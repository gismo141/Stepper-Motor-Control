// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VFj7292BCuB15bckbBBWbHAPazMdalEFRsQ4JN9ZvnZpP8+KZQu3aAg1CUiQMFfaRs2Bc4VjKjrV
2o7oATgdX06oVZR7DluCcFrGLHCKINGMvgShG9UUiwN1MvgcVIZE8Afzmh20mfvyzIJDUZhWwjDQ
lq8uKq4bCQ4WEKXwWv2T478iUNukkD6GcSAhri96jiVhxBI1gnZE/N/OfQ+mY2yWBnl2mjQgq9J1
0hHqZUaPsWOOJzeKFr0Ymmk0Kuc3mVWjS2bC1KAIXzHJWQZD1R2f86szeDKTjA4ogIMYOCcxGe2b
VYXEO9BomcAtrJ+8767GpaYjYBg0zji6r3VOxQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
3VLiCRKpnpHzEwE8YPZFxsnFZ9WRSpwIQFZOsI5q4q+Z4sXtIiXIFiGXM836ZCoui4OVJJ4xE5Bt
uFH8JDFCTxDgJ/2hlxJqW3J+19TJjrdxY4a1YBtqvezY0B+4HPfOPAE1am0Bh9k31egN5C1CgWjk
xWjlvPiFfZu8/Q+DY8Y6BPnfN+1vIAXEjHoSlrm0t6Bhi/p2hRky/Fp2+F355IEg98EKv0F7HJ5Y
pCxZm3hJVXCZ3qNSkiwbc8aKF48m4w2N0Cfw4YhO6Iv3L8C5hb1UPCBiyFVHG01rvtUF5Zg8nImO
VPP8pFOpXYI+hC8DDlTR5kDucQXZEWKHEWXgtCj7OKptDiCpyFS5ldcFsEeNkYouSA/Rp27Aw4/0
6xQdhvurEMLlzR8GEnHPJpwKlqOX1sq62TJQU6v/EcN/5ipo+1m5mehB9jrDuQyhh4udDzv75eex
FPnFeR6/yKPJ5TprVgdFrgOKq7QLoWScnbbFwXQtThOp+5tW8uKijxbW70bvrvJKergCOSVsf8m8
5NvY5Tj9iCl1ur1yyY/+psxTzdI/jeVbqE8BkzrmvuAl4pmEuNNXYZXmYm1kWhaUiLOGFRsBjbSb
R+xN2XiqhO738mrgpWkEZngrpng0hIFIt+liidDRkQfY1olle5afDl6VddiQjDGsPcad4MGJLVD+
6I5XVtN2QhQhrblLPU/yPPwfJ9AA2kFQWRVUwKiYBkjDuUCX7IhBTiGa8UW/oMZZu4B/73twXJF7
kVDPDADQv9ImBENTjTCUD23wqeFb2IY1sAPnoyHjuuhqPcNXbhREnlbA7FaAjvgMIpJccYlmY1Nm
sGz3vBLzbGwTMsdTpuILsUlzd7WWV4HQJyklzWIdAtWll33rJtpxagZMq+jKyKiPoMJgJOXvCZv5
6AB+8/wxnwoJQc0foMLSyeD815Zoz+jisP5/gSd5AWbFf3flfQ7o1wieF+nlt1VeAvCOHAg/Omk7
laDe6KqCPftjhT4CVjvbSvUeywFKaNwHXDpMNYDzcVS6ZKJoT5TshEyb1VETC7xh8+cBcs8Vfurg
72GQipd4V7bfhCO7V2jCLFJBEr5QCM1paa5uZCAQGWnBZ4HUeedVvdkBB7jT+rv4JYnH/7Wqp+HT
ifA0d242Ouo4GWvPi7l0smRTvGXJuFYrZjr4jX38Vmd5CD1DK7AiGxYyBpUyr0EMRhPi6rMO2pN4
rOeETmsT49+rJL0rqjME8OnjsBvb5sVk32HkXtMq8nRQpHwFgxYfrwgc1z1PKbV/NNCBa0JaHnni
GHpOT4qUEwgKXrL3x5UZoeSPeZmnxk3HOQe5u6SCRANeZnXH3/ZrDVhK2HvJ7HnzRmlSAKXyoHVv
FNItOAeWjUSOiror3k/ft368AcnLFBUz0X07KIh0tO4nWXQxOVn84VYrySmeyyb97RSMi0LsUy9p
XYvNF3VFDJiz4dWm/ACdrNLZGfGWfVgD4EdXyBg3sV3zGx46jNkASX6ihGU3RHt94cWpLsqdIvIt
zF1GuJ9h5R1LbNk5kzdH1Lg9CX3tHP41Ib6R4IyTW/ol4bspw+Dic1/TtTrFwiG6hpzRqDV4Tr7J
8ZPmLuP61MPhXuc5Iga5luE5Q72LTfuJ10ucINLY/iPdElxze3lCQAn+ytUtRMmUGlpTcO1ojKYL
DeGOagb+vwBcXb36RikM6wx2dWExmdweLFpnRQoRilomSG31+W4sTEXBE1h9qdDIxwy6/sC/Dn+L
cAT7dA5EuYFfxa7KeCIjKQhly4pxVPVgiUzBy7iKBnWAhk9naNOv/obMlDMN27ZCVcT9H/HaCmpX
HqrSBmmWohiWviL0fh9AvAu2sFF/GT2OVZ6UZpGVJPhQCN6g1qDojp/F8U/QsrUderedL231UO9R
kWgAiVzNjkKQ2z8IkNm9DKZPUYDym09do8OW8R9ZV55j/4IqGElhHjXy4t+1WLa8l9tRcvq695/U
hh/RB3hbFCkKWOEwhUzHb/N52a/UvTl4KnLgK8m42a6NYHmG9bBmwUysGg6JYZT7j6NQhqiWcaJ4
O6gkcjGZwfKLp8uUIGshdP9dFgQj0ihfark8n12VfKgdBNitUjE8LoA39/3Wks89Q5G1fVKiCsy8
XLS5oaFJdtgOpU5kifHZqO/n0JBCdm8wKfLUQLkOiNyfYPmQ+Oawf92bCTzxPFcyZbyILuSy9/gB
jX/i/OsgrF2ge9whDgFpvlweptuA50Ct8PEnHoBEiHSek42VnxgV3HbvysUW9VYCqnAILCoUeEGc
OCiM8ZoDdPPt2OZPzrx5AkxCkEaL8+m8D3cQPBM5JP5ais8H0dmPvNnp3AMX4qL0sKGphYaZqaky
8hb0Lx5I/bgUhj70iKetTbIOUelIRLyvk8NUHOJrKXxkNjPpl+l4h8/6UlKARv4GC3lnnU4mcq0h
FssxhCT/fxIf21fOelRfrfTmpwZM3QHLU3QMh7IPvbjbSMC9UBSjRTmZNx/xVP8oZGDK5WBIQGc+
f5fYmGi1/AwwdYj2IttTKLhEapDYLNzpaLxIJy72M2+tLVqAvELLeB5xfjLUNWyBJFiUnTLLI/u1
d40No2EP4L9gNN2z4z6M6WHWjP98yjoooqxU6A3gwpNBfQNPl84m8DsJxTV/MeUuqf8hj/STf3/s
4neDQvnrF+6MXAeu8J7dSycNdDhRwtZu3gWWdjHsWFyq/iOZHAxALbFAlyX8JDdXwfVNafuMK1xe
k6P6jPDQsC8J+Yb+AJDuPZYg50L1TkL/h/n5hC0AsZCUZmuQRmIw9+UBCyAjFOfL2z2PFk3mQF8O
K0VAwz1I+0oIAwMdVr/iDikSJ6Jer/4XxQIR+Xk45AdozRDAAYchzFngcQijnq+jdFnGWfwDMJra
TYnwnIPS2stEuxiSUY6YKbonJz2yKlVYVhuilJlBYG7NVYx1XyHQqbm4cDWv0FQetIbROgJJ6Vjp
XQlJc4c1OdsQsiQGjMtvBSybxjMl9gud0VpHiyhejJujRXN2xbAVOAFnuNoPIpcXkH7AUTZPoO7s
Hth8fdefQzLvmqusK4oMfC1ORc6cybsN2MDUV+uJvcbqqieg6NsDW1rVK4/aTWZ+SgqcTyEdtMJc
AnK0ltWsVyYu3McRf/yy7rw97NVv13MUZTcpLruniWn5XC4c4TRw9eL221UNT/eAF4rOQA/tFiqs
ImsPcTk4GyVm97LrSZ3SMiLOeUGpw9Wbkj2R4F2KWJh1ZtOjzgLHxHE2k9dAk2ZiUapAxTRtX/I0
i2mQUuXPXYSHM2oA8c1c2XCH3NsfwL5ccS1J5D0xb64o89D7NeYkejDf87KeHT6ay05fTlk8ltj8
uiaFpDHqMzQh6dsNQZt60RDFmAbN9HeKiWHyAP4bAa4aUCo876ilow2JBd0yOfVOGEUyAV+7odA4
j/fYAuLI4GyZWrKsu/XY12d9agjxp4iia5bSVtonAA0N+cdbGhr7aFZraiz8JhtZPzSDfKnEMPiT
N2CRQ5TuxruF2CrNJmGuNycaM+6PdaavMrD6nOlzxIPdgfl31dTNiE7cvgEBbgu973jIiQsvQMOR
acBYqmjJdeseZzaSCE3bklnxeyiFVjp4AS0X2G1NpZKfbRbd3NHg2DIaVFdCiRxn16gbMM8rfvHn
W6OK7u7PR+QOu6qjDMaykRqpufNvviGvhZZSam7rdPAsIbi3r/N3ED4nmoPJWatJsyQuNs9DvI2v
UY88K8npAhAULqGgtdf6cMw/Qypd1ErySDAy7TQgZj569W23cWM4CqA+b76pV8vt4jfYgl6pnNvX
NotEHIufay/N7dkXqD8sdYucrXug/zpNXlVcS2pDcagseoirBMNKdh/TiYsad4JgPoE6FO4bdgHL
xzwghq80ri3h6GWrdiMq0xYXzLagVdbTDztgkLzuMYLEdP+2E4rY/1NhUVg2JgwgRtWWZHWCNRgP
FoXRUq54nC6LGr5/UVLmOioHKbOdRZ+Eb0rk6x/e1jFUo5FtZLbRmB6o+w/SqQCmBU+rlPpjXMYw
Npg1NK43ECaZrdFcs8w7K+aHd8hgMcVD3J6XIDfux/5F9P7dhHsOUnqrM/6KUEvYK8OWveBTvqKw
kFTOQY2mKz0+ltwXTgrSus+xv6XsJlilukvCFsrkOiqgphfoc9/yz+z4FRjL02SJpIGVW/4+2E/i
r1MGRqklEXDkCUOAsL2f/Rxlwu6btPe36+tX4FaibSrOc0bQOFh3vxmVqdbn2Mkfs7Y7VOWFaISZ
dOtG0iXeOLDW8qRa1+Q5hpcIjsjMvzQMedA8OQAl01wH7WUBYQQvc1eCENaSUUZSmIeutRLwnMD9
puS+GAqkPIP4yPA+0G5JORhwT5mYC+PvODPDDTW4uXbpI62+V1jyx9uNUHkKeePhomREco9UC3WQ
BYV3y9G2eqxvuZAKYCCHSzZf+RuzvRPZlUIEyBk6Vcvx2tcli42vLqVucd+ZYSOcD9ci8r9RtF0R
L/qZDiJ87X34Tdil+T6PU6IKG6LRQq0WzpQ9qfm0FekGuAsuhbccAoMEin8xtfuedYhqoCUDUZZP
lZMc+g0429BdYZg61W1IkpfSv05zgaZrV0Zj6D6CZXCQO4C8n3pONzU47CruNnuKQkTO3dMmIZn6
C1u7uObQEEhV/aB2MP28YPTY9l/S3FB5LfusuuQD3UWPNXBK4EZSbtDzZmjv1hC7M7Ebz82Xkj3R
qf8I2IDBgjj80Yb3pfJ31KQQkBypg1kpZQ4GbET8KPPLm/RmIrIzVpIb7z6Ge8xXWcrPt6rhtUPF
+VOnAp23HB0KA1PGW0qwYF9/t+yu/uESjHjUTO9ZwHSpyvtGOzTJHtlL781F5PWQtBmiTJOieENv
6tqiWGKRtsNlkNfWWmHsD5LcnRHmcc5v/niGhv+Tzx4q+aQlEhcs2E4/T8Xw7vIZ4hPaRfRxH3Ir
8rMe2WdS3YwmGRnapk07BeGyHMowQRqSRLm4j97gRWeGg11eRr9gU5MNymFjmOqZ4isChQJiZL09
ADelLPVW2s9yN7cNtpq0w0MloLOA6o1ujp+/cZZw84Ne+KY4UzhdklNi8Hhtc5nHMeTXwAmYzbeL
UFdXvaRKqIn5+rCqe2zpL7Lhq68ApIhz1onf5RZX2crJAtUCsDLH61rcURgNjLZzk+8GEzijOI+H
7UOsqvdFgoR26PFWWEXkBZ8R5nbcFAdcACspAyxucJD3hcR28ASepwoMXyxdsIISfITLwXIoYcmG
tY3zOtMF/nqreRK0iwIjaIDk5nfR7x9JnQCkCXpwC6kqNoWlvrMye/GGITYCpoE7d9uWwg8YrvZy
ZY3S/LAJP+yGipo0zFE1Wr8eVV7zCwNw98y7AyuUJPU1zV2B2HsIX5tfc0zaynGAx1XsfIe+xIyq
N46AGRm1ywEvxgzG7jGpfC3Rd7UfOO0foOw3bBbXu+dD2R9aCAYIcLrdfRl5MjslIlzqkZ55koUc
pImJN/glIO9xQefxJ1ik6Lke/SzRUqhwEINOdiSXVsDTjycY3yJgu5gq8N54cmtrPT/38SoA2kmA
jhmtvQ3kbUnPDDcsq3JMErjG33ntg4VFFj507XWB9zLSSPuCPbpzoVSB1qPAAfnFXiT309psa9Qr
046D0QxgIRSFA6ZP1dlZ6NLp95NPwb1UScirzWE8rpZOasgO0pKKNq/be6USMVmzqB1lGnPUCrua
VUKjXl/sUC9pm/XS7ylgGg+Wg0iITjhScsdrulCpkNpStuQzxUxEC6h0pFaKJCgI/YO4q1K4s014
2fDi0gSG58DMufai+0ao01Do8Q8fsBo0upjaqXXxbjUkafk8b0N1BL93JVlBy2etwcAyHIMuLaWG
6bVE2tObiQ7MOztGoKzwiYT4PomW18aZdSa5weGoPhMpqqovmcvjt9hyLnUyrS1UAb2yEhwhHGUU
DnBcTyy7VsP5lPO33MyI+SZYEOKPxF9hYAPH9FC0ghndcps1lILDZUsF0ov+tGStkuEgovXcFb8A
9vzzx05xjs6ILYO6ZSacq6MfYQNGz+UMJOqRPANLaImhtQCI9QCoqnBEuJsH+PJxwezvM+mjQGrt
AKXYRFvB3QQQvumw6AetW/9qI4GyPjaYORAxxLMerfwdi+UYwjydMoFspr7KOvNSonlXmO0Zq8wJ
G3PZq5/+r3AUC67y0TN5bSoXZpKnmX2F+8EQqz5Zfoj6rZFH34K47EwwXIRl+9u4kr6taKaZlf8s
0ItL5D9oyNdCZ70oguD2UJ73OzZLGxuTIio3BXnXRi2pxZ02kylNWur+tWHQHwKnuVFvxFtY1Jsc
p9QdVzz7+3G2BtD0gWjbpPrVzAFh/iExDwK5e46lQFin+iUlTg92O+OwYaG4bcrJiogPxr2Dqonb
kC6FIDffPnjpUqN1FbCTXw/uvEqKna5G0S2Cpz+58p4WprHJKW4Cp93oI3gVCe//Vfmlp2Tymg61
zZBkLYjpBL+DxW9aUlxj1aVFVS+/DydIMArECfVw7YIg3fxVZadCD3R169ryypqwA0M8CuPZMK9O
v72bPvnlqazL+8lTaGbIQs5ZwpFuXBaV98bH9PsX62kPU/f0AYo17cuQEBvddxDhoXYK4t+6rsLD
Viq/NgrIgeF/M9EpaMlNKqFGlVIn+cxLO9BvVff7vrwBm2sQF+qLGTI7QTO8S5zIuWqSwZBXyyt+
hhHbftAoNAVbTD8nZ5psgkUFM3gqDrg93Jjyxkuck6XdOcMuWaSGZCMMSfZfBiHiobtgyPruEAxD
5bdqRc/rAGIGdmeG6QPQoRFICkqIz4rPOCHST9oobkBuPQYLrhYQFrR7yHCmDuuEG/KuCU8vEmpv
RC2PrAGC1I7wO11uXsGld1jTmLP4yXR6nBWS2vR2tC630epmA1euIuQnW/a0xht5Hzb5Oz/o8WN0
MBL4B/POai5OVO+0SPh9A3Ym3G2azn+H5KTL7Lt29nCzk0gYcJEehFofNpjPR7GVthlT2nZjCEp6
PJFhKJ9y8y4rozeBmLWjfD3+oYlqs5W4yeuoJCN9oC0+lwlwZ1sefhvBhKsY0W9Wra7mYK6DF+NI
oYZN+V9J7NlvfQHUgQ8DAJVTYyfketjW967mLukDRlFzXpC9OPEejoPuXX75CVwhEfYa/pJz9msf
+zIs1YBkM6/ByErxmS81hOEr9JVkfD1bstYy9XiQxmOK5tkzeeS2yG7GDb64xsRHfYto3IICNSk/
ya4ms+r0DrEzWeOvU4fB3XCWGCcIjicOxFCbeiTb8GMbR9SRn2D8izhRR6pcDk3HgPMwsMunLw7j
XgwWomL2oZcjRY9DzUVlObOFOw2qbdf0OEN5Qf2eqo2to5pqkuTIb7vQi7BReUAh8K3iYZoBAQCJ
HOzqG2GhPro7WLbL2FyMRs84RorK288MhV2pO1SFpd+265i6ygHGWp6lTgIMqW//8j8l3uA0+EJu
JsBfYJVWo+TiWR2/2gRl3O48Vh036LPjqKHWZNnhgJB62NW2LklajOd2MvzxgUnqTwBU0F1W0UW5
7VQmc6Dv3luV7YZJOnaEqYvc3+3ZEZ3vy6DALQUdX81cNHtInpmlr8SCfIUI+v/VoKAiCmhyPB5z
LSX+iyM8x1fmIx8uxEHpfYACFWr9QeiF597LJSR6yf9DYaCrCskjX2XaY5OlbCq7oh+ZyxHmRbaI
08NViZfanTYX99ZnoZ/R4eEbQ7rzD7rGW8CW7vGuQo4mS4xXycwR6BKuVtE28dcnf4qlNSO56sia
U9o+J+yA9lhBa8LQyeUnOgVqDWI++XMnDX3Z/lWCa7mN6PsLsm273ranCo/0zLb0zT2PMKKh0UGU
GLyu8d9Zch83hMYGDL63PbbczrSd+iaXmGR9TeS5ZFBy2QsFEj6HV/+HRVFvn6k9h6Wy3q8YCLNm
I/aTm+lU48+U0bHzRvk6jmmZzLj2fm+VWNlYoSKU+ElEIz+7huTZaqlfEhgI1eJt76KiXtnl/OSW
84BT1x6kJww/V4+vEthuhOeGtrC29f2jUjw6luIrU1ZFTEGWc5fm0dcPuXhrKuFSvvt8ncbQ80f2
2yAAumhA24z5UVXyFdhbIJ4S3F6gTpQ5HWw43/nX8BNByEYbdWowNFWZjucfTwCFAXMsJNDfNyNI
Oh8zS+XGCj9wcKgL5fEIbVcdOiwLhtVKl2BHwZWRZd5Vb4qtBuFXc4Mf/YZYk9AloZjACj7L49SX
8BQSanyKSym2mEYNajWeqXNSG/F1NY4+xwBeacZVKpualHHuuesSAXsa6iYLjPkXA7JUH7hGNTlm
4IjkbQgI2VHEP1IK0kBq7sqJMl9h8Y0fs2DMAblbAbVD3b73k+FaQQ6AvY9O2jrB5rqp7XSly3p/
wb19Le8oB2mzvpaDv24T49YGs9pVsUoO3YYAPY2icLwLpmC/in7d4liIuHCmAdhB0xmvJA5EIzFn
cBegqnSDFOxc7BfiB+fvEcEc6TZ9gpUyJXgVrEv99Wi5TrR+bujF0BSwr/tXvwiuHyhP/ypxYpjB
hOjJzOUIE7Ih8nZH+YBiqST4BPvYDsgtFiaXnEnMpF6uFN9MRJtF+cDPpDPHSia+5JrUqoY8v6bl
2xXmbq/WeELTHfKqrDWFuq5eywca9VfbL2wZKZWrRpN/TTFu+Hs6sxQS1Si4H0VHYIh9s3jE1mVC
Mupozk7ZBg/u/KFgNhc9qEWitb1f7QLdzls++2dKZZYE2aYWvTGRKFFEx2JtKD+odrUPQiptn72y
Xijghoigfmml3vKSPo8FI1OzAwkWQxO3mz0TTgliSYPlyFNPjA6CXRCobGLXcVV2lM4dRok9K3lI
sqkE4nWrcn7Q9lV1i/EIvmn8pEwzjSV1CVNQicVdTozdxMnSCvNvwJxdBkuAcciV+C0B5EKD4q8I
NqgWWjyFbM8+Mj2021SxwMBkRtXvhXxSZpeudbyNRapMNjUbcTqSvFCESNyZAjNQAnjaF5nlbFGU
YwZalqJQ6+p8GjlA88L+VAYHobpYYuodHZUydi+AU3s1yurnVt132/nmnOl/8UOlq+4U4Pz1KkI4
f/CArLQcHmbWyFGkXjfiUDngxLEKc74RhWaXnPPCK5mnKyDAM4daF1k3OKPBkwX6iVe9EA1BPwNW
GwlTAWl8crh0YLSghQMEj2ZcsvsfSW6jAoVWSirX4X4CzgJnoOi5BR4LlnLtfdlt9xGT3B08i4l7
d9XER3L+AJe9oWVtQYKAKoKRH+uejYkHDjoEq4bosQ9B36sguMoT535p/pvWweyDWSsgq9mVv6DM
F1+9mvPdLXKFU5s9apptKNtMoin8veyLpmCHOvVD89vX7kwJjnx16T+OeU/sHVACQoXweUJ1gnSh
dEHH0MDLK5YSHyJSdDHhl1zfuP3L7RhcilagjTh5SiCrZNaIwKE/dbHT/nZTT5OJX3laANXaRSTD
TtfcekjYcRU2WD+jktJPlGVB5lfcv5MeH4v1f44Zn8Tx0GHIiabqpibPSMqvzwci2TgqWESPk213
G7g45uOXPAZWmZcMToyn3ValoQrK+6I/PCUd2tBJYeMyv+Qa6ERMXDZKVFkW99u5ztsA4Er0tpDg
yIMXj9WquqvsQLC49Q9168dlLH1t3KIgB3Kzx9fPKLaiRClxwWxUl75XzSwtsjqOTLcw9azmWN/N
PhNnEd4u+VMIHUdl22W1IwFX2G0yaMUdbPISKLdAE9zXz20iJTinzcM014Tu1bc/QdquTEKGF68H
MsKFBiuNJ7wXHeZILqIQcZ30avGfmWZKkoTx36g2IAEvqlKlj/g3k+TSes3CJZh8HYecUvbGlwcw
ozUF0LePNLRjEEXa77og4Qgl9jFlt+d15OGZgHKJZdZj2mC4Y7TvH+MDp2tPeBZ11J02f1a/YFaq
+fzC8+FtKOGC/nfeiJUYB+z4/47R6O7mlz2/ZgNltO2deAhkG1vy/HreibH8bjBcSRaY7nF0L/uT
wkCw1BF8fLI16WP/xv5CkzQ1YCUq0lFWBEohkdMGGr4tP7MolW+RCw3SaihoWfRBtKsLwXfGL2E4
gtUJwxylun6CKBR2CDe6nvZ/lA/6C2CmNYjwkNASz2QC61Z2St/NbiBOoloDb5R7p96e1QnR0GMB
kYEc/WP0jqEPvH+0auppWDIzKyhkn8j/Ncw0cMaVsspPhqkA9yx1DzD5GBzjNuhj33a/weyTytXb
JEORqcr097T4oCiEQUxH5AfIXLfTcGvL/UQ7x+HqxXJr/HKZi5vsfwmjoJjra7LuYzRZuyz/c3Yj
XZF/bqtcaMdif7BZswiPjpplUrl6WfiExchXXOmUVxsGhg4hA0PZqDPAM7VHgpa6EwMkliazbmYw
ZmRTTVpHJ5tGqQ4KLL5IycjdJWarQmUpXBG46snpbWBSf3bbdOvecbq5YDs4GOedt58lyq68FlkV
T08PFWJqmCb5czdFF+fm8TqP7+JlHvQHUfbDysUKKJNvUBt5qbLZPLCsrIItPPci1twNn0t2Grr4
5vm7Av9Juhwjd3nyF54GUlUD4GriauDWQxGgf04z4OpVxGsbSTbw9xLigXR/ROi9Ke+Wb1Y74PYB
zPrlAMAqi90+bNs1AsDwq5jE6Gu276dHFhYUQW4SsKjqVEmuDEAhJKGau4YNAeLaZn1mypdQuAta
IIQ3lS4W9lrdbj15E1FI+f1w7mRyAQzs4lHLEIp3eLnGnQi0BUmu75lV8j2MmbAGNG+ZVbahq72a
PrO9Iv+oB7yYpxYcJF523fKYYuCpO4XI129gxJNtMTgwSlbAx1RqpOZBSLSlPzz84Gxg+lu0itZe
5fWYlyurGNuRP3gBebld414tur3zyAxU1rhkWcfUykFcgFOoJH7WPiX6Wrdj7q8U0f6DjlU859EM
4hVDxY7NnvgXH3zzliQwJtkEmk8PtWOjoS2CfkL3wAKoQ98nqybQIbnAPbpUmGeSfJ7XcNM938WP
9rbL8jMXpRrpdzWNk2eviVLepw4PLrxFpzpUPgSphVPdVnVk+BdXlJyNPX50qGYf/+aP9jpEzFA2
D0DwyZvohKYIjBS/oopHMeJiPl3GeJ0cLzlZX3SBAGOu0uZbo5IO/HnfiCVECtqfxBc8hARfinY8
P/glk5El+O6amQ6wHSsy9CjezUqmoD2GjohkezbhZbdnf/nHNRUjsBjsU7qBzJUC3qyhsIWboz85
p6VEqdrD+ncRm44tHeHr3xI0E7jy0SC8qyPkE35lyyFx5lawQS72Bk1JOFPSwnt8+qlw4IjjkTjB
apWj1O7rTDB7V8TcYlBfCYoZ3/Sk7hP9rs2+0m6mavbv/0XBCd+t/SdQIuizIEcPtYvGwVMNge/f
ZBAenZAhzIqBPtoSOrdPKnpH1X8kQrCJGpwGaPiWfc9dAoFuCqaUA0XI//hHFJmslMWUkflxnZcd
Old6tlBThbPmxsY/GyNnFREAqBW0B2EyhK9yTazoI/tXDI+3g6bAulhB0L769hdaaAwWETZpMvER
6u15+IbSEwvCIiyfSnjxOKp0k6WzYPt5T2MpRBXXoHs75vt0eHZNFvSEQa6wGwnRjWMlA/v2A6C9
lFOKVZ782PvUYhJuua+qIyCRwtGbhHeWC1Oiuwc+8WTLGqBSZubS1OYHUqlhozAQvxOMJVOB9peO
Ne0/ESOLbrMsXBQO4C4a3SWMMrZ/bBJY6KAmEHcczPY1HAoSFm0rAf6Ybf3pyApy75ATL/ldU+/U
45vUX6KpWorVVyDTkB1MI+WjF7qDgJTneiSVD8MyRLYcX7ccK2VU/qRHITzcvfPK0vqCtMQf08IO
ldigqufbJkn3MDt6fyqJvMy+uyUNDaIf6ukGiE9IqKooOlf7A/acKPzCTPRk9MChl4opgnql26dK
9Gv9EaXmT/Q61oXFoJD+CrqiocHQ7m2X442GMklvuCqS8KvfgvZN5dbZg1fbRDC9ZsJH2NCeBQwI
PKRDVOHBRVXdL4zN4PElDiE8fsWo8gs6dOkXEi+hxphji/U1MUxbS+NiAHxqK4TKV1ogVLBGB0LR
oXOdhMqGAtmzOkM/q5ev1Rg5iTzXmoNGc45CUFmjwafCSTu5IRvvc7Kd++5KCxwALiTTy/lJHput
suD5KytphrTY7bbPiWXA0csfrD/Tdqh8GbgxtMeBP7egwAbr+LuGjwsmOiigT7O2jAPtRj+aLF1V
cENiO58mIWKjMOw+ctclQMWHUJqiSH9Hsxy5BjJ/heWtKkRLnxilMUW3+Jd/9v2xDyzr/BhONIoB
buUQT28FfdXQ95Sf4aUTYweNMT17XN/8gC2+oq/8Fpd4MovL1rFPzio1/UT7bWDqGdwuyqxwz7GC
HklGaQ5a2yqwy8j5rnJHnvVeKNGOp5LaqpQxF0e0CfyuiOzvWQIJmG0D01mJKAd/EU/qZfvomESN
b4qL4hc8zzPSofw3j2BGTiyJUKsmQ4B5DqxWOJV1l+Q2wx/bGkaoImjtOdwID7x+F4dLVvKf8Rnl
WGIrXH55JQrLvQGSUZYAjxFoJ2R2BF9WK1ITe+AGSOcbtBXhRQUmBV1FVhoB+1Dhx3/BLMCFXDP2
pRQ+m/JpIUSmjD3Tev9cx5fQfKRy/TeBLXeZRUBCY+VfMHcJgz93kda9/EMyrc4SdLU9h/tB5Ezt
fZ6UfO7gReIWCiD+OZDrSk+DmOXrJ2KzOCKXxe+u1EmShm1shTjaFnGAdzCho9w3jPCtcCSq1cMM
o7Tha7dpsXRnlortydy60E4lHLrATVToQj88VglGBTQtpmUYcvMxC/ZRSw5Alpd1XHX5/SLBIzzv
lrDEDja321vGZJoYJxYewxoHx9FsPEO3H4sPyFkD8U9mawV7jneM4s6rnKpqP0YU+X0ZroEYCJgI
sFzRY3s9nyf2sNWV0WxEvei5wyGu8puynWY/ryg+msSs7Q06w9gOMea7TPcJsH7hRR3J5kX2SHKb
AJx0WhMNQm5tq4cC0YwiLhXqcHKuzZxAgQDXC/Lc+XS0x1BFk7M21E8YUi1IReUDqto4Vr8FtumR
iOjdF7LPXu7RQuMZiXjDdrtEPFtQxCyolmYGfrsJYv/aishmrXVszu4ruluiDbUdeD2947i+unBR
CxMQBoj4GOQw3u7UrUrOECP0LGHpI9oYrQw/rxdDwyMAqGo+O76qOxpZc2aagodBDLPtwrOV1smj
A85ya3j49nOMOrnvdzMbeWvhCcP/9q7fJ5/kYRK12ieLfiyqio6esY8isr2U3gDm52sWZM7nZjW2
8JWDQD/JEgxkGcGPQudU9f2FyVxvFdwjB9E28RCi/gXoSKps1cyPbWdNOhKkizkIHzORlasE2+7U
iizMlwkyvx95x4QUGD+6M1k8+gG/+XWAPBjRL5cHyF7OZp9jEa3Oz44PEQHFTL1xGPfjLHc+Hl9X
dLAOdpMAxtGbbCEeJEJxWpQeGb2Yxno1Utvz5evlHM0hsTZT7nE6kChIVYWa6kTcl470jqH+AsVe
BkRd0we31CEoCG+1nnvQs71fevgmLGtYAjLfXjqb1fXcXAPm3XOYwuTlBVw0SiX4LVNbarM+FVXJ
fO4W0cGClOZXBXUrKJGRUWKeNDLPC1x6jyR6TVgnImopG8sE8DhwwByO2AZcFAV07nogibRKlFXQ
sPWpnbHp9o6giH9Vz2Y14i7NEDqx1N8v+ayl+Au96zU3p+IEJaHkxuWcD6BCp0h5f4FTr1urQ2GL
B95ektW01h1xEu1Yo5ncjgCfahxC79MBJ1WQwdQCGjGiYLAipbWFKLPPqOEUuuPSetU82n6iajbT
7r3VhOv+b1bzu8l1k095j4GNTTe0nZWZ0pUno5Wxx1Xor7dTUDd+Zftia/FUhHl5+aJmLSMNgw/E
/BlHtOCQJgC8vvFDzywfp3u0mH09tw+EgBZ1fh2vg7iljGUNF9caRFvYni/vMDt+cTEBZgEdvGj+
TENhlYJR+C8MbDtWaLVrAVwvfRDPFNpAmRZZNDzgFTYSuqfehuJAe1Jpdc62oIu/SeT6HwdxZ4OD
/xZPMZQ/m1DtkmT4bX2HGlq/5AyNV5meu/ja5jOQl8Wix4jh5lTCVbQ4MsAuAN2FjK5K6FxfbY5/
N7xVGXU+93MkKg/wMP5iIb0ruIsubp+BIbl+L37dsLy5sUBgJrAFLdyJXLNWUcW0zzLq2jLk3+NA
Zo+w0EQFlnw/hQHitDAgIoJe/fBHTviYfs1hve9xoU5A9ljlhrvHIVBXXvWdQLCuJpKbp3cDbbnP
BX7E/+PHmUJ3FS4Qg/gMmOYpKkmxPxJ9AfXpWYjaxJxOXVUgUDn7t5FyUpMmBnTeC15PCIPiK0zF
+I+Ez0DxZjv28hy3D3cISx2c9P72pB5tzTF9oIKLNud/Wjs9GeWMGV0A7kgxpa+23DI1krtILf3/
flAfJbmzi0feTc5FGYEi5AUnMOp4BAgCSaUBtPeO4os4EA42/nGcOyNDvm/HmXkWIVEQ6jdT+4FI
8RYxgLKry7+yVf7RAyEVOOtBXEqhxbnSF9LZVZHJfZNBM8nsJxIfBPl58tDi/BuGt0FhyNqQwBMe
SgyyLNCikIiD7EXHLrlLgsf9j2frXGs/twaJV13pOScRodfOdo3mNwFDTZ/LOVTKL0AZySAdOGc2
2yqtDdMMrRJkylDVu/+v0MtgnEprVF/djtq4lz8gLMDP3lh72L9+BfGQUXzNqFdmrK7o41exAvDs
crES+WVkY+bpEpn3fjCxV80Q/dlOjokzpoe/3zvEqSKJlOJRt7RhfrADXlJiHyq2qPek1t+CqBBi
NmeuECG+DxVm77lwDerlfGR3x8DNYRxppB1+Y8ACeiEbjgD+GkwGl71aJoR6Wl8pnhVcZUSKt/FH
OVfuEgy/+2Z7bCJ70JmUp3AGSXq61EoOn0CQ+Ip6nX76oChRkDQxaWVq+uz0pI3XxOXVay3TdVUf
vGNfC3ebkHFlQWoK9ADhapqSprKJ5M9uqnniWuC8dzYQ2oQUzoYK3DDy67Rc/uoZtjB2ObxHVERC
m0PlhpHwZoaabrzUJVvdz86ra2SsmWHqVjG8Tl9E7QXuUk0bsEzuoQUNM2HakDOPz+oDjX5cVyFG
B4rA/u5R/dWsQcxEecYh8hiZtxDuW1QHXa510SwzDDtnmKaEOCSOrzRx7x/pb4YiSRlU8uCkJfHr
5wXHjJgYQler1rWKH9zb4ZRrnMD8R0vbauHlxRvdWSJ1+g/t5XV4iNWNgFQfkYjl/phi8Wxfy54W
UAnhIFWKfWzpHraRyJjIm+xyd1ZTqBBqUKz8PIAsIpLxG//6y0qH4LFasUhTAajcyPYBZ1sxuuK2
4MXhxeVTj1LRyMS9aGf3PcwE9MWVdTRTz2FdaVD/xmStv4/WeG9Bvlxm3+0K2pvATrBNWUGIlox+
MeEbzL/PL/Gr5V4U09z5NqwVWRIdWkuIUzPO+BwTW8YYTKzJyXv5zK5H0Bqnz/Vsw0kOy7R8807K
JiMCeu/cU55keeZVWClfKhZo6l0gWvxfxpoYyhxmxEOb2t/jNLLXshKGyIqVY72CGuP0vgPr6Z6c
3gwjSFsjsmIqCrDjwU9rClwXRNfhxuJcegnMbW9jM7HVjCqbSTSAevNR+ZwfsTwv+IHNGeo2LV+l
szbYh566r6I94M1OTPxQGIC3eAg8zT/RGGcJHx4v5XwhsCjBohYF61akGTuTuc27h5wyZga7lIlm
mocH2cK157jIN858AhmBAY/SDj8RsbkI0mkJZzemFtjOhXGGPzkq8CWYhOIGL0eymm634fyrZRGd
cwveOmmSE98NL22KHmWVv+QKckB7XosieBroUGgR4sEE1PchsMxJIpd+C8CgO0hy5cNwpm2WMARd
fe55OqsYgqPnzYrcLSy7LXybdYnN6TkU+SfbVthsGwq3oEAA1ABsOGE1ouswESgSokRpB6bxkFvO
RNLO5HiSt+se5Tkfuj3xMVNsAs+5FaAxdwdwAyniC5kjuToRa8OWctkldQV7mjIIE7l2TaQyaHu0
dK/XQ25ZEhZFFKN5qe/BOg1VhNg/Hh5KGh//r4jhij+9G4ab2/r5Z45hwqqAu9/rAld3lB2xj+0F
5WUv4m0rgHZavWpGVXHPYdr1bMJ6ss9rFiAsaCVQX8MLry9AQvk4TGjNgHfiFDiRkPPRzzpM5GJb
lyraSnZAw3KrWkIwxou4I7o1QE+1XID9wG+9/1ID4L021CRlAGqHfdgxRFlcCS/J8ioCbXidF9/3
/II0V9AwR4ASdAhu4HPVwv4xa7NXJ10k7Q03UBDk+q6Ns1XGLzz4q6OPj0uwWfpo5zcKPJRsTLik
oZLjthvuCKofV1P+GvRaxlfw8pljt6Yypy+nN6VP5tHRVW9756r7mCpRr9IvOMXE4hUuoecHRptW
16S+Yxd6MXdyyFAhEM0o2dVa0hKetpdq+oMbniXSshqnAGzY9D2xWduKL1hZji5CdeNOKvzzrF+R
HjTaZqYCv0IhMfYWGfO1cTvwyN6w7qKkibvQQYzMNo9vyJMHN/uz4hv8cFIweyA/3an0/kW+Vwcy
jTFgsnyHQS9GhvonijtYrWZCiblwZhdmtDSHzrh2evCcexxz3GshcXV59FHag3O53Nlb1T5ncuuT
9I2W7MqPJipOHMYMW0O15RoSv7fwDovKY9oSV/RBtk5/hwUaepSaPW2hw17XMhF3qORZs5qq6mM7
8ooxD0fsy0J6CGLJDi4s5ofTAOKvMds/uI0RkRQw2u8dh2/kR/Ggju7a1BCWsHK0bxslx52Qyb3I
c5zGCdBPXLdiIQ8mRTmPm6wWTVgWi9l9G68oX2k9qI9fsSq9sfqaRcJv7ayLwK8jeVmACS3perR3
UvXCEoVC75Yca8+mEy7bPK2zkNzRZWKxjT28H8Gh4z6tia+XJaoYsTWQk98GDbmWfprTJhy2/Yc7
1LQ/JlMsBqyY/L/mZkOK5+l4qtZrvihnSaLS3qjMq9eksxBbOQTDsGiXoaCWTkEat1TKFQJ7QCpd
APWqZz5+Q7GxfyFNR7MQAAWoeCqVrqyKkiI+Sjy+zZu2K8NAmXc/vFQvatvge4yfvyMnmb5eMer5
xrQfqf6gGqnXd9g1B2P7HZ0iP8Kns56kbnv/nMjVJQEs+0QJnc4+K1YO+SJWy/GMs+fth7w9pzC+
0XoV0W35F945KTB3MRh7D2TRtMHJ6i0DqdjhiX/m559A47A4vWouUilRTl7BCLK7zbvKVNQTQOD5
9YsolO9LiA3Azo1HSAD/FKtgOj/4l1IDlZmduzadLjp0s6Wl+8yhFNpZ03WCW22tSZ0A+kMXhJj7
zCCmTExIIpuPms4rt+p5t7U02ilErcNXInVQkQBJapzsg51iEA72qaNEW4Zd72dLVE11HW+tovDu
kp/gaJdJ0RQF9NNQ6304T5YTJa0kYRKU0Tm03s7pCa485cFLlM5u7VamxsOVd/uOyoBEYHEKYXTp
/Xr11u85hNiZmDp1IOob2MaURrbGtxSUthVwHxoBgiPaVM3iAl/L3IGLOxwPAYb0TtirX9Aah4CN
zb0nVmD5ewaqOgCsjBPsosBEV+w/++/cdeGu+oL38ePtFedfhGCIG4hsvesPHEYdNUt6bupgiPvy
+LZ1fkuW4APBohdlPOf7Qw15G/zqhi+93mNXJHyerB4feOKlUQ30NG1kHd1LVyCgzujns0laBKJO
kSzzUnbfuyXxNGPnw5CDaiO+GtKN1KcjvLDLySNxp2efiEfivHLWc20N/JZdQnk0CQPwKK3bOxem
Qtbq50gAb3s88u143e3IWzJfnwOetz+xxhprCvzUUnOE9wQpyWDsFbZsVQJ7c6KuvA56Ec6EhO+t
1PntGU5BCKy0ykJTCVJyVi9Z/NlEbYH+X0PS9NLkiaYWmIHgw9OCIiqj/jq8CUnJCvG0pNqlubu8
q7MjuHZE7Td1DWEM2lgXYSMYqAuZL1YXVeVJSHp4Q4ozg72vyWzV2GLE9CaLIvq8TjToiZF1LI+n
krGZgERxAnIDU5qg7ZxC7eAUKa74orV8rUAK8kPWs7FjsUmlNp3aebnLv6rwhc0QNQUF4e+YxBvJ
oz40VrtTotUsOMaimyQbNoGh2j3DnL7GWF0qhwh8v+UQZZJ+SUVkV5vPeSDbaGqYSLq8pOBmmm+1
ERQ0G4i8YA5LQ17/vRguGzNZ3HQp/Y6X87Cv6qr1tnb7lrSKCzVlT1xWyePeECcTkbAxOyRlayrK
X5X2uHzkO/fRC2/2eO6uYqnGv498w2XHt+nzZjecpGlQGDrDXok04TPS80WX9lUKBImG107cBEok
f0ft0LzTW7BkMzL5zkKOHcYBoNZBu0SGR8qrilIjm8zwgSKqP6XG+nLx46u5td/UssDPbfUOOpZJ
/8k8cRHk6k9QPdGzm3/WN0shrRykfiY=
`pragma protect end_protected
