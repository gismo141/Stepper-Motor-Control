// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ngoa6zcPZCb4gV5zHMeHaJ0+TJCyR+HGrdJYtu6Ej9qCNs944gwiU52Lp/+sutDMiqCH9CnCSktQ
gaY648PPbicBqBccaXTeeKuhmOpVQJeJ7oxMETN/tt/5TlTMTPti64uaBxEawpar5R5SPEJ9UYna
VJYr1qwEceM4OGEpSuUrRtJjEIy3QW6WAE8nsH4ZQevEUdmtPJPRKICL1fuC3z+fHCWxBFT2bRV+
7CBX/Fe0on8xI84kdvy/nOk+16nm8XWB8AAE7+0Q4lGAfn4gOL1oV5+1WCfxfZZUATCKNBSj6ThP
dT/jmkBdOYIYkGNjPdfPBAUC3nDlmMXlpfxVWQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
jwSK3TfUkqkiU0EBrVNnURqLzIiZaYMLvW2x30gKotdN4WXfEvvuzN2os2ohavLNp+ZqVp1yDtb4
w0bw0Ekm9ekuBaElHLGGiG08U6YGYqnh6kkPecheFOXRqoAtV85N63zq2f53mu5yd/gWqVgzlUQa
bggMOqVFtJdInGlwyj14Wh09SNluCmrLsBLQiwaCYtDi/6nAe4MkI2LoFck5dW4dN3kVhBykPuWM
/a4uHrVGOMIN1aJo8O7l76DuoubmPrHvzYUBShqEhfQ8GEsMtfAgsAaec8rxRqlEOyt7smcickFN
iZU9/ecsZo/if93IbLRrK3aaNKDdGuOaEt3hUYk+XvvefCSmrRHNnAA7oYBDOeTh34dsZ1WZWNqI
58rVHi2ZEecFGHdVz4+sDUA/jv/B4IYiuF90U78Fc9wZXRS3r3vCenr/LoZPY4Bdpeo/r1CCAIOV
EEBdnUkuiaYglQPAy8qVBPl7gIHUT0k6UVTj/BS1o4l2WXaf0EAcpL8x0tZW8S8NTIe1H8lYE+8A
f8vPSLMVgaBH50kKLVvOEcptA4y+rYzq2lY4peKjdcCaEViSBrwsSaWuVN0AReDNlMUoWVKX3Py4
i5RT5OMFj/le1amIudJwk4k4CtdP5UPOt6LrY9ZBQOohm4OQkC7/ddlUdb1VMa4WXoyS+B5UkVxe
8nIKt1UJdXkzijB1DB4qDgrca1XhzId5dP/XLk9CHf0stdCasjG+aNR77kgcZHy1uJXK9mO7S82a
gzo+AC+YKU1gDhLj5Uc8HZfB+jgs82Jv0tH8Not0FLNAd/HfUf5bazrAiZWi5dTGDl3Pax2phkQz
N3TXagYmFypM7uycW+zbblXexoD/hGihDC3NXDT6E7QzoSprgeAQgrAUTsTkmOsYvMoiWROuAdY4
8yXRhTZ4jufRDyje6nNPal0roQcD5rBiEIVnfMfgNILEX3PqPt8Y/MyLon760THF4jG9/hPzcINw
vGIfG2NiIP9San67zOEnPhhuEcgj86ptdgdoMFtX0+lORarW+eaNu0Qv1ZC/OauTwZYK5u80H3gC
gSl9D/TrBaZodMPKG0tj8p6jFK6EG4GSnNarvVxNvrWfxfjl4iIYEpmUoHfeaU7sD4RvHtljfPDA
+fjeCSrSVcRU/pFZBY6ihn6oIQnEE02sf0ME6viwoNccabvRqczobDhtMpOanOpT3M3ejSTK4azF
f7adHnfSr3Rnah6jExCVDkw+bZLoaFhejkXmalbUXEOAbTtiTgr4QPtFDDcaiefpEJNm1TTwiMpv
6dZmkis3xpvH5s3CxENkCUMy9eKzmSXO/zbzLTEJ2rvjxs/wsaiatYT9L+UXOpPulSMeL/RQDk1A
ub3jP2ZTG/ZFkczyet571CzoouV/an2dmn+Aht5BviiJsxcq4ioDv47fxKQXnH8HmVBL8rywIo/7
0w5mwxXwJbSTziHPkL9yGnLL5iIk1ou4tcV0T9zVjcuwmqp8WLw/6CksSumpHfIx37dvetC8E8hk
XXxNbxhuKJ/uKeED22/L3POYOP4nous6rFXejec/72T6QN1ZMgZP9ToBxDYwHy0zutLqZKYFrNEr
0ni0+25xZUcMjBGOjZDBIHVFNHcYRU30kmpUArw55q5GyKNWC7nQ2kSPsDmpokpT8ofrLiykVYLQ
VUBpHpjmQK27iRth6uaOVuAmuZpHTr/i8n6fvHbQq3UzHHZnc08pUAwAG9WwZrB2b97y6fNxDlHy
21OfN069NoX+5lHOUAhvxez/AtopTh5+9RaJNVNNLhR5sZBCsV+XNkVgDdi5xrMCcOyqsX8xkgJe
pUVXz4amov70HNeewqdyz+eiGdP78cnNNLSLnxRAlzwk296Xlrt4Ea5IVKZDO8y83IofFpBNLvsR
KPdmih+w7t2cBwGLpME8Os+aS233Hu+1Jod+hAboCgWimeKgM2DTwIJqyDocF4QucziFBXOGcH2R
7o9w/8LortsjVsj2zDxSidZcNbK6zrc6VFB9Ic305k0uNFsMIqXpQwsJsNcT49N+cxTW2CHMOzmK
tcLye8sCyv1NBivB1TXIQcSjKHhJe61gKjRGgOM4RKm5Y+g5KEEdOLts4t+c03CfIrngXcyR3jAn
cQiR6ub8WFiXCNWMZf6EouT8aMuPDwYehYW5+WFKMsTMrlZ+AjoCJdp5cspTfM9kT2YB6Y7ZsH0u
oMsP5gt0zRYPDiwTBsGjnFCCfK7YZCKX6i1K/ysehdwbmdtHjkQ/Ez+punPWlOVlQiAqy+k3JkFI
XLHR4qbR00CzMG4CCrdEwXO5KbMdowv8zkyQf87ef69r6QcRr1+bx0L7zu/N6WCxYL1f215MAnpO
haeEasoPfArsucwwDXOT07jA8cb16iI5LvCZ/ZvgqctUtBSEtOur+xfrzCB4OHb0zPWNcGmUTHho
8APFN1YamDQWj/UxnqAxvMkNbjaYw5YxBlhOy6YTxRp5yjaQCBP2LnzNCCNDZwMf9/GNWSGRzjf7
9ZPOojmyPJxauax9AjmOcghPgj5H5rxQZ7/ZqkfkCqaZr7k0+zZYIIMDAsXtd1grBFsyRgyLB628
Qb1ls41xEcjViSx3RAd1JJIe5URReAdJcqUhTL6RfN8bOFT4npAMUP5nssaaf8KRB8gevcpNMnUa
/61IFu4Ui1Ka/zCoyjDyK8LZlkmcviM+6QQWXnv7MD0BgeH2Li39U47Xfw/MqPHnWGTfdpH3UleJ
+UXAFTQ6nLCibL0zQS9Je1xLIPU8JGPLcgjEdawT011Y34qtGmcx/oJb+b3T/ZuWP/JJ3QG3Vtur
vjkVqLXy1wRvERg/A2ojPl5RLxPFBEm47su3SLymn1LPe/E9H2xwzKg1hH2iNJNPJfc/cMkoHQm0
GOrPGvkK+pciZr7JuHcVP2Sq0kIqFJMJJvaLhpWB6qTbciteRtm4ShwMNKsOB9d9zLvZqm8br+qH
4sbR5+XHw/4f5pwm3Vfv4DvYbLRteyJujpewW+g3MOuE7rE2wNRSIK5ZVCj3TYR89dytXi23+RHV
a3LUQ1rzPuaKSnYRRHQrbe4hw2y4iCF0NmSLFegjy7kg9Puq50Fr5rTp2nQk7IyIiFLwEYkFOROy
WLp1dQB5sJKBXVVXce81QCw7Y6rCvSuxuhXythtvWP5X4G5wAtW2dnB3omcea2cn4gxEbGQQySkl
pArTr9yNk+GzQTe/Sr4wDiTA7JGiHhhCl1C2ajR2FohvGVH/Lov3eA8l8EYl0fsDY8A0fS68FDrh
2/Jf987TI/CYvGDbSTgDPh5lAbMq1oh8ZpNy0eN7hpbY5pOTU/5ZFyONsrDi5+pClCFG54G3zZtu
POwTZF3MTD+550anz6AR3JTCY0pn9exX0pE2M5fWWGyg+2U91x0BW5Dvucpi4O4s6G411/jjONE0
3Xn0ugxoUS/I3RF+S+4zqYhKB/jBT7WUEUHmV77dFnmhTIwdW12yLGzdh6gG/2XwoEckNFopC5R0
3XTXz6iPn/hBjyvD53+Om5N6Pxnbqs4yNCtLv77i2+xI8b2OcIM98NASzcpSsTjqYYhzp/ywqX7v
xMId9OOcg+2jsDI9mvmNElrvHG3ES5lpDGABMkV0coFNM50wd7VbLH/Alxsp8WmN58xRoq/4CKiz
ei7wE1daIF7TiCxmAcrKSiFfWSOa89jtnHZnoDQmJNkEjSefRYzo2zq7bER77oKCw+yhgKIZsnYA
DvwcmlRPJsUKcPAuktZcEAV6rRg1QlxVi7S4lflARn2+lWKVuw8TA7j62wmCr0WnZChfRZr0eJ+S
dbPfX9NZzVAQswfaCFlf0z9q+bKM+IAmoAck0iBxyA++2uZBv2p4rRGQvO3yEsFc698lU/jBxvLd
YoeQmlyn3jzezgd/HyoTmebqFNumqk4JHOvSXZv+X37q70YOl1rIL5Vwe5j+TvITSa31Q6mWOQm7
u5u+EWGJX+L286NEin1fKxWYf8XI8nEovUF+HBUacoOff/1NF1v+3skvHAlYGQ1cvK6eKNyNTV1y
QUKi4BBG+Xb5HItGquKHi9j8CVebxf7CatRqRqH3TWR2zU+UW2ADeUzzuVUizfmWPtmaMJGkDHqg
qBR3CSmOtH9lniG0uPrvayGfqkOfHBu3yFiSTVoxW8j4mm8qYZdKJP2ZqdtAaXojZd+yWBQHMoh4
CNnCnCI9bSMDa82TZf0BTeDh/+JnQ1ILvWRWDUvkTYiY22HPGIfg75YyC91skTvTHcz6cmhVWUbA
99yAh9yVuasGQkG8GI7GHmDv+582jtgdOyER2wC6FxC9ISbspOGYh4bKDkwA6QB0Ox+mgycUzlZy
4SQihrKgkDai6W/+Riy2iC7MxChOD8MPeZDcRxn4dxmd6SARKJQLiP7g43hVPuiPSOQtZmrsmegk
lD21U0AkKgmgacM55Dmc/3OzFik82jQ+9uI15yo6CjqVGD8wl7U9UZY/uqKckMg8kjkofDRGegJE
TMULTBPjTuYXCy6PLwyhiAsJw/BVYrjy39unUR1ndXrjK4DEff0G78ImTMuPsA6J2GpRAr301yKm
YWefMiACryoiXDwbVinU4ccicdyZrX9RH0swVPtlATWPV4vU8ndmc3tkPMAvozGSHBqlp89ob8cr
1FOzD4UA1yJ2pmZ9MP2ylSe3bUgfnVQCFNq89NCuEPE6tXuL4417u1+MNm5xWgS2Bn/EMjVeblL3
G+BAxrek70rbQhYMC6etcLRNaSwxnw1hUAqSN8fyR/xSYcnQRct2vMR0PCw9LQHx0tTRSmsIOP2G
1sprkoK+6b9ftO58hWIR9OdfAL6SkibbFlfVJGfnyAkhPHlxa2758cYG0eXPL4WMU3YnmsCnIm8p
/y17MonJ2pJgSCAvTGmTFfGUsmsfxAB4DDQ860YTnOdUQXCq0QQwrfByg/7RbdK3Mx1bRySb0LBT
uLvpbHu1Xrn6PxkZA257Vziljf6tZPQltIxdeLAbh9IPHQmi7mpd6FJqXL6jS7oAQr3UtknTdmss
w/McuieKJcBWdnOfc7Nd1V/lLKjIpn9zF8G5Gk6CoM1Y9/wSCD4KK1KmCZPg+NRu/oAyk+a53GQy
WO9wuDgw7jvCyW6svbSkqPqrFlByIS+zNeqqa+5lPZ9V1jEMpXxelmS+co7e8NdVHsorvv2wHgeh
o/ZHT0Xy8IstRhEHYWs8AkOvlL+7qTKjmltMFnSJHmxUzer0fFW9G7AQYCAsyOnifotGb7jsXhIU
kyPTgEotgOKyQVyyaFs1KgTx9BqpVzsawq0eH0dRqYNbPfOwSTVIZG7Ikj53dC4QSZ9BakvQczfB
a8rwmB1yCFikRHOvywDikDD3XGGoOK1bqFCSZclEa+eDdSA68U/KMwzOzSUpF+TqMAxuO5nb948Q
FNeq+C7qKial+MmOd1mBnBdo7JAXjTkVyxuivGONroTPcKPYygM8ZF0iuMiK7PkcaCsFmM1lBwGg
auw2ctXzG118iZuBLh4lPT1sGOPUiG9znHt6/yq+fFZVTe3w4lHcR8t0eI6MLtdTXpV5n4+5z2Nt
6lrKfwJjVEpSMHO47GLbBmSuJ2eOemDig4h46GXFgvN5+qmmwe75+FbLJCSbwJYarck7lHQLOhlQ
J9qhu0Y9PXFRnrFcM8PqMcMMNMU79McjJsZ3anAI5jcgjfE3ZnZAat3vlh1F0kLnbL+6YvFj9yoB
/1/tn8a2Xgrm+h4sTC9NuRZ7We2NkD6/wviStC0+HnGMeptEA0p2CTy01CfpWVERhCAdmBFFpbWX
XW4nl9KwkXCEVsr7Ue2CDcsUu0xbQOzyyebT5IE7Psm9OqubI2qka4iVnaeMIiTCBvBe761AWT+J
TszSmrg65YqiaFra7ICMRbfOTK1Qf3pqrGWLeLSndreV1/8MoiF77ummagH5qkWM5iP7REvW5tXw
TvPOZE5B5VlyNluw9V8jKP03poMnPnOAKwM+Gdi5Q/bRdpskqlp1TNL7+aTT2vrPRi6ksvH9RMr2
TzecjM3qOEBY4SsKIxxfAvJi3uKuFf6p59X5nE1An2eFI7N2j1dO0+d5I6oSPHupTvoc0vbM7put
IfRI9Gy6Lc/Fhm4oV43LW4pfdmYsp/leFZUp2FZZhZDQ1UpZQJ2Iu/rFKQNHnn46i0C6WrR91ucn
3Dx1ESqle2qyZX9P00ipyii3Fd01mW3ofa5GmKIUgjty62HTUnonwEz9FsRhsF1zk8UFNJyYnEFN
eHlsQPbi7V3GVYqjttWd7FDI9JcGt0dJwZFlGwKOXgoSMtXx1GN2P7EOdB0aqiUfYN1ny7Xx+Ms4
WAKmPJD7nRUgvXiTyG6bc6RwGc8M3p9WexsxP0qWrCpx/JnTogrJxfIBHqCxK5eXFZ0XEDdnvYoh
t5++jOa8fy9mUwyF86DfGem17hSvEB8Xqj1lGhZFCESM2k7OZAOUNvyjj/YMD0Z3Qw85FY8saZFq
0AcUEUPoeIoWx6axW+0EZ+PJoRUFHZC3oqLCmvvnLvLIeuhbmhTK6/LuJrEVaiTiRSrQBUktJ2Ia
sHcNazV9+7Deo4wx6/enjlojXemRTt/WcnYckNER2NInU5gqdxC1nOivWl/gxmvZDNZjrM9lv73W
gq2cIv36kF9BFtboWWFXWJC+HSs25sqXrrApCx8dQZAZ7cXxf9iqXgl0e+sVDO+sDOt9sw6Y0RgW
Nq/1LlMfbcZi5riffPwdssMHKTmdw/SP7aoWO/DAleIkAFltEMTVYc0/abp2jr9VvFTWyniAiM6J
lsSb6AxeYq3PA//4mDH2szbcTqMmqJeYbjZ7eHZ5JB8wNQJegJdU45Hrmdcg/5XHZY2Wciyp5T3B
3lod/UYS6UkBDNVzWYElpQGbcFz2y2Gb3ms6RfKxiI2kXqCn0HfXML8mcOhHo80RSS9a70tHEI2i
OA14lmw2HmkvKsP7GfyCoyB737ColPvkroU42DlSIWkDpz/c5CNjSDifopcG1esoFZU2n+7PPTyU
4PjciNkW+AS7OVN7atxV2Z0Ls/8X4N7OHZGWnOEt63vJiooCIA92xT8PfORUqqlWqliX/aGxmokK
HfGiglhQKfP0Sy0C4niUQ0OUqTk57WewX8g1XRwuX6Lf1TnuxwB6+0U+G8K92MLf48ZWRRtoY7jh
rmT9j3d44J9td6zRFDFIs5ayKhBfzhfAKITzaxE0jPbCBlFsyXNUvtM8B0SYJGdiMSYkIEeRvZhn
Vr1ziSsixVxxIINEfsSO4171pKZbejxqzq5IOIvQSq8mhl4/OWJId5jf904vyVpIyyya9/J19/ok
w4LCxo1DcXr5mtl4Zeq35Q4HPSJQeL0v9z4D/rxaqIGZoAAu1u0ZvLb+iVYLERM6B19Thvlf7y5l
R0Nmf+Ej+v2RSqB3P3WRwRXoILfxqcxHQGrA9mpemjNHp7tZS91CyVUJVJWtdZ1nnStq90O0nPE6
i+hrzg/yUownLXs+josHdL0eMNfluyLImErJh/KTSoEZeQttc91F6vSu3qpftq4WNxLtyi0a0apl
gAj9b0v5ArQNUiooOSmiveztYmIZIaxTVJnfQ8NJotFucOXpaFwxpHN00HCU8uUKahhIsJVvN4rE
yhecYCMZW9pTnmOeWUoiPEkm+rbUQOl5aJIUKYKA5psvbRVpAe8tkTD1L696l/LNpeKf6fQZQtY1
wZkWHTQmRg1tCFDJWZ2IDTYsKD76Pwd8tlHpSERgt/UY9ubdpdn6wlS+vi3JlK798GqobU0CMxOC
1J+92lDxdCZ5AIpYTYKnQwBVmcOKymCqbDdijbQb5J/P4zRELThEpESBLj72Uu0T/PTp0UzYa+sG
2HxNMRLmJbb6vT3EPOqSB/5DPRCI4C2qeG3STgz4u87tnwBsqAkkMPomjBED13VpnmZSnt6tJffd
AOeDvQGdtfrfYWtbC2HJOP+nAuv5YUtOyf6kZY7DyV4dYaKkTv8mhwSlFZx78jkG0QeFbN1CVFKH
g0ftEvIt2J1jGnIAxqJrdsqJBtUUwFBCzTXKwlQCXu57wzvLT+bN8lobAHvY+yNalyDfQ3BsS4t0
XmqCgbbyvLmpLZS0tRuLro+UZa4w8ZjP3A3VKKiyq9DSi075EKuFGORZUZGom+DxwFu9T9QZlfbE
3o6aYU6F9z5bqvLnZPBXS/CNKqi34Cxf9aCqXanz07ek4/XrBr+XtIn0nPEwPT5m5q7hJGh5Z0d/
2ZivkpTcLa+/Rpe833ppXxk3ebDseWz57ZcLYbOiT2IABsb4C5f/pO9d++wAxBe74Bt/qJPhIF8T
EmlbkPyd0NEaSyD6YTr8bPmqgRea53AgZx2GIVvHcRHY1rTBb+zLrUzOzDRah9nxOJPGQBDgA2Kc
8uQf4oYkJVKWwXxX9H6p13YHi+zjzZOy91hvodE3uNZf8PcoDviOjMVL/12kWZz20GTqNJODBrLF
Z7jC946wg/45CVMm5WE97qbGXBREGqvqB5ZswyLlBuLl68vg8Qp4KlQ6gOcepGDvZ+11mdCqHzDg
EdusbFxf/q5cAtrmRS9UnF9No3nW0AagCTbTmxU2dcJXS+srwu0aQnYUVnDlPY5ccXsATlHvKxYB
tOzer7+fZDIBAQ+Ha99Bmpq09yJVFF2sjemn6DTtXray4wvuD5Y6uaPg79792M3amFCWqYjoUIcI
XekQAHGJq4RFpt2lNbJR76NGtyFlzU0WaigrZfLPdNfYXNhmTevOujS8qAez/6lAmyogivuRtDX9
3BxaHMIMIjKMUVqGJsGXsee4TGOQYZiFM6bNifGCx/kPClKU6sosgXYLQVgie2ywzhneXbH/y491
7i++0EpSr3IPz3hoBZcZ0ZFP17131ILWfiu5THeueZ7mIVSLKFIM8tkYDeztffSJ2Go+m5oC7UqN
EfFLfebsKKfDl1yE7HVOx3+p8s090sZnL5bMOhX4TDqSmrOeGTQ5tFDHRH235pCKBez6gmm/oAIg
d6gP6aGiBqRPp/77QHWOTt6Zjg+AyTzFfQJMwXnizFkyh5EjjCFlEbCBaTld7LJMKhnxrFGYMhwy
TSWCl8GpFOKprhHGtrJ38hvm8PlNZ5nf6LOSIh40f5Ot0T+8rwUf/0agbvByxvJKr6EraLkkTnvg
3dCha+O5hg6is0oYoRW4e6R54kIfMQI/YVI529jSQbKw9z92iLjqy9VIGhmil1+enKYuVDIm6kQm
2ioF2QOhdQuLnAD4D3/8JpD2g/9cX9r9p2WEpb72dV8q2QvtcFku6vc/B6brrESvE8flGe7JY9bM
AjPFPggzclhRkog7/7ouQn1Qqtiln7PQ0pVs+Y1/BR8WOHuvw18vtN4zIQsk5Hw1I2IQpFr/Gx1E
XsVMg2aPLC3GqhgodIT/+BKoyqKxkjpCQfenulNy4eLkDLQOSsPc+tQ3OG8mkVt7umKZUacJqcU0
qh64lmbo6xsxfD1dCMWuTlw8TCczFOC/m1VZZ1hfnkXYa0lM0sGR+4M21s332Ld0k5Il1O8E/FBM
x9IQbOcz4j8RMq+SxSGXLluW6qaJ14XePDEZyLTJbC4A1iBbFOROuPL4ow1gASVnFCjbyYXPPU3w
kY6JJRq0kAJI1yg2VURFax72EAXYcDsXTIQ9M0gmyZcX7lulGNGrNpECpaPGlYdVWXvT8ebhtq7L
26WJK87bheEfI1WZqniXEev0tXOQMfvR1H/kcaJIHIGBMCO0Xmn7tPJUawrG9Sqh4l8Fq59Xec66
ehp8V9zRth4+Tv/1VQLSB12tGAJd6LqeXqh/k19By3AN/4uGITEI4JQWQpQQFo55MphKf7r9vhPC
awbEwX5sWfXliV7T8gAfKYmSWMv+8GzA18dCsCJosfUllKMmZlS9EKNze/RzcHY8qpqCMHDFWZD2
otQnfOxbNUSc/aLTKmUPMhRSDPl1Zj4gKXyrS0H5YksTHu1feZDLAsX8gohEDLBaDzN/B1d0q3Da
EDESJeM1RHStyPv0Gqbxu1FJREKOKYmnGCmmCZQAkkknuQC4VSPnEJfKMSEjOcFJFRUEgSOyOI1B
nFWO5RZbz73fOqf0mZrcF0aRPFWvEiS74JuwgdqOA9VfOCXR34A1mzTkiCytPxhHGNRNqXPpiWWz
uV6hoZwafmmE5bCPsfT/pUIzoxxqAKmLiVIwijXecFDFBcTyaRUBgEHISHPTh9/IItzwzkVrWIGV
LlzPcH7FTpYPw4ihAXBccNaAmd7+JsE2se+gwbpmR0xYlkeFTghCN6emDCGljvFz77ZzwPlujpl0
ACfsgQVmoipL3kPQz3MSDSDdy6BOjoLDLAZvZCBZ5YXyw4i/F52l2bM1ZCiNTIotyPZbn2pBJTs3
4Ukw1coML0IW7ESFuYHlmx0V1FQCTOGnYXatEzSqlQHZ1nhhnAbfZ4nCdBU3Zz2aXhnyif6gD2mc
n7ZLC88Evxv/xmpt3EG9FY7xV856NiWZrsuAAF5Ge3xhVRnckeGkHGXqhtmmD5fPN9GqsSh78SgF
u96wLdexWrYbMt2MlX/p6LBWCqBE5Ki+sZENpco0xSsMcehgO2IDSzrKqY3G43ivHYtRrbPeXDQN
QPMPBL/Q1ZLCz3HRIzG9+CKixTFOyh1HTkb2NWkLlY8kC5O0RzLd0NDBOmimOSuT9QZdWjWDaWRG
cVbkS0OPe+J9c10ePyPiU0CMJqwaSn9872oT5wDmCREoicNUX3tJAF11JzmycH39mvaZ8X/y1/jA
9T9qP+HYT7xBaHRoSV8lRMqSgLrgRVqPwa9+WMzeKU+OG3/zCYbzJv+/5qgG5dsyGs1AdE1TZcEj
pPBejaNUwxH9sgWYfvpu7twamNJWHnaQHFfyqZTuSboFz0v2/BB1g/9M5b2hNHK8l72U1H7H5Dyz
mlqPnVXBRai6T1zSwvD5hEK3W4eae4R0i4rIScpK8vp+Ilv0ZI5tEtEJC2njfhXAT/lcHDe63xHx
oAzcPWqloqMG57FkZU0nZtdjRXctWHxgR0SUN6PbLHD5ROd5MIWij5nSWFVoPZIr3J/5khn0ZVNt
fkIh3BkMSX5myQjnS1m67ii7tVFQe6m45mCRaV7UftKqol0MKJ6zm8B0utvS6crFwCmJ2B2pf70p
E2pm0nrOd8xfi1ybzlVUuqSbuDgkTA6Mzy2S8cN59Y8P1ppU6tlA/JEbOD6Z2/o9aGt36JY7FH7z
M9P7fQM7VDOjTdqSyZURP1XBUBAEvH2hQ+Ojmt38uJyWNPOKedBocV8X1mdfgNtI/yKZ+dhvdil4
oOtYj7UgHWKHqgcOvKnD1SaN8/7HqNGcEWvsI/Z7oZUrMAt3qyf9u00zCRVkE0+ay8j+Roix8AL+
S+vdTbDxs3VVlFav0PzoNzRVFHtX7q+zVcJglQ6pDtrA8gOoGAhqbcmmf6u7Hm1vvfj3Rm21gVgz
KcZTViz1T+a/7P5AgiDHnB9DqcC5/pDyQQCLx/1r5ZJFcJ4HNP2IoW4peYlNUfwa7QSJKm3LlDm0
mkLcNcSDGmnkoJ+/sDH8k0HT8ZVaLbRhxm8jVAdDnZk5nwyKXQqnGKJqhB+JaiMFl02u57znKXkn
T7Y1AJz9AUQQRwLNNtWEVGvqkUkgwweXt3/DKDdA9mGNnqXPiObk3ttwY0cp+RePCYI+PZ5i4Vhl
dg4UfC4zHuqDwGkCEIbaUOqyOIS08IzM/eROefqTRW+jDXSqQy+jwjiewBYnBIBnhY+lrUlpq47G
vnLtV5zVflSfKV55YKEe3bHo30CbBLqLP1RkloGI1enAx7T13TYmeGJJSMuohek73Z2V+bXXN3fj
vu5/QZVv/ZSt3XyhUh9w/t+d/ixlFW1zKhBolf43kQ1MzcW3SggobbjKrIGM9bM0fkM6GNHDpodh
zlk5ldtz9KccGftTfAgct6V0HLW4n89rgPlAL5UHQPdfdr3mWNEjhVqj/yYn5tBQ7UbmzCES/CNO
GR0djohY2hPAmUo72o9cmLOugtMJ3lhmWPLRrS20MtyYMGM+lGt8Uz2S10jpiqFGl/Sr64by9Taq
PabQX7foV0uY6XM2j2rMwK8qLEfVEpSwpnnTV1/VGKZekN17D5tSpYu9QxNO8E7Veh8TOMolEs7w
PSKxJArXhMtGdvSXD7slmxTT64TyPXpxQmQ1spRylwuWByYqvpJpPtaOyayq8CukHhgUekK7hZQ+
Z2WNUEZi+9VvOt9bFESK+eiJ6K/fcV/z+qe03c8oHZ2+gBsIEtJUd2VRvJsCq74YKh1AAl7toaoA
WaIMRPJLFnEHzsQrq/CLK7jjkkyxl7ko9eJ5BCvckTNvpOgUPUWCsusI+mH31scsMUIRvk1BSZ/G
3MoghScGQpkxnquD5sA4kaMa43EyNrrbSIav4/0MXfQsrI5CAb7NGIxQiz3HgQstx/kfRsUYU5Oq
sG59Qo8gaiMX62pEiE8dAqQkjzU8sdS23cI3ewtFJslY8FAa/3lgKDFWpJRhgvG0cUSczMlS8dL/
g0WpjKtPEeroCo/tuujAAbsAbkYelDfW/hjcYBIUE1SgVBzbcvKAkb/4q0Dju47aKRJoaIhPmoV8
GaNK/nCwvj+gv/rgvc7H7n1eXPall3HXBJaPBdgX/B54gkn5Tr2IqAVx6eH+PsgtdDwypm2TBlPO
8qft/7cScc1C3Xk3fQasi7+ubntd80JOzFW8Eam5itR2/CI8uy6ZcGD5dWdl1Ey3yWAcAB6vRRhl
uW9/wScB7gq56X8WKv0RbGzQ3vnX+iTCpxXR3Q1KUscnS7xTBhU+XYX5ZwNBjQxr1+z4L61XnAHo
pj/WPPDfgn5GvNWQGEpv/Z523FFrbgVrD/XapxdAQYwb3nvkO/Fe8qnQD+Zg5bavoagVD0xyNnTr
MOGSl63QDc7+Tm5dwu/grUZMdDpr4U0Ua6Yvn1SqZWdMkSCYG5n36MAGggiq4qgzK0XoUrvw8ojQ
KYKx719acb6skuLJpC+iEIgsLnkvbSocNp06WVUo9h2H9KVdDpU8yGLb4jozx5nwUrJYR3CGY0OZ
/Bu4OTd2h6SAxWK8g3hdz9eDSKjohk19YYRvVn/jF2gjaPaolszDq8QvN65vyC6EbfyarqteHpmf
TWv0T2BP3JviL8q1v2/RicGHcPry5VaRNSYmP8RtYEfUMKc95ifumw1CR1pcRbDv99FjDc/UIU8m
9ChY9msaEYFmfkO/NliIpsUCS7Rjc3Nd/Xj+23kV0lc3mVWCDXheI7UILOdA2V4NEO/mFeSD8eRl
hhW4nUjkFu09ZVuVDrehqA1oFK92AjdLHE/zxpIC9MKaxZo+bJOU9U49uaROU+lXk9JXgw4sh3u4
sQkKJUfiR+OxbpUBEg+9XAbZpUl9Cdgocx77hfChg3PxAbB/07s6Yw0bIPecRHfmF+TmSDym4kD9
AXQ+A2Vtm2npjz2S8u4xTs2q5A/K1SKXRWckCXi+hTY+u5j50sJJlIbmTVoW+lWZi1GnzXzIdlA3
qShGYPcsESOPpB/bLEOsffYq9fdJZckNlH8y0W6Q5v5N3FRjc9C/sV2GgXyf6BOgIPvw+Xaly/XX
gw1uQMcOrlyIsIIPJc6GbqRFxlJsA8/KGRKjUArSfJSQOZZtVROBHXmXWS5ODlPw2IiHdNby6UCf
8T1L7P9Yh5vPX/gwVrQwcIGzynyMqrwcQs0EZSKZuvE0CwLTkM6VD58z/YFoZRl0tsPXkkhLT0+1
2yI5SKoarfqT9bM+jtmVUG5AIhlkZovZxf0eRF3FG2Y9uEj+K0jK/JZNXrF282K1nGducAogmdbk
bfnn1RaBdirIbj3RSXhPoSXmLgSCOhPp40shO8PGnsYKs2y0p75tPMLq/qC6I2iBtZ60vheg6kWo
hJfSH/9XMLByka4Pt9rYbljxVo2Lbw30krG0pB+JOZZBxo+ZtoKwTCfNr5VMJbwUPtK//cCL6lel
txCVxsb/ecxI8I5qnAOLnf3iTJ0MiSviV36rC/G2RdUIVQNGkES7+YBVPX01WwlzLubuulAJ3jrJ
udgLZXyJOpG2yLd3DCvo0BYZtTrdAvfQiC6DU+Q0LVBMesPV0u3fwN4DbfRG+M74GYDJ8lc/V8hs
TrbavvhMid7xk3K15T58qduzjZFCv50Rm3iH7VjO9EW3fmRfuqxGQP7O1r7/SDqBrPntCK5YCqcl
HRfq3SrgXUU4dLSx9CdMzc5yBbeWlSVR+YgoDuZxvko90EwUgHhP5lMviN/XnNH2kqBvBEbMIrLM
sT6FqibeUbfyYlYVLLZLjtHHx3YW3cz8ua14o5lOvIoojXAlRjLzhyWAxc7Y3tMj7CH4OV12dxEX
K2qaCGQbdNt2onwWyf6/vC/EcOslXzaLrl9w1oWGP+IHZxVsNzXajkTxLzTYI05O79Z1NflSY7zL
ZJ7WRX72yPFqhgU7l//Rv5PklgEPxyjIIh5plNuYtSNXfkaBV4hPm9awMgwLP70L5v07AN4OJcRp
7dfz5CVXHr6Yn2Dhg/sc3qC1MuNdkQQjUbcgmDBBOGgzI6JDOTVvWNJQu/KpPclvdQyTSGPmqtC3
AvN/6LK20ge3zYp5BjOVKndOmpvr3Pg1tP0VBmp3nD6Jpaqgg8n0kz57Jv1Vk04LmK0QljrJEhSU
bOC8DNhh8BbyHSTmBqhiI6uH6bliDUV4O5YljrwMrsEb5xDEUGoIRYTKu12fKXVD2s+HcOWB9WIN
BuUutQyWIuUwwUYQFJOm8oznEhBVMZSKnvyvsp6/rKW/KQvkQlPZDaZoXC+hfcBSpPTTcs3iGuMF
qyZeXCoatQnKgR3JzNTiME1xuhsQZRlma0kjZD+Fz46GzrRW4ZnUf+T+vfUupCmaL5zHkKDuEz/4
ihPemYl3E4oJAlGDG/XGjZF+dQ/1O2Qhb7Mjk2nRdIZcFXVEM0zcHy3vS8/4T//XTG90fzFdaxA8
wsoK8Orr7axpf/aEL2JP1ZHlajBSdGpNzYEDxzNXiP48oHw5KlNKfj3W0wG67ZQFsnM+yn7h9e2V
JZU1REJFzVaAVAM8VqY5YgOReSWh2N31EY4yFdXtKqTByhlV/wsPVfg8ZtznUAE6N6Kyd0c5oDqJ
uDnZv7UTvUDreWZccOu7mka19SyL9hM8lEVcwXgGWU8RhRR8JyCXUK6a9/tmNNfiDmLB32LoXwIU
+6wsJ7N28FliFZ6oZKADVvzEDjbUwtd6KlXfZVwN0LkykC/QlhCkOlYUauQq2d1SmOShvJ5A7xzD
jlLrPwRz5tlMOTJj7Lqt16maQLscuq3XcodYZNi49DPT+eamV1rO6KCgiDbcEGBRmlPOBfaYVt+N
F027cthGPn972V4+GhCc9n8eojTDPa9/MaYS0F9TPSkTGZsiq6JJF3JfHpWX5UWhm0upBAsYVNtd
/x/YxEXbofAUrU9pczpWS73eGtZZvkkbQlXNQUTIiQvZ19yO8GrIkyFOnOGgPyNvGiegMy6m7sPb
3i4Pro5u8UrB0FuPIwCCkBIXLGtQ4M6LNCd3X5bGZ7QvKD4BA+U1miyas/t2BrAdErWYABEi6GE3
48GkcLei1YX8qMhPtzFc7v7pkkRKaGoXoS+O0olbuEdh0WXucBiHH49it9u9GT0Jrpcg74MHii3Z
bkLp2CguSHmODdUfT8OAYdeZK5eksmNawNwHobnBqI16ZirJ9SOMnZgjLCTRlxmZLp0qZcZ72Yd8
J0578hxM3z2RrzuQ4iksm+DJVjPoHiwTD8fxQ1z5Dy96QstDcyrkM4EC9yTPcoVGeA4IvSadJSyc
/D8xGonFO3DVSjKqm0vok4oSWAXqTuplMS35u11NTTPMBu5sKIokOAjjrc//JVk10w5sKv2pLGvF
eq/NW/caEM+moFIlYEBkYKFLTLhw60IOMTBhW3ffQrWI+WM9/wBbaKO/qiwZH2hRmAlVaX/2ncA3
8Nv9rlYsZHWn06USWT2a0vjGh4zyl+ROQYjBHTnhVZ2hBA3iOoMdU+fzmlfQrh4o1PBJnC3Z5wP1
kpbOsSay95+7Dcg0f8OoJqRAdTH/8J47oEJAmJpWJOTqgEUHgw/qQTEJVyDEX7E3ClLw7/5GKSlZ
PMW7rTHJ+pxotCCZFISicZpjcb1NFc2/IfchVuWo+w6rJML+NTfvQFd8GRm7xt+eqNX+DKn6BBss
YfGh+N3YcpEfvtSsyURh7MhX4YLTdbpYJQTVONNe0ySse+MzSDFyw4e80ripyoq0wXQn29LmFDUH
jr7N7hKZjq/EAp3I9BmeASYVf5alxye5kdaVZV9PXTidaiGMzZB5tNkFH1VcocmAdlIXZ3yt1CS0
U1YbeUGUYMr/Ci5bVIxbJXDw0vxke7PkL7AnUfWC6JkAHOY8p0Fe9o2ZkkcB+RC+QiDn2r9JtlAx
6lqR/3X4cldh5vq4QizyN5KROJD9tfcKm8xWwLxoTzF1PAQajUEBuS4Vo3+2j9bXdz0uSMHcpvPq
iauvtoOH+uyemgQgWu4+yn0eXOKKqt2nYEhnDfCHLSuikDXCznlCYpTo+0z0U17WobOH7I9huWD8
jt5110/5T+TBvYN1GAvyCpYWNMZpGJt1RO5QOco56mZ7GMeTPotrSm6V/GC7XzMQ9D3PhTCMBNs/
+KFNhJ/bO9bM0l1zHi00JN9OKlfA6G/NgwZ0FG8UCmtTMLkVKqqZxSaRXMAr72FHgjPzmtDOvedH
4Jggk2gT/Uz1kh/EfeaxEt6ZL3RC95IWv8SI/++MroCYvsPpCG+739cN27Ow4sR+J66qKOa5gPns
2Cq06NsYzJZXmsioNT4T/Pq58P5KJdwGX8NbVy3ZkXxl1DCl3YjF2cy1A+p4xiRWl33nEsEMi7Yr
H1uZHf7OI5zliuTXDYJ5mkWX+shJw7C4PB4iLEgcdBFtrSvYQW1jjVFVb1nZApU9iqUA18CNElKE
uF4ApZRiP5eHnDWANT7U9iQ0aAaUbAizDcbyd0ehcwOc2mKEW6cAFZRirtXS/XDFhuGiSBw1DpGh
50B3wdcxaiKjWikJw3u6d40+EUUrgQATfOEHbkjgAMVSgdPuV18SqolXkYq/Mt8mrGYBxfOKvDdT
GIxZCAfmKrHpdEpg8f/9hGjWWeCT6UFGnmVA11yttb55k5OVFTWzDKw6Kcr86YPPVYm6QyImP2QI
mZFzyy38ltxgsrhJL5Y13bD0ycPJzM0vJZPsmoLgcei/n82idYkBJjAnP0WMdLIpSnaASgsHvfZs
S9XzIe3OGeYAiz6PS1uLBo+VuGDCwk+NNvVB6cwoE9MNqmayQ8G/WhXQx80KIKWQhkpUNRfOAOi6
IQc3OLEC/sGXEz07rNHK8FwUKcoaPpV7opMKosXT99tdkh7RRS0INRVTuJkK86JPJlD+TGYNpGBw
tTozfvFD/eURlGz5anZYd6H2icboeoExGy/d/BfklfPjst6hfJg/d6n69r60bLDU38+u66kmi/FR
0SRAbfU7YYh/dnn63grtfLriCgOn5usioGJ84uuNEVMa4L1zcCH2gZJDL3kURF/8bI6Hlc/jY3Qt
hTo05N+MtKgea5sXvN3cXrgGXZwLG+4DE8CE5cnf6Mc4bkwQvHQOrTJ0JjXqtqCi2Yqu4Sz4uAaM
Ryk60Rie2WtUnZqWHye9aT35JdFA5gp3gKBrVDyGoIRObxJqT4Tk9+qnAtvLQYa/8B3Qf3gbPrtX
h4mk6XT06BbLHJqMfxmEp9QA1kimszKZP+UTazHFjGQ/ra4VrTNf8RRspcNmLHS9S75OfsF0Ed/T
5uV0DrOLUAOSxjZKd0YuBheaSKZc5LAvFimnSgk59hf1QStp/iH1qxDAgKSJ5vUHu/mqCbR533BG
RTxI3l9q7z69NuC9G1CdX2wIVVkH85tOn3kiEmBH6Brtfo2U3eWaUl4kPutialmbLrCiyprQ2vKY
IT1UHaqxFgyb6sxoNxrTQUAhBK6YX3sL0R6/sBQjlEQMBgA/spMuwtb8/vYG5FqjZ6y6xmD8W3Bd
plz12qF73KEhAs1Ku/YDDTZMXrtn1qJdojmAzhu2CS2WZ8itVp2IS0Zen+sBThOVcc5uaZgeebd9
Wf42xfjtCpymiNocyH4M+HBdK/cTLWwjltFQVtcKUXUkOM+fKTOkg61AgruifyOD1CuiO66PIBcG
driY9rLQ22aHwCCc6p85uQ25s2Jjr4Ivo2edV+2GLm5BT3iuj6Oi7HXWmWZbgvze106InWecfVAv
TfURsA59IC6NQVFadwzqRXMZXhfcZ1QZHJeCbh/LZBIkIw3NEfE7RgSLxsLKpu9WmsUsCToK3vXv
vyZ5QvreD9qP/6wewoK4St2/FGFI7HJuhXt0qhQIrl7lNrw8nnKRo7slsGpl7zVco6ZB7P6mSkpU
HYViHTqCLYNau8EMguldpBdozOijz7snqo5oLSdlfy4OZmpaVlOIm36RuAna+uTPDCaAkH1+zVnZ
uHTUW7Wiws3m4cKLLVU2ktySPn5N/ibXCTU77MlYpe9kqfav65pH4BnH+0A9YOMnPa8XVQKh73Oy
+j3foThYF6ncQq4Wh9fFQrKuOJOM3E6/hPiDkh3kYULRpyu5vAT2pV8xaJ+4/CbwfiEIqqxO+Hyk
A6+8qJ36I01YQ55nrxb1cYOChMrlYECG9ldqCb1UJXEttmmsQCs3cv3qmEqvntVz5gb+7aOO77qJ
BhltdDhWsDhtifvscigZvrcJ3zMFtKXToFRcsFlgUuIlNP4c8/QtlGobBFfrrG6MncGnpB4JDujr
UNmOM0t/EXp2fv/BmKI2q7vwkWP5vlFXwtt8Vx9I9GBj21zcVKkDou1n6uBlfVjX3P+Esw/BsQUi
T81t+trSwl10wlY+HdhF2BFjqHlqV7HN8580FXogqLeNzfzmCfp/Vj7A4aIs/OF9xSm5WJt3VApO
yEuQ9agkg0sbY+f/TQQ4u9U9AEyJ0HlU8f9hnHIOeFy8UjAzZqCBiraM0Oq6ur0TRWSLL5BV9Iqk
M0gYf0jLy/L5jDa/qWO8PZA7CLx9Zy4h7eYUK/Wk9MpO/ij1YoRPjyCM9p3Dy5LUchV1lA6NCA/r
OtNg8j7daFQdpZ5x0w3fz0wjLTWLrjPyHTt22oi2d258WpZ277/DdnmcmNfJ2bFAYhcHFDG9rbJL
tuoqD+zEMe0R5JKs/y6L6TQpewN86/xHTxTaypzW3tM9zsly0Tn91OL6J0Q1sYjx6mp0NAcq9mqE
77pu+IPAO/89rb9uek0soytZpzcu0IVC2qCleS+mr0Z0amo/RJtZP/UJ+19pUAvx61VVJo03X8g9
vrkHTufMkLY7WPVCXvnePRhVpKYJyQC2Wa8zaKkCQj5gJrUDvNHT3cXkrmsvPM5+o7RuAkMOUPS/
z1WHA/eLn0tdvaDT+QS2amG8MykWA2OiqAxecECg6mkanlWgWoUzcqNEYoIIfQOkXblQSJd0PIci
hp4cQZZER6vd9go708GjHaIjg9X14z/dgTi8CZY3ZIDZohN8q8ERynTpyYepVLclMkPpqMJnOzar
elsXsEQhy43wKbpo6KI89tZ5lyai9ZZlNnIHXf0MKNoCLPYDwLg2/5RCvXAAnI28svDFcNTkXJxs
SKCeLL8kEa+6X2MJZERs/uX6agTj+Lu2/QUdTw6+jldN0r0gVPtKXrk3uNlxzofzQTpn8tXs+Vmh
QjgFHba/1Da5HFA5lYfyen5+5QGvJxoMYKtwZ84YqgaNJjdIKNkcqcIDT7DYXPpZvrWi9RMj/wq5
V5w454mYm5h+ORnqhC/geiIvQDuwo+fkSx/K0p2hu0ucNSYmCdELwaIbjTXLDWMO2F2D2pdyePWe
f3rmpfTjYVCZXVS5B4J6AY04L84HZKqKaJb58xuDMmPkqCs4x4wc3FPBzhgklqOzFYM73jRasMNf
ps6UC/Uz9TpHLVfbEkaksYN9YlaHKXvSw+N1sQZShcDEx+Za8GFjuZ1+aMaAt7gaOG6BpVBFsgDl
B6Mg41r+nVI0nnyTQx96uu2ZHG5wa3UXYcJWOauLz6ygNCR29U31RxfpISARJ9fl+uLRdir0soH2
BFcJsdLIk0bxHH/FHRz8wThBFwQ5VEdgfHNHsCEyONKmEC7rg18OjzvGvJZFgaIA53ao/0N8gC2Q
0+3YyYaQi0AY9IEDya+K9wQ0R/1wJttoVrMVE8XH6xPscpKWNOk7NTN18HgtMhFgYxLs28ZFvTO5
xNY+5Xo3PLtyvVeNW38opgAxkMuXCkEI8sx5o2BJCZZvYSdcV17IHZ+ZUmAMAjBO8q/n9juSuneu
q5HODAoYXs6JpCxu5SgdhgUzt8GYQyAkFRB25WMoCXw09Bc0Dpcmb4dtaCFZ1ia9mYpzJWJwsluD
m5WigG3XnkxC6Ve9saxv88rQpRwrQM/g4GXWp65mYr689vBZ9vEx8mcnpUZH58U+CwVRxIAZkvXJ
b1OtzAEI3GAVQ1JzQU2HC9HEzFfFeVPLK6h3WTTdn9Jx/DfL2ZKzykLmtgtcIHL8mlqEB6eW8LoT
tqjaK1kX9vYtTXuXSXuwzfgCjKEj5Syp4j+oOtnxA+7kHYA+J5t9yCYQTkYk7K+9c/v1V5L5/ptN
jmnMsFKLI9to9mhtJk4qol56SgWOk+BhtBqI/YE7MLDROB4JwGkV91DVsGsee3LehZ9N7JeBS+JJ
G8/l7103AWYh3WCpWlX/0P/UqXDB4S/34/vV3W/HyczYkK2NgRHXWCQYHs/VBYKBiMhx/Xpk2C9n
QpqCYKgt/878thDYmrdkCOkMC5ClqsWuI2DZbCnfy60362hn3L1bZrQA7nATyyrUZ80yVB8Ti/eZ
+tdqTuNjkrlDsH1YgT7RLQy8xFi87J8kjdLuk2cWM6TCxM1Q3BB5La4y00ihj685Nz7WVTViS0+f
XS3zafbwtqNeigB7p7A0IJrAgWVbYLfWo+9JgVtcQtdm/LYcgSDnx5nguo1n/Af3EVNFRjPjTgs2
T1DB93dV99HMjABN7HJqkCHKAgN8ZZzeW1OKuzDHmiARZ38O9tTUqtkOXT086gN2yzdY7MzYh2rf
gRZJcUKPkO1Oo0gf+xTEckAkrwclV5roXaTahI2phhrI1CoQv8+ordT+zkpkTl7Ju+dBAqkMlj91
hTloEHdzAE+LVZaR9vTgandwEYWO56Map9HMGQWGm2eAniOfz8ARQMgLY3RyXL20xyKsDRCn4xdc
OLQg1ytfrfBcDm/7nbvdkwoVcWDmkORSybidjpxPSkNZC8obsx0qEl9eGuPl/zzZY9Wf3qdmrNke
XMJ35UbY8hd1D+FcpoBsOVLa4ZXAqJFlTemIfbU8rzM5fiIAfzY3MIKKkbS6YzwurHfxHDqYt5IU
zdhMwKiWNLBY0yaVhLzrjj9KV88s3sVfA1EdnTdEESTkmYsSB9ZBiuu72yAvoMirfO2KXeVjaWpA
S/BseO4P1F12UYew61OIUeRSp3p2Yap20eyUGK2WAAXpjM4awuz4v8ZkUrYJx8+FikqEzFqa9dV/
HOlRyOTKMDqXrn3caTNqXmFnj3137qvylv1PxRPP5UB0NjZ406axne7X20m2GKecu8e72JmGLP3T
0fy0xUIQ7lmSrLv/L/ANZbayp2QqQzJ3yJInf5V2F5r4PyvXWlp6wuCEOgTF+dO3SwI4ozgAGydi
Dbc82vj/nZWtc6+fZNUm/RXIixFunFkiZLtDXgcY1LujBsECoc7rHEa7uU0w691YTwoNauRF/84/
fczVQLA5iy0tpo+r/j+DD5/jYeH27XWM6WvQ+C3mQupxKjXL+lLF5JzIilk8HLZE7tv0J7Lx8lU9
Qp3LvEK6NJAXl8VCZ26A2QFkrY1OsR+Rbu/JcF5rPGk97eZW4lqTGzQCwhiAmK9i9ZILvu/BQMj3
YB8maFdl/l8eWoKHwRs9WT6DrURxtr7AcmzRTky+MxP9/ExejGyKDA9ui3Njsi7O1e4DiSLy3Jbb
ykHMFcyQhVDrt+bbPq9EU5qKk9tI7XI1CKh1fPZ7pmRSON5BtFCOrnQkt31jJ3BDwWDjaQ+iqdqX
ikk8R4t1fm1BleprGIyNPNCGELz08w5y1DSS5wjicVi3nR5upJvEaeOLaN+33yuW1oagIuoi5BRc
RmvnvVHwQHYzFchQr5Jy59nt5/f6IHbg8//PmWeyXAYaj8RQY3eJoZO5CHHU028Wf9FNCq0kGdfw
fzSS25RH9KxHrnE712VJxWQJ/82BadkGTVQmiFHMRLzc41ABsyNr9f9vUWNxfX3EBDh6DA845KYc
Ul7i1Q/g9158ejqRD7xPQKX+HCsK2iSQTJYZj8fVbEq4OoXaan9tQacsYtQJDihG5m+iUsFu8Q0G
kffP/KnYfypqo1XHth/CABWHzBVh0pkY2MI+vq/2C366D2w24a8RJzIIkU0h5dGSafXol7k7Iq+L
I3EVJ0o6iZ7thADJVddPYDy49A81OS72jKQy6V5aGXGZCK5UnVeAgWr6WWrfVu3hzXt5Jy9TsGE/
mTCuABOcHdgbiLblw8x3/initbL3boo4kDdcXVVIbzOjX2LFuBCF9pAh/HeTyNzLHw+U1VIPhd0+
CdIeA9qYQ80FnU6UaOPp+NLB95yNmCJHKnEAxwe44tWfRxg3y6QvtSqTx61/9QBqHM072DSW+VBB
abl8FElsQxz0XY3KCHFzjnXksKt+12O+lCp+yQXZhhQeHB+y3DOoEne+TGYJLEoOcDKJvXv6yRwh
m2g3OkK+U4MhdN60m6dfJRMKG5uSNXleH+u/16pAXLOepfbTDc7uKpViTKeq36rU5wPkde+MEwam
uDJhkLfCG/kTA9pMNYvZDGvT2jvumC2X1B48gBqa9crL2zc0NcTeWjsEaNMATDdTBewvWsuF6VTw
T6jVKOp8yzew6+K88vZPIfvsrMWaRMCtchLNZF8i/4fMoD3hHInV/p08L+zWx3wpSH1CY58d74oM
GLgpX7rxJCrsX3JZ+m+NqqXGEEB4k0ANU6+JkKg64bDbcKOUp0PZFO6nSqGuCn+cg6pJWqkl7+zH
BGacKneC2atVN5T0UKEDx8GZ2j4X9iVNZK/NhmzToHIV1OOeCt2w45jW0dBwSDLN9a+Bel+igA04
SO4w8SCbM/6IZ5K7fvHSA6KoXMafuFdOZNlZ2vaq5usccDOM1rg2vG9PxeSxKGbWuB492g881Tnx
rZU4kIsdupElexJQH3Wy4lc/zSb+aKx5h/Putfq+9WPzptKYcOExshXVjYz9AaqZyv9shHBsQAhI
CeToXt8qUSFmERlXuuSnr0jKP6wUidSIPDvlMB9/4P9kIGyuFNM4KH9e+mm/tc0ZufzfXjhfs4eI
3apxs4awsQOcp9Qz1VCjHSGIq/AS2T9LV2a4QF/0x9XQT/xj45+Obhx9FdFVPMPQvd3/DOYsdP1u
s+VFQ/7G2CjuduMEfd2nyYWWCd4wa32f8GOuhZPUP5bszxfx1hURMruoFzYNh2HjIwL/QlnY2Yj+
e2rUAKdedn0NjKu/8K2fC6eRqPfakhACOvNRA118wxByJYJOE0DNEg/XJhwWPcFfWiQHZHaV7YaP
RYhBk67thIz/w9cJXPIMVJEXLrgcFxwfbcafwNNd74NfFp6bLOl2KixpGXB+e4nLS6zfvtDgln4Q
XoYaVN4cBNLYw2gpZFVpPc1TrKFgNN5b+uXBDx0Ra8KJShuo+v0IJ82djSTTyCm24nF+Dgnix9pY
GTsfNqc6esbD9b8DhG+sKjERYgtRbTSRDj66nH0bxCOClYFcEpC/LrRnHHnByVYQQ3xBIOSlfu+P
Q4t7QeOk0HIseuukj0XuLvOKXosknCtc5L7trQXc1T/YsNHma7ooARqf0dcDkHwpAdGQaemloIZM
/SHm7KgrE/b+JKfwtYEsS9JH0AVdMHlf7MBrureaUboI8leQUfZSW31EIOv0ba7yehkuABBL2cKk
Mn+HGv+vgZZ8x5ajcqF8GlkxokJW8rD43J0RYdL1TIirYV3m8c60ZIXgAvWURkZbFXKH5C7hxrXk
KMwZtFoufPiO+7+qBO8u0T2x07k+n327cjthbmQNpyPxuBfVfvGvZeC8csEQocNVTtIezHnIeUgM
Zg7RhS1wfTtz2LSUQ6Vc3r9HB67eEThZVRRvbGnKHGpCZxD4Q+wwwefPqsGjQ7tJPsDaSMhzQGVX
fJ70Jo3z8BFEEsR/ShF2ICWh1WIbsQqpgmpb/BW1T3h9RB4AukoBsKgbDXiIMTnQWXense2MNWiA
LoYkbS2mPx+hC9lkW3LPxcbSypCcpL9Qc9F+0lCCpXx2nzusTWakAmoaYGBolhZ+E3yEDa918zMX
+EGjGeem68j/Rt3JSmaqw6osqSI/FA5I8Zjuaibw4SaUNTLGRG5xkwYWS8SPUsbXXQqYXiixxFQy
p8sl+KvWsXQIXhQDP//uv8/OusDnvnMCPBSBjxvPZu3TbH8Eo9N9BbASQ7z38dO0PXRh5tJwlgvl
V22gMPUoGXGhpOZmaEs/hRNSA7fP2Jp3QmV4TNTQJgqZvd7/X79QejyfKR0S/z6CsXPcHM3tffTc
W9GSsmJ7lglr7MqtQc2sx4+VFKhQQW2ZMjFb8k4zMp3EloxdJ/Xe2yHHsi8EZXmWnBOnBn+3TBvC
Jd38kzmDBqi35IQk5gDeZ5H7U9uW6e+q4IDvi+6//bpXMxvp7JxQcfPzzmDUiC2Iepvbq4+tkEMt
VLSCkoeCgLNEahsjmQX/EzKcAbt5xVmKjBverF8rYaxcev9ANmUpmGLUM+u1w/J2Wm7xPdSyc3X1
vw4bpI6mNwpxiBjfuYsj/I6WHrTR+sPC8RrSCDWm4uKZTn+PLkQIdek/dBWr9WZgzV6EAIAKQjNo
pZti/gfZTh0liG7lyCiPJapv71GwvOLknws3QhBgMFEnRV50oO/dso2U29yHRcUu4Jo8mfs38Bfi
O2vAK4IBNK4rQnREcvENTKP60AVoSu4WpWmIpOrssgQv7JVstbQo/qQEFBo+j9pL5IzLST1vIbV4
PlCddiSSoZaXymsvMC1C5JVqk8zt3wTcGE1r6y16BbXkWGVXhsXd0mW2npitBLn4ugyv+qJslqsB
AV+C2RIHAKKnubQwldfKAQVFn/frH+vKQ31210ybscBeYnESb/jqna2oJ49ZTIToRVPWipU9sGKy
XBs5IMAolayPvkF6mZm31bWd5Hfh3Vh9R4/nDagF5PMt6Tb3BQrCt9ajXXjqSF8Aq6549xcvZ/6Z
yVgWwWoUxtW1vWgpMlmUaA05PLhKFBy6a3m00thowls7iDNCJMBfboG4wpvyezLqZ5bx1iVDDBJg
NyE0plXyB9iukiAQJhCa3F35gQmXvSZSkEqGkC8a5whsX8cZwRE9dfRPXKADkqj7vCDVG3+pp0Tz
BQ6oHWba+Dcei9FoNqaeFrw+pmTe5BVap2zZUZSuArxErvOW3BMpTaAyAhdtmaH6akTjBUSkL/64
K/aWPe1tzitupf799F5MrCP1i0zQs11epzBKamOP6E/ig8impkOQqrtPpHhYGmVwj/elnmjoygBI
JmyYC/dVMS4lK2CF2IBeTmpRHnoSbkHdwOC+QKqPvflBD3OLDPnd5T/liFvHsDLJsZfVIBfVFX1y
pIBjny/Pos3/MdQe+k6jpRKdmEwIXfngbOnm8WxndZOIZzV8hoswFb0G0i0shYCfABGSjn4p4fDG
CTUvtNGddiDxm9wIRiJXFQ4MnyKkHQtkpZo4+JxOLyL8gZ9gnPIIdLosiPKqYmpfEVronF8exCYT
72NEfiWfpWybiLQ8eIypaRKRZ7bd4gVEJi9AxUCgqIzZsnwjIS4CrOCScMgRfxvyocE/o6YfFj+o
RWWl28GWtIN3lqHFpQssS0PRHFKxO8CtlMDrKvkchRMqjYLjc7QR12foLABx1IfzfzLXEaIQrGop
ukJHujAD9PZmfcyCGWt09jZs8CvKX3QKy5R8pL55KchUo6yfHLoZqjBxbZOYoSM/zW8IvfaPq9aA
h2xZrsyhhxoHJsT97UEeaazOoZA4HLOLPjmu+AkwrfucJ0ShwzSb9nZg0DA00zSnSmMj8+2c1MvC
bYApTJO4T3fvHXd8qmPPwrVdO4vWbjvvkG9RS5AZWqzpT+XexBenOVulauyoNtulWncP0n2+GxYB
fYaaaaokCbY+Xryrr9gEKb+WulIQbbeU3QZG/z2n4DmBR8bouUDPth8teuaGzc9P672AlM17aGdy
oATWG6H2eeCmJznU80UyufbT7hUyj/lfxOwMq6WoSJYEWtRvlrcGyPDBmeLVEMGgyQtIVgLURvAi
R53Fi4JPdOGWDfrAkKzHO+1/z5+VjTBSY6FozSfWaBUzBIve/IjfZlWYZydkCktYAq2qhXprB93i
DoZmIlJgA5TsFOusPpgwJY8YHsYrUc2GcEjnZwSK850xvpzZbQS0myaTlZTOQEv5nutPI02mDMU7
pfxxbNTa9WqKh8LO17/iy+X4kJ3auZjGMD+wNDg1dc8cWEWhA3Nha45c7wOBy2VD5gbf2PnJNqQ/
M+L9zWLzNvk5ji54zwkByvA3jz4YjkfLiPOyGUtqO+yvHUj8oLDXmqVcT2VKyIeFhwLY4Y9lVvTC
8junUgPTT3CG7rOxpDl12yJ06HXPozlaz/fWjdQAL9ugf0WdXyBzjjS6bCKgrsx2yhyZnZQdsLDN
O8jAn2lGgRP8j6X8vFOLPxLaEr1dzd+uACA/lYMvjebrCXqQcFnH3IDz0XNx7TuCKniqvr7A+4Vw
ScR9J7vFmvNXLcyfHYrqKqhBDLNQvxfw8u/QTUHpro9UKA/Ld/ey/3oc8wleVFX72kK74+54arrW
4odJ11T19zcez72VGmrfhn7QSrljv1ZxnlHyYv9VnIoi5zCyAQ/ddd7yLZlaHY/Z/pD0AK7sG0DB
bffq47TVQYPwUmK6TuOvkvjabIcAJLl65lVOYlP6fMT1WTZMbUdXDv29GMNLO1Bt9obE/7439NeO
6iJjD7+eA/WmYcKOPA+bvxgrPDZkpHZGit/ApyYK652PvKpMJ7Murvktry/6KVsq5CWHKksT0Wcz
PnzR+fOmMjnN/+F5GwDFzPKxX4UdLdEsRtDfGfgIIDgTXP2xr0gN2BzjPnaGXB1bbPztytbzu+FT
42yfHIxQFODf9/hNyNdJkig660J1DvDshDyzns2mPtUuGLuUmuFwUUhx+kYV7a8skHxXwTK1EagO
gT9an5JzwdhmIaW02IaxprGs4MAylQwMqlsJVwbsgoaT5JOVkhOL8CjhCSv0jjWgRk7K196UvXNU
JvD+FCAIU4/f9Pc5+gG7yKaDxpLPn8bXksOU55iM4wZI+xtCWqc4feLn5X5NvIgYQubdy7bnRTEa
AM5HzMCzb9IYdLSjdz7iRMRQmsN7QnN6hTvfO2RZw14/To2muMnvVydSWK/vSHeV+hsbRIsTW5JU
kak6y/WwvNvPXIoX1nQpBdPaxaPkFNqsjK7y+VgfnHH+GaNae412cN5kpclVc/PhwxK51h/wkRpe
0bCWsbKIyGF+Q5NHbjStBi6FPY1lkEEr/8Q6dg+BHzR6pufg2XAi7LWwLtsiAUUSN8ykJYa013qG
priuWl0vUBoDQWU/nDFriCEbG6ukIcpcff54KY9SISKHCDqqP+U2qcMXEX0mC3tmhh5M8TCnjMDq
bYtkj6FTrNgKdlpOlBlZjb70m/qDHUGBNdeX/H2hhcE1Pt6cBz29198str7h3Ltnjk5zxDKl8Bw1
D5lyK/2FtSbltU6jyNUlZgPmwtwyD1gVG3GGhMutitcOL59eUThOCxPQ950jxsORY6m/lCPmdU/k
31p8hI+7B+AqlO57rRDebGvs5iK1DJF5pJRcUPvbKzLwx0oHd49gbfVmy8mogZoPKcHwlwDb8v2U
rRFYEm7XxJOHxxvZkFgE55K+acHGkTTWdmagnNbTTPaOqZ9fF+IGAvn3mBtpwBe/8GRDZ3chGMQZ
yJ4AiA190z6JtQnOUOWfO4IuMH0+ibyEeYy3wZh4j2EM4vlZpiGT0BOlPnxHBwxn9D5nNR8em52v
Fpk6fMJu+thNBUH6D7JqdzKIAwkq/briPCaq8mLxUcF89gbK7QsKBAB6Y6A39XB6roF2CiTBCXUB
bQaCVTrh6OKqu3tV4GyrsUsH6jiDEi1Uwf+z7LSQaGuZMlvAkzyBPfxHoWhs+xgBFbAz+Za3vo/O
EBmaU9tXHSrWs+g6d3nZEea7tmlT9KrdILIpafl2N8MVUDJJIkKjI6ZFuAzIVfUGEuBr+Qk7Kh+B
pZ3OxySyQmlrv4c4H/Cgdl3GNXjspifHJdF9Hx/woUbxO0eLP3d+78yR+93FKbZ5veSGCF4t1jcU
cwnQXQ0vnXWXabqCYov1yUS2MkCiRQZuWNShdnAIdCk3dpo6OVaoNrOk/YDW4uA3pMeyNYUh4A0e
pnMYDcMwy4TDlWKH7paiUXRwR3tB8U4MbTNdp1zC/R7fO4o0v5hPtgqE6YTVtlnwAvKeWgUaHnE6
fuYg5k4smCpgzoXEYiX7A7slHGV0KAaJD/xT1aYDmPjUWvL2zUvT8E8VOVN4AhbA4p9dZmk944K7
wiZw0fILy2vVPVLY0OGOFMRF8eE71gYvmG8iVeoUjpNeJZOwtkb6TAlVmo/QWll+n36eD6ctKnY3
HyM1AJlnr6c/lWPOZIqTWHn1/44PgSn30vbw4mDlGLv1F6vx0Sm4qAUQjQeeVQlVRKiLpx2BqmAb
6KDKNm9vDFEhMyW1QwA9/HjrJmrIH0L3rMijzjlKxpWSJVXwpo7duV4k8386ULMj5auqZ7gragzM
XhzLD9R1Cvzu8bkjRNmUhaYC+6eHCDWKBr/Yt3c5e6pZkz1/xTI0X1I2EQwJmqK2jxL0ah4uLZfU
82t+c+b0CRLDYiDPfcr4JryPYfgZC4JHYNMFb0cjl2cH0VhOyjGo9ceqqS1hjSfBfTjnKz2TpY08
KVgAqE7emKUd0vHkSphNkjf8MSPNTpPRlFzOM2FDCpT4Lu1t/c/3uJ1+uWt2zeMZj/Lh0ab1fUU2
ovPFzk2RXyuRMNV8BI/SuwvlzY5f7sluZ7zf4h4xzGdKkmBk1O9yggYpy5QOeHGqIWBXM1ZAo1UJ
QN64VHXPC1MqbD4Nsy7s5awIBrBZD11EJEujNCgcnjRZOsPunvcB/nt6xIQrLMnACYI2tlIdZqld
F+srfORF8EE48pnD0nm4pmP3OQTbV71GIa08D6WKE4Z0LKGo871BEbPlfMuxz12faRefIz7JB2LI
kccM4Ns2Jbg8xft/8/Ja4bWeMQa/yfBFj8RxyWampmJGNDYxoied6cWbollxt1EM8f+PdQw/8/IO
pSsNy/IXJadZtjdO0Bzd5U/HWkgq3WzmdaqF3jMzty+7r3MKxNI3lo6HH3Nf0ot0kTDGASWlqD21
inP7kO0nv4ZaWyQxShhWLri9lPGqIGJnMFk8dwGGXhkZ6UWNsPUFB7PEnS0Mi4Vzc3hnBrgoxY8x
ij7q+mtPL0v7XnabBnwK5WdPjFKJEDaR61ndMzZYwAJUJuHzuael+aqKHswM7TEBxriYz2O9eLqq
PZM6vYaFFu1/p/A/ZcUKzowjmy5Do5BfmWtDoIt9GIIHj3jweIqMQTXp5hqzJQ0wkozIIhQlmJZ3
YiqYFdyAeZ7nj+NgVJ51Z2hmLNM+ZhLa/bdZQlK3oKP6h1uExbsh5TdgChxGjHnIcvKhht8I3p4h
lIQkQi56IEs9arY29sH72O/Vq7Z2hsdMZWl8v5rwBEZcoYMTTcXqF5m38TxZsaLL+U3h7tUJEsAx
Tl2H3LctRt5iSw7m/w7Vg957vDvgpwXyx40fvlnzrPAr2J3HnBDvs384LYkw2ilgt2mvBZvRXUxr
chkImAbIJXnf0nsS8bwfN3xHsXO/+LRaqjkLG+SaKi88c2Rr85G3sW0cVUO+tOGtWhbcZuauKhg/
VEmVBRPoNpdNSxkgl7XZkHnegeuzuQC4cx93ZmgWOPaWNcCLp6bgNE8dj21WOrI4bdRWVoEShevL
0S1pauJBZ/Msfu2UfD0kSDwBWc9j5yyvQWEveyluqGv9WU+qkDCo6YuyBAizxSU5+ZCXvNZNqAkn
m9C33aIBUZP5r4Alga4PByzCrVLwL2wby94f5GVAFw8uyQUwaPttIBub9OgCLTYanH2U5bd/dLgj
5A2i5OG3tIkko0eIPN9POGceJQM2iFX9CBTWPsRkvd2sEjkxSzrZdaX2HVwyqL8Pz3c+mEk6oaSr
ICQ0/sd5+qHYEXSqExbyMgipmQbeqf1nyAzK71hnfws5b1f6SH8//zbZeqXlo5pZMQ05+eu9vDi2
sFQZZzUCOVcY2PISL9n2rFGguPPchhQJqB5BOuqGsQm4+q8jBb9sLz9Jt+RvydcA0Ptsa83snswK
Cxch0Xu76LhNcdVtL7ZG4XD19/YJ01YE+Ns504DWCzmoI1OJfouuTf879Bi4wFO+q/N2DMcEz3h+
hGwiP6vwefE1GSfmfjNnSyYCqhEF7sT7XD46bfQ0L1p17ux5gyLIDIC9zcXn8RUG2dMqSqAa91tQ
sUK2Mcr6UjCI3bsnpBNQtBJhTamIWLy2Uq04vSuhgIYOmW8aHihfbMTh96w3FeaABbpaAr1K2XwZ
aKoqgtEJXYR8DIXg+KKzVt0g6vzlqv8UailmbUq8bnWRb5xqmfQGlJxl6rJHtkoTO3586hH1u0O1
EJ8NsSZ0+Lim3Z3MTcL6mkqY0246/t/Gc39pWImDzLFl/r8Muv3I8/Jd+j9bF7MFY+NLBXJpkKDS
eky755Psg2nrqLqAmM7oaJCMzafmk7WF3aS+oTwWx+K3HuFoYCNF43gIH9RM9zDXXTBujup4m4zC
iy/ze+YNRAZLUcvdQn24IpHqJr1BGPdumZB8KNDzyk+OW9QYq7CxAsqWc0+cxa2pHPVOkoMHSl/a
9syf/k2oV6R5dlp47lFUJuZCnEtKexSaI8/s4mAhwsrY9EVpvyN+p1BcHosMRKpySKTmOtC+e2WR
nMrpPpf+l2quSLWdOapDoTcgN92OYsPSyQfcSkTP8f3ipL/Y1ryvAJ6ufzcdtdBaH33s5FKOwtiS
2rxikju5/EGW9f7c7kVLI+oOFv4iE7gC/F42FCu9CMzNsyiGzgCzOYJJBt8mCrE9kXcvydQx0KdV
4gT7ynbgTLX9XzFVSjQHORD0lltPpogZtW7q+Hth9NTy2EyRz5LkVtw17ohI1MrObwzSdSgE4wFk
B6zr8dvYCAMlFBSG7Euf5B3NFHQZ1iK3PniDRqk4no94UW/Tten2OmGg+szmpQmgU6O/4GDuoGqE
KyZDKZK4vc3puthL0lu1EMrK8YLgzbQqry8djtjzJ6bHEnCdx4U5CCKsi+f5BhT57TohMIRhRmHF
81z4tbMHqfpzJt896kHkdiw71tcklKuwVX16tnSlXeBVb8wD0R8eIMSlgPmUcMHNMrcxVy4sCZir
TsaAL7Ic3homNnE3e6jh2thQ4XZHdKRbgKrP2HNL9b1WVRUj053WyIXAA3Kb29hkk3z6dlHh92v6
4iBujaMw2f9iNufEwRO+qPcmotC7UqcP+4uR5MGQmk8UpoUTB5hz7vPUsKQkr2DdJfeGXqFWLcsy
EIwY7pKw0VGBK3H95rnbz9Ywb1vnoA8BZadjjSgw6h0bt3LspsLd78uaepdvcn2zDIa9EpcGioSB
vCP71KHy4zijdu+gbHcjqkPJCUfdT/1fdGS+elvrVcx8cY43tTxaQoiAosNIDQ4fTFkPthT4xdDt
BmEVV6bFqy9TtdxBJ0VlD1W9d/i7kRGw6B+9twC7ltqePIlvJ2yFYfVjgmWXJzpg0PNCnwVyx0pw
u6wt/8XxKZCJRkiW3k+ARuFkSS90rA3kw1/jdSXRVjh3rcR/2KbS8OP9uA/pmtpbE0JYeP1LDIRL
3i1/XtBtohNAhoH01zNr8xlibTEooiwUSh4VMbEXjS7jnkIWnaLrDeQNvpp0p3rAhvKAYO3sPFjm
o9adycPeIpIhXpAwBJ7po7MbFUDG92yQgZcjwTHZU1uJBqCC2/X30oQwTR73zlym71XThND6dMyj
O+/oJI1dAsVQKx8FbVdkapDvjYtxWwdeEeZ6BWFnw7A+p8YRV7jp4YPDOtcpU5rnSbbIQVJ+Aqn6
FI9QZQvBgItwwvgg6adXKVrpEsSEj8m+p7HbPWrsFp51CUK+Cc4YwLN/MkkveyWf1X5DZt3ZuDZx
Hz2aH8M/xEVc8iT/Trp4hARzH7sx8aJNt5uE5v6634s04DC/1c8YkF6M+Hg33GYxAlsLdiS0jDL/
seWGwDAH0UdQAdN9WMWQvwCTWqPDhZIeZj+qHftbRiA+NDIIx+gmIN/o7uxM1MdqSOrrr3s/Elhr
6/X+t+kpZ+le93qwm7VLxDC9Jfqmf5pveGd/qu8QLCtS6iixVrIiNWKZ+EH1Dh3yUoIyTMC44CZu
xCCxIWMWCQACLB/TRjVHJcWrsprKFyJjUohXI2xYtwhCSgg6YH7Iw2BTgjslY+Yxe93e8aj8L3W4
vMDf2hWDssNzvLM3555y2j4RUAL18/ypdSzmxngkZRY0M9RHF8SLWC4QN2hoE97u+S9RVGJ65DRW
dRSO8QPBfCe+H3Jd/zW+FpA++ozopGYgLTmKq08RevHJUQLpS1KrP4WSlSlMMguKKCTC7A6SLVD0
/dsy5FhzEu5rzACElTUcffPzXZXzsUkgS2J7fMh1pYdWRZEdvQ4i0nB5Z7VahTO1OD+uXhVY+bxW
hI2OFYZgGnM1u9CyKAWZWwZ9sSkNx8rWhT+peV67RdWaNoIMK2d7Yf7mupaSm28F0LHmXfKrNB8Z
L0GFygF1cvg9c+2iqoKnHVD+DIN2rs7tmOghSXhpPl6eJZk9quJvYpU5rcO03erNZ1+AtxPAFa64
ZPcwhM0DXSt4CrH2oQ6rIqE6GlLfTIJ+wA71x9ytJ6T+HUwQV0YnjmKlv3Z5PqSaMHhkWwAppzTC
+Sxoz1HOsRG7MownEJQ6Yx4wbLRsBG28irkivNe3Lo+WqvWNXHYZZDlrpv5aMJ/dWEHwabrDyu7g
gXbGrMUuxaizfezzwZgdYISp5fLKL7R2eqp9/w247JvpfqXbmEqOLTEIJ8ABh4InIKpKv6uz5u74
Er/jHHrKoVlwKZQMrB52oK8NsXfsMJibQxR9B/64mrxSjMelV+X/pJC1EzMLIxc9dq47BjfLshkb
yuIMaHm6//P5rqL80m6pDej1wM8iOiFm4ciK9R8Y2sSf3xH6MrxMPkTQV0Tt5YhH8OhFWyrprE+D
vlkneoTYKOEhYs7VfkDZKBLMCBqg7LkA5v2QjZfQIdXKZzu9qe5FbVOr9w9uSRnygJj07uz2dH94
lcDVkwk+JJ/SHhr7VzqfPVqH+eb48J/EuUdQpF12m6zJ9oOJDTX1eJvKxKoyQXkog4nOzpJ8IQ7o
JOkiTVdQkUPPFJTkEzHE+mYHYfvgld3aD+L1nyuA9xTv3k6nPgx6K7YQron8/bNhRkTj5wXKeC/Q
4UQOXue2dgaSkhIYXiYsj+9U+dot+0CRede3RlBJaPLxqL+VDoU4gsJ68u1DzzCdlZyFDvbVoNPf
ikobmLOGF6nVPQESwe0IcnP4SW5M/VFoaf+OlBZC2qCz+iigUgsRSYD+fNmBZpCSgBcum/K+pDsi
3kwlhKIaOhAdqj7+3Fri+kCOLqP9X9BNUdPX2wdB9hDDaN+kkUPfaDPMG9e9Re/lMek4vwuajP3O
KDFTOG+lINDTYXCKwXpWgq1HJN/yW5gwOhtibGdf3RmmWcOFxWOXrf4hstPDKSG2WBZSfCs7cFFj
nzwzqE1AQhOXXGrjAfyLnoLQ3gwUnGMvMa12Y1BgOZa7dWOnc0GkZk2UZOiz9t+CE/DCN6XRn7OO
QBIi8TH8dSMS0FvH6MmQsL0uwTXmUwKYl4WEyANd5ISZxR3hbnq0p7f/KhNLrrInOq09EI0rpSJg
cjnLRGkmD7p3+Y0kJTOdy0DvdHhFsJstJxUdUgYmbGC/j8LVWG05aJIblLovAidnKOmCCq3rSamQ
CI7AREbo1E/xQhcWio1t0gefqBHvRD8KdwrutBhJDr7U2inciyrqnKCvfg4e6AYHyCGOZFRGDbOY
dIkocf2MgaVPpAoND/eu5CXuaOdsBM2LXHIGrHcSt9a7SvIJO7QmMPIA3lg8bYVkAmtCJux3nAZD
evBzyO4Pj9ftyRvLgWZvVIMjgQu8Sw7y/jA7lZF71ES9YKIDCV+Y9HEUMeR0mF/QzYZxg8TKJLqb
nkgAEMEz/Zz7pZ6iLy8kS4I7r0TENmDm26F+aGB+ppnZg6pLiJUeaCRQ5krnBTKpzVV9sF/gEu0H
kT6v4nYOD26lHNRuifIF34D8tI5//7dpXATSZQsv/BmJ6KYYYjbYIjuuLyoyo0eQfzRofzTduwf8
5sQUwX4w1cigbgjzwjw/zHydFUw6vOWIJBeGTiDkCnOVn+iyEQkjU67tCGQ56MCXfRMDsaaJAz0E
mxGDq3F/sGXsxtQ5ExVTSaCilfD1gbsfivy/U0kNX86hvJIRcoJQlPsJ5yVjmSqrIgqgv3/idxJe
QeFenHxuC/gUYAzuFS6Cz4NYtRcoxPiJStbxHHzwFPIe2+NA9yYzNfNWwEnol1yZexiSuFvXQXlt
OkC2B0QeKKmfisLye+Z59JMHTXrxF5boBz1s6rjLE21l4Ato6F0Vx0XkFcptTkGEk2jpDwzl7vG1
+g0jeTcG8Eyj5/gprJ6ubgpr/T+Pnbk6YqzKLgcNuz20bWFNMO++f366s3nLFryoTqNw15A0x0iI
8hAdO+ndQ0o/jTAQlhjFdWvDqYFMgMGCrqBf8tPLuTQT59lPaViBDhLK9fN+uOMHP5xdk4tF1cbu
gHGjmEzNqaBLqcMj2i277Zj6mV7zV/9urG9/VsBxySv47oYYsCHdfOdKHmnYI1QWLZyNOblWj4lZ
F8+epw3/tWMhvAixZc8p07fLUgZ1K9jn14CRSSGWaRNfrKfvIk8ywL6wB+GdY2nrp+r7qsA5gFNr
0fut7+4ERYG5Oz3NunaU3TE4NtwB9rGZ3h4iA0JOSUYoUt1cGdWj6JpO1Z5nGIK3slyFLTcg3XdX
3MeSQroioSpCU2M7ea2bkwVMbeBI2DRnNRq8GO5RztZQoYW4sVcTCbx5e5IMZbDTm7tbXlLBqCw0
yC/bY8PHWBtuFuzC/DGMAtdmUArcjNsUvo0A8r7CrIiD5qsmr1N5F+t3OZ+dhgZi+xbpiUPED5wb
grtYpMaG5hYYupii1gypkUWoMVHr3CeyQjuUP+nZWKDWKggGoLgpCwgpCoT8yPgH+vzl/DhVCSul
HHP4E1R8Pk6DCuyC8tzWPRsyqVnYxnOLM1fG0tqDm2oweEc3nA8bEXTVM1EPFDVvWddwG1Svuo5W
TmoGdbteUJi5EJrsvn3glVK/1ErTzQ4p4dC9YM5TtW4mPM4kR1blnqSIu7qJJuah76Kkd7UoL81q
BOhAe51m8Yt2+Nt/Ak9rySAw/OoLEYwrx6MXo47YdtwIRsGDttv4YBr6WE6QlzlZOtkoe/QAhxmY
Q8Y3YhvA6B113OnAJzsc/TtMh+sqPmRCNbkCfWlnGM3g1xKjlULmE5CshuYEeK+jNmanKg6EdheP
X8tHRI9Rsr9aD1tdwBiE9P8PPJao/lCiQjT+gxCB5mmL44ltjbGT2goT+jt6zjoGxvAGNV6LBo7r
iHEu7hQ32ukOtVINuajUfZcsAWJkunkQ76edWTDMBaMwhRAbGJzlAHd/r+HaDJN37dp9m01ZLUXx
JfRsIQUdjIXmLKUcWQbapyV4WH8xVE0VD9E8VFMDBTs/lZ47J0zGbPQ7wbeR6+yQcL5DpG+H/rz2
eAeJ0UUB8aQUGtr4M9h7Iy/Lbz7T6vt2EJI7UpcE8z82aFXV9k8GfMQRDX141NLjIzSUaC1MJ2QW
gEzoozoRi1oZPab/RjzrPwvPsZiQrHQA2eamzlOD9F2EH0ExXfdROdEpPLYrQg8lKght9KpLxQ+/
whrVI9DzXc9JBRL0B5j5DIMVmiun7CtSGzh6no1KqC7nVzZ501jqtGHBH77oZj4AeZ7niBAAahXF
IrODXBkx4PMV0+6GfYRxO359EUXyEPbG26f7Lk2/pURvjlWtQQDIzYgCKJOLrrmc+U8lR4qUAE+G
Oj1A7Vx8SgBtaX9bjPtUV6F4y1Ey2IW9WVbvNHxi5ZPFTucHvu5rQ96hdRTaiyxS8Tl2+FJcOOQ/
EAd1aM8T3TLwspWcvnBiuOttEDIwp8N5Jm0Bcy20d2LR1FywYJeRPOs4hOGtqtDzGCmlBfgNVNL3
Vm6NTjHP+9c60tuGn4G3H0eicrnj5b+AFzPA/dkO3U633vbBdYI60mZVvhlrApf66ht4cP80W0el
DKqKEw8kIbW9XE0iblQ76yA1sP+Fy10vsHlbdYTENAWRbaErlg4N1UW5yLpetWpP70H92qXWPaPY
1mpfjIgyJ4E0koReVLzowMk3DqOyqlWqQhEW72K4jgG91dH2QEiogbe6kYoDaR5xv6+o1tF/LlqT
IRDXgT9ooLk3IDL+snbeyvC0bJSfawGIpZooT5ON0n2i0m7gqlXW096+sn/SwSUB6XsJT1G0ka/3
uL8UPswdSOmytr0fyl6V8kc4tExItuwESe5dToWKK843cIOpphb+XkmamnX9kSyXhw24ySCc271Z
9AbKvUhcQglWaq4GJNknToRE0SnXjccRC4xtSWWbRdio6OukD9hNTNIWcr7UTRkE6qz9MF4fWPw6
/Mk6nybsjuuYSp/zNS/e8fNEOIXXsAqaadc8jwvJNy9EpwPysg3HGjdIlMRzdM5hmeUJN4XI97/G
/4exyfmmyY5qBbJZ6nXyvcADA8F9YaqwNL9osxUb6mekk7bRE+YfFibKYwaub/JkWlOXIABSyNJm
OBEOjJdi7XZoqvg3+0MLTOG9vdWsTvXZx9ke67XlWISik21byDm8ANbrB3jCPeS2GgSwDBt4vBQh
WZPydaUoCq4o6lYBcrR9ZTJM+QDI93G73nYq0dKaYI8bM5FVgtkrVsPv7dK4SmOMemIigR56J+oj
QnrnkYJSYl5fWoWKz7Y+XpVmYVhqFKbP1ftDJg/J5AqSPutOZpzh58/flrOBOUU1n0ohHbzdAqPo
qVUH2gEyA7FOazht4foQgH0vNJQZ/isycw8NFl69ay+TyNzkjyA5j2I9ci7+9m5YFbFZpva8XgcB
ek+UP2+szbgtP5M9s5WQywvCrrw7A3T8KRmidVCIZEsoMDhlPzJvAVCsDnL55uaY80xPhFnPOpjD
RIdGtQlZED8E0A5/vLb9pUt4Xyeny2kULztW4YrAJGMqaj6Cy3J3jAAl7l1qjTgvYK1O8NJ4rFJZ
iL1xh7BOn9ym4rXGIeTPBbLpuroEK9KPGa4BCptP6tEQzejKiU4wpu4tZrC/Wx1OpsyabDxyDgfG
5V5xISxMUxohK3D9aOvFmo6rWj/NOvCxLXwc5fdLjAq9iwqWNC0vE4344xGoKIWyqI2WpGQ0imc+
X7xJLaaiTZCI6jB0d3vrfF8stzI3nEqiI5TPnxgePmS7rn0jfSdztrSkfV53DPNiqJcTx1oImoxM
Z+goZNAqgCRlBhu0cnxC4VAEqlrFgsQaNBO0G5K4IWIAKXPFK8pMvzyvNYWPbmyAfwh8nfxfDyAq
ylKfw6Y4IM/BbBrhshEpqGs4k9xRVWtMSIt+rTeCPkslt11xP1I2CJip2jb5iaRhfL7BNl0tvutA
Yx7QpGpxRaxWVkVC18rN3Z6rj/U3weJUUjKmQy2LVOtal8Aj6cAvQTmQINyF5lsCV5Pp36FY4Fmj
yNME+w56j5bpqfDsa7Th/AFkTbduCFlZ9zeRJLYL24jHBBV6RjIm4gcQm1pPCV5WvrlfE76VOPlR
SNW+2Zl889mJrYVHXqG4QZnGclvYniA9QtU2G53RnblWRZngHKby50L6Vp2uEAMNG1StU//oI6tk
/etAL6mI5YsOF/3KU/hVlHCCtmKWmqf2hT/z/7CwahxkZnVIcgSVZyoORcKyAr0eBHSLOjuHoIvh
7a1I1QztaoakPxookwJkBu8kcqhQX8Rx/P2BdPqQeYgFt+4YVy9bocoMl97chex/rJgGre+oO0Zs
gtatiUNB/23JCrvw/l7w7YyUODdAweT6gGH/6uVOv6HZIrJ4awhqKegtlF5JNtLhto2IaVdKje3K
RvFnCBFyaM2Z08uNVbWI+Ga/oFMMmMSlcQR4b1iJOZ5X5vwwr+5aDpWT9BslIU8VRkN9k9r5G9nu
pZiE6qt9nnFhVqt1Qwy7eGpi+hE8sXtG+CoyfIo80wEgZL4gSWS+jWSRd+0IgrC66JWdfJUpNq9H
2WGhQJRdP31MSjrA97LVqyL+fzvJEMX1umQOvNLpF7iS2S232nog5bMq64rTznDxso263L68mcRa
7ebrrTJIfZC22qleX7tQa8KXbjJWh/NEMSzQ2Fmj7UmdMdfYu4LZta/3iXyUBFlbcm2/cCT5aKVR
m50r7WQ+6dzs0lELg3yT8PoJ2wB7wOQ7mzSr+MQr11SeyhlBg+V9EuQhScjFZkNNlorigNtyQUZS
pUBaPc8t+dvYi8HTJyXKm++obNNzW3BKtdFJynGV8m+CwruGXsvSXD5Y2On3rE1FBrjUbaC6oRxC
U9hV/H6mq7356euiFxWWXfaN8nDupKulBekVM/tHsIkDKs2D25uLfrnyvAR8faiKHeojginACpso
1+XJ3JR6G6yTZAJxJja5sMYbKtlx6poO7yYyQN09nQtfoyS9+S3tmjs6gAiD3bK61o5RAITwpZc5
M1YsWIrpt6BpUZuMr4D9Ixvk+pWxhrhU05Ke1eAP5Ohhe5slAUz8jKTDstgjpWOws0HaUUKHsIU8
Z1FaPHG4Cz5m88iFnwM96GHn/77OKgnCIg==
`pragma protect end_protected
