// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
N5MQFoqJ13acI+TatsrnfEWC388fQbhjFUAbDE4moGyk9XQ4NDyVNpcBWeEduyUqNZIXhSY8qDti
kZ5AAFvMdiNoxiIfmJY/VC3ZW4k5h7kv2LmvQQUqUIEjo2g8mH6n5aO1m8cpz79dcCrGEZFvB1x2
5i2rtO3ZgGvmKQ3lE9M1teXFTYHSxcZXuX5glKh9AtFpy4eJZqJbPELDQ53p9/Dmx05+5ZZMSbVi
2+Ygwx2/a2oGAKKqCwF3CTtqIBQiFz7cSZmUMZvxHyO/uu8BfmB9ypM6U69tQah/OvDCfKt0Eq0R
u3X6Vcc4mVNbJ3G/S1FgNKE6DxraDD1XiJgG4g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Z4YMnMndUMIL5Vw0mAF5xcgBTVfgvc7WQ28GB4GQ9Ku2R5B5KEGhXRx9I1YsNQviwoujbsb6XHyC
EN+QvjuNGWEBVBR04G+B8HSl3U7e97LZJg2An8fL0sEREtSsxsFphFydijluT+ilF/9qW5W9byh6
8MpowMLWnBhuLdvUKUQ5mxA8yoT+U63sSsta4J0b3x5k43MRLsz/zFwBcPnXAZKkz8lbwVQWce17
un3eGfnw24TAi5R5c+xZnoqGhWJmY/+DAvMb4N/sg3pzG1FhE0hh6V9U5DeTDt/Xe92fBDmcs8du
3uJVCExODuOc6mBedbG8APlyEpWQzCHEJhQ5ZAZbxCvuURCkDbb0eZLe7YXmJTyHuRDsr3kroE8E
s0e+fE9lFjasS5X80+4Wz1KzuWiMDrCe570/hzQQFM6xyPeTUJ0oHvIlMAT5Jh7efiA7OXbxFLa7
9/nDGS3WSpN0zpCiWHYnTWMGgPSc4FB5ZtYtvMrjRPYnzRsWslljRz8GbJix3D+GtJBrVfY1tVje
8aOCu5KS85XPIKv8k141x5WxLXHmzayQwRdi/QP8gIKTSQg1r527DtT7ptwSxGeo1atIXPMK/INs
youKcrViMtWUCpPyvtke/H25cj/mSal4PX8PnLP14vKc7v7wbDTvvCbXeZh+VKVrl39xAZin4mfV
Zt3nk3/Q7XzqASThvGaQ7lbTZdFexaosk3hbBiPWcMRmoyNdxi3rl8QvmqKfDO76M4OdZxoAfJJM
wOtrHxnaGhwOoNdwz3a/DhM9Z7B/HEP/Qf1RfPOrjTMKMRouCfj2Ujnz0WoENw8WtigTrW7eaYtI
DH0npVYjYX2E+l+EZK49YICjkSI7CIsRA9HOAiLpuIl/YSjdvpsKJbTQ2lZieTXhF0Yg0IcwDxIE
V7RSRGV+lKnbT0gak/YOyq/4RBLbgcfowSVYECOcOVpxB5bBGxIAE7xw+5lcStx2rO7U/1YYBRDj
hvBEAcXBfIAqtyEIjMs/ncOoiv2gyqmf/nXDg2fkLjCPIyxGKdaebUqbk0Ug80EGFb18aABat2kz
IYXweYc+9G3KDii0X33BceOXXW7xsP4kXUSDeqT5F+3wR9i8mICaCg9e912woZINcUb/X4nS/qce
ztpiMJh6dSJQ6xClPbY1C8WImrcITAocvgtEHZ/lDDkJ8QXFEAMGpDEoK3fyu3P/k2IJAM5syP3Y
nMX1bSIHrdGkAvSVxeNjTixBDpDQGufGWBc3PLJnjLxodRe6TuJ9qkCBquLNaDKkCJIeaY4Jp9K2
PB+phYH+hu9DhCGHtDs+PpXMks5IpyiAbR6ajsltp+04F5CUmqSPlJZsPGQL0L25KmeaGA2WpJhD
NB8ycSSiSoVBXv7RlLTtL/DlRET+SRsRspP5zGb0QFyvj27yhQ09NaCS5wyveCUDOCKsUzeToc0L
2aU7/rngeQHi1Hijfs2ppLGtxRuFCWtHWFXzzhWdj4ah11nM1jmuiYmdWukF0yRxV/bgWpmscAnH
eliV0wh00SNgeBp8jDAASG/W+L+oA0FXeEqPOQw0Ayov+4bAGDcch5StCForjSuHONEp4y9Nt+JK
3m8huXrEIco+5MNUYD0OXglII7WcQTNNzy7wpYZ4iDnm5GnShBf1ZKZrbpRcrn5r9+x9o/BzV8Wx
MODXMln46k+Zro/0z6Td4e7UzTBjrG46mgQhsEqdWqPQQWC9/VYjszwKjG8eTdIWvnntfpdIgVgb
8ugN62B+QG5Xty2WbvNFAztouPirxEA+IzN5WWFRGhW107Id3nqt7xSEtY/B+VpuVq1zyURTY0rI
hSYTBv+z/dTdCoaGM4lAAyJRF7K658klAImZ7D5f43liM1h9FTXZGtldL93Q5kNYsbh1ik3lMuuY
JDKhhDxoZBf8zLgVa5O2J4SztlzE79BbHzuz5SsrzQ4iO8jXeOnqW2RHlgCL5wnvCpDu589Rg24f
IWAFw/bgfsGd+4t9wymxrm2IxRsDf63/3s8fysZelOSATIF00Z+OdmFCZZoRmExvmOzMGrRSzoxX
APWARyolHVWNRY8MTKGxOjsLbc3YFeP0uuSKCarBtrFbIQiiGCUkvQAxym+I1LPNU1J+zZk2LAT4
mEVUfF5huyetpYReEfQQsZNVrhX9ngeegApWx+FPrFp+8R2ZpfB1AimgFu6es38AK00UJoAT00++
vpn0Vaw6weIJZaPP5ulYJHPznStadYmzme336zulh1pZvQHMX+kiZy2Jlmuk3xCNPaZgPCTgE2vn
LIIxqThKxKCcqogDwAMorPlNwuiB3YAYGJa2wrOf22GCC/+oZHonhC0r0LErWgoWYxkq9jiQjt3b
6lOetPxoD8e5kBV6EbkUWHXHxnpPjc56z9p9rYpyT0T/e4s9d/aREK0A7UPdZEWllOiwHBQw8fnT
zx5EWfg8EsFsrAOs46vFCEkM9z+k+DrDor38u7fRRLmUgND9irZMxQVxyxc5Sm58qgUbtcxxaOVs
DsXgiwkdH/lNWGLowfp29seAqqTV6uugKoDr6lpcVQJ2BS3sZVWlNOpUKmNmI/4EmAXcyeIJnJH8
lzKqm5kdqiBomEDjl0GwmSngM2xiOSP7AtL0DmJEHKq+7RJx+AXyXmc0reJREktMg3O9ix5iQlUT
7wYdqEaKgIsPMEDQ9WrAV9V2z+InpBtO6X06UKhRyu130LptlDtpxe88Wut8vU5uZapJOjXv64we
AdglE56nro9MGy3TUJIOnQ4g5IyfpcAx6RX94MDrozSWkqS5H+pjxo1zKwoG5YlkTp1ROVILpcYx
roRlPi/DU9L7GUCjsl4SKsiNccx6/tWW1IL9shVKIebrkh1DD5xznXZOb2E1QOeBuNA6hvNs64N7
172jwvEBIaAVgDv8KR5V+Jdl4zkXntse+uJmkWDRJwRpXgm4331OG/GAfkg3HEoXBYOdwDwp16GX
HSkdTF0S69TCt5XwM5KUoGQuePWS3JuArvhbhQih5/Yj8tAI2EJouO5tHzSGeZC+O/F7Vfxw+X7U
yNQ2WaPIJhpr0QkMHLLqKMvWmjfAhfMK1DxrqQHJ6ikWibRl4YVdGc1eUYLeXG4TlS/tC74Uf8tZ
sOVlbhrikZhJWVlNTavMwuf4fj8rdEqdSTyeF3q+ONhYW1gzX3W4LNkdfhP44cGE48iUPMrXDORF
EnsBu4QeAKvnJ7pEwV08QBALCQIPJw+fXjicgPgJ90aC6JIOuZYFuERePGdS+AcLTc2lEFI0EbSC
ch0xwNmxZN4VxmalqalzwTCy3OmvLwIQENTyqSZ51yN4KaxcXY2/+CwpX3WLqYdRT18A+PAYl26Z
LR67ttEDlIVzd0slepmn236POuyEAGI4eSHNXPfFGPBrdiC6XdO1tPP52VXVrbvP03NnS78wLlp4
7lLjjHlqcUyx3xVpRQLPZKpJSTu/5tH/O5bAJuEc0Mx7jrxKa0UREG+qBQ74qBVdHyVdptAXpsTJ
t9BMFYyYqbTFUq9h+c4k8yJ7et86E7r/0BZMEK8VMD/aMQKQXna9F/w3sA+UGHGQB91TGwrlnoeQ
7TCE0S3pF7+EWmJeEwFbaa3EDRPUuqtGHn/WcCISrtGnqxlj9tPEtf8EpeYi2NRo9FEUL19phmXa
DBbD9deF8sRJ1HkH92rlTMpbLZdXi8IGdHvDBVw5RkSFxgkmS5siyC2PcM34gzeAu0T4Uvmcwgbk
OJDhpIhwsirKIYXO3YFBT3cng//GiWGNV8iemlMPcKZlTBNYRI0Gew6L1eCXol9H1RQ/Wc3kwRTN
3OioyVAzPh8kqPivUjBhBO2v61YJaF58U4aGSV4XBDUfNgKPqmZ6Ouw38Vr8tRqRqhEYGto//jwe
uvcdTLPysx0binypYPTBFCI80qipdh9Ts7/LvebMA23K4E+K6kBEBKInzC3Qz3JOXfh0QOmaQC0m
T3FNColgjnE9BauWCLHfsKZ8qemOe1MwnfxLeEWaEfwBb4tW89DiUYk7DtFe0epYvPcMjR30OwXg
P9DC+9MPtTQ2y3jr08Iq3fNa6iVX+d3C7tkIMpg/STs/oxU02kHSyp/0FMUqodMnk+op/4v9stQO
hMD4/YtjAv6OzqcE70oxAI4M/xKh4Afg5+yif1MkRJ7giTs1YppPzWOnijdujg4HAE5p4iBSND93
kXtToL8WwClxlNLqYstLeayJsxE+QFu7go1nI8E3fekPrKo/4cIGDPxm0+kV+4oy4N3Hq3UQ3ADJ
tyZf7ORDpKQnJbBZ9hr1FCM5BgccUJI8cEM8Oag8RiWJV9NkXouXumdzGiQBFW4phw7L13G+APP4
c+lZ0wkzUqtJ9Tp1Vyuy6AqtJdfBEmhvYyldcZ6Wpju2ToNaMJLNA8OB1Xc+NnKkLUipd3aKO8a+
jJYcFUfNSszY59qAzT3RIgEhBQZjrZIZ+ObL8GS038RLEgLHavVS/XqsBsDVAvTmfIGcho0D9oar
Ive8wRdr1MLGNIEomRHCOKlOwK1FXDAA7t+WrTbqUPswFOE8vlz5jG1op95VVdFSFv32Jr9/a8Ql
6sM0wlN4aGj69IKr80OIzUrOqarH/1Pkf/RITwsFAtIFfdQ6uvKfwI963V1AW+iZEllU5dW3oPOi
6+1OqJnqSU+hGR+trI8rIcuCdyx6xXRaC+w/pCH0OKwgR/jtiiddWaFkSizVCpY3SJjJxLutdOUw
f6pCOJBbmNkvqtBbWc6qYpXi4t7h1lhn7wr7k3HZMY6LYChMQ7dREVFGZk+OwTevlUwiCDlPw0i4
HFNoNQOM4pSsrvGuwKCtdvdKvVCtfqeaoCm1MRXxUC3MNm2gypCV+9v/iB1p9obyNu2FyDkxqNja
W6YkAyQvyzJZfLVyWwwP89V2HC3hwyPY3Qr+SeuNfAewJOGomrOX/hMyQGXlLPZv/H26GMerCeug
HpGYkVVkpBEfO88iFOJe4HvEsC2WcSRU+68fED4E39DKfTo5LLDph+cCzQqnRWPuP0CagFYzIgcj
wMFBAun7FMaQgyyq+bMrbrMoi9LHmjpTMeZpliCgxA8oe+GKLwyZa0gCsvDSk35Pv5DuXb6z0MzZ
z1lH1fU0XMQmiXK8bRSLd+4/bgZ5INrwZtiViNidVC0gKYFlSJJalkJRyqM3giyRCHF/sZZW9O2I
GQLh847U2x3Vli6X0ybavJnMgRqWlLbmI+3XsapvSYR4Yn+BxauhsdjpgWYez7Zc/tkwXYMcN6Ar
t1FXYatOAKQW3fJEhsv50jMMU/oYhsRZ85vu5Smvgeygm+Dha6qfsd7ovFW4t4Qb55x7zjFN5wFb
9OFLYVgION/kNx/mWAiPkyo7jzZuSHwfj7cPy2Y6GommZTRpWKPwpq9dS/nS+ha7s5ZSV/k4H54Z
d1bOjEUUxbAeaNSKEIdNMiE6qi09Ruk+FQD4GfKNxPPWsqt1b/8KZ1isbp+MjyQvK880TwRFM08u
FJPQ103GSvBuAkoiKoKrvxvxrn6/9SFDQFVOV8eNlajGqMsMkbOOrwsinF1uDJNTUYIV/S4pc0iW
Pbc+Y1LwSEx0xb60RiUgz6toJWnCC3NGY4lmN22CoCnY3lZXcQeOGGLO7cN92YJJF4I/CdKgLGN/
ZDiR9o32c5rsyb4qEqjBXq+twOWLpOKK9gGMjcUEce4JsGcE17r8jirzf6uFT9E0L4141E24kYrN
GQH/LoTviCX01aWzuh6DWJoL1tNv8X6dZYaSLhYyEx1h/GFLuiBPagZrseI0qiz+y8wozvSxx2It
3mEwG9uSbgD938kGF+HEwwJayKdoHjV6eEmDbJOM0w7anYq7/WogRalA9zP9QF2Ua81ln045zBFM
/5LzrG+xG93rIhLgMfX7MVGP5KMDtRBR45Nds8F23wibmWo0nCK1+/QIBqyR3nr1KBgBrYErkTqf
zdl/gNux+ZWgvpLBPj1QZDIYl57X2N9ZeJq/dz0lpQg9B6RHll9zBDEPqnfDJOrG5X71AX9W3FGS
2/ENrDtsqdh2MkKHRGs/MCIBAxHqkw2zNL4uKOGIIL7IqtomypBgn4dGGxOP+qgRvkCpQBzetgEb
Jko7opdfwSAaLaSwwEE8Kn4TPMXgKNo6Fvvxh0zefeZkTBPlmPFV6xf+ln626/QLDT51fehART7x
RpA/WblZUnM/hAsw8mWzJF84KkLAPBK1OHQ9L1PPNyp1R/LgcjmJf9nGMllU3FEzjg4JCJhJVMgp
U+yWqZ8DMkGKMUld/aktMeb10HZwySvdOl8DzWuxBpFZoHMwY8yAqyLc8g9NNirTrmJu7xImHY71
ye8Z1mD/c2zv5LcCUokLbHErvM4DAqJ/P0wwZ/6rqbsn1kOKB51aBZShbbsbDLJtuiMjHC6i/rZP
LGLc/WNUDVISjLV640FtXN5x9lhB3NCMketrG/NEt4EFa6OuQaZhR/SL08FDKhhUykZXkbzywfhg
gQ01awoMbv3/MyK6vu2a8avJw0semdJK+SPOIIIAJWXoOsmuoc02eJbocmlfvGQRPvSW7+aawS6b
t01he1aRZC86O0aIo2IaCjB3o6KKVi7VStxNGAhn2z6UOwlxnuUf7OBHMEXU7iRkCysWjSutJLjp
5Hp8/sB2fiDfDkS2PJvbszRe+m15t1tNCYQ4AHeA62HA7YVmFhmRTNpKPVDxdcGRR8x5zA768Kqk
2x7mxg94Cdlv1BZ9Yk1EM9+VFsUWczEdjPz4jFyCvxuNsKRqi8abzwswVj5ZWm9abYN0c61s6jh/
X6tEETlb5qSi00FOVVGc33b5y86sOGQQuHbWFh6zQ987K7eEhsY7aTiUcOLQbRpjXolBsAd43bR3
b6MHimDnk3x874FpmPmv1fhqg5sL9Px3uoPSghrsyqj/+p220y9q2MhWXGDjnXGkYdHiLGmnnGqi
1tA/eGVkeyQ15YC4UkXFQlSOwhA2PKKBS1kl5/Bf2MQcqvFdp7i2l2YeelXtPSWOk5+cyptI7k2V
yF+8IHKugu0O7c08OYbrtIdsPapEvvyOFt10ILQRiIs9PPpAiBdF1Rgz8gcaf5aO62k1/m6zXs91
no5RBs0PhWJoe+YVpFThjIzgMR2+Ium43GbefT+J49b/djkRhH6bCcWTNwYXUHwGQzhN1+QxU2lC
U6Pf1jUj1UsI+yrS/ZMiKFdbEMEMpM820uTGyfG9uUaBM8CFUNTxY7rxwcBt3ih0i8RqXTOLiLGc
5/q9q6OLHmkSMuJEjmgHS1dYQJb8rBvq+kPPbTIHXzgwj0O3305kVZTjwMUcQ9ZQTFLA1uA7fpRC
hKex66GCstK2D6y/DLBJBlxoYoTGXTcaHOu1UEqAYVgAAqC+N9jsIrRrfdBRicbyKziQB9orieFG
W9T1iBRTzs/9dAkmObkrvIIoz3auvyGPXCG3jidDoDoZX6JGtr55ESjUeav1LbQg3ntUyUp0ERRS
XPVaOzUm0Q1o+lM4R0bzrDI2TZiUVCOvVQ8arcyFY8sllxWs7UKalB9LE3rSS6v9p9ulCauyZs10
KIk+PjucwqgdU818yaCCeA1uhbRdOxk6CaPVQP/aZ6Owu95QptOkWreUhKw8HcB0wU57KiBC8eQZ
ir2cr8j4FejORAYN31Q0BVee66+ISqKGluDfInky5vcq4IhIV0hsOYYwX9fMcYeA8OTSTAFVtmZV
kOVd3VNh9zpBtLVS7U7BBi3umeasdwWj80u+8XPZjRcuKwVJpOQEjY4PfhlMgPIBnARBRBH1Q2s1
z5FmhvECGpLkCcbILe4n1cdBAdSEb7nXYf+u05ouH6OXiac5VM1g+Br1S2vM20wMeMjHXlRCnrq6
i2xfIZlz7nJJq0CLfiQdJx54a6t6dLvgNuKEcS+udMk9Wg5/e5SAOZQ9oi6iJKPoPksqYh+Qp3JL
VLIYrCAG1DLCxAwudgCdVSF42mHcWOB6PnqAINWzfT4ixw/RI8mH8UO8JddagHYgc4ScCQneZeQ3
dj0gj++dzU82hk29JWbeONT3GpxdlSuXZSTCNZBPfxpNJLc9my7BNrnoIV784eHIcZDBygalqc4u
POuhw/D0NW+r1VISNwoYG7+w69hNBCRFL5u9Lg0Q/vSSEaGXBkgiFLgl4qo6GRrCX6Rom2nSujDC
mZmjFFm0jr8UBFlCgmSb0vXv43YTzAUgh4837Zh86Y7jn0IFMVbiF26xZowCNWoWqEXw5ucf2O73
BiqRf2aRBuTGQN1uhKNjyu1EGCIBjeUqoDx+Us3GZGin64fz1AlRv/NiS6+GDNi1XpXoN/cg9Ahc
mqmxp7mdGX68rMNLygkjj8HGAdoO6ZGM5Y/+TWBMCB0mQgasvLahZoM4DRAyehdQUQT4rVEAbrMm
9FCNaOp7uZD9cm9uD1Q/Q11R/A15axJpUPbigKqkg4Kxqbzyh30C4rFt8RuguHlRrp+qgh4Q9E6Q
OgMvjKkdqrlGsYchQd65SlNDAUUIrwuMTsCL403M/dXShcfltsLGj8nPqUnlQi13y/GZsH6k4ES/
chM5dcp9kmfLKaiqQazIguaGgegXzRecD4oxx5Sf3MboTxSpOMUzdsiS5KDB6qGxw9qMaQbY94gw
IXp2D6sUdmLksJNZJ5kj4rp0geW92E36Ukw+Dncwn1OnvT0XPSxa6zTGiIz7SANLPpWjGwXmNjvU
bH5354oJXvLq0y2UUVwauGY5rv9sKZRgAo64lp0+ZrWFDv94+cwODLsjfy8XjgRZJILUyNm2CtFK
4RwmiPSRk6uNkxZpG11dfXxUOQIq7lS9CJmT07RiXLoaHBHdguXwNKgmPuYaqX5g3NchIA6XrrYA
UdyY3EO8MzNTDN/yEDZq6wSq5pGHz9gE07n91SndLDvidAB++tr2HcaNgTNxvA4YgapBAjcx1B2o
6xkQ1wV0wYyzlQrJDrNWy7mJpx0invVXa/Qg8kACHzPCctku6ullUwU2NkEkYpzv2HZ5y0ZT12qo
h6YAmcdbwpCf7M+XGgyIyuAYaT3W1V8Hv2jB4KQYHLL/6TrJHuGhNWLUOMxXtwzVTei27bc9x1i7
v34mxbY1bJhq2XTKTHTSHQdeOl3Zk3N4Fm3K6ZoABAbbEFOXISe5HOUpsKIAEAOxO2sVsXnt7a/w
AZXYRkR1iorRrBZcE6tFmyRs0Eytms5ubvrNIztbwTLAWK+LR34bl/nR2z6S19o6MC4sUFn36/0f
3RYD9bfVDRnkfh1welA14+8l6aKoXtN/xtB4AahXkMRBSQ9w536RbvjjA0e3xCJgoEKq3HT8aw4q
zTLlNVyouvSbKm9goI+lFF5vC8mQRpwG6XvvcpYaRxAIYF+4lNLHcLeHBfuKEL6kypdz+tcf+EOQ
kDYCJ72aMY2ce3sPhO3mxzCtdkNgc+oUtRvmZs9JNgmImwNm8kG+NU3q5wg8bXC/3bIQnMEaaxuT
LBQ/YbCOBPoIvnBiHSc1ucyuN9keGBzfvWp6ezS61eIhzoh9vYskEDOpMLRdfJ9EMYmEw0PhT7UF
pRobqiStqeTF+4RfaSLeP0iHoEXOWwudhgwS9/VO8dK4NB4qu6HU0kyCjX4khBoR8g65yiaydcF+
OPBr4WJWUZHMwzNtFM1mWhJtpWthPIBlDFhQtdjC7h1ElLNw1kDOWWnG+hbSyTfZdhje+4WNrByW
GHzUeVZgUP8sGX0vOdG0bdgee5WFCXXNQpuuE7Qw3OnxKkIR29sMln2vYFe4qNX/8sMjM7+L/vWL
rHotv286hQ0ELMfDKAl4rDTxs9u02qHbLg1ThnrRRctqO0TufYG1SlIUwL2ZV+xSCkSO9x/iwJax
jGCjQIMw+yeoR3IewPekEGko/Nyyt5vlLsGFPMASS0UhLb1Cs8duPvLsxVyh5LaONFm3iegDKetM
THO/Uh8V0uz7MpdQCa8pnNwfKgLMpTjBV4gW2X4tr0KaM8iKGirxq4fw1graYEbM8sXd+e6h3+6+
LKYGpKhTd7t+abYy6HpNEjDzcPoX6IHs5Sv7VJcXfCtGlvvo4cnCi1j+PVEETzfqvMN4LY51xAm1
S+xQ2RQzjuSwy7kHXrMBAA2Td0H1MKrV4kR/N9bYBXu4wWffDEeoS2EDafKSx8QYg+xlf+W0B5/7
/46ucxKox+433brKGEiWQYLFusppXmCrWLV+IovhQqME6hgVEstndeCZ7B/LqoYePkxx9+7/Ft1Q
ibzWv2Znq+0DwbMr4++NfxD226jbUSomhQSnDsuksRW9e0rKEnze78dUr9U5DV3qkXuFmnQJlmIF
ZmwWEbgGGWpLWSmtObDrac3njeYrk57HYSrtSeNM71Q8GvmeeQc1o4ei0+v7s8475d4hUYDgON11
3ClZAts/LxnXiNrYjhI503a7uUhCmhI7WgE+SObv1VZEh+xTo+G432Y/3/8X4mU+2r9Hr529lPL/
BDJTS0dp2YH4HJTJ0vnI4GI8JWAB1Bq1TQoSTqjeTt6annyStMr5zxV9YvUyxbcuc6gbJIhVG0CZ
UkGtsfAyph8QlaTeo95XU6n6YaLl5f7GKxBZsdtK7if6A7oS7WO758CB2jWnV/UyWxd3XohA3Ddi
xVF4W0M3aZbBh54xyQAIIajMgezrnam9RU5/Q14uacZeMZMQ9nvBEEuIoNJiYAOjASxRNl4zDOHc
mtLM/H8v1XE7d9ec0OEkR4sZQ6GTTilTljP8TLbU41aQceZUXRQ9hT0apA3vvKegqoYSTakLnXSB
X0c/eywbzBL2lE3E61ZRqwlITLVnSJUt6NO11x+hzZiiLkXzUsZ8YimmNw+2KNgPXbilD26g6V1E
9gtWop2auFV3Z9djDz4d7ZLUg+f9r5piUKp/ppAZB3S1u18TsBZjxKVoqg1S8XmeoSo97qNuZych
tozL1p2cMl2db/DpnXiFenhbbixyFjWeEp+ZkN5xw67uFIRMY4BTbVkv0DgEK6SE+aJy9/7Sf3Pn
EyoAAPulL0viNDSSSfDr0IosxwoQJWPKjcG5jRHFCt+dCtXseAh1h8uXpoOS9Ynguwmw6PvQ9AgA
sNLT4kIcFPVJljrx5H1yq2SXmEr2mxiMHE8lCeQvJ90NZ8prt8nXZD7tbQR70VbvX+ere2qJUrVv
Ks6Ja++TX533Zb92qSB0hcm3BG95s8WPBW0yLpG7Z6mOxfNWEFJHhc+i5O0pDgx2+TqaA8xrfsEB
kHh1Ax1S3uLAjElQI9KG0FEHptrcEbrzQ70i2d1KHImfl6edqMbMlGh7fHJIy/dMESwVBBwOzxpn
Ia7cb0sva1u5QqYxfDbcp/mFPEH6r+pKLrmbMb+lTq+LESE5vE6h8bgUcje0uiIHE6xFpLeI/QtM
Xzo6ZRMoLdlOAjk75PSH4IfUpTTB8rgtTs2fQCWQeLicxD2qmgP8FMxI1/mdWtkYDPzo4MGmAakN
KhO+7hhxjoBozc97Vox3kl0+i9JHeNnDAEbdDgBFr0ryHB6SuEF9pmy5fVOiW0qcRM+CAzLW39uj
QG2vrKxxeCr+e9NwvEsyQpYWTrv3pklEAl+L8ElQYZvJPEL4vDO46XX+wap9ZSHNInwJ5wP8R3sZ
AsuMBNiKzp7EKWj16AQRWpjQH3XEdJb+5xG32TH5qBQCXFhq01FLowwfX+3Gxp8QQnMdIlLOSNne
Aa+H8wIyd1SwsiOajwQQsGn9rthqysKsTVDbVW9rg9ZwzQQnqlAm/n3CYeGnoX9KUKiZ1GGYukDP
tjo8xW81Ec8tWUNBP6nNOLcrzwyrSzU41XYRsXr4Rluv+e2VgxvaLIUBbSDLgqunM3wayHZ2ABXg
60j1ley1SQU26yhNQGX5lK059vgGACJQAc0natQiHoRvRMybChD9rHV3jw5kIllCjdW7vaVt/4+p
difnqlPg4jYt43y2+0/lA9fMPzHvJnUqfkbl88TbuN83HHHFT2tfr820oVEWs/4bGep7b45Chi5k
T6juq6cTntgaultfBtOI+dMoIhqaRuBvzgljoBzTWHWz1+GFQSkov6bmrv477s/+6QEUjPl1g9SH
WnbFdOt049cv8KGJI0zifYgjGHhsaYbYSVWZexCHnnNktrrKyeAuo6KruId7KMPi92vtzennZ5Ss
kOKfKv2fq4wdZDDS4DFZqYuigKSKBvM0iSnXZwrysUkRwEGkVLGQ1ENbY7cLq2Gp8PPMZN5LetM6
iHZMKQg6g+Q+a/MdXJtCHZf1lqMMLFZm1cy10Bd46nAxdtQm1agXQTWqXhrkaVxiqMzfAc8bCTJC
mL0H8ft8BQTCLMqBk0wj9b/HOeS6PlnOuFqZGy20a3asp86jv41EEzT8OlhY+AxCStBfkapyFJh/
BYfpm8i6+S8tQsyk04FepeY5s9VqyBPRN5QxJHsmkmKDoYpyfA0lJvGhJCQfVxdHqskctpDT6v8G
Gunyf0PQeiMR0XIxx8xOgcC8EGe4nlcpNu482LLVwkG1cLC35Ncd66vEQJ6rOkjWDZ2XnAHwCZV4
3RXrtlubVsKjA8ae1iXat6QNuvulVPf90X2saYQnNqauYGdod2mxy1krvOblmI58IgvWvKvh5+Rj
UdjDxlG7jgfzuJkzhT2mjI/oGZnuIfGeBBlHBV/iQyePADBU+oKe+TVxs6RDiJOs0UIps0x5Fn0x
+z6vomkGxB6DN6x3nkaQOl2IqAONwLV32TWj1islcYEGSIbqTGAS21hDOLLDHTsRsF+pWjqcf1dl
4ZEY8VieKjTpuoesza5vomIFwjF6XvV7mkF/DzJdHOPeVPM8Tl+60qbjf3wXwoRWE8JsFe+SMai2
JYW3O+J7AEspqzjpRDrXUiSCZ4CrfZU1HKwIoohTOjvIuHqgdqJwhOkTuSvDtlIOpl2fgim26PXi
2C741goMxstS4MGlxg7n0Ku8BksV6tkulohn0ogwYGrku9Fqzi78cW/Cgw3kIpaQ0hOxccFAhqWR
ykmS/1RiKWPPbWu70gx7kWWITh5OTwmqVgqvLb9utElx9W1cFLAaui9GQIEMs79IxMyjGXA3EFV6
ICh37KTcPs/7wtzTACZjTp1P8igHwWsQvK4s2MmyoTF89Fpob23tx3plILUebtMvUnUY2LDlkjwk
xB754xb/GjH0DOPsO6vMq55SxNUd9bZOqXhsleCcXQBSOclMxIH7yBE8GXveHPwmJ3i9b8hKukmO
T52YuxiGfktzcUVZ1UXVKlM3f+fxoD7aCDmx05438gUhmNEwaL3D4yd1cmbbeYx4VaFH2k5SUvPb
/SoEvxdYu1ElmO4Uhe6yIBo5eiR6sEGAGfMoJDEztOl7lDOJuVh70WnH7lZ6dbYOcT3eMgrxOvCM
SX73lGwwR+WR/Cv51/qXT1e4vU2glICo1CJzQJcAqGjvkZKIspNEV07k/hwgAM4J/IuGdH2gqRTj
0duoOiL5+t+mdKxr8vIEXudbs/GJO4DyP8Kt+s4yQcyyTER5DL6Mu37FbEjJwSeUVzR18NJrgMCU
tCPlrU3k/RZ+D/DzihPgPUdZaz8z28NqRay6OleiM0S9PfTU/6B1zj/a8WiSBP/mgus4Gtq0xOp8
WE5qKy3Y7WjPAurXcn9T6Qi0Dwtn9k8eCyfiTju75jyVhCAP+BWo0ZrJ3rbceUxaMD0RZdFSEk6d
0wNG2wsVHIyqsRNRRxbWQIj6W9Cw9vs1y1Zbq0uJo77HCSJHOFqqf/maw/LedP4Hcn7nA9gldSwO
pnPditaUmNsJ3SZYwp5ehrtassqMMfeEgM2fhfA3ncU/6eonkJWvSM+hsk3wlVbttV9cMTWXqzHe
UEw7bUNqCVzO1PB6SQ9VPErEu3epplJe3ldE7ZuqbUTqGzCEIFwwevN6ILzmCkMw2P/0R7Kn/UKU
eOhCAKnLYBR6b1QhcOhqUIeaOk7azA2qbxEXobqvnRGZ/5nVohEN5qAasKoz1ePwyrcx12I33k3y
0ian8fVNqTHMYkBxz0cKMXsMy1qwnlGTfzWC7Bnhz++b0+bSN2fR2Y+GwSuwarTxXbpk3sbr8xfJ
1HOg6bcseONjX0krKUyblQnWzGCEn9mxXjQ8kA+3Yn4+j0UN7Fk6RRbcjFBnpL7B1/JeG7/XWa1T
An7A0y6aVAJiMI37/JE3w7lyGCiKp0+n9o2Obv1fzxOIsBgrW234LLo5XNUE+Y6XzOCpgMFOiK0l
9Tx9xSp5+1qIWMRdVDWK3L08gAn8CtkQjJ2weIQwXIeXjQPe46vYdWeNEWdWl0bcVHyCsk1RsSDi
drIkaVpV92nFEz8a9mlJnIuWcLyb30OTioUbDr1Cm/I08iVmKWPND0J8+M9oqMk5X3VMyTdyr21y
NOeYnZiygiWefPqtyFdAjpxMBlMkrCp+T2IL5I5ELJa2cmlK8QfWK+Hmty8PlAXYFaxIxHZKzTnL
UltNMXVDu/GVbr6Z5dPKV7vdf6beiaiZt6LxDR9AmqinK+tOV3pZLuC0FcrmM6xXP5ckRY6pVE/+
1W1iotch/3yFau8o0EndFXTN0bM5sPtHPMSD+GnvV/i/qLB20Qty5Xk+4UB22NVBVqumNAla4FqO
ZaCbNQ7s3I28sZwapOyi7FF4/Q01+VSo3W7HYWrXyKxc1QP8McG3Rx8jYL81DKPQd5sfkv3qgRYq
A9O9HJ//iw0bBsf45YDc5JjF4lezw48JXck8YDQDk4BW0ZVbzes2TCGDu9b0n3opW6lGo7i8bWZ8
9K/DfeceHFbeZRbEkaTWqcQo7l8gsbEOko3ueHsXWG2jmRwV9tRtJ74lQEMGWM7DVRCRQpio7xav
9zvrvE+xojZwhVC8wXKYJzywTBGAq+yMplQmq700wCxNz/eL1DPG4WKzsZy5cR9mm+kLFhM7FAyU
Y9b/rnF46d6KwR+9HlcXZFyaDUEF76SpF4OrQf3SRDCYcW4W74LTnstWfiFMjmb7S9yw4sM/ZRmV
Ws3VAOW+yUpPSma8+cv0UxW6sjZz+xLT22L4g2iHS/omQVhcIUvp2aasHdbMIu11HYAS0+6TrB+h
pWKf4WE6Mbe///lWEh3lqTWIGvhGhlCYVp6qZ0VDbJA88Ui7Uxmgel02BIyYJg3ZY+/Ch7y4cvsl
uJ5tifXlWWtlMhcNEwUTGBGjanJ7/D7Wx/WHdklTVFFMtWaQoMYxNV+91+jx6bl9Nm27QTOnvjEF
tc6ccgOegk34Y4ElxN4Lp2hgibPD+EdDPSdL7FtlGY1pEkkXpBtjQ47wST/Lza8e9lLlFFw+MZiv
2rsVjZILcOdP71R5IFLaZ4Zsnsc00zunVO7cs0LPlitELpmADwjpWpe08ShpCOEM+xU9LzndqjIT
QXkgLHkNPD8oM5aCG6jMso4CUsRkdn6DHTV+b2HeHtS45fjj66ZdlXqmNEEF8YEb7CmE6j1zet9b
Yt6cVK/49cYYzPNMChVcbxcx2leoGCXQBxX+o/Pu3MrHz6bNOMXTln0ManLchmpAr1yMVKWTgWGL
fEnWXgVyAWt4HMcD7D6q7N7RwW71rVsVLZX21PNDul+4SalKIMfqcb4PWySrmCH8B+SsgjwWRvao
41KuiaVVuEo+eayk8KDd3zo2N7pwivedgxWKrfWjaxc2LfemAX0ge6Yamc9EjlRJ3nuMgVkFn/vj
gRwYRzk2P4+buJEIpUtcunc0xpPFDYmFMAWEaO7HZmj2thEAx8tdcyoRinvE/uDdtOvkN93WezQd
daVdppNicksTa4vIqJV5t01eBrg/IMDRNtcPm4tSld8la3rqXXvktBOw155JZnKxBWDpDEgwRGiZ
CIgbzjQBH7Dd6yviTE4dZN7w6Wxom2XMXjFi1KEQNNRUpl8/2HgD62PKrM0EywDf33GHpljvyZxx
5eJa57KtA3s04ZnYUXVny/buDRksrIbTNamIQS5cx/3nAAyTcMKWRvjnZkaVGVhILZEKlbPPFl4L
0iEcetAPmyk2KTtGudcHzrsYsGHHtEUtRy5z9WbcHnvChh4xLOduSoOh05U4z6TfK0U85YH6um9F
9YYcOstmw+EUJ8xTNvD5OleI1/PShukIiQZTmg+RqHpZMboAEGBuVeRnGTdjG4DCf/oH3QAPZPbU
F4ud54PHTXw4Z6bRZX+1ba48d47vTU6J6smrOqUFI+o0k1nNY+RCw2o7kd60eUKXgGPOiKOiwmWf
+y6zIuMFj1JVfvzFVXWkeEJnK1zqZQo6gIvDqpBEwu8pDy2idvrfTB2EDhCo3zMIkzmDk3ptE+KG
vjXOXjHVLPWjIxqg1XrnapEb3WCtvs/hEhd9QJcQ7wKPDGcU/CVSJjAsjMxIkUnmsuw5rR8C9AHT
obfMtSqsKvaxpU8DQYv+g2OZm0cboiZ+mwswVPGGA1iZQF6aZstVGL7OmZJ1gGTzidJIV5/EyDYZ
HAJfNEyi7ClU4P0qp5OEDUbrcl3lpsshDCZgrJql1NJXts52sERHpte/as+boFkHWJ5uZGSndFph
S6B5KufOuMY/AOvB7EXqOA+aYfQt/WUFquUBQ5X/CGNT76nHskP9IKHvnjZZU/d5uqa1E9g8x/DM
1/Xw7KJFtbr7mMysyRjWWd7NKFjid1MPD2/p+8AQU7kjYOKqDo/6UR2N5i8kC7ngznS6Iadm14Y4
F4j2Mf7/nWiH/IMSOSYu+5IoMw58fTvtbElEu8EczK/RaIxiXJ/V86hTS3gjiPOFJjQT4nvlb/qU
FoPCYyBJyIVldxkYSkRcqi1lFAjacHPnn72lY4UsKJXmrgwYYU7BthdLYk6UFULY9b6/UJl1F/oO
AvdLqk9uW16QkLHPZ43oxN63O+HXj8LwnvNhvtqkzgIRNCZCCINIkF9Qh6nc+YoPGr0GrQ95DhUL
sGa/HMLven2QhK98+AjymffjXiJmMD5juJuLDk20cvCSisLLfo6VUG/mbxDoSjvSojkRv0Oqx7ox
Ais1OwblbXzYZ+PsjklT9SEA8G6EaAHZNY8G6yyaTp+wMO1+DFI4z7GcjAOIdLTzM1jQfrSvzdu7
BNa7prFX5Fhm38CyZrmoQsBgD9KoejR27NFy+wf1qQmgOlsU/eOvK2lJPcZr2+c3R4wdeD2kgnmQ
jDNOz1bhDtt485YvXOCeX2cZVCawbRHGwvdCaYR6S/i0oTEppkasHj2vJbqexQ3WcvTqzRJuiAVR
ohWcIb5YoW7/yVX9Nw9akNVe2QkY+cMJck/dd5hSZxoYQTbJeJLdRR7X/VVxliIVvIo1m7M90dWg
T7SZWT6ynSGEGrEom1NOn7+csK+JMUujZmBEEg1Hw9eFpDaOLBlhDfULykEoa+4Ey7HPlWAWQSsI
DZDAFdhAxvKk//NmPc5TDqT9mGXqpYGowiHGvvqlpr5dTDGHOujs5b31/SlLWfIgUPA5y0NnlHG/
J8nPy4teuWRgzCyJZBBdOTlbJ6CaTQ36wCuLU5UXMLoWOtnKYGuK+JanNkz7KlyPEEN5sjMEl3pl
PLUP7fOIqBm/UfR9QB7AhH8M2Tpn7UTf0RbjxD61M3RwtqINa3kkLEf9n2NkWCcaCAZNTfnr6V33
ZEO/Yb6syswEulrMz0j669oyx1UIUWfyXE6yZ/UGMucTNxcSqrz4gDLjvMUTN32ilonerd5HHNgH
EtqH+Nk6YMf6BmT/+GWhfJ1vefYUxwBooB2zZKkYQ+Nn1JfAodtf9cR3tHMkHjf3SjvtG52IL3P6
k6iShG07zO29QR57YnzHDl6pr96S6l21mL35N9IJae0eTuQWKFj0lPwJa8Hcs1tjLEyW85UhdaHj
42TYjP6vZMlJDlNfEs7Irh6IpF3+ZIJYpzLJiZdF5jSgae3QWPUeVW8i1STRKjVgnwKn8ks0BVHj
Pd6ztMe0AVbHPDzNdRsCfudObSpYJmK4PzxqSmnXnWMccDL0uCFJSJeFSU49LlpogT7GC/PjCjgv
xwwSe1g+z3jm25Luv4JthJBY3U0n0BrDpngWOGX6/j/SYTf51ao77GLNFUERIs2WWSlfmfPBNtcN
uLTpkEsgMIhQJsbuJcV4KIEfM/43bhbkJFaraW9Ss4XaaPAWspFQEsqw/5kXYV7bQBwjTenj6SCO
77hOwPaM2Lb3VJHVpO3djTHc9lRigCg9JTAu5dJZOEWpZ9NxzjmP8OKyPtEbTcD1Zc5xhLvp1uIl
5v9XmyVyvuR2fveIAmm2zG+nk/XuvEZHWakgUbUWvv3FxRz6P18qCnbpZCPmYMHw4s3RF06y2Ipu
gD4UrkymAkG00+5KekWELoObOOKjWB4Sirn3wpxtNojSsDQD/Rv3gSmc4Hq3M+/FW+nnfw9teex3
a+rBlOrvrvNV2WenOh538RVGM+xwIZ6E7NbmKaFyj4/rD/Z2xYzALkQvr9oyh1V1bzDK3BcHmfDZ
ln/sgunO5jrGK7ek695oNVxOX5RJrabPHfxuw3cfNp2cYH1dsHpmzMcCf7HalVDAr2A36LOQqzIs
r7MThzACAYfb20o3ALauLDIEDbGITs4/miyU4HTfJiAaw7L9WcDZMC4Mp16DgA0o6l5dmIags4iQ
jvS/poDlwdmilfD+Q4vH1axxStSaPOHlWBCm1Ryxb0h2+0OJJd7krraGuwt1Bf64iN/CqnNyU4u7
vegp1T/tzL8NUEmAjKkAi8QNleP1gF/1N2vqBQuk+jbNN+RoNuF+3G6ybAdTi4qNyYS4mc6zh8S4
AxAe0YKf77ekei4Z3W2niOYFnXmNqYQK/Rncx2TPjn3fYL4PWAjYGQIMM6oGeVw7Fj/OL/Hqhwr+
/SbXuxCoYo7uQSYxHAoSX5pGVc+S9cpIrrzFONu49LhKlByWbNIVBxLWoQBE6R/S7xkQYLo68h9e
kWDDhiluz2Y8rpIO5oWUGo3heOzOVahmDOiYZZTTYvA+DXQBxDCCcFpDF6uVS3B4s6u688/vPl2S
zMPcaQxZazvDA2AX+AZXHbAAn4P/Cp+NwIJ/GP2WcnfePqMLfV10gLuB56OCLSIp43gyG6mkpshD
Wc77fkmspBP3SKsaU0a4POCBhdoS9EDixbD3kkkzbY+zLQEYq7fesWDfYLsKO+PNQZodCkepVIQu
2v8YQ+LknUSrZ4fW6fLE3XC+a1CfABAXpKTIkagDwD450zpTvf2u8IMk+NbEB1E4ILs4XG4T28V3
hTBS1QnNFekYl9JaaGT7blUrwt2ir/Umf5xQSFlLfhus7bAYwLaQMqfd0hiMEDXHV66H/wIiV3Qg
stdTNDJqiD0xAwVET1U98ictb83p//UNtbZ0e8CEXwRMufhGDMLSHZhd/Qfdsyyl+9/x9ayyD5cD
3lmDN9XpB3WFpLRj1r7kTxg5+4FsjEFviDu7NwQ9+StXVvZNXFN/Y+7wUo3kgMlXFZMQlgqxZbVg
L4AjyHGIsziuvzac5ft1cy+d2spDEakG2ZPROn4D9iL7oTHi5JBpE9mo9LLHqINNfRKcdrFkDmHY
7ZoucG5kEtT2TMIY6slwi6lCToxQzXqjYNO2OkOyQkl5ATm9kExY94oTupioy2Bgqv0a02Tnjkwa
mOxC22zJbi3XsC3pNtkk+CjknVUxu//6rNWG8hOl2TBWA+645JpR/uk1z8VACQ7kYw1uxgvvz9lm
nNYjaHmQh0+nbatP9dUHOG1BUGroMtq0pdgqOrf02DPTkzmi4uVJKnIaiaIR67b3BDu0MCBU1gd3
xtVerGruQSUryMifBsCSjMyjVx/mEDvSNluYjz+g3H5DkG57TsUO6UPS6kgybRPuoBUjGyyS/4ja
LyHDOxSzSoWuUn94PV9K9GQ5/v7EmO2vg1ebnE1nkOWsIbZNoIyXrZhd9VZVaE2mtoSOPrnNTF5L
0Mfckh6+zbpg0lA5kcKuqao8LTQuSvM2tfcGVdzfl20+m6UMMvRjLePpvat8GDoxQT3Gk7TyUvSE
Z7XtMiEuAw/zTFZaKcOpBbx9j83N315whaNdQ7hha6h5FjblKgxBAVNHt6VVbxXiLIcKJcn4kMks
s9XWtJktYRamMmbjSmlJQtIjXuyOmdmulcY/QIReW5pTZEgKODUQRtsD1dMBfoCgKcXOz79oWQ+Y
X9g6SxHlHKYs64RlvBq671Lye6Uc7w7+cqOwsBX/GPcgSj1c5/8tLzp6iwH6l8fGH85yPKZ89HYB
GTAHKwe2ec6E7vaG26lcMonrViiYaazgoNdGiPHp7hH+3tO8SfsE5ENJK8kBaNm4QnYMFjUM1/Vh
8vYV6RiJ/SWipzCo1Zwy2QBb9NV8LQv13Ek0cRXPU2BNqKaY0MnyoCvyYJ5W7f+WkurN+GQcidVf
h75KpJHYMe5gtWOuTRI5mai5j1bkg3W9stspiRPnWi8UfFhTZ9xikIZzx0Pdqrj5X9qMyMzWhFKK
mOKBqk8Pr+VoIQLtv693+i8ZHLrh7LmG8P8+JFoAlzrtHpZIb3WPngyyogjl46j0bk7cEzmDeKGz
xcB7e4NFr/56zqzkce/Egph6rM81ip03LF/Ao2NEkY49N7JeRcYi/C4AmIYsQACgB+V3nOHfsq7Y
ptFtWE9F77PLvji7JCpNDvbC0+BKwzfHM+eQoCvJ2XpQ4Y7WPIdNsf6lxhwSZOYALvT2BqSbbzbB
PjQI09l2BOz+CASK9QYMeg4ygYPHwQjyklmqSpqAQ9pVhcJc81sa+h6RTBvmyw7kFj+EuSO1OtNj
G8bqN4LcES37XNuQL6iDUcOrSUbbdzUWpTVeZ2aaBFXhoawjeVgB2lQ3IPygLRMVlSp+RignYJuN
Y1agjGm/Lt/VAe9FCAdZokC4rKbz+kTfRh3GDRlmPPrfidjvHhF2eu2Y8ZLkSd8ysSxdMxdgS2J8
lpEN6FkzA2UnKAXaJba57y/vp9BrpmCoh+/keACNKvbVMGsoAz3Iol+YVSsjSmqRmdW+/mLXZHJ+
ESeBU5kWVbEhsE0NSthYkF6bTeh3A8d31d5dl3Ibb+WxICNaH0+b2Uf9WL7DVOtR1CvdAi9kPEFn
gZM4XGZmZ2yTwrgDSRVQeZs3KDMGDeeRNi4T0ed09QAlyRbmF4pJy8toaS79aVzYpR8T7HnXsCsT
MO9aEQyLzU3kmKl8+EIz0ccuUeZ5ZyyCLCOwLmPhMCAah+dAkKldsQy1TS5gky1P2Z7zXaUdeWOZ
bEoYuQuZ2ibJ2OnankKAxn/v/O7fAmvn2nVUoVydvS4vEVoUhSOnCUg236qlp0az0Qid/nYAo0HP
5CNE1OjPDnUWAoGhR0p2d6tT10BfY9ic8qV2wUxBv6MdTKgYIV0pA3j47Jpe50rsiw3xpKuTw0at
T23RAH174N6Nb9tjboQ8iUHPL7q40sOQuNR6IaqQvnzkixlix9BPT6fasZunuE9MhTdvKl51iwCc
xDDqu+UqT2C7GSWh338HCKEu6dJnw/w03D7JfO9nVAbw9KtS20lrgSg90akvHIUJf/gZSL7P/NpZ
+YolD6Z2oZhMFPvArezrdmrJVG2QMPykVOTjyz6YI1yraMLka3GuTMc0R5Hgh/H3oRpsUPDZAZpC
cduPXtOfgvLxKPlcklJCA1OTUjRJ4/F20LMoSgz39MAM1IN5PL51ANWs9yGpMW6kU5OYPIRuWTyC
IcAnXYfZGznRA7Yi177wi3pYnKHrJkOqhfQHjrnMJ7vRfmM2bsD/7L8KkiNYV+eO4pc+nRUWb0b+
24iq/5L0JUbyV9jUv+a//y/BU2E16OQNSa7I9vGGPS5vhH52nXHSbbBDu5Xq5NbwE2HQLLySLPN9
BcaG0TRIKcgqayvLWz3dg91HtRh3dsW4Q2LWGO+POXqyQyNp96R70STAwOY1j6d+qi68LiT1VUAS
v+ZjP4MlrfPTlh0ipiPZN5T6LjeksKltKXUh+kXChJsTO2CjcbQYF8buZ9XalNtNXkw5HLFHYNJq
on2pfrfdAAXN/kzvdohqxoS4BIG6tiMqXWZCFe2Bh+KnDrhnz0jpznzBDzh2LuDajv0XPH7PbjzG
cD28DHfviZ9GoFpd6TpZWl1B3uovzVrqtwyeD6XH3QtVrHZXETesLrRj8u9N4A3zmZHbdc0RbJU5
UJFUjG/gNug9biVWRunOySPeGRDXOewB8dM6Lg8LS2kgjx8ryBLlCuOHHXdU+yKjNVYo3xYLJUAt
wpOhjWOKjPnQaE7y6EKblL0v49nz8aPn3F8ddi7lM+/HyHH96D2UUHILWgVgTA8Uc8x0hOcDGjoL
gmlKSV1mI9++vAjBQqxEo1H7JcuLgVoxnQtcSO3g+pG32sc3uMY+D1xnFa3DyAxCqGqZXZuLJiBX
xv3gEGeLebeyZOT7+nC56m+fT7M5rucXKDu/8hx5axzU/PSiI63JNB3ryQJgGX66Uf1iInVxaJtF
3TsMt347mc0Qou5yHrIVh/EYGNwhKgjZ6pr9ekXm7O+8He0gT60XeqjjWyFtXRvw5HO5X36DII2M
1Ub6XkM0bkcf9mlZYEUNdjAdbCz1bRglPnKCiBOcmlHank8B1BOqQeqdHETrn86MG1Ye5kDdmtgf
1V+mkpnzKm4YuVGHWBEiRBr3tkJWVfs5jURcqHWKe3hig1awdNlZetWTM83y1Q1ntgoV6Fy/UNsu
8LySrh/wQ9VVwnPcLxDkeNMuYeSup+Pu5cK6FeiMYTfCfqHUkzrqkAvFv2cb+XVkbwUimJkV2mpY
67btMC1rWX5/QAiWnq3/pPHaYekS0+XoOBce4IJKeKzpncCDDsjvdp4NE7LTv1y0STmBfEOD5JFq
VpXuMUKlbDZPmvYBuSgGJrkOLHKnB461q6Q9hIvzB2wZ3qBKU2/l1h/dKBT/K2miQ7h+c+d8sWTP
Fa9uLtzcaA3im53HfPfd8PcETv3fr8o3leCIQE4ESFFahKHrIc/T1RCutSaJAlf+T+hNLzw8S9HK
UzkOYBm2RueRzu1uVpbr0d/bz2Qk//CMa2MjwgRale04r5FDG6xZhFHS5ffgn/a2L12J6rWUL4rt
uQ69yRwPurcJHOw1Q8xw5cH9IZ9PgELGHK5nXaGohECBuSaJ2CWC4PXMFfTk3TudtGB7Zk7Klwxk
S5tiLKQnzMPPqDihs9EtaZBXAApNVfhR56aWyULN2MZNrvzn1hXCuPuL2Hh4f4lYi+idb+nrx2em
HxeFUs1e0b8iuhWarAEQ8M2X/2ktiuo1LGNhrd6vCRre0HI62ew95UD0xU5A7jwlalFesqMgwRC5
FqIaB29sNtLYpVP3j2i9ffJ6AQOJFGFRThWrG2zIuUnY+PAtL934G63/r/Rwlp7XXvQ6qNZUSBaA
6nUoAzxBL70FtTgukj203U3Ikez7ceSTef+7l9Mc651e9W23lCRDYQLeAXFc0MVJNkkJ/XJ/UMId
LNhtLtlqpd39TKGepTqGV2dRZVsIUr+I0zQ3tbcmv1HTDJowwA75p89AaglEnrQt82dP1CG7mPhX
8rX3XbhfLYxjgR1Bxh+6H3xkBc25QLgfAfyipfeRr9EvuRJGj70Kk8aeT9aNMTE0myjvVP/4FXeH
6Llt/iv6swvxf7T3+SvYwtnfPIxsqxOnykZ7uFyUmDSJ9DNqHkmG/aP447OR+pv5u2QWBw0ZMHva
o1V1/oWiV2u+QhhLHiZdzmUw0BDiuAClc0UABdQmu71OpVYDy5VyQfNdjItp5oGcOdnHO/sx5LHE
ukSoUkxMQfqh4r0Q7ih1yRBB1feWbJFtSuL6KAF0OtZMh0lO+m1v9kcKdLr/4SwJsbScZghGroeD
KRjdzsNuLF1vbQUUnGypnTZj43YjUSzRGx73OwXPjI66pLfwO01pHe6kmVznYBnfm82tg/St8ffe
rly3gf9mlaWwWSDqU82vcK6amocGhs3JrVQqZR88dtnlVlbaTQk29hfTsYDUnXiIaC567UFYTPxb
u+jptfJs6zdAXevRM6BLbpvVIC1sGBoKhjk2ZUrrm0SjzrXObdEYdBeV62yyEk+QZvMJLRAdvM4y
TcxG7n9SVzTnKh1zYsmYShqkzbBFb7fO8Ml5sOFrD2wxKq69pteQw5hWzaI8Uu/retzcuQRMGpTv
3ehAUZn9LmFFvJjgXnCUG2RYXcm4EF19OnLtwi4NgzHr2XK/HOWyVbZYaDZVri55mN0OY+YWyG6B
rKSMuJZkuhu4KHaUhudU/rOI5EmrRip24qq1tUj4NGu07v7sbfU0aUMBJepNslfe7RFXpGYuTsHB
d8yA+4Sc/35+OQj0qx0pTP/WBcI7I7gbBi+pXVbVo5YsxC9xEBnwfLdphgT7EEz3syXDdN6ImoTS
wPHWNYVeFdflE0KZBTtV3N3VTvBswQuchXLIfgDGs8f5A8xqKTmcp3LVyrqDfYnMGVqL1Z6i7NQK
XcPsvU1JG5+hJHdeiZrO7sls9+dzGp0e37V0sGqeCyNU66gr6aSP3QkJumIPDwrhZYI+KCNSJE04
a/R5/PfAJ0hzKcMVDO7XWvkfdPRJ1baTycXzlbSvLuUyiIGS/O402FmW00c7fgMNv/jJytyHoOYp
0YvCkQcowTtVct/e2HrfCv0zUXmT6u4p6dlu9jJzXgRn3zEjnCOgHeJ/kriOOb4UwrNhb3GgXbnr
OTUFlhdtadeUJ+MtGy/i52xK2bsnt2IPRJJFCoR9Luhpg3QMd88bqaN1FQ5S+XpbMaj/FA27SBtQ
IOGdmOdKE+aRfLxr9vmUeU7RklQCf8v6w6ehKcfBlUSvPpWB7VZJOt65YFm5WudSCOLyTpgWQr+5
o2NymQzZR/rrbvXZyn3BbH3zG/4NHLctOfhuZuO9uSnEJPt3azNWHzEyH7yRZWSHZk99aXzJhVBI
woJWyOdI3ZUA0TIc/dlvtvKd6oc2e83oZlYHGxIwpgCRpUoc1ZNWzGUgZr9a6DpWq561iEzaAK+K
1JFz36krnQEsEBP24Ble+AJ2YlswM2k7alzsgAL9TjcndouIcyhm8S5/L1mIVurtMZPE+wEX9hOD
o9xSAznK5Nzm4jdX4wEsUcRbSo5qJ9N5DBo9P6hPuoUH4qapw3JIN7CFZ9zZ9H0A7IF6413G61B1
0CKtP8b+PdqNBTiFmWggvAwhFP9zNinJkWuwbjQUN0JBd92gOA2GtggwYgPsOfp1CW1ISeJVJDxS
FqpDwQpa3Jy9YAriKhESq/OeLKDDxM40N3ibLiCLG5hmhIKOsJruZ8iyqM46mC3lxdCLViZ0LN8/
Bb0wNy0O7maM7aT26Nm5Ts3l+wQEq9I5/YnscnUAM1mOZv4UsvcRbwvxfyAbucMPsr7TkElNvdLg
UceS6JMwN434R/2U4KBs2PWFJdwhdqyLh3ca/VGS2VCsv1TnkN2F+syah+zKSzrX84/lNLw0hYgF
4Buy6O5izEIlbA1Jhfi+MHBCD01exHo49sIhffFkPDpMi+HLb5icFnqHvgFHT1iqTI0q8mGx31T+
EJKKhi5QCk5BeAksy4uGpRRXwRqAph05Wzpez/TNE7VuB++86gWjBlGkhSyUbZRF6LxlER9yLvmM
Y9/DP1zy19r3EyCgCghOJYuHwmAw3kNuTiwqQg9rj2MmistFsBlrUoj4Qn3pk6mCbtCZ58Y0AUsC
fmJ7usjDGMUAljC92qFWJdaP3g5TAY9GpesidpABs2v9Slqb4Zv1ATusuFyAmKuzTCKW2/+fMhpI
rW5ZNrGq2GnUYxRIJ0wKU/5gF+tEPSUC38a+wyTeJBU+EgTO9ZsnHHvENR9efwuloBOOFCDvMxcv
U2U8OIHN1Td/AzFhFnIC39VZXI4phFYhxOt6msMESY95B+7Fed8kQkpxuHKIezhmN47b0AZiyi5Z
YgrgPLYC4egQJ4BU2cxi2699U7NYP2frNnc9ljtEf2k8vGNTUOLkUJgOJuq6PSVV8kD9oRD4CkJc
Jg4FZCq6e5sCMy3mIw7UfwBOk85Ke1GLt0LnrtLc71G/+38FvupzfCqik4sLTm78rID3bCFG5Y0A
cwoBnIue1OEdp2zY0N9k5V25CRC4lEKXwDx6K8qINiheQhNNwu91Jv9aPkN/K3iDMqzqS5lDfZHY
YP55GzmyyFTnbWtrEq9ON1he/2NGFvGN9nAlIzQLM0ihtmgMzTUtgR+Zxb6qW1c3GC7PD5aVMSZ1
K9ZBWFsbjc0PCO5QnB+0oYtfTduqwiDofXnMyS3rnDWMs/40g0CW1GgBAVWWwrhN70i7sQpWaxgr
roqs34FawDTt5MkNLUv4w8BkZHO8Oi8jqvPke964GmOaTCM1swv/zl0u+OjYzMfq9JqjBLg8pSII
PV5nSbHlg4ylZHQC6NT7XrikG1TnAoo3g5NxecxLLrSmkTdqbeYEjes5tLIxmvxahLrX3T82E9nd
jS5/5VvKwKK4dmkS0h/oJcisgrcjISSA45XRq9wOqe4zpGpw68Ecn5QHOOVr36ug0ealGrrIa4Ql
LTq95iDZPFeSXmHrfK8vIeTLhfEUyo+KG+891X4ZxBjmXD7PTDhIgnkoBhtxhvJrPnszXPjrzKK4
n0/hP2tGNi3Xr1N1VOS50GtHvnNWnZT2MY9M7U7sUW0swPT0N6tGNalM8Rrdq0lzyS6dYUTs7hIX
ZtI43AkGyadDaARSMAVb/JP2+45eWsEesA0+jxHX/lQpSntLsaslOPmlcA8Vx7QceR0N5cUQ7k+s
O5EvRQGztm8VXWG1rK2Rs9woHrnosFZM7efWGN0+ghDlSdt0gXBcONuJ4EDbWuqF36I5PtiMRknh
XeKjP0xbUfMAh5+YI2c8A+x5BgUo/e4rAGIkzRjI6u53ycVdqn6g9NywKZ1WtIhyEQHF5xWqc5Jz
o5R4sk/YfDtmsP2j+AIjmQ2J0i/GEVz7ZWbztuf66ZXn3u1DPPtE9a8p6PtlcF3EMRtUkyUhL58J
HctFV8ioMVeJhJ0upA0E98g29/3Mlt/k9zkB3DpqyIUzGikF6PW5Un5gqFS60Bty7CpDB8GNf349
dhwP6n6WRugg1fgMKeSg+JL5fI4SbAH3nMotwCbNxCaVgMmNa7MfayZWAGuhVOKsGKZ+Rzwz9mGg
y5qKltdmObxLXXg7mOe3WPRPbBMq2HvF7v9Tr0XhO6C2Ycz4QXoQ/f/h5j8zsZZFo/RgwpuSheSC
f4cHO4XhT7LlrezYdFFbdZ3revL43M3HP5F+YpAiN//pEjnpbhRXA5x6iUKWDVfVquRyiLV4NGo8
jwGm9FDuIEqtnuloby3f2YJwca1xWoVx1ZLyi44DMox6w2fcsqFdW5TfeXL7pJGA9LRfyPDcO44r
ka7qtnnHtOFnHqw7YhZPEZtztEIQ5FRL9umO6oSuB+TH61x6s8XFONvFMfsWxuw5afzdMgO7eurR
ZUEXc135tRmrZadvlwhRGYgMOMgAzcZ/BZ7xnU+JZjXh+hI9Ub74L0N6d9RXsdGlYr7DUHR581Pu
wjGPgqjpUR/RYxk0apkvO44b17dazOr2sIJ1Gf6J4tmacwO5Vpuj4yHGA1TsKqyUM3idXptHVliv
JJukdTdBhxhEB5+x4BVQ7LwnQ35IO4VQRk+q/D9dnTLFJRfKjtTg02zdSgISq1wxP0M8rRSWFFQZ
XJ/VrH/M7fOhhrC+EjWJGZbshVrji0DyATy4KqURnt0ucBjWbfMAOCK1JTNit7HUafkGsIFBklLZ
9JReNtxr5YsfiGSKYhDa0+Ci2AgDtqwblsCQ+QcdDn1I7VfDMu4TV3xf2DuJuUEdFFZSNWxpfFkE
Vm0WR2PuxaLMc+dcvwWIpm03uPAaOudHrWXddzSs4+YX3lZbmB+1Yxg9wkOfmbaAW7hhCa48YNl3
+YliE3xVGYhI/NrWn7NKsR/BZNyXmdyKrmXiRvHboNuH7ZAQEV6l0lANdKHCPB1I6HjhhqJxNzpl
Ffxs3VPas4VFpNJksy0utSyLqhDplGNjYNR3XlxpijTIPvess9cyJliQjuLthAJ2+TfaIupwuPNT
PieptAw8cAWr0CFxIy3rHKSUIQqY9V0Bl5iv7Zgn1eaBYlukWvn2YmLxVkwePZUBxB1juzFaIeib
KuT0csyOhcZOcVPaTGuk8+w3rxWv0chmRZpAqufrhS5bd1XgDcaOMtXCnQP/qxE5LNqt1akRvPpm
B4ZSHcTni+6MntykJfexy1d0XdOVl3bQvzi78cU0VkrrbXxjmelG+pZTFSM0xEf18apUGhIWJs2Q
twAsjpgblrgQ2hwMu4x3bw/h9tqHfCdKJ6RFSsjP4USFqRw6aJtRImReCkrFhTgbTbUPapJcQkk2
xTO5qzpS7T0Eu8gNDUJx3z5dtuJ/S3OkZTb61HZ3t1BPMIp7Hv9IxrgEh4mHdahWp5CbCqSXISDV
0OnoPLzcyAC4++BFcRrLMuN8e7BbnxvxsdnPdyipQ9IKz/ucWKMCo4nJ5jezGzaZiytXpY2HpUsk
/KMbN8PIaPRmmBi9DlzCLYqJQshi9btQJ6c+Pt30dkzBuJo/JZQH4sw/soMMH3bM5xUATsJ6Xd1C
t17U90yVkuuE0Biqegn2QUQtbNnfNtBlxpGIOP2PcJT68BYkct3begkEiu+xHiroByTHJ5gBpjaR
bGhSPrxROgx+QKM8tP4pcrNsdN5MHH6/T5EhoZ95JcuNHxVdzVAhS9EZ/I6sZq/s9O3w27gsZxNZ
CECnRm7V3EABS0KKFE6R9cozcB0xRqPxQDdoxO0wysyT0q5MjtW147s0Dt+/pBDZtfzJ78h0b5U+
tuwun0FgaPoJoTjKETZSQ3EWgRas6XZaXrxaiBPYTBOYbUks7nzV9gSCvHW55qRj9r0LD1b14Vw6
98BuVGjqdvi23QPN75IB7sPtXAHZbgSOVJD5vccnTSYm8SmRZrfVHpFy2R2LGNIlNtCpTri+0vEb
mvOL/duOmejUUCJhcMFOUJgBmq9uRgS60NBmqyj/nJxrWhp3bNnlxzU5fG5bkiOYnPoHAiUYstTQ
b5r+VYx5pHx9kHHF1t6yhH/ssjx+ECJOb/ut0MySQLrSvgtGtKNjkyXLz+jwhEEYDoqCeh+jyPXx
3PcDNS5cjSmy/9T8Iq1Jenub5FuXa2Dc+YS343ke5ExqwGDkdB9ePWRePJ3J9gjPzfpxpPhfR3yU
ejlGjVqzlCovJW9FZOX2i5eC9W8OOMNY15mZ/8s+RwyDTUNIS+dewd9Xptwbwcp1NjGBjEQ2/2q8
wJyUo19iGFucIE4M5Z2ES347R/zmum2if37QG2Gvapcx/8JwXaGLVtrw/b06tAS2Q91OnYJz+42z
a07HMFJbGrhkXlW1ZalyL/ID3hPNADsLzTw4BYoe4eSjU/iZMfx04Xia//mPsTSrz9gaKMaSNni8
x+jSTFzsnF+lLGRJvQ9c305wQBt0mCKkCX5wkCKCeFGOOZYuMsFnUcYWGldp0bGXTBA65/riJmOV
Fm3AjNyqpRmgiMhc0h8IEkjeiu+AAeGiALW2X55f462uQ2OTnDoKxS986zAZgifsvwjqyNrtezGN
WH0wrg0eGvTLcGNcwzPtnrR0cBKBU79dHjv1b6hEZA78gGVpHoSxeRG9VzfdjPS/SZb3USWIEK94
fa6/X10hsGkhx2vLgVxgvoi0IG4bBf4W29oLPZ4B9gG13HK2fBJ5Ke8wu6BMiRvnKBCslqixHoTe
JjNoVbxrfq2oAO1A74YukIy3G4Eo7rqGHC6x1Nm9TIHSl54lLCSZewcjLXxcDGOHfttt7Slr7XGR
OiZeso3+vw5BOuArzcQptYs9SpVZvS4aDpKUpQLdk0i312zyIF4yy6ygNBE90cbNpeHXMAi+vF48
Ube1hELDpy/cf3N8k2iRp4wO+nxGbU7dHTCBVDuLJwxdVtoNnxi+4wxA+vabgMHow1FaDpwufQbP
mbdaCGd5oaM40smyhHFs9vF2mGqbI3QhSH2SfxgSM4LaUvG+pE3gIbepS/2yy3z6u2Qw9KeXPznA
pVF7BxGWonhQyzBLONBdfeNvwp/sQpEJpEm1xzqK/j6ygGtJGnTZx6QMw6jVRPXgaUF2zupqQcYJ
N0aNKU9uWoU08pjAy7xz3g+JNLbUltk13tUHT/yoHJBkumrVEsTZ+CtBI+SyUEDw3N9b5SNsN6ge
2mCjynGeXpxWyMHjzCX/0MUrjQZRu6bmXY0TXGdDIdgxl6BbK5P8aItSOm35EXkBITXiywfs3tct
9WZqeXyPLF94i/g4BbnyeoD/DnXC+YE5WiztqmChjAiCMH3Cvk6/7jPxzfcU12mSopT9/Jv7W/Qs
hiWy0gpWyzjJcJZPSDNvWHCMrrrNubuCD/b0eDGv7DdoSRYPNoqLUXAGiPZFXZp24jiJ9iVostBw
M0OM7i+1xYlyfYghJR8ccOaHhSkprcV5AcLESbJOoFshuNgVZaVaieEXk02ZHVDIhFNgrzlfMgtf
Wl4svqn4HbzurJemzvkAjORGmQDcoqwsxSrGRytzyBv9ITSCdWcXM9f5Km3tUmk5GDFZdP0IXCot
l//VjxUyRbl7mmNLLhEU1pTXafO9BQBdhlHHH+TYAIHjcgRitGsOZM1wc0MUDkeL5RFo0GBGofaC
ipz0MPJjVgEtKhoJf9YUlW4QpmPAnriEMaeG1VtmililrI2NEagnbq95ZKR+Vl2v+YMYPSt9BU7U
rvenVoB4nLKspNlzxY6f82qFWvwrp2ZWbaaeS1GEaJHY0cIBMebueQjWjkJimmkY7rnc6wxm+hkC
cs4QosNiJwWMIrFaVYeIO5cZHn3lLdv6V6+qA8pdv8WK8Wc4M4RkOpiaNgejVBJ7p4u0iKkI018W
zkNHpfCbRH4yHZoaZWSmCrv1nVcgFNg+wesElFvHl+Q2KDaYaVcx+z9scOslBLyUCkhUtqlw1t2L
xN5Wbs+VtnNYmHRZ8qcGVl1y5gl9Thx9cNohsQvD59fNObkR6pbt18In9vkFGgdUwKorS+sLmYnC
8o7RIyk407JpqBo2EoNfXeqoYplLpnclrwjqTKJ7tiSfFBrrQJIZ118Jv39zT8aAip41vUM70IAR
Oqnisvy5CfFVnPWWmp7nX4U9TZgCdSLomIKhBE2rBLxlp8CuZ5LVmZ+KlMOKvmZbCRq9ynQqg9Mb
fRz64R8DHyLXtRmSm2lnczYkgbRKg1syO+H0nT90W6zptYiOkf5m+FFWqdIf2IwsM2R/UeFFSGu1
MufPXiqAFYft1+yuYps2dVBTTfgMWDkcbgHYz1b3JcJkcbm6G50Kxng+m+BT2pM5+h9gLoQArIh4
me+qnGaWYWgcQzyPD7QHG8cbnAPJYL9YlrMpr+65ptQBdxBXHN2J0TbHPXQT35iV0YdtQWkEIddF
q1AotZV1ipQLH5+0r6NkvzDkars+HqjWiEGQ2MGt9QzrCRl12auLoSfHZhEyo6fcbXjfhBG3DHxh
HPvU9VyWcsNLtFxyb7jWXN/DTzqcIuRW1sSi9eWrHcP0wTfZv+nuEAfIukTXTm1DXqo8ESSAwrbG
PVgos+iy17H67qv/ntH8m7gicAawg2rHvKwR3KsyLY3a5s3nBwOgz5p5jJoONS+f4Q4BzbAKzTcg
MV6XcFPmacdWSNSkI7YrP3kOllturCzc9Meqqs0OYHnVfG0LJdljzw//dXO6VeWDlSulVmXbcg0n
e394+uechHjFFRsSpGH1PbELbJ8YhsspZER1Z6vZ34Adkn0sTM49kvXoq/LIdyfzJhm5s75bPlbW
BG1ymTDJmqYQIJMlOJuD0/COph3gtaMJGMa/+yFYdCQyY+5fN/gyOazwUQotigfLxUhoIv5di4l4
CSWli6JRN6V5yD5oZeUvnBIB6UerMYnggS4bOL3tq+Rajexw2H9xUag5ud2QBmxHNhZvYzQ4kIPs
wuzkq237wYCcxHK1vNoui1Qw8FgpRoA1wMJUHixP3F7ljDleMiSTXo4Rgmwy9lVXmH1sIpU2entz
0Dtg/9wLV0uDwCTj77c1dWFPgU3NTSJ8ZcMCBkO+mDRIm3ULcNSe+PBIPXFM20ftyF7mDgTOCUH8
9gAssOd+QRaQ2D2Le2ytamfHQNk3RPyrrnIG33xEKRBnHpIP1Bxrd6B9UIJf8hDkrzfJToox9Plw
pubiz4IRFotF3n5hBeHCTMvKQ2Nv+riXTSWBeYDO0GsAyd/v3U5XDQnnY+Fga5Lo+f7o7JSzj4IY
HcHKym327Tt+04h8Gpw07fL1hPrbicTCRpyeica5jz/ihJMwf6v2s9TYxmtR5vNZaPM24b/Lf36i
5+26me99AlYLoB4dQ8fevFqoxGxBDIpDRn9baHTK+2xvS09XQaSZaeZSIRm3E11D3QoHV3Y+gIJP
fmOkAewBqBIr27WM2IR/v/qDhiUwO4tde8T61rHCjKvN4muX2++q93soWwpAI7Kta7+8QXigZy/b
tDbo+WQ7JY4Z87+NGGsY89oH2RgC1NysRXF0muYS5lIaSz8E2EbL5O6fzmh+aS3IFH4db4TGZXY8
mKnsgaqcq1mZzo7wFWB5MmGt5SU8Xl4+JSrMJWpHCgEZ7cWorUW1QwIJwgoMjtM0LhwdAVBxSIsz
e+QCu+osTw8NLVTXwwvRUFpP3ypZwBuq+4lnACVZzL3uKEqIDBUClUTA9SXwsZe5nD/dcbr3qbnW
3x6OF7zSFYfP3WmofijHoioaPSbcjJOXnMduCJIFwyOFjsaoIM+SqRX0V5DP84SmfrcSW3kqt3yk
+PY3Fyjv2nLdyaPykpPCk2cG9u/6LYqGz0NfUgLOHmee3Z55qfMwEMkfWyIf4ToXc1N/DRO0ajjA
nz5eIx32Jkhl1YP7F5baH3syh7KLYBwdi20KqAVvKs6fyGO6n1mA5sLLyGJpVTuqUGUJmMccgg4F
VveZNW01fz3z3ifi5DmQlOA/D+kONSpJIG/tLMdia1h6zXRjwvkEwqgjBILWsEVtEVkkUivc5U9B
TcWRsM6qLcbOywOAA5SZFHHR32S1SaSRCPa6zelRK6V8RN+/TcJqlMXJNoA/lNm5bTiTOFoodP9J
1KkPjGl8H6xAAIBSpV88dWG0JB3ZMz+R0eIFf2capzkC5BGghyIcW2sqavZb8pGAOVeytY/yM04n
CGJcsQAFO1MgcBJ5jh6eF/LGiR2fuTYrNvbT984kZUHLC4EjlmEx6GNylrtkvk4s4+hgK/Cc2nOm
pds1tBiTEhJMUeTB9p8/SFesyFIeDqXOsKLUZ4yl1g8IC4nKM5qWcJIZoUaPX+kx26HHBRsjM8fr
pmY6Xc9uqCkh52M9C9cnAPfPXY0jxfUNMfEuQRgYJlADlzQU0M2LdENOdEF3V+trTWc5gGHYJVry
CE0quLigGxlJ+ZfLlvRAz2kenQ9M62eb7PpKroUBxgBITZGGJX3kug2ShpJXFsCNszWpC3U74HWF
fXTw+ZIewUNEjLYzfZcCehIZXin17gqQQrM7iNZzC1YFz0Bi+ytNuPh75fWNcOymeact9bXA7cc4
tizozpRUaviy7c0iUiB3kBMVVljRuv0TWonr0al7IKoFVb4CVn19PZC+zHKRl1IbnhFprwIlJgNe
/d2qCebqfo0dahdgegEncSu/QbnezD11HTkusNRJ9b4ejsq2ZYea3CHhSVvdzmyTEviFOdcLmjOR
95py5FdtJ/ofFI5gtCeEwXZ4HCsj8ZamHLmPMPUOfZ4GmNdB0SqIgYU2Nx35rilQBNywfizBJAzg
FnldwYJllKIqyp3rSDomIClYunq5g+ZV3AMFSWfV23cbuzgyk/RxxVfKg7YToH481O2oPqlHHkAP
ebdVwKGNl9PQgvQnBkwHrTTRFnOJ+CWcy+YAq7F0396uJ3xsUBqZehg+sbrSghbuMStwoctHVUBx
Ws3jB6Y/uh6K6JQY7IesIFvgqXge5kqSG4Cnix819HcDOpOeSQnedt8WGDp2siSCWpZC0qzFyEay
XgkgBX+3SO4uxD4zlXL9d0MIMg9fMG+ZfQ2qVavfGAUPdOVlVzuXbJD+zSDa8df/QOVSrI2g+RwS
+vQK98tDf1F1FkEncYUl/2wSySJ1zqpAYYHdks0auQ/vn/yt6tgkk9Xm7n6koZs0IK+ID/wFhJ53
VtKKiu3LhN8h6EosKXjiwvpN+T6FMRHzkLCWNboYX/d2s4MUg1C+2SWIZjqAOL0//wwwSqbXD4un
mem+gEmsLnLBlGMd2ZQH6jePTNvqoG90yIED+I8l0EjD4ezR584Hh9pTLmHr34lr71yAfHfPeOTh
uybmXOYWlf/InBavtTHxhGioBXD1jSmdPxJ0hhmUpeBFYwrefyQ4crSQG2PJWaAXK2o5p9vCIuy6
u5imrz2V6OYkNiaEahJJlDkGB0vQLUlqbt4AXktZupbBZeYCx+0U9WBfvkrywDY+ISqkfCc6I1rn
nuB4kjYbceZxPCITULw7ozej1tFWQbPVf7G+Ts2l4yJKUBfqx8w1SgHFlbeBNAXixfOascSuE7tV
eZ0VmjpOmxtY6maghFaidS50yyubsRMTJJ1n7+GB/jwI9p63G1UYaioxRx2Mcvn8IKTmgvkYPe0H
qiWVX3Xfa397CwPq6JNC8wDuTJwMR4N3mFBkjKKxJsw4uAScbJmoUJs2kwpgiB+1cr7pY27vc/EL
wg8ZRIGkpiqx7xjOgkeVTuqfkPc4oNOKGmUaRTlzFohTVs1W62p9to4mDHe89WEa/lu8AdVpUS8E
Esot0do/VUrxX+BKydv38LrY0F90XvlG35Yia/0w0lvLCiagWAWJ/d0Inciyb7KpPM60IKlZahQB
CBKE89+TadxHOdGnhTBvdLVQ7/1rT64eniB/5SGjZtqCeMVDM5YH7pCXic/7rm1P2kGRzVHv5mC2
lX6B4zByzSt5GHT2BLYZtGiuuyEZuGrXS9b7l9SQ6l35oDl64z1zlrY9v5Bdzp9ZAq+woFzp56AJ
MMPV/K07BUXj46Puqjt5Of1yASVH16UI+prA+55z7x2MdjhvSruW0tvb+tsqBWFMTBustqeh1xIZ
AAIBPs4rHilrdNz+nNsnfn1RxukA0JHzQMBWU/VX2+l8Yr/+pRYjvSpla3KRZYFcDtmU8+hST/I0
vP3s12ph3XKF9g9Z2nyUupqkhgdXz458b1rsaOH+kk7Y7SDrB/9L6tYgG69nmj0ttte2F4p6Vgmp
GmyfDN2BsqUhpoFjMKhWHpgLc1Oo+vRRdhmiQlc2sy2UTBlFIH7dUEUwVdKzQwPabV+Ivq1lTurP
U7Dbxcg0JKNd8q9+rrn7FycvC8dyp0a3uGK13+pav+p7uqw3zFIrGhpqehf4yMujzwknLy9A1kF9
1V1TTSyj9WhDer9A+T1XQ2y2X89TZgpxuIxC1Phrq97ZVxysCCOMPJRa/680FlOMYR835DrAjT83
v32PrTvqyGdSWxiH6U9gmQq0bU7keNbwvh1GhaNRTIJwlCasugkbyoZvqeERxtltWAIt4Vxw1etQ
jZL1dDuquqWU6CCFWvTgwOHo8QVElV/+e+teRrQKtrYIrWm7K0eS5SQ40Gy9l1x9lUnJzv7owYdq
R63+F8ojlTjyNFPgdROeVGxm4CzKXfbUmS0qEP65U57LUYRNDam3AHnDrW6AaYm0qSugt13qoRZf
dyveA2qA5wHIRiU9vRJOiBuDPK67Qqkrd7UBDi9itmCJoOlE7pJgbIiCJ8Fvv0aWo15O0qNX8xTr
7/V8QzU3F9gq1QUiexXkwo34pTj07pXf6fXXkiEF308K5uV0o/1OWWpfls12x+9qsg4BzFzDB1bM
2ZszuQoVQgU/lU+BJr+zAP/NdTsoUGx6ThJvA8RK7Qcy2+vzT4NphArLpXikzUJDq/aAj1mkbLEV
U1tiUZwrYPbz0V7rNVSHVgSxCqWamj6u0jPcT+UeiDfYSf6uZYfkMvG/Va97DJqHbCes8Eo6x5Ih
tvi0xrFG1XkkLgf79ZlPS+Bqzjkb4m6r0bHUlNDA4eATvbCtE+ZXWxPQEoT2YnvGAB//mR/860ma
Fk4S7gSW2fYyRr7jMeO+HuuULvvyuQKroId/JHCg+6JaypbPWnpAfBQGOSxpzhz3j4hgKl+a1E68
LXQqXFTr2JbXAYdFyBbNtcI8m76loZlWTV2ZhQ1hUJ3UnveErdGtNHUqx5MiAPp6ize3HUjrh8fc
AeSAMfRJAMai6zUneDg105iWC6urnepBCkIcYYy8wVoCqGY3Yxb+A2mdRJkGzSXEKfBoVTmSjSGz
TggOa6uuBxnHA6NZS5+y8oE+s1h8yjQPRAWQDcEUp9CFG3j75S8akMwg5m0YMRWHS3ZjR9b3NRfr
AgHbcRjWOoVMvLrtu50F9z8wm/VoJY9MjpB3cDTEjMUYpwV7YV1R1suLCm4R0HhN/gGTVOLQUeeq
ig2GpHMlD9Jg67pjFPDSiSXQ6Eq+cg0KUxMur33+tt9+fQSLsncRWliClMqeCOGy5vndeUfAy+vz
VF2V0JPk1gRgyc6QMw/Sz6xFkaOVHbuVadG1u0VApGPSfZqSTsWi5daoth7dVelAVtt5AH9wWLYI
8ucf8r6GD/YdeL8wmIk5U0AXZruJ0GqjVQps1QW4aeG+FLY8F/T+pdlTdNXJNdEA69wViwZ1kK+E
n/jrwHZ78HGug2oA5slmkYVG94cPMR/HMB8vmrBerusp3A65UsKce0ZpDrb8MECZw7qOZGB45tt6
Srhq2IyqOrk+cJZiykQhfgA0dIdFIbUifhu+g4sBoDlrABFbrL0sH+C75Amw+uHW7fSn1oifaQIV
8pfz1pL/fluxfSVY4gZhwZ294e3iuyjszv6N/riFyGv7WmHlKpgFAvtcZTD3SxGB1fJShhpyK2WM
AXpKVTn97Lh1zuJBcf3Py3bTDWo3UbjtA0bYbLBYSsUGKOYSspJ86u3diKlUkZoJxPNYxBKZhYYL
8o0ByVTfPWfh32xtb8ZhHVbXt25Xw9jIQ0aAkQqs8YVHo4ct1ybCYtQoc8Evhasb6fYT2PMehhee
O7urIhXd/bDs8bC71L+sPq5nhZHLSPGBF32lkaIS4Py04TnNSFoYawFwEgcd0WVbZ7ot7NYkBs+R
JVFn6FT2o88sU09NiMwprBEZZwdaoh072Q/4VreokZTZBmQrY1DEKzBCNFNKoNF1PR8Oc+aySug+
4PZ4xbnidNjp330LhCd8pCNEnVfKTPL8VLYAVFL/nQiVvWsw8oRRaqXRtivsbf8o2KTYbVH1na9t
BqeXoqDfPaxUM9xVAmkRrrO7VXWDwtAFXDYDZ/32p33uBznMCjAjDuBnffnV+7TSei33gxDmbWgf
K9NIrU+dzN1DtRsnxczxHqq08Jamt3kTN2q3xHOE/rl2ZqhERtWvoC4BibvF6ndLOXyFh3uqURB8
nfWlwEW5SHZefXX0VhE2/o3UF5GF3C+Y6EroG55+K6UV7pquBQVhsQIDrcwepeO7gg9jQxAuqXlC
L4iJNtIagLY/nzBfwyarnfNzQkjlR4q2TqFCun1JeVk1KlUlZD1bjvPMOwEx8vHWJMfKCMvc1kmG
SDMYmvGztYtET6PyTwaGKkooInpadJ7GHJGZBkacN41eMGFmcPbXD5bQV+1qWUzgwJT3gI4a1m/O
EPuKY3JbrwWVsUDo/O2S9Rd7Rz8X1v1JfVDz0VFKEVGKkxsr1/REj6Ffy5urW5D8UbfJjkrrafge
PmbpZENNBlUGWjMmP6OnbyfKmHT9Ua9wu+JvQ2WuiTrA4ZfWfECpf4r6nq9+Stkry0A6lNihPa1A
1NUMhnFrfbVkxVW9M2ZxWYq+KZBQLd8cqeB3PQVEs66y/GAes4WyPWpPv356zMBrKeLEdpvweQ7N
biLNmGQYGof0YJtGWsOHEfAeawlyQd24F/TANcMzuNQWfbmi8fi/O0j+y+udLfm764cW5RzxDdei
xxpvT1FePgTx2NcGlE1OT/dTukzXg0Cmszj3MYdvRupQHS0ImiC8lN/tlkRSp45dnbshdEegiVaQ
Lac2PAwYQcvNeGUE9+m4o5dyjo6PuJsZVthMWZgP0jQlGxwINBvlOi3f3who5SPY0LoS2/1tP1Ed
PV+NSpo23fxiqgZwMGjU6KbBOdsyEAUNi0cy2ZshZz9Rev8c+4yCfqYPvz1+Y+pyOS+iHVxf+usu
tiUlH5iAVWA+YS9P9nvr82FSz0Oshi/uh3/Hh5lF42838rrJFg3LT+iZXk7WFxHu/FBMkIi0emKj
jI3VXD1DehKacZI1/mCSvWYBrhgERBnsPWw8Rd8QQnOYxnrp+ZSR8TITGWOpZrfXwkbnxKepO2DH
iH+pn56oEWhJll2YrnpbHG0Z/15/S0O6ENI14pPNFovcsxElx8cgpuS+cXv21cld1p4oDo4/9uC1
5QcRBRZmPNscMkRf0Tzd2upcGH+8drdunMZWRodXzAX2yz9YbeiNAiiVO2XUSLx8mkXl4FnJQtj0
lvU9y/ePi6EYL3jkgkj5rCkcwDDYc+2jxVZ2PENQkIkzmz0q+5LnSqFWi/tjHQ28MvbgSS9dM+0L
WdtGJMzdytwKLZBe+CldIUL62JLc+v7UcEVg+EmV515XHDbYx6/jbmvlrfOkVzh4pDTa7T/o34IR
/BxIp3nKiofMWEqU1kmqlEhrw5lwMIfJ+q6dNRKatirdEZTkRqFO0FYP2VWTvciArtIsTWO0l+TQ
TMi2kQPTCntw+PyUGdwuViPms5pQSHvcq5jOEsNjef/Wozr5pliZGn9VM3473KiosyxGX0ylown2
E5a1qo8QYSnZ7Go2WaI0eqrW1IK4/Bx+/wiTGaBzpDFXy2W2FXHpFG+xQ42ahWmFSP/iA3kadtEz
a8DfAP78lp/exLyU++IVIHjdYVrSktgVCYK+N6PPg4kpYa8DWFIYY7oST5fV3uk+KYDrAVvGLC39
sL4l+quTmpHVRkGLA3FmixUE+JJCOvVezYf9MM7nA83NZsX4tu8h8+QQeLtSXeadfCPhuGnYhibz
qwgAkLAKgJhPLBecNalu5xq3QHC21u0QFvjZexZL8jMD24biIctjtf02Aohi+FFVFH6yUqwyyCbu
swNdTIkteqVRQx4KpAhfjqXCB0mwfabKBA==
`pragma protect end_protected
