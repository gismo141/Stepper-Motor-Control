// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
kr4YCcov8kLne7yERU8tTjYp9iq0d6/WL09zzqbC1a3zt7NXGpPfn7K6Lr0R/W++FBtUNRUZEPmV
HK5fAIqH+VuEkaoKUOE/0oSw663UWvQxxlKrwzDbumo+gpRkwZRGBViAnfhWfywA18kx2UrgpMPh
8J8VpZWwnvlZ0PKuVAqlUnumoTckk3rI8YzewT3GlfwXddH8woFRIUl3gq/YpcY5syzry9EyfIir
cMWs4dKaqU9G7Jf4CosRVjjci/OUT+7wnABA3HuA2eOf+LbIle7fcTTMnWEtYPETF/GKTIGVxJFb
tiVlk+cOb+0iraIMsTVCaQF45lRRKdHfKVRAeg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
J9H6LGJOx/k12I3iLrgMHG2yDNIZYt8pECrXL8E3DPM4sa7+/zBhSDNn+CuMG74qRPj259NIyrx3
bmHbsEqp6GFbKl/n6RO351NuW9r5aKNHE3zjOYHVjDQBdn/V4i+6urI8IPsI3zcgPg2X42vQGLw4
HgQKh5Us84QWA19N+KmwsbUVVsZdVdfJqz6zDvS71pegwWWGPhitOrf4pzLimFbsNFw3GeK7hrR9
PRLAGs0D9dxR/fMDTyK2/L/Z4tsZUDO73ZApLGE+QMjZSv09n7S8LBMDvMkgO0mmHgida4HLaE2+
IWexVd89Km/ERL0GdeHg+4/bR3fCFzjSwCoEzqVA9HINKs31ZCPM4QXiYJNfGdY6xY+KHS71O46p
H4jMbp2LjOb5GH+yhtx0+7eGGWXc+7Kb/p0GX6p/zYFJMB8m+GGcNtBI81xDZ8wvsqqQ1pK4+JGr
gvu7MUnqCEee6hiflIe5Q5SwouuJCnhB1dYIcFSkQYSWDr1NzrwdgwPSy9YfValv0MKGkFs4Zm1T
7M/iJODoEbtOvRrtALJtS3Qug60dtc4qrpkZiR/yF2FjCHxVA2e57GbCkBMvt8yHE660DKKEcID8
I1Y7usjbpEkfvWKCVe7PUAgAUYpJWt6zfPqSOfVTyZnYbU0TInPWcQplYf7xCSLh9EKR6Vp9tnOa
VIPvCxJLY/KRQgMJbZPz4ZlWBTWYSu+lHyhDAZBVcLvzvdnl/93qP5DvRIlrJhQywwNHYiM7rqiF
qhr/hu6ObsNcmRzbTb9UQleHe9yq/+saKiLreLpHozQhYuZdJBimvRWRBsghuYZMaa1kuL10iYbT
1lb+OnTfxWD0m3YOHcGX5tcy8zK4fv1B46Jj27rlbAT3QePa249GHDLtTgoMe4jnIUtm6dnJfsmk
D8BF8ql8MAd7dqWmCRRqVpu2xTWBBXkPmfs/b9ygEogV1nLe0VowDBbpJFlVfDdNm5QatDMssdJt
bfhC7xi8go9tZQ/ab5mCY8HV5QogX553aX/jNKiAtjHH2yGMufzVDbbvKky7kiW8FyXUH18Z7ocg
4OlGyfX0OaKo9sjjuN5aK5xgo4UfBbLW9Ynh11PHe/CadL7ne8Mhe2sZw95I+fcE65FuY8KK+Lsl
xLOZ8YNYFNrlHcb4YmFka96f8LPeXarVJJL7IAh5S6JpVElFRBiqFs88OlBxJ++wwnkiP0Tr04yf
iQCIYhh5+pOTZ3CejfkH9wrc1BNk7Uttg+i2s/i0oCsGBywmdQJKu7j0xskp+GbbL7Q4gds733lL
b31Gon5pgPYBvoU/YQl69f9g08C61V/KZ6bSrc1LmaQdxsOXLxsF6F+OMWPm5+kKoZG61cznIZ/a
ZbEu64yfIKWM24APrqnOioRkJgYZRNsf6ORYT9yuASR5vH1Xi5gMGFdKLnTrZaZPUI7Er5IyuPa/
QxMkFzPpBzvTlRFOURyvhOFiAjWrAYM41FY2wpptLXT9i4XGygyTt4l215TUFAnITyDBP0wxszot
nllaokbOjK3+N3A+EXlC8laGLt+8HUeTr2yTXaSwADRo8kPoMIEjEpg3iijhVl76+i/Xi5OcuD5n
PQd4t/POKfH0AYdSm76RwZtDIlPCIPstU51xM3fiO5+1jknsIgd6mx7Nqn4vZk63qzgorLP35x8g
BhOtHqjdzCXz9f168+pVBTaqKd2ASXSDzEf8EWNQxLaL4Rx4NzahGM33UC5KwUPnMYLNKjp9ueUz
P0I5kmq5tZCUJlPHDmV1wEzjcMK4KSl3Pzp5bGlfu7eJh51LjyZ6z7T7tsDs7/63RJIAsCa+tASi
p51DR/6rlYAa7CsKU272iiVfanp4BvwLEBn7g2rV5dWN2WypP5LJU06bFmoMiu6+wG9x0ez1O4Uc
eAROfXozAlWiJRHrrw5mdtoPpcGtpZ8VaHKLBO+d+h4Aw7nqT/JdNCHdoaerU4oWCAWtKlC2eWMA
nArcOpzOkh5KpZo3um9w5NgOEY/ymmmU78edTNoaLF6srEk0HB2V9QzyjruAs2OgZRrCsUHabzKk
FBolIzIsncoSALHxRc7Oaf7U2zTwFORysxk3/29WDMYIW/pjE6MGHBP/XVtftAxLJE+C4kiHRdLb
AfBLC1BAP63om6PFqY6LpZag9PVZhGYCMpHZ0hF47BX58Q09Qi8gql15sWfYV6eRFGMXRbGx1aX/
Cgsoz5Y8RXbgmjZDLvRxEuiQjFuYZQdAP9Ck4XlsgOaYpXvrOIzQgFam/ODwiCQwF0St7ACrw7Sq
nXGB/pDhyF8TxmVNQ4Ho91YpXhE3mc4TKp8jUEQD1r7oY0f3aECbYnpVmsojNNw19dWB9lFy66X9
2+DMC+sa4k2tGP2l2Ydj2ibjbM9E5fLSlK94DGc7CgHl4TO6ULIPoHwyMQZV83EWnize//a9ez+o
dmT3P04663Gjm4NMiRQ3eiNSsZkvND9f+xC+6sla85R0o8UeGfl5/w19aDE76C8tHrU/0PNiqzpT
CF2CFBMX6/EBgs3oqm8qVnqvjFZ76c+JvvDDFhi2iMwLyllVvqV70N9ZtUKtzc3awaR2EKjVy7Lf
NFOLLZzym5RdRQ9EIOuNQ/VWNvCe+ly/yJCZCvKbsJQSueAaUSqGQurHspuLd/Cv5nKEwSLJ6DNU
TyGJfhwKUOYeA3zIN1Ifp2Zm9o02vS4olJC95BQn2QdcLarKtRFxKDqrcrsVgNvk1B/TfwsRHF8o
dzRqjW7as1TC0/Is5hWkewIBeCCOI8MKsur5z0VWqULFegCDLyAh65vsO4vYWZQST0on61qO4nMd
plRfva2IyvzbGurCODVnr7FNFGoSgnPm4CqGm8+U7bqNnJrZHdtjGQtWr5+q9ZNAZrYmiy7t9bJX
BFv/qizxAOHCiG6eRB08VM1MwicsBHHrw7iGdSalwRpl4iwoPyjEDUhAh2fU9dmrHEIDEQ7w5ZfN
nI3QueXDGxykKuQms5XDqMV0nUN5+ZEBGzy0qrKf9LM33TIkFrzQLyfRd8YcvaA5Ke92LBwXxs0A
6TSen2HuI1S3QDPoPa6VEp11yVQevWqfaoTLhUSkW3H4YFrFeNq8GO/3Erm2UIdPd/oi/zT73Awo
5mIll2k3+yjYPaxPm+8yoihNJeLn9o5fOrCt5rhqCbDbR8Y4s3bwRpKw2NHsr8ewjq/gYxitwjx6
ED9lw7wqcNicX0TE5IQer7Xpn80ZxjHX3AzFzg1iqP14WfVdx6n2BCLs7nsJiElKtfvRX+7paPu8
dg3UR3jnWt17FYMh0z6pRUXX46bBTWQeCWAobBIZJ5adYIWVRct8O7LWAuxzV+eqXei4N52pVIeY
OAfoqjs/p1xn5LXv3LLBYLxcM717d7mvwaPzEdA+03lkG/rtLwnd7SHckEC6G8VYuVgeycMXN2pr
RgXp+UWaL2WqxJA0gOM6MydEVxCGvHGJ19/JDp1e6daxE4eAJ5HRUV28VjqVEmIWIdWFuK5owxme
J6xsKSnTv3UbdvArpFHGvTzi2xHY3TcR7335WBCaTe6CrDYWPmpfyBdE0G612NyiHxPYzWpcPakD
3P4kzfIOfMBoiG1uIMfc9lCsAEx0t9iw54AOG2AA33bimYpX00e8dwjaTCIH3g9PkkD7x2c83/3f
zH0p2eGMUJ6qBt3hdj5GDC+az3B0tr0dLMd7BKVMvqYnrQ1CwrHHlatr2ugKsCmbQIFbGLhOZdYg
+aZtknTvYCtj7wJvfOPwQKdUc2gNFtf24XvwLkxC3EMNiHsHIcfhy/bIzfhi/bUfpjhLleKnTWGN
bwSTe5yuDuvhKJPdd75tQj2w9Rl63gfmSFhGB69USPmV9vBrCgRQKNQ46IxWbc8YgHKajZPKV78d
oT772pCwTFb47JbY9GoVE9On2gRvuQ1ZntXCoOl3EiLbn3a5XZaPF9/KBg3zO3+ItSGaXIRxVsRg
wv6N2cymv8h2GBIFBRy0B6vXOmZC1/nfJULwHusOmNc2ivXU90jVNjFIhUTE2h1Pqd37vlcvBWKB
wqRa1cgPshN0ZSC7b9iDLdxk+nMhLyMk1cjC6JeVUGc15I3iBCbocNJ9aRBZiuLf8NRSd4RvdLZf
sFaB8xlUAuZwdIQvHimHrlZcSy32lRcbzcUap9kaaB+e8P3Le/hOZuk6KWfjA6rf762RH2N9+YlN
YiUctsyWKC7lUWS6AGiRiZR8+5PekvT8Xj3i1SYxChQBumXlnvHR4sWuRhgk8k+D9SoyalIAfujz
ZsE7rdYNoH+GijQazAPzlccjGSkgjg7X72xNoBBeVdrIEXeUp/bftqctsQRB5+jtSon3HtFWxfol
8FaLcOzsFTzO3m3qLe1rLScKOhLf7aMcy6OGn8nPR1A/pSbi+vjGRd4Ct5o+IJL7j0xyXPPlKa5T
dDL7ouwAeKcYB+v7kDsEzqnFCokHASStQrYWbMN3dlVrbNbx1pZFf36XH9/ThdAicJstr5mamjMr
+LDv4IN7PmzhpxcceMCiUZJV7d3beI9+ZVwspjdIpVu+BDtbt/nQBQvDi7sUl3OzYmla1bgbsf9S
1lv20cl/zTyjsg7YLFXQYtQzMuoZVSIJg+EOAEJnSxVM3T0X3sBPRosbEJou4qQbx2vKoIohCz7I
0UUIF+ZNB67Z7idHZmFKqu1Bvm4wnqNgLCUxKQQLUIuw2+dS89LX4mndYcvhw0MQInEUcsMeSoNd
zmY29yKeJstLzx4V+l9lDH2cVR6dTuwu0yil7rQ9KhlH46nFGxNjsNTmygQ9yb0QJV5IiCOkwn4h
ncgexH6q6fhVHMQrB9CRLM9Gcztj6oDRrHSHliVLRIMww+dyruD1U9wfeTvxzEToePquX+8ZC4Xx
/u/ZqeOJ6tX5aLSHnpOXTQ+8QFq/89tUBfPg4tfTfoYCwOdwkTQYsvBUZ9iADaC55kml0qo0Yu9I
jCos145Yd+P4Axyd0xDhrUHBBMNiwcdg9f1g0UFKR/Co9AnI4SCHGGsgU/Qz2K0oer3wbK1q3V2F
Exv8dvjyINk6S97uSe1lPQiaBCA5mdRTfyEnHoH003u5T4+DIqA0+lRv8C5LXs0JyXtf3aG48SUv
rdjERimb8xymc+oNfZGe46tHpUy9fV3QQzCRJ4Bp1i80xeVIoUxinmXALZfaPFO+qiADKWwEbQj+
ufVNrE7ZlFyYAmXtoY1feVUmJQQUkk763VpKIpCWX+3MygqLra7ahqXGDnIha4BhF21Ru50oftHa
XIBBZdGcLRA+Zg/lY0RkRZYHHEsJ2SVBO2rhGL8HMnPuY5bJaiZQGoPDlYUmGovWLfb7ZNKJ3y2b
+x5VGf8wONTHrDyd7nIHSwTkwIgUWxHDeuL3ch0+F+DUtucz3ebpPoplN/cDVUc94KPQKewiHBL7
cbAIcjfx3oUF9KRa9pocUZZpziIxmjqq86bycg2AGCYDL54yDatD0AsracdXA2PPNiF+3ZKFLLV2
WkXTHq0zHtUe8Fr2Hhhw/07K8D6jRworjQCg/g28X1w9GNCCIXpl55AB6vqccqSeQPgSodXthfa0
T72RYWFzb7UyLCPF7iGUnuAVBY5ADVVmSF/kcfn/71yfQ6urAE5FLr88BD5HTNMEee4eAySUh74r
twHNl8kauSZ1GvHh+JMbeZS0JJFRsZMsEnlzaB0I5lqzs0Z5cA/oTkiKdFtiLPGZuLh6z/WFGasx
OlkjHN+N+4G4XcvLZcOk7DwHXuGfikLqHa6AWtv5vV4SzPvsEqavQnvoBCvcNQzfw/jgTb/P51Ep
CSi3dtatNX/lNzEW6ebB15Q5I33XDnFnQ2+Ap5eWEoD5DljVp4HbisazimZZS5wsna0lYA1Ea79W
YwPli5CtpKqgPbKDBIdwbRVaKfNkXFS0tT5H6UrveZgB994nYjAGDMqa6JaTFCwdk1JQxnzx5RwP
7KBO4VNXDw9Z2nG0slx1Kh2AZWjB2h+MDGIAlfY0BfD/vFepNQCKRE8SXENq850XZjzE2qGWdMlG
UUPblnarIRzkuZsIH9Ki8t53lyiqyKtRgmaX+A4oXNBgd9DVaH0IkBVrH5OjOv2f3045ZrbuEEjB
cYEdRTxgrhT2kQaJcbTTuOa1AkEZzk3pnv7c1ikTL7YhA8UwVy+fF8kfEEyKSHT25Wb31YdYnjAr
TZQWXHJhYWk/SsnVLdDs8mfO80zCBB3YyT9YtLSkZ0tDtrTPQDwuPtgp6vXJxc/ubOr0FOxxAZPX
5bwBLqMeqoFKTTzSP79rQD42GngQVJiWo0czM/sD+2HwBJ/idybz61EUwHUj56MLRDO2DfYm8AOp
+I3VHAOnp5v4VeHqVfHRpCxnoy63GdH9mkrnO2GQOKgLQAox8Pun7hkIcsoJ8pcntf3vY9ZhFKhn
wVsM4+btbl2eRX9iA07H6IXZ2ICWgt0FiiqsygHGGu8FxQ2ZES59NYPR0+1VNIf7ERROXHHXu4nB
ZDAvi4BlGhaKvntFiX/q3ljsGQ0DlrrPdr14M8XUwL+caXyfwdJ1fsu/1sc/GKctboMHM7WiAKJg
eDHbfwF3yVpEW8z+Z0r23L243rhBDldd6TMgTaVwkzZNVVI6EH4wCs1WuB2RGKlH8OwFj50iTqKj
g9020YtQYh/+2kNOoR3U2lVi2lzZbo0X2Htlwo9dOakbzHcM6gnASnrkyqA5qGVmo7od1A+tjoH4
t7ob+kAo/Sk7/8fSWQaYhlruiNwGUvjgrmebT7q/+wVF/JY9EBlBHF/oGFK1NH8GBzsIE0q2rKPM
9klxoWwZPyUfP+ir9UcbyS5ORfa5itzTeP4YrjuqUgAsvugJTSc2q4PuZKyXBAOpi0M7n8nMNveA
WJJwELE8NdrwlSI3uxWwIIRch4dGaBlnQs/+etWMH3abVUzdgw6hGxaYg5Rq4deDbN+pGDpfuBEv
uMHFegu3iPrU37mV5wbGcPUrei6aI1TMqtonYEIjVHk4b75MxXzbo3qBIjTPFCoAKJ8C+y8y75/f
LgcwQ0QYkd3T2gn4Vz4DPBKyGLQSHmlo5eMta6bLVOqfSzk9mtLNtMzhXtf7MwnIpTdgPRRp/4az
APndcsfeTJ4C4oEfN00YtCJBmz+V6WLLR94up6Ywe7j/2q+jWzq5KAQr6aFblEbANiDomXdcZv6k
QqCfzNvuDPxvelSXAzUhtxEybeGZ8DOVrzWwDWJ1WC2kCEYdqBch1vqYUjTqgB4NxUEZVX5M6xaP
MBoZD0O5L3LNnyisd8muO6SZRMrFi1B8PNSStYEsWrOX3dj/zrHiny8wD7gCBNRzHx9bZe+bwqg2
0oLmVmzxWk9Q5DUMCzir4ZgtfHKiD2Q5S2FwU1yM25ayL4C8reRQIOXmzjiaea+IfLf7ynt5gk3F
ZdRFfEJP0eZRWVN9hmHyS/4Onev/nlnLcFhUEZfGBK970aNHrVms97zdvVXnhQBaEP/O8HRwiVl/
o0HKLo4upLRXrw2TuPeoZw05h68h3k0n4rO6jcVDIQcf9/GNqKjuWzKAecswGXS/+J7dQXO3fpNa
tSyGgBYdWSzQ8WUX2cALPPI5WDE9PeZ+G19GjJ7uAaF7yxSQU1mzkt/fUvFzSpoc4agQv6cxv3jZ
cfA6BaEzwp0KJbRCQBFFMFgnE4GRaJSUjv4VJrqHlvKOjOFAU5DiZvtVKDRreim3VEBm9NwTj2fu
0LPSS/e4PdzzSrkLz/anU3Gpibsxt+N1MLMfzHK5ofJg4whfM8IKXeFZK1eGZ8jCVzGEOs9++1Gx
rB+/0lzpiMZJZx64K6Kp6xZf0scHrbDP2lpSqc6R/1DBJdYqK77ezRdqxmE3TPj1FXpMNDcxmeZ0
OPV+VnCmh3m/CAunaozo8i/uIJ3InYVCnTYk1WxU05RvFL/BwknW88VzTj9PVc8ahGXVXhVLtqOr
CwfQKTj75HrMd0v41OtJ4IlqE+9knOzZ4owB0W1qANQhpxevt95FlcIc27xDv7h6wC33O/H2dhD/
L7qk82U+5upEOsBbgLzM1/l2pgpPw8RAHD74VPQA54Pw4FpF3A8Pu17IzTm8v5m3QqPp24OP9IgJ
N0x4MSFBsJICpqNEIz7w+4CU2U0GpkjKi0SY0csld5i7ZlFyWrmUsyFzVpeukb+ETLwDodEzyQ8Z
CUFpJ+yw7ioueAQx0pgWlUukvnZwHna8iIjEuextQ8lJuDRikUYBnOukP9vif8FqIVO9yhdAKB2C
7aNDW9uQvn4O7RpQTEc1cHjA7U8Cq8yBLPFDyo+2KR1gZAMwVNY1o3qkhcclCyTa9GR6fixRGuPm
xte/DfG4Dh5dM4UFlBg6PbH+RAIWNKXcDuOaRx9YH9aOVp2Sa5ukezBNNDUusyZJZ2v5N87YLfEt
1tI6oJ0k04WavrkUCKkSpjylApCE5zx+L95tloCsiTUZG5GbjvkChcxtino4C0UftN2VNbm76j4a
wvm6brkCdWojUp3IbrdXKbVcQMYbeBM2cQlcwQHlfB+xOr9ZGv8KjOOToIDNL8KNYZqj8M8mThYl
fUCsd7l9KdzbiArXez1uS+2/BJQ3SAdJpQ9h5OzyKlAuZmDrfA1KD4cUpTDgNJPeof3w1fcg9RmO
NZRkmoD1z1Vl3Nb2nkCD3LsbpFIh9+Gnxupl1T/f45KMVgsNrzq4YgJQv1yrNOG96XeguUtqFmUQ
drpmA4qPqYwbddyd3SkgT0K9CHeqFUTp9WNt0DnEGaqiAN8uH4A4ZzbNTvVeZqq+VDIOhApaFpEE
ewNdhWEc3WUS00RdUCOg6dFVoDnVFZGsdY7i/hYBQYwr9oa70x/WN0ptGRYOALRsFomYSLRv3HBL
jwS8b3FtVHU6DTBwZiZILyxUB6vmMyfQeoyhglJvPlqVkUzVIZYYMQnq0LUqFvKRlKV/J/U5gooI
oEtjqotyLm0kHBRDp6SMI54jFS+UvK4ZmGe6P4Oopp1xRotAEFE2fe4HkCUMg9TfUHaE5KAoFubn
cVoB9QJnDI8FxvuMMoYn8IHg2/zqYOqfkz/vIbhhbcZCU/9h7QqRRmUIIvd9n0bU51cjsnG2xddx
UUbalAVcOIl/ZQ8+r4wmHv+DF2v6zad4/7lvDQnc1NMkjigRZ5CvYORGwBpDVUoy7fXeUS+7/pDz
fqduDhvvglIcx0p3so5t5/QSfXF5OFUAVJm5Gd3rT8c4GzzOCQfZbC4uRm1+19RnNpc/YzrLIoKn
IFuF4+qG/q9f03en3hD+hsV8CCWeB+3eusKLFHs14Oy9oIXe6W6qTxbKpRxwfFoQluJBgfjvcEwY
T3PfRNGBb7mHqOcvpFYn4VWEpXQmuN5bXaHQl7EaMK/6JVd7rOXJkfiNxYOQxn2aQP/pC6EK2ToH
a63E56ON58CqzewCUfGPIp8pxXIaR00MFkYaIuVSgM9daYc+oGJlmStd4P78pywXMunMPft1iIM9
lOR+Mc0zU5svO/aU4cQ30WhGz+4dUXdlQB/Fhv5tcFw6r9Hec6Ff0TNYVxqRWMFRv7hVmAu7VLpC
x//zNoEZEtRGXmjdeTQjMRYYoCkDb9fG2gtWjjEsGQhC3FNSN//kVWb0yU4Lqxp9sZ7NSIrjQZtK
98MGOilNTTAu+sDbXz2SjB8Ep2tBuxFB1RfGWd0jrOuvWQM79VMyJlCu02TJrF+HwUboTJggvokg
WTANy/mHo8rBp6YQo2zB4pS4mW/OG8j11N14uOyw9ZA0aHDtHP95jAADn24LgUK2TW/UgozvzW1D
erB3S+oTjaVOdeVDvvxM2Bz3HJnYja8tOgAwLB1rMi/1c9f5SjtSEGzT/pKj25rNAB8JVAcP8UmQ
qjn6uVrc23mrESXJj45jKE0TN4CiZ+Sn/xvwFORK7Na3oGYdw6KxMznStF96fkEblUxmia0ZF3Tx
3GsGMM9Vp1e+2tIf2kpoRjxSE50MPRJzt6b6vNb17iGPkJk60KJYHyedB69OageQGhwdiMlbNap8
y1XcYH3GR2fsEgV7iTH8Y5IsKotMZvHYZXVBagvGzVHBNiDCvI2gJP1cdHuY9tJme8RyKt+vn0/o
e3INrpx6be2PcKhvZzlwRiYkzo5gr9QM/3+7HdS9FbPk6+g9MSl9XMt4QqluSc295GV9YRUwBdMK
D0jzXOx9DEEmX5bBKVLjOA2X/PIM9XJ95TrofunBlPOfbZvLE3E8a1OPHGUR9cmY1kbV7mvNUX9t
V9Ib5Al7Tus49CRKSxz+A6nyWkEisOgX7L6apmbzwrJSJ26v0dN5nZbha1KnbSuz9NCXAvphUH4d
v+V3dvrr3b+pUTo7jD3hE1vqabnMx5kW6KyN/2VHpOkDKj6E1IMJksTwk0VtDGzUvjPRxlXJ0UxR
LCMWjuaJZfAomwZ9hMvY0uRXg+o6lkaSq+GSFjE9dD1eLikgnX6OeKZ8fY93661MHa4mzzkOIkDB
ysb17EfKb1GeuNIkXKPJn3b3Oh/gY05bKfiQw1Zbo5RQSYvvh9oOl4iPWQMU7Ms7zZtupUY8XASp
nKPfJboYk7om8ZaVBYHBopJybt0i5NiQ+JTuDcFBoAihryzD6uHtBAFqfOJGgBEAP99fTraKwnTR
sKcTUzqxtj17eO1CKz2QGBsYYPOX5sGg7bGxBEBWUfG8ZXk8942WM4H8MOqPCCRVzoUZ5LqnzVFX
2F78Imlp130ziN0fRG/7ycOPDK8DEQPQve366antgQGXtuAZfjF0BN7FW41UJ94hjFHIOJpXE26C
4i9Tncky+8VlHQkMlO5mzJvIJJ6g2Qar7palmaVeiwNLPnsUzU2FXaXB8kuoYmmnCxuN+3Vv0w3p
OZVcEEF93yIJy0WquuEXSeDOlE+FZ8dpoSUq6BkSwSldygithwKVr4REJwEm5hbU8cFrc0evrdoH
h+JXQ87+d2Un0l4QQO+vUMzLqEDxOlkW5LCH0RGmTgieSWviFRWC0VNIIjYgBGPbNjiKRWjQoABt
qwBWVE59flU6Pnslu+QeRtWy6AMU2U/Qa0oWroRw+EWNQpkuIGFrieGKDmBovZE3d4hTXE4appUk
RYzP7yxlBzaoVTOm8Eupzs0C7ef9ptkTuZBRr4K2no72kNDzX5l1PkCvoLfjbRtIpUyPNQc898SG
aqCs0Iu0sBBsEphai7NPnt+KJBDZPJvRxc5XU/xJl+Ki+LPX6U/Xf9MBZVxdeRAlitL2YkbxhF7+
JnbSnUFzMstjPG/O2h7ZXHPMJTZOzfditzCHNrU+YdIEisFUnX9u9Yz7M6Nz04nsh14k8js21UsB
pmnk2zlFJiTl0mwfwqC3uaYDmeqmw7aHPjBXc3uQ/RxMYxJa6HEdHiIbzgNDhrebSVa73GPHTKV9
pZIMUyHRtxUH/PwQz+aRXkofYPqaxgPW8w9dcw+EopfpmiJV2j106psNxJG2SQpyKJnoT1ShguE7
Th7W5BF4t1wapbmhpQX1dIr8Jp35ZVEOI+nrnfUwCBZ3Vu87LoHlQ0ZJVHp6ZQUocLoT+k0DNXj+
Ge1nCC7MCBUmNdGQ7E483i67MkEtikOLsV7d2CYiUwZuCHnyMvHsUx9Z5qPoI0qZate3/ZpZCWeS
NW1L9O9dm2NzphfcbVPHUyAegsLVRHHEE/cOgJKfa0VLrvH8Lxcp6FRMGk+dc7nmz3B2lzNJtZdc
VYEb4ZlgFEJGLRFmBuaBcYddVbj9iDX4JW+izY59GkmM7kX4uVUVsg/0oCToE+b0fHq3i8G2uoMx
trco41P3lC5fvhEvM7xBGgpLWyTfpHnNi1e/kTYhztF6Q+KNFGNO0P7GCPH95NGAdU4CqBD8z7Tr
XTcn+6PzIpch2HVAFnHZRoHje4Qw9FYe9fOiSLLBmIzNX/y023hyRTrgXA1sjFKlvhxSnxKWIlz7
QmSAB5e6eEYGg3mkVPUkcx+/pkrnE2Lwdn5QYoPHIjHThePkiblwH77fpeene/2Gz27jABcTcpJR
8DwZqYCELuIZNq+k4//KGpZf3IECErrboaE7e5NA2Y/+zMYLOoAAbYuVXbNSF4C1ihqIUulVQwRu
XGY5ifZ9+qKY1H2RZGmys+pY4nRgwOuQ6mjQDo4NuX0aUrKmo6JKxqWBWAl+nxqF8OxhhIIAc81l
CzYTI6uarQlxIdMXeNp9f/wUOAl/e1ZP927C6BtX6SBxE+3+KXHOMWVl8nMCMv5UB00klgwudGxM
mb1kyIUUn/QBOIFIpcVN+roeF3MNrl+cYHX6IoicHSiRcGYvRuKrLpEqvoCKats85OO82jcQTx3k
UlbWZcKSEIfNpkwB7LbH1/pR+3zKgvLV3YVc6lny8/ITRHJelcZuAc1WYFpOkneOYuRKzaRGZysi
zWvkd0Ih7TL9XTLJH+SuWS8nBeqFWGu6Yd/bRMooAS4DKks5UNLOfJdUjW8GEMGmc12LkHQ0wMQ+
185ec7pSgH+y3/gbPq5aUHNYXYa6xezlZ8JeLee0G0NT2yj6OgsGtyRUn7QLiNYN1LWKXHv+ssX3
b6xIPGwHJH92tYpfXk8MYFQBr0Jfg+FQ9m/RfcUrLT7+mCTx4KZigc3QgbZcrDG3AuoZa2I+4/TH
KNyGYXNWV4UZ8jpGGqVrB5VZiJ03NhgkKB/pLL6Pci+C4nuHMeBolzC8mxyhYPinJKGe5JmaBFGN
PG+fXmEQ5pe5myqMoDbB21+QJzDjxRehqa129Y08JdhWsaCMc41EzXCZPJksen4ibKaqOoIaxPME
TBN8C6EqsJOTmoFk3F9lefgxXuc25ABLvE3d+HAkxtTYu8Qyf63r49Xpw/vntr2ibZxsKItINaza
rHO7F57+PPUo7/IkKl3mjm9ExtpO0FHykLApiBx2AvJDw3eH1PWLuEacHRB4HNcZtV7HR+vPn5QY
uwXDK3TPNwVsqZHDPRcMVhKHXQOiEm9jPXmWrzVRET3n6ES80qx9r+LO/QxQyk1W0DjG/8Qeky0Y
vs3bdr3wPTphvgBYk90zYQ72fB0hQRjsrUCiEcCh8zLxsuY/Sjp2LZwZkJ1qVa0QcGXBTVKTnSeB
868MGMKUzOhIu0S4Wd1ptE3l7DedD2LDouduZL6bIjd4w6mEqvrgXtdTy8EGV+JygfxZLOmJ3dw5
3EyRQMIcECwGRIa17JZSR4k12NVE75Gtt3BZDblfxNePnJbZOE4JSZfHBoqiZX29wEc8v6mgsen2
snPWy+Y+H+20XTc4cKHnmoEOHZGqLogZRJR27w61eKVo10ac2NUZMzsfoYw7dsSuhiVQtvf3aOyD
NRZjkGK3X0prrgEVMn/FjfZFRVjMsXymlDORxGCwjjSJCY/qeBlpWV4s7GiaTu/31rmsJ3les8Z4
T4v3qtH6+YRKCQym2Gxq2k7iPhBTR8EZvxFinNSTbntd8ec8umg31a64iYNSrFHneotthLTxpo8+
pokvY/9X9w737xX9b5/wRIXbt4HDEBTK49b8mR/jwC8p62//qqNPZ1bG7y8mocz+2loFIEFA4RK9
4Ajjw6IplSFP5BoNxXmz3dvXT0gjBOwvveTgZ/0q5lSG8ATFrpxS43zIudtQOGh3XdZWPB/qGN3i
ypMpF7sAGducnUQtyEqr0Cf5waEcng79h8ExOx9PzbLP6iWP9oNUDDO9YmWaIrjOSmKv98tad461
WucwyZ9PHsWfyy1Z5QyDEPXUMxfv+cBxgw7BS/1iJbvF9cO2EuAv0LZzpc2MMyKHBOL5oBDkrAAk
8CWXKhfjpXKmqbnuuw2uGKqEErrwvz8mupXcrRPQv6EuAjkVhBINt1LHVKZEANyGDsoRRlbKg+Nu
uCYWwxVKvfDScjV2zWsBQmivB9dx1Br+UuT4/Yp25V3/p8r2HikYvV0m8+kNMqZARJ8oiDeq2CRv
JiPvnANLLhLMoDD22MusOKHaj8kZpU189LOKNoZ0rgh9HWCXZVSPpEYC+wc1qXMZOjUVqG4SXh0n
jA67oiQI7rplhtG7vlb4HNFEC4HUtTPZ7Jxm/Kc4mVSkUederoiXkj+QT3LOgFbBRWKNdsrKZNw1
AVWk46DjTwGkxkBN5KIlvobIKO3cOOeiv3YbEEYGICKvR/D3fk6Lw8fmtuVP/aDIoy3RkHbJ7lec
uN/OEXoN6IjgVrVQabJeF+3wuXz5QGWcS9L00wCJiHQ5lQy3uusmTMWR3VCqFE3xSy9lpB2cBQE6
dW6UK8XWu7unZr39Tnk269AiBkfpWd9zAIgGUTJytFCZNtg7SpObkqQHLsbkKxG91qHzxpEDbB/g
KYcOxDZW2rqc1nlG9C+oOVvoLcW+q6XERatAM8wSqiTWvIwLAIy4N3b8nLpSW94fuyd4oasiZif2
eEqZAV6/hTQ8TqXqTnbkibeIVtTCVhdSTMzfNmFNyPl2UFbdUsMR9Z8uMNJrp8SFbVZ3bpCO6vAi
4OmJVUk6bKD3bhChK/aXrRg9EiOcRMggyAPJ3pjedCYWnFGNl8d8xksfAZAYMtKogWMIoDZiVvrM
ngfbrEzrwspyxa0Oluf3K1VBsElGybV8+HH+jvujkw9hRrBhPdrfpOkM9HQK9qic3tDZrIFeWk/2
nDNonFsG9lGBReIs2TztbUIjugCUMYHWTKYultz2ts2fUbf5V9ZazJiDV30UZq+EBGAhflGlLN5F
a0bKK1iySQmFT6QwlIwr4Tl1O5emHJRhsQe21XTejkKhhdfBnAX9R74NcRAX4mo2H+AD/0d+N7ri
80JuA8Mt4NRvuBsKgKMfv4WJ+G25dhQJhlWg0kd+YU6Xt8gcjii6gnAtcKAXg2c6jYXFrSK+2OKz
CuLhUYkUAxOzU9TTMrSZlJcNUjDYSexfLeuNG5VwpmlPXORWaw+mHtDhWNaSdXVPETaf2EUaAdRf
IwsC3sDYCiqciWYw0gXlGF0P88KFglkgmkJVPQAb4ecsUSct0EQSSjJrAgXUSR2qRduiMzLT2oo4
nBIDgD+6+z6dZ2907bxuNwq+NymPGInxVTA0uOPW4Qvo5sfupEseJAecyCAgSUttXPfMYVKuzhxo
LTOzB7o6duBtWZ4zvELho6hz5b+S+K2/RK/hfU4I5ZWRX9DEwoSYPD5AahR1uBJY/gJxfOb3haqH
9X5YpSA3/NGTOsMgKw3D6A30PZ22N3zs5lS0AWuMPOZjy9cmNUdZWqpndm9r7NVh4rtaCAo58ADE
bh09ryKi9xYuFqxzbKVViUVDwFbfWv5oGIqjphFOtU9xgBoN/cjH5eCvfxws2Q+sgWHUb0vKKe64
Lr1u2C2ydhi2OzYgK/Z0C2JszZf8T7LruI+DyHdNmAUAI9rec2HPBL8HCLxk5/4+2b4I32Nwp1VY
tr2dgdCEHKeGLbUuQV+SwQiifO6OwAB5+oSuWnq3UjAY0pU72KNbFgC7KNBuDGhrPXcP9rCk3J53
L5Fhxyct/jtZImJy8OETS0hvg4dy2ssMmwp5B5KBWrEwsoGNjTBc2jDLJTbvppt1bWQdme18+GOA
ZdVOeKoIjkacfsgLKZsrWiJ6dVBmAMdmL7AG+LwQL69Qk1bew4JsyReif6rSDDFnxVzoJp6stp7Y
bKI9m3tF2LDF7UpAsopYfHh1EbIMEHhpRcig6Hy9+3wi8GiM/YNbxFbWxc7FkEx6ZOWrPgxDHWjM
MTkjmqaIGR9CVV4QPUQe1IHQiMkOTFnhgFU2eGQ88goe7G+tP/KvRBSO2+2/wbBu6TwhR0yyEdiz
17wrYhkmV/SDykucNNK4v9CGbi2Ya1JAI01YvigFCo1cHCKOBkP8zF0VKnDzaCPGSb8mdXXYZlGO
xauAvMkvGWDTa+CRJEAhvzwPKPWrKBERHSGMwadZT2VWVGSm7TmEwcZwdwV3IEakaeo5CUZ/y11d
mx7A7z6PSihqbDOX4Erb7iuY3R1l7lLmhZ2VT76zJw8lGZKqkadmEjrXfeQ483IuFq4qRTmPbWxF
/6Nl+CSq0RcqRoGrgFs9NURC2nTCY9NTOc40M/a6lZHCqaJWgG+CAkj2NlMmb5kz+AhAm7dnDJbS
yuM6Iadsj8bJXR+ERlPlIHVOGQUnPDWKyjPsiXZA7ZgXZsH8czYzlFbEYK5aHMRNv3ZL0N17GB34
SCa1mCXdD1JGGpGRKuFpQADCtI/IGepYzYmzK6wLvDSeUJY93M0kOZVBYudoRX8/vqHq0C2jJpzy
mukGG1KhF81B3iuGqycSnraqE9Z8GndJ2W9d0VMSAZVkt1TwhEg7ArWGZnZVrtz80dHfdSAgziz/
Zcdk1G/MRTap/sO1nM545jqGP5/teVJCGSz+FoWb6Jz6ClH/hWEGQJ3GU1SzoBdGnriCv2nLEn4Q
y5Ba2HVCTQFAuv0GrHdDy32/3urwQtJiaDMcQXa8wgNx6p8KMCIbVTJkZafHeH8aTIocIcSpiB9P
g68Ugxd+nFqd+3sjDT9qllQ/6suTEUKurjcvGBo6MyMsvcU/BYX/L9Mkd53u2PRP9bWQG7LCoJCL
Jo6qCw9kIC/r3ZNOVFfEdKdFg/wMmk270mJpjmDNNBdZykl23/8nS7V9v6Z241g03MRckr8wzZwt
R8+WNIEGZfkZYSWkClMFGGKUKMOMbg3caYoX079sgUGktDH3szUsLNZS6ZdxiWq1XcXkUEu49pSL
kI4KCYwppGus6b7Fg/K5YGbpQI1270oDY9JXnBjI/UBPiVOKAVoKDaYZWuQ4cwN/0+bwuo33R7jJ
b1xdNL7HRsBuZxrsWOmr8i3G2mDmOczCQZKIwjbjeUr/vj1rm2Qf//8Fer2f/GHFSZUXx5sANBdL
BukuHyDGoPBkgaK30cAB1qOixIY=
`pragma protect end_protected
