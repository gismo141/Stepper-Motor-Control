// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Q2zd2K9iIFXfvn25MV+WtJSvaCH+1naeTcWVGp03C+Jx+d1gEOkzkVdm3f0MXf9ANmMjC/zhU8h8
cu5TrjmrxAlMTK5jZC4+j6xA1ITFADBmo94k5mqRe6SYvh8LiSvZbM43XcOTUQjqwhNdXUdNd476
yJCq7j5gjWaFjUh0cFrxJ4FyFCHD1Eeg4hDrd6hJMI0jnxtiA0FfJEXPRVvwe1gIwzNJUUnfLv0G
umd0LPENBTA959jKryRY9oFZELhxaWCKSG31O6wPuEO3pInFELsZxC2pSRQQ3HDq60DfLzc5GTxm
rn8sji+k65USLAeQ1sCPFwaA3tDq7l4YlCIR8w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
3grhszvQDNeoJV1WpNNjCxPvHv7URcp1Riz+Abzx+wAuVh8BP3ZHbAXi8VYIBVQyD6hVvgQ1dEiQ
QVIVcUI9KnbzWA6mQlhMnmDohsH/lQC+ekC7CXG2iIW+V9OCn1caqTVgrMKDLyyUasbJ0O0uUkPR
LhBW0QEsjO5AjePwzUq5S8/mH5BNQqc56vd0SZfVJqR/IK9jjVjG6j8Gid2lDzlEVDp72KxMAgaM
0zeZPnA2QRpa6CGDL2F9GFiktpOKGQC6uCpm1pTcdiuha6bmBDkSVs4OAsSGV/4NJdkxHl082FVI
i46h+FZ8+Ky0vwpcM9+X5ibCWVeSj4gNSbS5JwRYn2WJ0ieNPfVCADWDFRG085CY8m25y3IG+riy
8t/BIPDf+37S9X+mMvEPh9E3u66/7xKvaol0doQpBNeckHsZKdA41FKG0c0sQQIumG2ZE6KldIHw
dLNR7V24vth2jdafqPrFfIVu6N1FpOs+H2pyzi0H+zI4NDgKVLJut1VBS8oymfV3+QtF4p1iKyLz
kX1SnvXASSpyeXV6iHoPptoxWNDzr2mgQPPmU1IraHa4jkHRvn1lu0iuXtiw6Kl325n/PNiKVK4m
11mUUdOavigsj9Bh51zbSDEHwkEbR7mFS9o2cRLFOhpqL6JENkNnGi5RzhRDRiXlmGgvvKvHTnKd
LmbYl5GUXF893tQzWTpsdJ1T7jnmoZRZQ8WyIBBPh+wIMGm+1iWa2SNMisodGJsFYzhlV7lazaQq
XlLUQnttytIYwX+6Rxb16GODBGrBl9uJP6n2prLHiNBfHLer5ExVQA4Sv3Zm9AzD+xIGJTE0eF2o
4Ka8a1UcPdL6f7oNUigaylkeYtIbd/91g8hz70ieUVb8YmoC4l1i94G+yHcC2ggcg1eCFG48QJdb
O71ie5e+Zk5zhszJM3B373n1hC7N5QAsZio3DD8+T0j4F3QRVnS1CTZ54ZtQYBwL5OfG46CK8wja
Vuzpi4+ZMAtvDZFvWVTMuHBY2rKeS2YM5tTMc08CVPXhmTZ0iQoOb4YHMlOntcL5FAz2xeVYyQip
UwiB3KV8+eXcEp2HYxvFphnluuypHq0GeCG0DdhVQ9RJhimRwx/4vWLQmBLjFdUtD0rL8crQ60rD
xPgqF43jL+4Aec1jYZc5d12Gds0j85bt1SyG04jBFTaR1bNFFdUDHbthgWivs/NQnhoShas9MQdz
5qYRu8BcFSnIbOvyH68Yg8IIlcm6UUBIsfQhZygPb6zLWKg4gpUupMplicnelsitilFsXCJDGbft
K4ZCsS4p7iN6t2rtX3iv0WDXjBWYKi7Y8w3mqnS7hMx7U2Rb1heiYnlkr+fkNUHgvC4Q1Lck2k2E
ybiWMEekLzOLtKTFyZ3DUY1n5ZyVHJrfGwkQ0SAB7jVssuU+6GE6/DVEUsUULu4ScnanKFqxq7pY
dEQaaiPJ+FZHGsIye6s3fBzQHfyFThhB1h3U6zn39m4RJrpJaSoY0UWngJ1U1MYJUuXOHdfe/Ag2
WT/t6X7NR7GB1wKKOU4UzxpAF19wMWZIN4TYhov9AKjawZeAcMop1hN2iqAGFVPH2FmyGYDpKU9I
nDohhtLtbfP1PsLgB/10tPp/Hth/+ap0sNah9ums+yL1QGEfFWlAFmWL9O0yS8b3ggScN/A6rXMP
jkWlFkIbDv4QLhgbczNq16Xb1lGa5Rnx7p7q7t+SfbZO2vCZQswT1gCy75JCY2Q6F6JFGV9Crh4w
VW9Rp+JWYotgRkrK7TP9prMm47f5JZrumNM/B2s8yonn7oeP+dHVXLkjGqhZjcHodDAi/1lQHKuM
iUXRSW87Sd5f2IPdCzbPOIKygLR7mKouAI5AbOJ8mKobwkWbgQYGdzRfB1hUOtAV7UUdMuF6KFGG
2WCmXMw7b6elbJUrnDhiPT6QW/qyIvI7O9CjkIClTHTGTO1PxVS/GDiVUvDEpbGwrjwnKF98vDa4
yt66Y7dT+zyWK5GfW7SpKzZ6JOT+1szKToD01V/w40j8UEoMzcPD7XQGnZr9UJyPU8guyoBLlapZ
EwR49EI3LshTONh3+13IvCWmXAkKIwrNoNesuSMb+jleQ903qczmd4vBDrLefMuZYEVGj4wR087h
z8o/ZeLW1JkB9zh0Rh5FRThBabshEMpQpxHIgv0l/oJCt8THEiunuqGqi0udA/hdPmPP1XgTHa7C
H7HObPqji6MpEbA2TVM25w6CkdR3LvXLtMPDIUIZOHcB3tKthGF9CsW+rO/iglilGP5MoHm6pvSB
yl5cP4+UAQjhUlfU+WCR4+uadsRzigBjYp9yNEYgiaPIlAMMsfeTZxZUcZLHtDPYvUx6eHLd5l68
PFBa7Bf4a1cUWLd7UM+jJpQr12gIqyXfAij8Xr0WlebBC0/dJ9M9ym0HcC7c9NB/jCLa4AZoCUAv
BMcJyZ9iwsDt04aQGfbNxFx19g5aHVcoTy3/MROguXiQTZF8B3vsO05BTRm8yyyUMcxw57rIKglA
kSYGSfBTJMpowePVyao5a8M9E1+bLXZukpwyfAm8yRX83o/mfQ0Lt7VPgfvYDfxoLnZ6FASuoXK+
6mF942a8eZd9YMaYT51/WhN3b65u51V+ooi+klrSogJgVc9/s1Zw1Lr4GsCPDreNQHUAxHvFF4qP
JsrTb52rXDHiGfaxXZ9YYYH/uzYviaocck75Rb/FrRQhLSH75WOElhDrg9BYu8gn8GgUUSKWYroz
svIIIgakPS58imcW5U22VXXfwaD44djNXmMGZ+Qq+iccLG/22AJ3+qs9uEt9bK7kJlyGAccQ5CN0
Xe9QsqczY+EMw/TrLYY28xaFfd1lHozBOe/8qeMGkjHzECGdg1pbo0A1qktn9yQzL7M3W/vnteTh
KN60GEmD9E/LZYn/Ju8rBi9kulJffJ83NrjWUAPQi3xDvE8+Faty/eCdqao0jWPtlU/6V5SPaC1I
gMmNsBQnvmoagZG9LkLVvWVqfHZtzha2Drd7/jpG2gU3QNzaTIbwY7FR8HX1xXuAYf9O5hu3OLd4
gGzaHFZqx3ZPXn/QyOPVA9Y8S4JaKwjd4TfwwlrZc7K9YTZ6yHj8gi6jziH/VpXxdlQfx/9uH3IS
T11C7T4mUwYBgrm5OS6gJlFefR8UyC6FD+uxHPeEkhKhJ70OSBgEOxXLjV0gfizCMSyDxXb4dH10
+3G7HVxR+LiK1+3LqchgyieorMCV1Ls1M4oZKSRZi5Z+KcA1OBkFx1N93qvt2gmtSJEYfnLKF7OU
5FJm5w4w9In5esEh9EE7CkTgPMec1vJBJsXRGUnl2rBPKr63mQ0wnM4XA5zp71BZtQn7mrALBIjg
oelLe77Go7+cPv8AbfTpSCCg+5dETlG6ZDevvCjn5oBoX9i/XsINToPUN7ssi1ceZIEKz0aZY0mI
/4pWUQQFKXqEW+8IHkTfHCdKzD8W/kO8F55yckpFBQgYLiDUNbMaFAtL2nJSejh3HDt0znU/239P
UG9jaZIG/4Z+V2SgzsUB2f4GFblb6FYxmqzhDPy8tJWxKIOpipsg0As8XseafZaoZpebJvGyYVc5
soXj3hcWqs+bMGf4mfSZqSQbw5np82NIMjVuI8Z7M1DNigYYJ0q4yaD0oPyvH+k9ZDXYyZ03qi8V
4LKgKpr9mABAqlpTx0SOCr50qwaNcjF+m5iD04F8Pt36qJ7ovvrjaEr+I3G+4Hx8ii6wGlI3iaGG
zS389xWLr7Z8pLy0O+WbJ/baGojDDix+Pta0mognUH454Bb4NFgb+tSQUs+LyUb/ZyEZUOgBUjYv
ni6CZ7LP+LXMdXH+tL2GrDpClY/M7r1pSxB1y/gQbaSXCZ0A/+eScx/eVMf6ImZGVok2giBNhyKl
526kXM1zG2YfDD+npub1rxVrZ/F0ka8Zhb+sIJGDoF04qU1nwbPfSzRzfjkbwcrlLYSQiw2wFPMR
338VDCqcX71Ksf3YAP5qvGuf2QBO0qAjlbE2FR/wBV1wT7413YocFws9NYBRoyel0CgZ3y83a6Pa
/ahQZ4kgJKQ9de8wijLA6MRwvtzepMDgN7gd+FhNwDFs8XuQO7V0vrKVXFqXoulZ1lBgHCAEIqMq
l3tRmxWNN8HVMfWcXTozl8psrEtFie7S1vVG5Ov30zUFzKdfYmUe/K8Wo1iir1di7hn/mwnXXLCb
il+pajJSNU0ELZXWdCcYDZpHNCG4iavBU25gVU3bsvIk7pPIuheQtlLeTFoVB6GF0f9mQs43u59q
FVhiIVwS3IkgzHnkdlK2NulBmMVU5dYvH8ZYRZAEfK1/R6wrwGsUcCkZLnfsV/bf0/1zg4KZrBIg
PKaC2KiuM0Jsg1PSy7LRzo5/gWADeWCWSHa09tR+SvGSn1TAxq7709RHAWMfjBjM18FgK353mEBc
RAGqXtKmgepJWwQZBpcKRShl4U1VlEqyio7ONVAqKnRqZJIxvVICJIxVGbrwncxk+9VqSOxeDkv9
VbG/KmWEJjx425haXchIqmg1YnhzR4cdYzOZ9rXv/usRFugHHpdg6eJs2T7BK2FVV2uL8PyuKK1R
+8wCY/wml1/Esu7FpGAqo0/yB7sNiN/Ptuu+T+xRD1Hcg1ubZrot04CGHVb/l9IeQUztyc2cUuhU
0yvI2cAStNAW4X3erOjM9qkixQcWmM/B7DgJ2Vfjah7QU4d8n5XTErj7s5mWmcn+GeycUKm9PAPW
Z/QAhc4sxX/zs5g8/eVnjg/w4vB2dyA/caZK3IIkmxLuynUo3cIyV9n1w2ePY9zOrAMwKwqNmSPw
ov5zoYMaGiS+NzLAUq3mfk0UI4gZbYjmCFLllmud7lcTz9S+QD8IbbQkz96TQ4mHbOyumTZP1t/a
Du9M7CAPZPfmqIpeQC5KRDKoTUukwXVXHSZ45LKQLc6RHJJq04PaEvgpwy+GwVc4rbPNX94fYp/Y
l+JECUt+JwE/Esyh6RVMmqfCr4qhqOYlSErqvbYNlRp9hv1nltVUJFbb58oqQV7iGOrvRBsCRUxJ
9ZyfxoEkKbdLdHUmgHPfWhR1Sh0ns0w1gcpAVfMm/92U/CxAr7qXCWtmvrDk6L07JYAhHuQNqwxB
syetrp7v9ml2RhtEpU7fQgaMOflZNoZN6huLlkdSHlR3XpBn8qluccqprKRvpLLRVGQreY+gYLD4
kuayxzYgdn2qOfPttUDQZ86ki7hGZSCiSoMf9ef7d2vB6ewaORfOGQgbhBDh52RufiuU3EUSAINS
ZEbyWU54X32zADfCZ7Et5XV62gsRN5RKqEjm05fIDMXVhpMO2joFfpZWWiZBfR/YUEzQOV9P8xOA
/D36ne2wQ5JoKhSxYUv2uvQMdH8TB+JHwtaD1A4X+mSd1CcHOCZPxvRqA4yxvtdx+Ee1WIJ+imI/
h1fVOBFa2G8DHImFrEy4qMGve6Sff5VtOrrGX4WVblZs6xRUyc8tJvjrBYKmiBXDPmEL8X144SHQ
KwHwwSkCI23KIO7RwGyey7125XWpiikZnD+24YICMMIpIef2LR/Z9ZOCaDAM+do6ABeChzd0w1H9
nrY1HsThPMw3Ef8utZBdoPMmzqStLYYv/8qqPzTw29DuTzNrFqu6FEeviOK9c8wGGBEX+hcyEcTz
yLipJvarmGadIDZ18VoG5sgNHyGOr9sphdITgwyScQYJ3DwAjfcSytOYbQ49z60pambhby39wiqG
5FqtF7mwuHuJ9F4hhADjP9+YkbV+lSVjlYEDOx3d439yhWMDZkQnjCO1vjdPoIpj4uGVObbNCxW7
jrOpDnjPWd3qGOTVo39OYYiVcuL4rrdwh8alMJBMjjVRsSSEg3cYK9O6KXqbHa7vZEnvOZ0NlOjc
i/0mjuFBhxnnX6Avg9y3BS1Q7Vg8rUzCEfmcadS9g+9rZQDtuhWPF9D/3f7NjOEvI8X48FWNqJiS
RnZ+5xCGvLRU7rqEbD4ILfxL92o/enntPSyoGlLTSrILA18Act1hfl6CMSYvBW+Dxt5FgXgRuEJR
ZVqyZUPfkfdkabubYrjd5pE5IJHC/Q+94kZcKzm8krK7a6jf449/sznpOAJg+e/TnZ3W/Tjqfqcq
yEraG4embEUqzSBgeLAgfLeBPq7G6+Zl+fMWnF/eBDFaKcHYGBGKqUYdqtjH0Io4nzseySFTcM/4
9eVadwCwZFs2xXNGXNeBOft0ozMnueo3dXZTBObsNmUdAYyWgDlYmFHOmYDmE2N0SgpxXc7b6pfa
Y0qrF3s2f1lTvAPJY85Lwy+YhpIBoR1cAUJf/cD5qH9ZYXEUxZ7gE/ArDkH4BsNCYziaX4ENCHTs
rl+Y4q0WOTPQFq2+FwhKxpAgfcwfwlOVM2rIxlq62fhcDR6eFZ2F7QM0RBZi7BELJ9s/L0SoCnOj
5vECozih27vkCr8b8IbAujl8X0pHvtFEgZf68DWc0pZJLL6GW+mP4a8uP/CDfRR9uOZBt51xfDqo
xuRt8Q44eOwyIsXuoqT7792jL/de01D/uALT026R37PAqWarClwCK2Xao9gjHtR8uQyu1TZA+0rm
lbvguMQe0mQNeAhdRGZUE/G126UJBJNbj7NMCsymSXnU0mxdfuQENdcuFhj+rhvsJ+ja9Z1dfG9m
RXG9oPTBCpwdCdOLn2s53lLQNmJEGWWVQHv/yvplnzAQnp8/vgJiEwyWY/P4k5Si2anGXjx9UR53
7YOEUCJGU7812BsaBhbRNxqTQPP7jt1WQdsNPnqAgiVNO6fYeE+DMpNvmqANE3IUCacAlgx8X20I
UZW7Kq35LUwL+8XIQR/MK+4iQSpsjQIgvSODHpNly+coYE0qJ6v9MsR9SQ0ipS+kqLymBHepbb43
2Zi5KWf7H7lriTdFMJbKLgDBk/CRNDrgxvb1X3mu/uj5LPfKe9x/wdSozWLrFKdN9DPsW7KqcSZS
ehAjgekfA/qnuNF9ryco3mQrDu0hkvVKxEl6cR80I397OJpPKDjBAPaN6uenInYO0/4+1vwGQL8J
3EHC5KUoZVCkD7nhVDuBkYgyMfficMCDDoDlXnRExJh9agiUPLYl/aQZe/rqNksaCZY8GpIBIPwc
lcK5N0egsVFYSX63rLQcdM6TjumHNTWfNPuiSuNBNoAuZaDuWSM456+LHPJ5n1KXN2ven8XFXdwg
UV0PrUncCe4y6pYhrpnai2p49VBVsjnp2xbKqKYC2fEj6Np0fAil1O3FcUOaYVr7zh1iMCOVXeKg
4Mt6SW+cg45eVbzuez8vNP9sQEMvbtlX/XP/EVM8NHxc7rReWyLwl5AbJSIXeqcubsyWpmxO3Hfn
i1dhiacQcLi03c0P3HBrToRMVf7Rdw745Rtw7oyqDan7NsmAXtqohOJ+evhrqYD7ZeMmSEBShnf2
dvqZtBKXumze1158jdjCNTzDW+JVZyXQVbqYN4Y79cL49aCqth7/sWI6fe7m1DFmaNAQZyNeU9QY
zlNWY51pTfDRa9uY15j3REOqS6zCi3gZoeXbC77/c+VvIHAMjJQLOJQR+xUKIeLO69v5dnMsSJW5
sYrCFZMvD2f13a9pXBljWyk6gDUx1hJFx8i8/WOy5Lfan/rCYf5k12ksuz0sIynRqcVzxzBJhVzI
vwTCzhOL/7H/vy8jJtKWDKPuO2RhtD/atfJTVTZ2ZSf9l3mj2pnhNHcQPpT+1u1jM9bjreBk82/j
L8ns2JzC1LSTMOpRaK6s0CG+IVn8d9TmQWg8uJsblWSfd2x9d29arCMUvQTJyhgLCWGoai1RzK3y
ZyqnXFZm+gT+lGjh71/jDQVgyvbUtUU8MvKqJhYzGfFgrQyHE1byvu8Vucowb7wgxyW58zHuKdYs
PYgMfX0Y5vsv1D48L3Wkt1YXfC1uTyV8eeC6f+D2nHlqSQpZImmuGNvPemvQFxux9PcZw+4F+SCq
Gjn4k8gwiMRu5PN1KC5C/IJeYDgsGKrHwEWtTblcsaAdU5LosewsKIUgvKK2tqL9P+WaaYBza1/D
ZUC2R7O9Zb/nGxzFIElVDE1oUI6Peiyufxrdzkvm64HaAWQqHEX+xUe4mRFr9EsHQn9/DKmuJ9U7
JKad14GvFJ1MkFviDVN2POxz8+hlnOvjChvopMXkypnVsL6qaV31q9ZtzoRk1E9U5UKdnzo3AZhk
WhOf0bR2lrX/m8tsabiccQN6oOHELNqmOdNXwMyom6+p2eTnTUa87aEBc+2i0W2N0YTBDkG1jOU1
29SoJl7qDoUabXgSl94GQeyPHLF+iFOHZOPqPZESlqq+kLu06rwH1OKpHOse6xKnem3fDumk5Xdt
JtKl33bFZjpjT+60VmhQbrXbYwmcSemNVUxhyedNv7qR/w0uKzs487DVr2fKy4G/svXyoD86JyAE
rlQXYtBxsBg3ZPmpw6oKzNgwtCrqlHQXAEyLqt9thPkeDzs0OuKuxx2nmVtJK5uCO671eZp4qn7X
jxZORjABGQR3rxEQJ/SiARQDYZ7JCKkzWkKgbtJdOpNeRAwle+kWdkysMZmr/f12NXBxN3qQhglz
YDX3AlNwLQ4fKKLqDqIP+qb6Y8lvFnxMeZmIKZg275kfYOvk//OoFWo3QOZ4s+f7jfpQYs+mP5+R
VfHjqciTqxoc4tqUV2mE3RF/7mXgwTiqSffsTEp9MuY1SJvDLi6HDk0TWSMVSRUbIwxHTaYLSqY/
WDn59drLLJIDWCuELzGsbrqyI2ZxagYMei5yHZP1+lIjrwfyeItZuQg3FT4Y1+BR0kHiD5v8807S
5CruAdMgE1xMySrJPzZxVet72pf79WXKS7fIVsLyJ+Xc3KiTQGq0c7ePI/R1Be1Cu19ACBbC3vvW
M49fnabjWLZ2SRUXc6dDxi1+8SS9QZXGA/ho7khCGGTajBNEiqPWyfoTgbk4IRlI8JnTPup68gqs
j2qWDTWgEVHNV2XZWRjg+gt3NnMpIljQmjgmWjFNi5qXYxFaJ6ww9uewA7xFqWEnRMh8KVYptUTg
gMXSvqdRe6/cvt646NDCZ6jslllh/d1aYyv9gUAYm7dCGFWZz0LCE5yowl8/zCrDit0j1ALgvbUM
Z6q/vDv8odOlORl+Kw4S8miEAlsGuVcutmhsKhkfW0Z+ViLZgWv5D7Kt7JUabrcWlRf70Z8Tv3B4
nCPyrJEof3vMp4XA0vkK4+aB6mhWWMRoYMpJF1umcGc7N0sF1DcKjS1ERc+bBT/3gBxT91ATjC5j
wBug3dzLAQCnzEm4ERAW/9BAuZAgzTkAF6emm4LUrVy+DtiP8mGNF0rDxjTuuFJ49e+YHGcuQRKc
sfuSLc09Bm5zThsru9qEnuu4c8GeYzQ055boadgvD4Z+QFThMj0RawobuR/y1GRyEKYZ1wKkMVZF
qyFLmOadeXz6A4OERXIFjXDBica9md1mtzctH/HRhkxvmUXwbvsIH7pw1371ny4fIyjWiGWr9Mdj
Rxp8O2Tl2B7nBlMhSVT3NH2105MVpZq7k2kWBnvhZbw/Ae/m6Ssqa4DV4DebDer3b6/ZPb9QhnXl
uRlU00aV3d77inlWUA6HLsAzMM78OeIRmStG7eT+QzOank/IXLDj2LdOQgPpk0iYR2osYj4wvxGN
275ArrGtgF5JL4qA8qfuwJyUCFJk/NHmgJe2+yRSGZziTWTa1uBd1XMxMXxlrwwwA6B32w9PkRKl
dZTLFYV2uP+52eaUrLRJinfsfsW/0KO08QGzpENz2f3P7h2AHzJTD06Aqo6njABb6RJZmleIWkvN
EuvT81t005RntIjoN+FkponvyEmUtEins6tO87Oce7ssKR25pW+xv6sOBUf4mapRfpc/2kt/CtY9
s5FRGlp9pcf3aBl8hU8BZwfaoAETvC9wR/1qf9dhLDSDFWkfzqIrN5FjGOh0zBcge/otAWoitvek
GjOxLnhCT6KmHL/K6PRwWJ9ivxVjhSvf3X/IQ0CEp+3zpbfLJxf6LF2WqNUwB5h1+4H/UMlF1ckK
ufB1EmKXX867Usvrgmwns5mFMJrCL6VnzBCHt6eFbJrtFS8wrhNkg6paHAa9q9CcoY0p5YBuCGHP
kiUkyal96Wv8VNb9DJnF4ekdrfnvquQYZ9YTAk+QSWYaL30iH6ISSEYlidOrSyjWQ3WP4V1byKkX
64UVqaqyRDylJEgq4FX+xOMI0s4EZyezt52vhy/Ov9W+A2H/sG4dtOJ6941hsw0yvhUpg/wqNvS/
ip6/jdan/os3QCv2136YC38eaPrtFr+sOCT95NyOiXidM26pCxpeTkVUSAa41Kan+wRoPLN01Z95
UJWbcNaa69JgeJZd5MbMG1FH+HQwGX8MzSwCIepxFdCT5hFlFJAo0apdlpJRGxTDAlykC1LTDXx/
RhVZFK9YiAwjhW9IqelL5afIkicmY6FxtiS1IMteDzoy0eHkHHc+YE+iU4QqZcs9lo6aONiSimrU
WalaxjbMCVblRvL6KX+m40JbE4d9YNltYbPrzZ6Bx/qZ+uI1bVpEZrsb0dYPjwWyKyPk/Klzu9fg
+izFallch8Bc47BHPzKLvLBR3TZKckaocKw/pCdyZtJanrImCLOZIVdRg8+PVZ8vaH27Ii0TOF8c
7QNZsqrMHiqNXQDE2T1PHEYxw4VTzpCxxpvyx8mRNlEeT2MfENAXukVkXxfBUuc1HcKE6iVHyulc
cRFqUKwCgjdTEOHDYnNrCR7FloLUgJX0yrQHsgEwjoEccEc1wsxBslFzYYZslM4nQX9Q+erSm5CP
p6HL0H2mf+pSGkgY8d7NDiySGJz0Hxia2EE9u1YmNx3k+eoZAYqcoZZgnzHp9G1hX8WinLgrAD8d
cTTzJsn7kxU1ZmKo6R/iUEdtLAyAl+IK0sWX4fnO3vDoyGAtEr9jBGianpiBkEtiibLNQA1YK2el
9zd/UhzpV3K6tA8F7b9CmMsLbpMV4d3PcZ/7ylDe5R26dHD9Eak+vCs/kNvnyb4O7RILXsatC31A
HCY1Pjx0bdY12nNFk+sSjqw55K7/aKrjLfblHvixrmGw+hf0J2XzB751rHPTgHhJaHRjWz8DcZw0
+EMWB2RCbw9S/IQe7A9kY5rFgqOU0IYJpzYdaRt7TUlMJ3Y90DW5t49kMpmgAYtg60btVfO+IHc4
c10jVZi0/Y9X7sxYqPZZV5e/DqbNvLr64KXyi/MbV5qI2fAOQczOntkSSjurk0oGqghh1fMq+rBO
IcU6NSJ3dmAQAZ/aeayWDz20Q8mQH7b7QB1ZuFXPQJR8GaCPbfcCUffyEJ5yEtkw0rTz6KziNg3e
rW2GBpNJDWRYLQJ7hDq5bPH2/+M50jVkNiRNyCLjZYw/YRbnUMjIeSWbsPi6PaMwQqqvuUDwczwD
I7MFqyogf7ZHhY2OWrp8JhN1Kx9KFcMIn+lwxkkca2gTspSsk1FPBMf5gxLlY15AUIz5Dkkmv092
8tLbrLmYaPBBa1Bzz6EaxlGRaAzseMkkmcDf6zOM12TX87mooOcMN23EvFsdsBe06Pmvb46VS6Er
C4KOwwScoc0j0rQgrCUmKgJBn5lEjv9w9YCPcV5ExQL+kzGuu8XNdL8sWX6iPOUUxLNqVOb+ZioZ
vy6mBFKUhYKP3iiNYTBquAvd90PvwlLaNeShjasOdzfq7gtz4BKrsF8k+lPj677i5UwaRDy5eZTG
kLFEHNp17GoKRBCYKUwZgdtUxiPcJLBG4i1ZhlIXh5DTZ2nSHOSMWZyov3K+CN1bo9eWHINEfsU9
RNQLOSR1u0WXqzOaETez8OQrxza03Dkty2D3KujIGdA3bsFWMGGz39+gHAVmbXHRYxMboMAWh/uV
lC8LPERsU8t6/s4NBFPwouIFxl7puPjnnHhr1IsJk5hRTeuwUmqs9FIEiTRcradZVkHKJzO9aGB2
qtfxz6q249v7K934m2+POVrqRBvb4Zcq6C0AYeAept4wMfx8fW5EfUvVOgZAYRnhjrpVNMG7CofA
yhkr9bvAKCR1l2FTV+6cWTidmzmNlJ+VrYZD0OrNg8bfAHnkwMFxZ1GJnGSuMxx0n23Fms5/P+BJ
77Z2FBmLTVaGBbvAPtggGd+jB9SL6bWVIvAXChv8iE7HxXfKzgILfHt+gEVjfqQ2fMVqTDTxwrwX
VFqWU/u8Q1OnrpyntER4YoMWrq2BBBPcHLvXd9kDzE6rR4wdrY4hSdcR5SxEU8kkUeU1kbTh0YXz
jH++yMjqjyCRWsUakn62WRpYxWnVx3wbGv3n+cNQ885Nwe+NlxRQyv9MC20d6DLV8Qrlb4W/nfqX
m75TUblbvPCruT/YkHxJPKAlEmHD09fx0QCIfJivbAQ/0+gua0WzgKzQw7MQxTdQ1SVi7Ycwt9ug
jN7D34NsurhgfmRR4mPe7Nml1A88w2A0aX1Pzx28gSa9uCiE6lFO4GBfx1RvVQP2aQ7hVgNeru9R
NmIbgjdpSQ9xLLfy+70wraj+mEWeKkjry7ymWxXfAxCPz56Ip1JV+XsMLKPKDRMB56GIGNhiBpDM
FdvEk+gXDiYsFBd5EGKh9R+otYDoyfp9H+fWQ6RltLWWW+iZnVPgpxV5LtZIS8s6BaYdM1lomR53
yTxRlqIpiWsqIqHUjqRKvXarRBimeoe1uJz6IcuVqps4tF4TlX5pnCkGXGvqA8fmQWmRf6hhWcpY
Vo+94cOGE30wO8EP1Ls4LShTGSai4c7jGsdHhDSgqgZNSs2nJC56tYY52P0t/o6kTcB50luA+12e
HA7cY5ljWRdv63WOclayVMb1YUMSRLRr5dtRiuvdsC29shdT6M5bfXYKnZ4KzaG/tiBmka+kaNe4
iIi6massH5gEWMAzF059/XCsYGmi/V3JDoRzYXdJJdzeZyXBojqai80fOBk9WJI2VEnTr9gIlGO5
go5V/jIQEPos3nd0ujlAw8fbaVmAd03R8IUf/gtKZPpgD4IqOr4HC6XfgzwSmVFgaNjjNe1aynEF
Fxu8Y5hVGrza6GB+eBUZahO8QQDqRGRyv5Pv/MBUKVFIgwMa/4ixI0CBKxn2tO9TlWelpXdDC6j4
1gjx0USq30QDzL3A/LsPM8Uc9g8gjCsCdS6hULH0raZWvlHGo5vqVpibkbqDorbOb1f+mYGzbofG
f83hHixuZPnv2ycfXivpc33A2u0cBft0TcnDJ6HDUuvlUiagygKAjWeKhrC7XnokaEildzyUfZm1
A2KXaClY24XCZ1jYRjkViiPotsdLtjxLRu0KwNDNDUzN9ghryzO4ot3+tA0PKDkV+zsP3iyId0QO
dq/4JvcWMnmE3Rv6mfynkXCW85O8YSPYqX3vm+nfvSnYgS+RlDhptJ1NOgYiFK+lKOjDdBMCoiE/
C0ynywyKhWIoDJ4Te5WReAFdRbf66GSX8Toow5Xie4DdzCJg0wqDAYANha7d8KgHi2Eu/tKlxhwN
1T9kGjw/hIq1mDkc1APMVx3/lWef/MkFy0pV33PYofYwZzYwrdQ/TK7LD8xk8KbbejUzc6Div3zQ
oyBYXvDmsnBmvgwgP+GNH3HhUop50K+4HXZ/LMarYUNbwG+wE4QyqyJbuGsp7U9iA7+awQqGdx/K
rxalHdk3HoVvUc53Gv5XQMXTuBqi7eS4ALqXjq3ZDPYHE9OM6JznVO3sJNgkWnE+1gzAfDXORTmp
D5BxHV4PVVRJDizlu0sR0Rthx1BLK4wuNuzFKKC25QiXZnk6weYXWC6Xko0em86UrxAD9ZlKeGAJ
hLHOP8MZBbSD+HsMUHkUPjik8czgVxdMFBSvSmaPy8AkETOvfhNi+cFkXy/Jpwdlb7ylIuvbL+4x
abJTgJ++97tzeNNcIvb7/OQohFYcMZeFhNtJnORcAKXYhTMn9YfO3tbH6E7RDGYV/PZFlS8rmx/8
pNPBZljwEe+9rVnshwRUAtA8IpPLIoXBvp2u3RSTBlTCt+JMIOIv5PUuJfcGxZWDw4S7VIUQPR93
yt6bzQa2j5tBhLZJm0/TWtMRULBwVg7G5Q/5xajOIZZr0ivFwGNwui/i8HqnUIeH4kWl4UHmEgk+
Fgj+yl9/h+KdJbJ3kdICXTJup2zj2lM9sP7u3D4FIVy5hx1QTQGYcPmxKpV+pL958FEPqD4656SH
ITgjimb0eI5axxUalCVfzcgIgONUe4xSeGeFyS7dEgG/dglswnJXtjgiol5wEZa/u1C7i6GLRo53
J7agyY4vhJb3chw4m/llf75HYCW2pQxmye8woc5YAmVgXOYINT0yxE3Mhk7kmrrCu2O9EsoAxYG5
iS5E7E/lhlsXUHihOVBlSqRapYqZa2UUjAjLqlUfUtLELgVLcrkedImPlOiWsy5kJIU7+ySmdKkL
AjNThudnzP5nlKDyPhUQFeZ5/1b3zIGTyMbGmKlRTxEXXGBg8u2BffA+brG8VaBt7ZFXmbldUxkb
isJI6T5C5DuxTTKpD6zO2qtyF4AhbvPovtmZwTdD3aT+Rx6gfFOr7GpE5QOL0TCO+NA6yID/SSgy
dK4ygemkeqANHavhEu7oQ64tK3hNubexbjFMO+YL/YFRpBNHZJ09CGFZZ74QqdS3sG7ZwsYcDRZO
2f5VnRGxsolzSJbFz0jwX3HVtxRco82cww9Niecbirq+ctrzrYzaXx9dvL4MqAgvn2/7PYv8LCB4
HYnMy5QrJTmIHwz7OnAmfYqxmiq9xGlKPYoml3tszqe83OabVSqxpgtytUYLFPKMx8+NfR7rTUcL
gIx2nyFAeVSoS56mdfIgeSTnn7F2Uc7j5VVGSgFtW/gLtEtU1avM2kDNCs4K4iZ+0MKK+gfpRbBQ
73LSZpdsExAbZ2FQTNwPgBrYVzEICcEwf4bLn3icAeYQth10eN8meI+lq1AKX9l4XTT/ntu5u3bg
1kBS6LXf08i3DSF8oJfCxv0Olkgh6UO9+6I+B/0KKR++jhH8IuUB84IgFctlvpVXEDoXSEae/s3+
BZA6iTAVqvDxHbUMeixfGBQkti76bTbZvKyymjP8PaWK+4o5iozq4deJo8SYaXDLmvxM5vGtIotw
2O0cJSf993iXRdgT4EEB0EFL1ES96GvpVvOlk87K/81XG+4djv8m/RQV5QZ2T/hrHzpelVpwDKNZ
uh6rpBRIJoyfMzBzELsYJO0fBNZQciGfA8WKzYNIbjvk0P/MFJQrgUagxqTN28DM8nnHnCIX3S4B
wR3T3/+5H2x9fcqMf1up+ZY4PrmKyjqe+QrJMPTDhAu47a9liWrsbRefcfj/CvStW1lVZB9Xt9SC
tX9f2pXjQXZ8WTbsmEM/nGT3qluGWYSOj3iqNU5SvHiuxhDH5ETgg5kWXBBYImWIAGGbC9hiMuQt
0If35ldxbjBN5CXCjyRTyumbyJVRYu+GecQyZ4zTqZCgmt/izEQIuNVaUthERgm2Yxler0bJwbWZ
Qp13gmHFpMa2ganl2bL7WoSZ+R5KwosgH+ZzE2dpmw35Jo6Nyn/2RsgRezzjfAMb0hpzTitIOTbb
Bk/BuQqfD8pHEeBbAyqydGkxjlgCP24XqaP2NvVF2GK2XIhSdmEzouaIMR6jzVJ+JSQTyOuVwMYO
Y9IU2BqbBEy9LBh3P3izelWC50qcLV+CMOj7Q4uVkd2bUTz51M7zqsuLXQsnJxwRNnJ/yDYWa4IU
Tn5bJe2P8DKmjPQxI21Yvrs67VMYzS+qLMmJAMrzMZVZthK22GkzZd6Gm6C9OPPWA3jRCtrsPgGx
03HYePzOEQS+oDnJmDDvmrsNVKSD5Zv5Q5YdBpfquE0zyW6IF+IACpidtNeT1S8KFZwO8hhQ6/9m
J7MDKf9TH2FcvimgY5O4ZHFeNIUsDhnNUMqfBe+oFkXVlKswpdEBRPwaZcMDR842ZqW63Lxw4Vf+
jrCocKRVS5mBJOHDw7ShgGvIwU18xM3WLlVe0l5lU9SPUqLouY0q0byeV5SA8SidManrDJOj/FVV
EtGtH7HuY2iyivLH/jX7i98oUu4MW9jmN7/4ZgXMS5Va9y+YgWNETrCzByDYA3oDMkIXBUnLumgK
Q94BGmtSBGBzhS/mD3kv2JCwYIYBkk30KCnLCymh9ZuyRRJrSpuw+6Wn5TsChlCsDXIZcL6wAIzT
8QG2hjnJOT3pMUhs87NsXXDzobNB6cNUmNlLBQ24TmkaakByYkhZI44cpaaP6J/V3EnlPROB6YJx
lHI0cugL+wGIA6xLMK+53sr6QYl5TOiRinx7dr7LYcG8ZkXHdm5F9bUuSmGGum6QaZ70yDPLRZFu
P7Uz7OoIiqDhFKJi6S3jQ/VNCqIiMmvR75wwP4ibyBTVOAnx49j3+T6LHPU/rpNvzxFG3hPoUvJ6
EYPqbze222PfMo7EbtXPbH768+Y3cIqND1YiM8gh3YzKAJzHRlYgMDxMiQZGZzmwxS8x6axgKRu+
nANbp4DCMQ+DaAnds5BAIirl9xc9K6sAF5eIfeqKaPDtGYQ2vZTQEBKyT8kseviKfWl8PPJfqGpE
4ESPwm9gDa2u7CLnuzw0fmAbjOvCaW3VCspjvK3SxoJoSD09IzJ2BWnboNNszjpafpXGuWqavbxh
PgbCzdXdMU+FMj1XUvXIWq/cP4MPUL4yxc3CdRAdnilZuNsCgbIjjvpZ1T/xyfcGHvE3h2f6/yLl
FR6bHFTObHPUnB7EVHUA/ihpNiJmqd76VndzMaSPtNwVwceGalfESEonNLdXqNJ4j5HoB6MwcJ8r
+1IaBgXewok5D0E8avsb3v4/Kk72TtJFMJnrUEbjJRR8uMqCTjJ592L70wLgLChdFTjEC4CdDVaz
JHkyS0N2mUCj7xgWdAg5got+a5a7B3RNViGk+kYHVcmq+H+/qCUm60XUBwJuMYVRMy4LqddwDsid
gUHzQmLguWIaU6yUwKNEwWqmdRe8LQOIhZeihn23HbEDkvLSGzgjDndAKc/pEiwYGlpY0e919D5H
k5AezdmwkXB9lqTmzACObOynwneCK9QJhB+RCF45u0o5etk/Do8DW0IQBG4LCaomQMV1XlA6xhHV
lYMNiHpWslI8Q99qSvzue9VURCzp+u/Mb86oa2Z94cO55eyhdaSQiroSt9IHQ+TxF6NrFNtS8rkc
fp76rYvff7mDYKjd9vnODLDnYFqKNcSBt7cDM9gYQGWfMvV89c9jqZdt61LzIyZs/sqlo6j4+au+
HYXHlCZ66jgC2Msxl9s04eqWF1zWkjDbkvGV7f7zuUzcvIlUXqPhODfNzFa3KLr6IaOrKluYP3FU
/qapbpl4AS97EpHOLV5lQTbHpwGppIqE9W6ncyQEz3IXDQvZWW6fZfNlm4APVHG6sIFBhWBQgINC
frrBvLvC+2aZYDMp3vzDHF9KFNTOBAs/dF/rtZDCybuaIhARsaOTl2eGR0GuiRsJwY0p8WpS2enf
sQ/Dei6L126nGqfvILTeefd6pkBE3L7AEruRo0fAXsxef7qbzDhcbYIGvnckdSoBPLLTXikdPml3
XKY8e+RRzjWMenSSFUX8CxkWC5U7xSvO5CziWHFqTOJR+xO0AWzSeU07w3SkhS8/d9km67hC8Cql
p1HNAhBjVfon+XGA5GY9WC8gIfSLULCqgQiE3Bhx3XQHlZnhiDAaZvxLIVDZyBF+I8+L6RauP97B
02qDmEj1MO/zY9cQ7f6jFAcPRneCCDy8us9Y+nIzjT08SP0Go3g0kcdnuseGAPB+ePv3feXY1q9Y
X8RVAsY67bQuwaZm9MS1o7PclDR7bmp0PrUEZW2/9SI0Ki3VaRwvoMM8AscJ8lmv1NCFAnTx/+1O
zB6NW2VKDiqFA3frn3Lnrk5rlSrsCmHjICSCMcLeU+MWbVKjJNofB6TNji5VU2kjkxPRiPcZH3CO
WsiYRsNqWMDslACIUfCB5R1DYWtF+0ZuBl4vRts3918gkiBvqT7y4yGBOum0CDrOiVXXjZRIGCzp
lzVhdn+XuLnm2Tf6sxua6YhDC+ern88cGMzMXUF0OWr8nEXbeEcgLoLciBUWNYMzCn09X6w+b754
x23ZfQ0RmBftOBG0VlE59FV8Lph0FgPghVExIvbk05VN6duxY1Ry8MFv/Y/gRrGDe1XivD4f5a28
/Y10mVxzHmUFx2wHIkxCztar7Xn6yhzLONg5cc6Q1mtkqkH8EZazvd9VgdHb7qd1WQkwiwplHZw4
gdhAMCHqx0a1KVDAXHs8yTrNT+ihm/yZJXhappc9T3nsQxYwx+mnfBsKEaIsRZKknu4bAzDcji++
fhBVbNe84O4C0XdH3Wk5ez9zbgq9cgUKZF1cEdwbuFJhJ5qa0wVZG8vHpyty79WOxmF1twDRSWjS
yX5L8QaYNGx8PrTZCG2C+/NXvGek4oxylYTNra/L7qfVE+1KjicVj124eQvCzV/PcuN92eyF2039
pEEeRrNUrKDNpWuu8UC46Y0b9ehFiPEJ9o8hWFTF/Y7JD+DDxPdGOxSvVKC0UcBdJPC8Fs76j9lo
aywlc1MjmDyzZIrkiIIO5O9sseYGxURuef+B4m+c3h+BmDYkZghPXinL9khuDD/jdi8RtJV5jWYZ
BFfQDhjZ9JQOHI3wEfjOVZ5N8Mv45brJTdUtg2l0L1elBtAUgbPaLaiSOygdCUrE7BgKghyPJt/J
QCuqZACdImy1JSI3EtGeoRDGl3zTCZSlB+8LLNaQYtzTRbF9O/cu3PhRY6m7tXeNdrJJvRDpcpXr
bZVa/XBrbE+SUtyKt/MXyFJTXSgltXJZ4x6aWTSYq7AO8bYh6DQ+3/hd13N4c/suwpKvHiMI1ZcN
bBAQYRIDfFD6pY8pjRe8ttch2HzCcfyJKW18doSQk3xYS1Y2Mwzx5t8pxqaahzF2sG7uPkJ6yv2/
sKtEJStSU2SrMswVY9fPnemyfeL2Y/RawlqMMpc5Ov6qBPzfpxfKFtNRCUDKBHfYShtvkuRz0N/1
4ydZ2QxHbk5Bp0Uyj95NbqVQnc7nXebPgqP2/UslMIM3TgKdfdZyJUbkmPJyhS93Z2/OFdeap4jn
EW9SSkXfCqhiW4ozvVtnpr6wP1uKBVNi25Hb6BLIaczh8TMHrGhjGgX6ppdXpFNVoSyPnwnPZcXh
rHZeEtbiwmFRQnyIwtTGNEwekscdFkcthEQ0mvxaeemrj7Ndu0cWEjKwVTkN9YtHDBwm4pBbYoT5
Hf0vPSXn6cqqrF0dOrw+G4ixkUim0PuhUMXAEsCO2vhJbn5qDxs0Fwp1oboMpw6Lo/pfaXU/Hf0D
p+pCWKtQw3FhBnMIlVE31/iBno56osM6mdP9mUsyLeaHqoxkVNoPTDmK+I90ZaDU+tOzIeWGjCPd
rQ/pVGjOHfh6NnSJIw6rcaHoZs3h+wbhl9Y8/QL0R9Ve69w2Vu/KdXhWALBwOdReP6r6keerAqI+
lGeUuCNbeMXkM2KjEEXJCu17jUxtSDjKC767CegK9p0YoXO3cLZxsEftaXpMnKCK0W0xpC1uxNAC
oH30gGO0C5w428mVtcqU0mKNi9sAIUk0C+5fry7feyk/zwzS0Z5a3V5+MXKawJfXYepfLHOi/CTT
nA8ymGPS9bVa0ahgkSgC/qg0+eL+DcMy/OlWXf8ipdwYAFZX1Xf0cfG0MdbIY/83+tD7FfHCSd6E
TNSFixgxBKoI+lXt6gi7fHHleytdqiJxT8OyTwoGGStBEoVT+WfsMV1amUcv5Xn85cbKyA9fk5N4
ZejtsL5mJBerjcmNdbNGvx2jl3tZB24pgLaScwy2npcyCS0R3UreDfkjreseSdQKX+FSktmVYt1R
fcFC+fcD5TZs5jGraHSvC3o4XZ2TR4jvf6Ka01k9oL+3d/1R1flrt6Tc/PDmuupSh2unqlN3gp2j
F54h2Uq3O1TXhPVR5t7n6LcJC0g4SFa6QDi9TqvpO7Cjktosu/Bz+53upBXVQ41U7zHA5StB31Fs
RusBtSbybg6B7B6+PbiAclXakA6WZ8M7YPkRxJgHzx39icIsyQoBByX+VUxn/3IO3YScU2BxR4Uf
boqJUeBWYE27/ZX4O88E8Upg2rrYHZ+l36MtKR6M7iSK0oph0R1qyCqWnEN+QxOVqDej/c4lROIY
3WBuAodq/J2XGJBwqWlI/Y/Rcn9+X5GrjlesmuQr0+scui062OwwO1MRVwib9UJB77TeEG3NQe2p
8jLYbH2QqUwn0dMGK3OswB4kve1IrNbS2KBfrc741b9VYMUQScpIjz/v5QlLqQAeK9Sg3+se3Awb
qLmSEYNGDWKpp1E71EKkofUp7Wi180mWciGZ9y4WwShdKaRyqTfwEPEFuomdxwE8dKUWSE6SKmBD
jS429MjHkJVtmKmPD1y65ZEOxg2yi8YIQqVvvUdDrEvqxZQO/EklhiqBCFXnysOPCPYhuM47b94T
xbzSdeO9txDXai2HtW/SOMPbh2hEtAQMjv3935nV84xdA6pcgPRR1pUjHVdKf7JuNrI20HZtsNBb
l0s2P6lVAquj7O7JwTgOw6Zf9GSP625Yo2H5++Vhbf24FDOuNaLIMU90mah/3h+o4iibiMWSredv
f8SP2zuLJ9dk/egp+9ElmesdQr3yh07GDlMm9Y2+p5nAkIdRge34G0D9f263rm7d/Hmd2MKkq6Tu
3uqwIhHBiUL4HeDwh9/LPMOJi2cbzOAvrnyWx4hROcc9QfgvmYaFrj1P9/fihXDsmXJMxGClvxvX
0QvRibRxKy2Rw79qxUDW+BRjC952ZbQG7zJq9JhlZNyaMfBDVqXZGt3+RDsCmkZ16NcKiferMvPw
HyGyc3MI69LSLUyXhDm8N4jxiGEr4Pah71ddIY3j3AwaZJyjVsXtlqcxzGE1XPAqvTHuVWa7IM/U
SfZWNV/a4iz8z9uXGCs6lqCZEleG1Q+jtxpNapazuEnAmcSLCUjf7NveJIdRnOuqWb4H/OT0r69O
b5iWSXfsQ9wiNgoQ4JJ9tS/LA+J5rLDbTEXjnmRK7ISikEmeMGvweW3n5nuFSCayOJmgfbb8Ttdx
1HIzA1f+a3hmKnklWg9kXzoIjieMDrSq5JI6n4aKsjSnH6qfKXy8rW4mvZJM4NexR9tz/xMQe+wO
7dsGNPj5OhUXQUrwsut2WrN5CUqC2ZsthJee2bl7JleLPwSUDnychXTJEimgsfnYBZJ2VRFCcyPP
DMI03bYlP2SumajhDBj3zXdzxdEXamN3kAk48l/NgjtbSnctR7HZ9g6PUGu3mmEFAltFCdQwThaR
nPI3g+5t0qr4qy42ICHuc4JskJF2uSB29FhaWVkmYYAz5JdQDDeuzrpNbODnjFAoG7PN+t7bPfIi
UyY4Vgp4SRytMGKs82BWrXh1TN4JGNJuZtr+BQOQd/rARxr0tVD4AqF+2ZUK1woRApaFK6qUiXn4
AbohGM0Yi8MSnasIQUo7RWr77r2kWIPwY43/W7TQe6Ozoj8HMNljapVXyb5rJl5/8VHsaQutcucU
hJ4hhBKO3Kit47CxXtyWDjy53PpzFln03TMJ4jkRPSOEc1e2atyQrBLthv0Tzyubag6drCaY5vKV
3Dd3sONMxUyp3lYs1AlRtUngBOh+PNScCRE8YNAmWziCNCNn/bvd8vyrqdsLAJJNzTZxjIcsXOiY
RhwdvvQaJ6LQg4xz2K4n2op/TjE9j7O9kHcDWUySQGSUpYQqDS0gw2r5Lv6bgFQOJ+FrQDbxd+/G
STyLX1joc3H7RHws6mctqpHBMvSmZdz83Pgtw9LSEwPxGBa/9RUThioM/GD0fYV6tb39KsSEwInw
Xh71XypbZXIN4wWjOUwuEB3v2mmhl6DvQy6w5QucWeS7kvD/ZmIMtTF8s33rrjLnJ2XR3pM40+yh
86YfkpN2DzY+OhZsbBoDXL6q8YipYosQrQxAZasuIWHQ8M4rra8UCrLc83qO7uQ0O59akhpgdzxe
bJ8Gb6ZSGTCxXFYAFy3imvfBmcdFSwxEdhHzJ04MROasnUS7QlYwah/y4LZ+gE2lgUwGlSJCS20x
ei97Er96NCUz5suy26xmvM/Ot/ZEX3UVtFDsgdVa4LjtxQLJJM2eLWmAkaYkNsrYXLRG+CQ+zNu9
bIlwUPsPGahCpXmF62OHXogKhY4uEVEuhZaJS7eGczSM/Wgs3eUktuKg1JC2xK9BA6OfyFYtNBQt
0Bxq+qCPo5/o+FCNOV1G34NiESdjFz9u+d25S+OqeoyTrJ+Jh2YxMBkREXrwcmnBwYEmaEdIH/5h
1MeOrPPVlaG3bcerLEMTHm39Ch4xliUszGzoeiGVAt8vpn8+hlfnTTWbJ3UVYQwxfarNOTTS9mWO
Ukm0CKzbhg4MIQ5UG6mLj+ly+StT1PsMJG+iWxBqDbkPwVpwiP1ld0FbSlqFEpHXU7J1Hg3tUMNl
AWaad0sFfuuyQBxRPooPBOLOy8EM/QGkMe+wsdc32hA/Nqi7F1Jzjgo78tBEwkxKPG9dIDjG6pt/
CoKzu5cO6RytlybnuYYAbYJy2PHa/UtrD9HfqetPQwIF8z+U2dzJG5CLJQYYqqwfJZESyGF6L4Io
6QWSmYMdyEy63yw86xysS/HdMej5z+8p3Z6rPR5cxdhGF9JvTSXyh+qHjkJbbsj4tUvbn3MFVB3l
uiV7XUep3fyhydBl8M/XHJCElbaEopSoq+6wyzh5nEQHc5wAUBaoPLXGo9d/w1Uh93bzwKGLZ9Va
+oCpRch7Ctsmw638iQskVal3uNqPQJswKkOHtn4yZ0UI9vBLFK8p0hLlhQgMCcRwB53jdjP5EYpS
Q8sjYWSDYDoAEqnUW2I5GmoCLgg7TKPyLiSJactZ8vqQml0UadHtz1vzWME7MlskYshHoMc1KY+t
4PMkxpFVE7JStCG+T/nI7Li/qBg37pKWGmxr7jciH2XVW0ozTQuC/+VoM51sT9YBUb1zMAwTPLhQ
7oZ2n6ipbxBC1OXIi4KIMHzdf24wls9kvsOFYBX4FxAnEcpOoQAMH5Pi6LZ6jc2nQPNz1aCQLohq
JCXmVnveXfSPVHnuc+AkcKCAh5p9sc1ecpgMatrPvnmqI8FLqeFRQXdA8ZuSMcn8TbmKDl/eAotj
gIKwUHBz224wJd1slxpGurHNLtRCUiv6B3V3YjBZ+2VxVhmlfV7XkEocFtiKn2E603GTafi9KBNT
SKyccGyCDdf7AovVhhSzKXmJygxpGh0hcns1CWnGoca2QiXEyOFD2NJQzSkIWXsmcTcCS4m+bZCm
Ub8u1jF9c//Y41uBJFgyH726Gz3ai6mhH/5OQdXoHHL8xgt40E09JSPJhaktnO1hzu7kh/mWIrd3
9IHvj477xjFaokiSeaDTMcvy3iHyRSxmE3+dEJwZAhRQ73UxPr8OFnj4Q+IVrKNf1AI7t3Zm2ZI4
ba/F99p7UsvhybskuubLtPo19CxxGKQ2ZF2F4e/Ld3Q3cv1bW6tlYL3qFcZmQr1CwI+idQ9jXFUl
onN1a8w/ZsRzHqZZVMJYSKBWaXPEaxWTBQZUlCtnqugcWSL4mOinI3h8zTBcng09pdVJv/jWvGFP
up0yOIND/ydqN8OzYUPFIitSE1s6gP7mrxzslItXtRvyrlhecmohcL2rokP9MouzJ7wGMwIeVeW4
pv6ydJthMFMiOumzS99DUO0etTcjYn/n5Z9IPkmPAEsFXH6SL8ruLs92xSFs3vHDWHRSlsozfJ53
Z4dlpJP7lGfYFt620tC7xj5pQgBAArxpLZGsHqvabflVFUGgSbn5kdQEHhfYiuFU43LhwrkJm+ts
oD7jx6I4vH18w32sKEBULJVT2tsX3lkvvJexRc5nqvcBg5l1lmlTlVu3LbcO7aEZUzEmWNrDx/0K
HFuir1ndQUhKbYyNZoDUXE86AzcFhrFt6qVzg+rcKxFDW6ceIJkZBdkMKDhyrn+EALStWmWwhJt8
TZYUmBg1e7A+W2Wge5HkJPjt+18opmwko2rZXzD4Ybehs9Nnaywvw1xrFyWbEcJulkj5movSs8a6
Zqr0ZDd3VP17JLAmz4VA0KaMxFvTyN5HKkinCe5/MV73td1xeIym63QHRr0auA0QyTT+9YDVQ2qC
Vxie9mKh9fCmHQ0fQTVx4mBAK6WA2Tv/QVifSF8AghekP2zMSfoIfxi6Z1cjl0BuF6mCOw42ENm6
llwm5PO1kNcL5WwCiE+aInShuCrVtqsPTMzAJ17EezbmfDWzopJrHbK8jK6P4zX5C67A396tG1ws
Y/twyc6AisonISKiY/zqQrOqQuseUEyvF56kqmgujzzrOyICrEzPNzSahRNloFnJ5iX/Bk/UiEfj
tTLbqeF6jSJJhjFxs679UsHJD/VHD/IYSEpduLkXDzEyDtKNjtTfOOB4dDYKdmHi4RKC+YoZtUsW
L2lABLsHR1lMkFLPaj32tmnNi6ABseOTEKtHBaCy00Hi0PIWKrmVLvV1fb8/as6MYGIcd2EqZOQE
mVek8GammgaJhgy6ZiiL77WAV6dooWSCROtP0Pm1RxpmWK9CGBOE1mOXc/B47grQqn7Kl0fweRK/
f4WU7oo5uMphmVBfMhBn5SPoZwY+vS/MYqNXhg3KJAhKCLh0WFV5wcFadJ7ClNXaarSCVmDruhBZ
J3Cj1PRxEjhcM7/SToELmm06Sfg3CEQY+kSy73+Hr8ED3T3/rLIxWZqYyH3Biu09N0OQ0UZ9AEGA
Dh8mvO0VglPjzNSNnEZKEsCcnFCF/M4ivfLWWkEwExOsheTuUz5/+99Oe0nmVkZOlYptOrfaHAu7
CSuWVqHRxsICTrFhL2h3kibkmWOadPo3WDASWiCWeuvf68pLMoeN5Qbq11+wxmSVpSZVAMVrWqqc
16FO3vFLrDiu9FfwA/2e+jdUUGkcl8RyzJlOPYWvGKBclhE26z805zFaJpX9nKjTqqBbLApGSATY
Cs/O4JADaV2Qklu5tTI4X2OxWcxAYollMvm/IxsKGmKRfsmCO9/ACi7+JPUUfrQCDobSDKRDIiol
dEDo2rYR3yLDOpLO/3OmNthUrBlP6A1hLmt9ECk4cvvsYrxSm3s4yKryNnzMZPKF0Vwu9caevyPi
WZG258wb7/tdLID9T7FE83MrJN8FlXCgFBvFDuT5BJlPIPoE8+DVY8DXIi67gTfwz2Fiz6rQ2f3N
nuZGVWT6p9aER6VNDc8cLW7Ifi/mT093TlLVYDLfgCcR9pApx0mwtlIsiusBHO5kDmiky+DMkQ1w
xRLyeuC3n2sA2TYHjOYJ6xddOYkSu3ecXfdDEIm3cQqVALmkphuPQcX6MBlXL4vWOVM9xO4k1kVu
wLnkv5XJN8cbEM/09f/K781LjmtAe0Crnrly9G2FT8w1HdW02yRJiZvlA1ca3d9+oDiVUid2H7RI
p3orBF3lbls7Q7UAEYd7Tb5LzBJDSKuA7EWqTEboOmecysml1VB4NFXmaLWj//MpxQW61K8plc3g
KwODEM+7qg7mEwK36XQ/dUd6i8lElN13I0xeIRyMTrDp3xTbhE7cVtEuwF7Dx7IaVd7vIfgvld/Q
bnTCW/8OICAPQzAIX1VXJTWMeYx+PIUBVMtxaWnFX7clpNmvA7N8Lmlo9bgK9ghUhFXyFtZ/AjnC
xTtYZZF/e3KBnYCIcqqDT03DaZsq/hwCWcE6vDdpJWtigK9UbcU9ZpE6apsppYn8mDyADPtHtZtT
H5iiS50OZYjLKT4vdwgeiLDDAapkEsmBEpnOH2n5OzrX5RAYQaHfPNvbbW6JRowX66z3ztebVaaO
whuiqBBvq5SyNnuv1F/n7fKGkZCtJ/vUzRUotminEPRpaOg8dB6RaI7z0IW92tKAYVq201C18f2S
8HcGhmBfMb3wiXHpWvC9+VCNoDH2ljqDNqjWopF7BCm1hsskC4sk+0O94ewWjuLcS8AXs81I9tbz
ZKxhcwG0eb3xPPI2I5T0X3yeKpj8fBrZz8Nyj5MjI8vm3lNYy4OY6/kw6Fi74FyGR/N2qYuCpURW
a9XTNKuPQlTyGmZzfI7VSDpx31kRtfcbWs9ZbrJJ4tUusuwef1oii0R7JLZC58o3t/xHGd/UGE7f
kpwmU/pkgwzmf/fwBzXtQSlJx+TN3THsTZFMDaWfgUmBvLFuQlr+byFsni5E2f+d9BPo0kDYkFZL
xvVmbr2WbSqHaG/2FLv9JVH/0ZqA8P/wIuUXpDcH4dZlRAYUQQmEjWQetJPCI3pUccIHjI1+9P4q
phPn0an47bHqhw65XvtWcBAMxn9yKchBkjjwyjvzypT/H7Wy8KXVMV0mWI39RskRMbStGMMkCOe4
n+nqzJjkHcw2jMSpY/V4pl2Ad4sb9Hu9L81nMPsWMjhpCc9n6rz4j5LbExc2c7sJlmQ0lXwRGQw/
XvDSNHKm9IRADHX/6QQaGhXJ8/sPI5QoVfsFeziHUMuSdQJ8vNJP0zn1J940ZmHnLO9e9sM0k3bi
Yc0/5uQ5Ihs2RT/WSd3zX31Pj8iFESET3+DdM+TjQhounXNN7Eq6G06qRp8b47q7xrkexkkLC6W0
NhwWbdMRtBVct+bcn0cn444thjnax/bat9eebz7enkY74JQ67YR7gIYMPCtmqdrA1CCgVNzea+4P
mBpYAyysQx31dna13coNfQcHYoY8l5f1JlzJxBou//Gi6g0RaZ2AEyv7gIwKXfDZ8PZjJ7Zkh31T
ArnR732SRqFcKuniDywXdb2FyPS0o/EE0B4GPkePyXKDehViwTNt7DKDTXXknE0NcJAjGkGlDLfM
rIPMfbjnLYXKvDE1dzdlrEnjaHj6t7/6FblL6HlrxvFNrqV9L01rD5vSmk/Ou32/wDyNbYfq0S7L
+7xvCBfsVyrDqqYgCYzxh4mV3e5guAskvOhRPF/hOqFZuiFbkzIZL9SadPCiK31BCNzJMd/XIoJ9
xNQQyYhTrHwg+9E6OZZlEzAnJAKMmnxZ8VrE8L03Iricj+TZ6R8p8GCTPHwwn/26B9Cq1R1934Qf
m9U0yFcLaI/T/RtqBzJlIREH6okCxzCoY+13noyQsZepnos7E34KsN/dtkv7E5EdqwQd9cU5J236
S1TwpV6kALEaDKNGTUp/nhmVDCjb1arwiViGQ2qeq5vbl8trHHYzk3v0n1GznezrnuV7dndaB8C9
HVWoUqq2sVtmIL6F0QDdGhyN2e0cpbFbsibnb5zy1dLRQnrmJn8YhoaSonUJ+yqc2CA3M8oBNfER
Pu92Qu4vkPHR7+cKzD0evlaV7XKmrM0QK6U6IlBn9vatjZupLvAzWrmSMxhec7+hGJpZ6lg3z5cM
m5zwAHy5jBFv5yrcRIMGbPpQhIEBceShDsxPpXbdcWOyUjQmMp3/brfVG7TNQNwRLToVYbeNC8NL
R76dCCBOrQKlR4AKr2Vt60iFWBoh3sXVC4Lz9r/g8iPJyfMyPNlSnhyq/mGpwBB8pRuLlKZ1/gOB
8ppp4yCSUe2mv/kW4jVcfoOYGF9fYz+1cujAt5POpAH7eFAc3lZsbdgQ3BXbA9WXFWlABjogiINr
JSgv0iO2LXxjnGWFk3pPH5ira2Sw8obN3ZNYtpPXYRaVknAFVoKoF5bmpqNcso39aG89G6M8tSc1
+OrSMbVzzLK6JmGQFKFSUaxsamezPsxCEUXjiP5cGBnlVqz3yxOsHUY2iFz2jnrquLORwa/nVWtu
DJmqeOefQzr0nw8cbvlDTyvdod6TfxHV//4SHulYIInR3+rfEzSyEZ0ZtlD6cJnyBkyQajJOK/D4
N05dUEMUX3XnWqmXj9QDfhIr67frKaV2iPIyXR5St+PLT5wTRfemXqZp1KLqdOVuxDm5/w7bBOLh
rwys2p32DB8S7ClJutkR0FsB2ghK14YLjGlEWcV0IW+mN9Q9AXR1k1P9J2hPTs1d3qbomxmR11v7
3FcBNXjpzLpnksb2WCKoooP8vP9IYEsLrHTJsMEFpWg93AC4UY5x7iR1jGboPcsAUpDEttgT6lna
iIDa8bMlbYeCPcSI/O6Igt0GUDdhISx6sth3xFVaUT4l2VL3SEPhrQnKjLNziibNLmZGIU/wBYs+
j+rG55InetiiktHGlBTTUgRhZeHDBfdqaAv9HoW9i6zr/mJ8gGoEIh8iY9myCRqkIWokVCLLZsdd
wgN+Mqqxl4hQur2Q0Xw7RrBi5d2PyEw5qWlPf/Mh4JVqz4MDBDMq/uQ7uqUPugmFaNeXh8/LVxHk
BVfvypR1F9pFtfQrGeSwli1+4k5tw9vCozUt8mXuDYIr9W4eJaH+mK0weA0v9xZE7S/wJmsnFSUa
qAq72N/eEsT00iyS+3ZL12aj2WRrjjDpr57MYnx4R6/nCOgph21f/HExzho05Ijj521BfgW3uzrg
vBmQPMWOddAvaDXNSRTnMpfHvOZbpXgeZmuoev3Xl+VY4a8nAYquGSCGo3iLY20qK4R5kLnYQb3I
2e2J1wnf2ZoL81lLokETtK6/4losTFc2LfDBmRNSoNupHuET1uzDRgSh2/WU5EuSP1adASAI/BcF
uMaxdj0zLkTMw5oH1rxlkh+eu9w7IMv+hMLYRM/hKP5G5bGbrpnSXaohXj1nJ5iwav/kT3Ro3Z5k
ggQbSDAEeVarg7td6L1ZNVPO+5xlPlMgxVU=
`pragma protect end_protected
