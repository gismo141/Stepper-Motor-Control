// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:49 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JOvKbgrgAxWSMtp/wOhM1Uo51Wxvk6Ou89LWNXH4YBpTgeeALVlZvus3WM+yzA+n
9ZlUwsuJxvGnbMn35/mciWqMlvsUQpCKJdVaC32GYbJhWIDEueH8vLdtKdj/M0Sn
cu+uDeMFd9OgxZ8BcFuH2OTgkU67Z9icuvROsG7wO3w=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21552)
LfaaPAHeBw4zhbI6P1lZf+vwgIiiv40qK7c09M4cEcObOWbbtGZZ/QhGx+Dmj1R5
Aki9TAOwzJDthXBhWGZoGCzvsktJbjizJDuNx8qbPZGT8ewmDNRLCwN/7TCFIW9O
Z3RGHaVAXOmq7xiVbaodjuB4G0jwqteP4NPzntIFlPZdh9B1K44GOaEv3ADvkHIW
7Yk5FR5VfPC3Gqka8loZd1rShP4bMm8xZF7QQxgR3u29avCTsWN5CLbBpT7Qf5yr
rjkAVSTxWEaJ7PppZRvxcIQrdgsgqCCJkBzmRS9deXfPi+ZuxL9eBUM4GoK21nSc
8Jjo6/MQatA/h/iSunqs/ALP0lUzxEpZ1rZemSlxwqGY9Da7trBeYODsxY7ODYki
2Je4v2cgteDh0MmJw1Du3XKOlmzhTR4enque35J0d2w2FnhzNeI89CJZ5/fAhA4w
8XpKMmhivfrvjUkkxlHDY2iryzC5rEufIki+1kjbTBYz60VQO9kEUZzwfUX3qGj1
nRiGVBByOBNbxes3LIKBqmcttnDtOAItCHzwBTEVDz/JQiUG8UbmK2RL8T4F8nHC
nZVIAGoPm8tNJKzDqwNXj4D4FZfWDGerlnvca+uqnzTv+vSHTyEoQ9vd+kT0Hw0H
ByyNKzO+f0jNlwZPQzLDFeiXwMzFj4dUw3ItI7vPzLLRJSMxwitM0GbtC5tHQMtX
vY3Wk8BoGZGOEZebYhyBofXwZ89yzLwaZ5RiexaKeIqu452RZZiOUHWZVRE+PNv2
ZGMCkFwhZvcRbc3VlqSP3SZCR0bR27sWy2OFXsA+xIKSLBD9ZeT6f2v+nGc97uHp
LLz2JjOCC6MsqwnFPP15wdgnOlyTBKv/cwKm+Sw8rQ28lSfbLhAUDCkFO/35JYIN
ivPIMZEb+EAhtaEpVOlpFZamYWyHvpnsWMt11H5UqEvO0AaGxHLyi6+b/YU/w09v
Za6DJ5NqScnQ9AeQo10BDXnPFnZu2Ob9Sa8ZYLO4mQ6Jf+HBF/L5OTmzi/q0TLJs
P6Msf+C7ugoEzws1IozusaST8q4tlbOL1ni2ml5VE22ppKShQsy7QS8/Q4+H1sOq
GEXd9yrz9lEtTxFcEgi04aOZ9gCDVWiYxKWaZryrPJYo9ABFjfIyVYmWOL5R4j2L
h4dnGS/ubqZUS8vmwtHvf/KqmVGLNw/hvjGj4ER85P7c6hwIc2YcTt3f1GqkTZMV
2mQmxZokxcPARYNh24EqA6OXQvWObzIIW+wHMl1lxfcdD05fCabOpl7EqJukGbDc
5wg2NX89Qf2/NRnACjwUF20VlqP1efUfnoMjF0WrrtxBGX58VA8SxLKl6wWBFi1J
VGyfh+/UHij5/ev5GXZiJ6+18wRvWGpANucMRLKjXrw4xyXOpvdQ5n7TS15m59hL
gW+V7wY5tcDUH3wKMR4uMNE5kfFaQRe1NNZp2pQa9hLlquN0jrkEm+4NseTx2Vrh
dkH5MfYMyjneJyU+zu4eMhQ/M5dTntB8oB54yHfnH6zykJHxzaZm4VWiyE8DMGXV
9zND9In8zpxfl1hnWVASsUlQ0gWbi4DsNg2p0SIarCa2zFfxsrNv+cExbDp5K9aq
h+Zmm5qPUBVBPedUm5WV7Ll8mazcSo4MyU4c8LBpV51pDkTsfCq4fg6sYMw4BPm+
5RvZ6WEF4QSwVas+3808l7lHQ3PDyNfjCCR4kbqsFGaHMleNqmcpr4U4yy/WU7X3
fv7+ELVK293kvuUJnmcd6ZzuA6IIxlCZ0w3jhP2dGhertK/iJf1y1Mokd5ZnKO1S
WQ1tVgq0D5NeVj32PYuAe2IZxJWmWKsefqH7ZQHcnzaNNjpw0blj+T38MEH68/XK
0GfJszeWeiJj1mTXJD34UHi5wuNAHv/QLSIuOGdsbA9aVjWKNbfDGqsQdPQdDf2S
ArYmjqc5x0SOG3e+L8pqVxI20CK1LAVMAeHvWzgTOjr3hAfg2NB8WaNrrfI6qbu4
XBYu/PL0hKcEfVVh/KeHpH2AwykV/ApqpBdo1wAeCI6jaEjMeHccCi8Lb4ZuFor/
yNJWfOwg/QoofKbxTDS/ZNmTFcm3AxpzlXCUCgNhy6oqr97xRXLTz5dJYDNms8HD
JBSi5AvoQycYQiaWLHAs996N5/ub0FoWM3UUbNlDkG/3yWaszWt75MyZ5tevbndF
qqn+ZvJSejTZDjIsuxpGL5nV9MTuLbbdx0Zq56dx3/makgUnc20tS+bGYwKSfQdM
w1dyRZChN7soIQyFmSpGgIG5Q7lOnVJWzooM9ftqpP+Ydna2d8gkHBN86fMDN9Ww
f0CDrVIbfypzBrReyFHTIK0TjEspeB6cqXcfFpv9bWBv5GbsnDASntuWGemtM6M4
zcUP8/Z4o4SFW7nGqkqwy/oF7dp8uvbphvHj6NOPbcvaLoxaN3ebY/rC/c/3AHhJ
R7H7ybCQbl4N50pNs4HvaAyL8q66i2GG5lJ8H5n7lyBI0E6su1pGrT9M7lTNTJQM
1r13+SUPFcYv6EUd6uOzdPZuXK9YmaFI8xFLkwoyJZRcp41dk1fht1ea3iVAdHd+
9hwr8LbIUlsfuwZh6GIZScxNDZwhOPPXSEm4Gg7/ShtJBjyP3w3wfd7/NwcMHy2G
piRqlghFRsfi9H6PIBHjRPH47hPNzNb1wH4NW2Zl5/aKgG9MRPFhW1kHA81vk0fr
8l6vJZJTRoJKIxv9q1j3SU9MBq47BEYJKTaKr8cRTzs+v0HCurCyD9opYjPubgaS
ykI8SbXq0JjlKSvtjWT6A7yKadJEzRjXE5lyuODbI4Ob1V+wuw6Cxz5jW7Q1sRkD
DiIKz3BZ51qqgb6bdNUj2IQ3JVrtBqjheUeakMdyi4wveQASrhWwosHi5uRfBGlI
o8aYUga92y4uDSSSUJ004KhBLUJACnO3E2Ho7cffhjno883LVJBiX0u2vPCpbuSO
v8GOzO+jRB996kKAktV5jDHtzr9saRLzpisAnAlqPXa98Jph6kTjrT1qs2KxLTdk
/7S99sOCVpNUBEtpJYYPIT2LJWnO9Yq7w409rGtX6cd4O2J+5FHVgAJnuYTZq9rH
grn0r6ueou92X10TlVhtBGqJjPpzqTCCcTVrqz5VqmJcGQVebuNsV/UmbqIeEijF
ZqFJitzX4t4FO+SHydFFXMPN5l2cHpwi7J2276Xpxb1CP2jn0mDaFtP9GSWTWKNH
6FOmLe17593HoElMncbsOQ/FcbCXjz+W0uWZwEDu2uP1A4A2Brhvf825qKCWBVB0
eIx0GGfXL4wTBtbi+nEnFWq2TcDAHG6FJ1FUsVb2+37BRPiO9eS/gjig1z/tGJ91
aBPGp6JgszC9XU+YTUy5ruSo7cje2rBlEvF9rsMqhvxzUV6lBRsICANPLYqG3ouf
mEuhwm1dFPEBpOdqa1cTBY08X/yoRpW71XMdRkSXq57vkqV1F8lv/RD46M27Tscu
mkUWRhr71Tq/DbeapqVcBoY37eZlP6VCE0dnHs853HpdsXMungIXlfbEH4T5H0Vv
Y010wNimfp56RaL/i61ktRXEV+reQsKx1FwV8CBksgPX3sy6bO5/NwtIDxt5njul
6ppYc4d8cMqLx+XELgsaZi2UCsiZY+yoxX/uxv/MMBuIfq10hJA1s4ACHFWUZtqK
VAwWpIkTFIVz63P0zMdcuU1Gi1m1y+kd5HEZ7isrQ49gUzJ572rPaYqHhiRaUeUT
/N0jeQkCJhQX3f+5ENW1ukptqOKnWErxT5i/zC/kAcgXbp4B/Eo9XRJ2A7OpdOOP
d2puw2whcOU4V136feXLGsgYbT02JMaaXKUNakODS4GT2fDHxQSi7rJKsax+rPwO
9lXKeuFXnPdQ+FIu4td865IxMxqFDQpgVEM3P2eamkZ+d7YZdnspRST9/dGx6aPL
pL5B16PpsuLyq5ZReLeGcZ6hrDKp8Eed4SwN6UfC8IFQJyMlWVsfkKeBZQdBpigV
RO0qADgvsgT66o78qfjNNshOY+4t3k5zhBB+HModKgqm3lhhCeBKjvBOPNgi5H7o
1K09yxR68KcXf6/VDzblN3RApLzGdNUoTjvukhDxfolGbhi7E6Ge43Z8mQDrEYxR
et8fU12FWuoyXTNgp//H9gZ8D9smnx1l1U8qSMTw6RJrhqhfM/Wxnm8kR1ZnUA5D
C2Fg+cKCH73lM2SvjCdkn4o5sHdMkhNclKPxhOQwxrHejidnm3HsuyUs4MBdAZaI
AzVe+C9qrEpTpZzMSuxHiYAyZIMsn3atN57qf6Rx3JKFNvnt6mhyIEf6YI74IJPc
PtTe2YT+BaIq463MiBGUstdPHO+IeN2GQK28y59sIzsylnELPzG/vsGD8yM8/Zhk
oXWGQLMXs7QbevcTkUIFP38hQU4Y/bupRecUurADUdROhSoY+nFgreZBbnrJf0L6
PNIguBdx3LF7e9ahziUTS9YUI9iJs+MvzJqGuG1FrumN5jQYFH+ag2EBx6xs5ft9
cU1qG8ByoWwo+h65oR790XrZHZZQuf9gUCF+nP9uEbz36AvwuwZGfB4GMcHv7SJF
JDqREEfNniHGqvSCvGB6myMlSO6MQgwASJIgD9c1AqGLd4ylPzpKntEXQ9qcJDSI
5xuNM90qvOSd9QUBZj2zLc5NUPTQ34be73HJJe7Nd0Vkc48oE1FcBj1DqNvI2RaE
i/HVSWTFConVJ9e1rVolPXFGx+nKoovPFDFvwTpaXBq2y6WTLsaOMWgXxmJcJg++
iqAs3e3rvyTADIXDUqmUsGmK2lX82w/49GYEufygFeATObNEsfjLuoLi25dOug5w
D0xzPsJB7eFtmvH0xW3Yf1o8hFYUBpsgNbGhEticxJJM1HWKTNo+UawPkEgDVVkA
mKf3FaQDOWiptckTDLJhiMdUclI/Tb5VQNVkWuTENEksEgwC0EFeZRrxstx9mgDJ
rRoWYkChjNezDlfUBXzNsiI/BEbZtuqcbEuzIa/LRr/5zoxZx451DSxjNjKpjobJ
6PBRWLLrJ7UcTgLXAaa89uJOF0D+wvksHkmsvr9naGWjdyxqlyz6nte/s7L3zu2m
TqESsQyTmDTSe/p+J6RotQpQQypocMZIYk9o+4Mn9O0aBuCokJRkElLijDkqV349
qCWvaOnbOy9KjVzNDoer/2mwwzVMiZNt8wJ3LVtw889GitJl0RIYrnzYyFbd8sVF
mXMmLu9jOW/xSLp8vWTiNa6f0JoPfU7KurCh6m1bMms+g4dD1fUnLijQmmx4xxZs
m9rqCFiF+iJjVa0+tvEk4McpnSTck0nnf1gOMqMrX6OjwQfCMBXwbhjEiH26m34J
NuTuQ2d0nXfVL7BG3ep/9vo0N41OdFtwzHegC6BAs04atrZvZ1z85afP5tjWyLa2
xkYAWKTqi8pS9/AFUZlSgEjhdONzsS907lQvvqL4tTMGnVuWhr9x0s9/0A646dTj
VRvxuOT9zNYesjegd9F3w1767Bbu9nKYjJGZ/xKJqhdhCNeUtXf80uJz9Ln6o2h+
9zE9RmD5bV/4Mb8ZiiwTI8jCbxkPX7BKlXPeRa+oNajuMUuwOdYKfCYWl8TFzfcE
cJO3QdFqZcct+WoU6b6yeVL2w1i2GSstcWgkgNj6ieZEM6ydtxu44m59jin4COwl
JqzCh6JSZG1vWEMJoVkC033MBqX5n/bCo4u8fgvWDxVP8gIwuwocLQdYJhtdJPgb
uwO/EdRO7hq97p3bsGcseIrcHm4rzlueE+DHyu79dzgspXalupVXkZI5v+HdPjPw
cLcsLWRznhq8BiFqCv3AZMsIHJQncznO3xJLWPGYUvpyndGn5jB5Q5rR0J8K5stj
675kAICDj5W0qVZYYzSIOsAlP0zz95kWnieTp3AjJ/USp0JDudjOu1WDGINIuL9z
0f2GNP9hpHZ3JY7mcNeKkwg02bc67IlfH8Jv/pbKuZptCN9dxUjO7bNZUw+G+I8y
6Dz0OWXspkUmWdCeIhW2b4WfYgsw/CbFQKs48JB14laHRu84t3sNW14tnEmMVfSK
TN62qZGETQR981EOH08LXCDF/A1E33xjbyGpVo9/nZg+OIhCWzNGxIAXouM3rgw4
UauswStG3h7AweIjxv7Hb7z6hGdaK7gmuIxNBhd0RT7E1TBjIgPoxybsBCsp8Jc6
x0dnJ+0ykCqo7rpfQnW3mlL9ZGzwGvvXDEDMyUMAUN759o5MOOjbTiQkwdxqmtNP
KGo7hBW/TrewieOKSiWNqUCAvomKj5jkimwPV0iPIhPMFtfpr4te2vyvtQ48EUNZ
tWHnW9pa6OsDl11YDfRvqkgOTKRJSzupAZBY5eCUaS92RqU6gllWZie/ZIzn2LYD
ukgI/im263uTeWCRUo/ISo7lrlbPRDc+pTUNRfW3UTQLe37XYqUowZrMPxff7Jdr
Fp1Jx1pS9Z0ydl3dm4MeJaqAHUpaYmCM5UvycvwjgKZtrIZ93UXUzISDBFEMJfIQ
/MlTh4RtR4tlKNDs5KLBLMhAUe3euZ7DRtl/PQPSTqkVCS/JpBQ7j8o+TSDdUPx/
re2dW40QNuwlw2D96djGZwHySwDPi/o0SxrYIEd5wbRpgGMP9KSVztNNz0zWOpFD
0l37p7w13LB0Mlh9unfZgY7yXOqsKupio1H5a8rMIb6bdFLBgs422mLM54iFMw2B
W225lw86kmakWldj0U1RwmxGUpaDMvdvzAdig9s4by2AjKT4rhagHEzfGsl7/4CG
P2B2CSspP5hhOlQDustlUV7qx2iemrZMgg+I/q4vWh2ZeVj8DU7bh23TcQrxdm+g
NDO0GmUxXNGpDLlYAtBXNCPBMn2/GDEiNwu+X8Gjn4sjTACifUkx73TdqY8Xggbn
JirgAa0KuZ4K7FAHbiiPbiPvDlQRnSKBUpmjEbXEa0qNSWfQGJj4Sxg28LZEriuV
AJirLLlkYdMlPmJOvuFSOQWumaspULSAkAQjyevJXVnLsSdog6h0qdUtHXNU6jys
8rv0my0YW/0eGNsx35laEqjca+RWU0WmGwmWNBsWhrGFYrX04ehpSs0xMDkEF+cq
3h8zw2kzV6UMXJ+plc3VFtb4Umk25LTlZoMvUK/JNyeZLJfnyQT+MsPz9UtWwfjK
j698lO8G00SGa3lAUaPmA4q3vF91A4RFnduvrolnD2UZ9V9zRxPdS5D7jOY43c1g
HN9lyMZ/iTFvKJ3pmuXp10SaJ3OpT3Kc6bBQrhBAarAU0wBL/LI/v3zdLSLOfaHx
j6MjcSK3HVUEqBEWohCc9DiP2ZJae9tk+mUpWgafGi+AQjFADJ8+sNNwlL8xW6wj
w2dyawPy8cxQL6JCCwkjDPROM/BYmiUJDNwxZvb/qXuFOoiZiEOBVYtGbUB3sJ6f
8zV0631Fa10F0jMZsS/CU1w7/0UxiKJGBja2oV5IBfnGa7mQMdrBN+So6OlnhWIJ
ZgoiJuVZOiJfduunr2auR5IYN37cJsHXGJBr8cNYIJuFOhlCYUQzmT9OkuWdYg5i
oXyUk0+5bCQmf3KNdLGsySKtp+SMwp9EjPrx8tLa+nnHL1D+f9adAWJLMlnC9QGM
dqxNO6QnPnzAh0KOwrjJ0XMi6qpi56KuHsKGAUnNZ+w2VIjBXrMWalWNMRI7D6C4
PSAaUqNZMP4DQCgeBeukjuWXFEECp+Y0FZAw/VF3EJalDDD62k0UOgMpbtUZvgnI
e9aSO9pXpqoPPx0Hiqcc6XuUikL3KUBUqyi7C76G/s2PuDqUy6768BdqLxeHzIXl
E4Q54zSgblYTP+FeOl40ygk8IYJWtWMWG5aGQODzVXn90z5y1YSPyPW3r1qGxSK+
J2uoHpXGgleeWgMt7l2vr3k/ME1AQmKg+4v9YbHDHeSuPeKpEi5jXzc1ijQWLFuP
USmi+kvUBb+aRjw/C+J0ghWvrDIeq9ASzM8EHMPXqp2drH7U4CxsmBFrwmF+qp0m
7LGhMgN597D7maQdZkh0w54tNSn3WBZkna5XLodQM3H1ckc9LrZrBcSsKlvQai9Q
JEA0Dji9gmV7lkFDJrnB8t+6/5SWtQu+EDzXTAtqJ0syC2QuJ0mvc3DM1jwr7MGz
SW1iMybAxzQEIOoSbEv4/FQhFvhXoeFKhgUcv1f10C56GETan3Ig+0BIYzJ071k5
zs6cSWsVn+2KY71RfsMFeLK9UtlAS5S3LPU7bbxe68SRURwisaY82qa6DmmxoyK7
SjR9I6w5i/vTGG09wgisY6ej7KohDF/qza2HkyHe5JO2BCua82o0Gi8k0DVoTxaz
fqOa4/MdwjqvGtnwLAnSwZP6Yible+Z3TNJ49UpRWoLhQuoxX1RJCdnXYRuw/qVu
TMZew5etyv7XaiJSVgbWTzheMWN+RGT4Y9JarKShONST4J3i8rCzk8Pg1GNkoDoO
CcJEDnWg+4iureIlT9JXajLp2stDQ7Ovl9h2oxv9jUDhM2cAWOY2K+9BoC1YKmDe
COxg+oG/j9Gbd26+E2DCFhrFpa4FAa0E9c4G7QRmS2AC9i2CB1nvN2ZAa9JbKA26
3alN/eBgSwPLwLLP75CJPaFcP9azj+bm+tF+gyIAqggmNmnsnhwcDNBcZImTwjld
2I6K88qREuTFpmcqlguieowTAWrVMsjsbON+sFWkZMoJAEIdqPfd+zjVDCmiaUSz
H9AAWfBfYa8V8fDycVWQPHFuLOS1Bubna/jJgqUGyROuuzZwTnP6l9y6So8fsUVL
L2XCbRuaIQwOVxVTL7Y8XjRgM1jngBX6DFsoMhLTm61iGZqY8kF8pKjh1rdYiphD
px2H3OwitSNppaQiEe2SMvZxyh75gKzfSqJ8yUjTn9ulws5efHZg+RnUxqux9tHh
U7VV98tuk8yAVt6/zljPJPZR+5gC3jUz/XfajMewOnWUgrKkfsNHgFhMNM9BN1aO
wd7qN1fhJ1tqEAKzAgPcyS44lddqRxg28SpTNI+15UQ1YRAhvEhVytJUQdrEH59d
TNtRL8w/XI9TTYRYCIvhIHTdXCTZqil+QGWPs8sbmdmRnhfZsqu1t4HYJ7m6ExLE
360XfKqMELi3p8yiYbjkrbodyVsxQ8q1GoxyFOv9mhXB8mRHeO7JWPPd2E4p4Cjy
QEPf3Qi2S/sIlcfsnSJWT0cPWSq4PEElbjrpdZ49SKA1pFMSZpzACbbORkAb5kD1
OlcN/eU4SFobxBQLtFPTuqP5AmZJ35vJmP1dRvlNp2JipSJIeF+msxXxDfGsU5kQ
7yikzRDg+5y8fy5ZSvrTtn9A1r5NivapNCZTw72fuj1UvToDo9y0ljw6iCdFEHNC
Y3mCaklfYsr5CJQWG3S4MLU1U2stLnKhh4Mj6wrTx9CUw3WXTXfeRC4OFV1HvHuL
SYrZS4ADXP4DazUCfoMr/5dVS6WxMei6QgaJlOPmdvH1fjRfJbw2fIOSZ5ICIFmX
xRR+PYrR6KGplQQzzVsPwJ0jAxYGBAcFO8qKWBOlkkJfz9DqY585IWhwM7D85mB3
FO8HhgGIpBiwLt/bVZsPSppn6DMe3AnqVEExQRQkcqC0NpC8MFa3Q61xlqX6cS86
8KqXt/qcV9TrKx6oleHr12QF4P8/vGBSKGpMD/1HL6gjupSPA0KjkubQbKkEySK7
qOuA9XQCVPjaC72TMI2dWVp9XN0dZVRnPvmXS873ivBWYCKqmdoFeBxlKbpwAzix
fpadurX1biLCa9zg8dq7r6Yj/PGVD7NxEsZ7r0512zslA2QPtgtomyLIqdFe50SS
z9LLYYXVT6Gv/VIGLxMhFpbTi7flnHIdU5Aaj7/T+9fEsO7ipCtgPtAFVJN2IdZ+
taPPJUPDKbJy9sQ/IL0jZhz9x1bci/s5PvPig1ffku7uA9Z17QAYm9dg7N+zFMFs
jAEcedprDAoMs/Fx08lm81ud/fRWxdoRRvzYWPc10vK+j1Asn0F5E0raTpKWzkTK
/snD8dcNEeDaFnHqxL+bVNIrD7+xY/3lSps8/djovCh4q4j3x8DrMM+CifC07lKq
rzTQMhJODTiqScX3oTP1R6/ZYws7xtDrVFrEGfd5TkMTv/TErL9pELRTIVgIqkYk
LEPyKN8Ydh4S9qYzK1JozoDzkAB9yaoi0+tnOZgb+7bN3ggkelAo1by7gf+zVy+L
LEfDIQ2eEtXWKil6lHPY/72+U5mVt9V3IsUTbLFHfOIOsRvZJM9UKf4rusv4D22H
wB33VzuaDVsgcJ/7iXkt2lSkWQbs3bUrCHfGgQZ7wdoQYNskZMXO392F5BWz+6yX
VvYH59o+0DnCYhcthldTfVL+g6jzvBCxj9mTtKe1HBqfH9QSi+14JMqXmNwWUFum
B0oKNV7ktr82VAx8ZQW8VXZYRmZKlkAajbkrn0QO3ZVGlBKoQhXE9iZIfYEqSKCE
fqDV0GXqahnv8TLO44rXBlwCFRlaA7qngvV5Pkw0mwdk/KdWi7CQLJ6ItduVvtZh
UVDTrUsPg9M2DeCde9rR4LALdctbvSD6RxzMvWparl8D/7IDLKT60hkiYvJm9pZa
5oxezzUMh+CfpEZkD95JG7WZK89b3ANJhfmeGve9ZzBXFx3cJO4cT2u7ZDrEl7Fr
U6hqjlYXyKISeQWsOmXT0kf/YQz7TfdOi1TNH/XIhGB/m/NvHgrvQFN6feKiBypA
91ukhxPX0jHI6VAwrIbcCr7sh7QND6xi/nPAooDT/j6JgxSTA1+dSgE/1EJhcY2a
39YJmzvNxpzOW2bpW11YEQ4VeRfUJT77o3MadFFhCMGaSq7uhnT99F+7NkecWu6E
oeSOmQmCcIEKPrvr88RBT3pqzXXRyQnyKYuAksnuzBmxauQcZwfXdwZ3a5KqRRJw
FLcdHiqRO238KrSR5r11Gp602IUrJdZiORBux4P0xwtxxQlizL1TKZrRrQx5sDyo
GA4ly2f1dVOvma+5Btp7M4ihDNEPJEGuMYdqwPWIer0wwDB9JgxFHJW82nrn3E1X
lB3r8nUE9fvhkBwf+WMqf9IEKypHC8Wsr+rw1C0nUH8qKD6vPgcpwXndCsqdTjhC
cDw21uacUlebUCcAVkYPLGKOVHWy3dUwJjOLpdtnYvidFFKIYFio7BAR43KpGPfJ
rw71j+HWUomq2gLUYhoevqlwLp9ox3mw39x/gweYygbKzk7Ry15hmlfapZ8+Bwjr
d3N4rJI5643Sv6DkAPuKkCGlnKF0KlXR6UIxSsDvkrhbCkzS/Uoiwi254/rdPk3F
oZ/7jqzK3omy/HZuzycJD7ncFGS3IriDRXQQ5KtRwoUuPWzk3JqhhIOMl68cQmyZ
NA6pR3y5y5t3abUYjnxcckr2/kiPXZmrWREJ+7BUV6z1IIXVmsb6YA1IZb1E2mpg
y8/BzZhGuiNuhGWfgN8AB7ndrFiamXOnz4gU3K4Va8EZab4qoCNTYAsPL57LWqs2
Q3bGctH3D2RChjVUYdrBsepu6LEm+SVTLRNnnYzLrvrE1U89YxF2MvoCbE9MT9iw
NVatNC8L6hyjXcsziCNDMpoTPtdVd3TTlJ6oCcNtJ91DL+VJTykiUlxn3MCz8t34
bja4g5DqPiZu0Uw89OoSk5Cy4MBj4ELSB09XfMo3KvKjNd1OK1b9UQ7AA5ytM3Al
8atH0ReI8GpOOsKvCkENFnB3gLeKG1ngHM+OpnP5nnLMxLYUq+pWU98BZIBtHnnK
KYJ7zS7XJaGvq4QQIN+Es+KUdrz6QzgrmbeZbrQtUVBQMKfRgOJD+mFFvPZsEJfp
iUOGyYX9l4bUgex+Xpkr6rcdfj1Y+MpdgGxJ5WID7rDwH6vIjuIJPv6GhUPWdJPN
EC4V4al2pJgDsSkjDrvPMH1zjPfOf+IOMkvmPhPIeuRw48z70tSLEsTPFcAU7caK
M4SgTms+FEL31cuDn3qfKj/TFwHHcYstB7TIa1dtMlt15nhwLVGIwhSTN9CKiG5v
96LrsoMqKmmxu4zAd8G23wVEZY5iqaT06AMSrEqx0exFeH49ULLon/MLpw0kDJsb
cU1D5wFDScjPxo1h4NreGuom4BJi4LbF8Iowbzr8v5WP98fKRIxMjQ+PawhE+wIX
zNPEjsVrPav3Mc7J/2j0qYSbUj20sqkBPCUHGF/YqP0K4XtZ3saWCiP4bIh3jPV0
7A6nlKfYRdQnqm9fUYtAZFUju6o4QPeUyam+lPy4kShUsyQ8l1wqdg/gA6ZUbK7T
5GmLBqh0tw0VQfVjjX60SekvvqIJbypfMKdWL/U/1INJ/M4GtSul+/XQnayWfcgT
ajic4Ptk2oxVeBypwkpSx8W57EKppCAi65uxDvkw7AAnbOfTGz31Rt4JLNTNPI5y
sWJ7/NCczLihAXtR0SYnUY9OLFVXacxx8s913P/Ok0hgcwJqClKHi79qaLH8V2an
XsiXwABN76Cq1f+BdXtd0pQpckvdMuBOX9JDXuYLXOQa89iAZraE/fbIVlKM2Ltq
CiDmAPo+OLCYRhuj1DBZcO5ak60MsXjyZfTWGtrkXRNb/nRRKZK7b+4gf32+TTCY
xbaV3hjL1/+OBxzselWfUEip0ihzf2iP3A8UVhZDdDAOfyBgbSL61e9U3UMXZw65
5gKY2Hpl2HD6g8TrGyxhyUe7OYCB0bH0CJ3Q3jPCw7h9XLhfXmcsS0bH29kTYQNU
Eaj5amLV6NQEvH1mdVBEh8Ot11ZVot5SdwJ/xK7ojaB8XLYEUQibCIOXq50CC0QK
ZwU3v1k1h3DZtJMdoRd3EogSMqUYNhmiI2MPvOO8ii5mvhXIRYpk9/h9hD06HMVT
OXrLHMeigT6SpM7KNJnF3Oc/t7GEKBepradrnZmeMSUOZeIlezx7p71n4RRNP7x+
XsCayvjvO6q8o5MDHfJ5b3ukEEw6ebYw02YDjX2oq5Yj/McD7zL5dIaftzzmeK6C
jZ3elTnh7ewx9RvP6GVs+EVBee/IMzDGSQ7KinB4njcQKXSp6Sn5k9IzPovn3c1n
JZEucuJfXGtc0/46iEcIFyV60GmJHc2KymFEjzwm7kkfStT2M56zsc0g4U5BtA++
zIFFxGIKluMJpi8bnprOB28bDZ2Jt8ugm277Pc3WNqyGOQ0HGfELMxWAR3zVQqwL
86bsXcHiQZkdGSV7qYR2Qrs5bwYFlXlQaajt+EkUGhEsIikhUW+HKyM7J63fU25B
kszihEamwk2Z1+Du6tHgu+HN/2MJZnlFPdpZUy4SQynnkONU54W+Ys/VqJhZXYlb
isGU/DZRlJPnhsrpe9tbcMuYkDlrG4ngx7458U8L4tGjVK8Gu5mAANLYqo98cHbt
/tzIerO2QWO9bCqaDD9u3koKaPno5JN79VSO9tFaVW+0tblrRU6Y+atc88uIOgjw
SV1dR6DXQddUjjcAL5bSNeSjocrT12daM85i47ZdZHx7wYhtSSS0sOy8NDXJ7znw
/XnuATxU121eaklXzHRGz3NLMFo2Wr9Ke6qe+H6PwDJZ0DxA7qEdvP8/tZt2WkQB
AeD12QOleicVBBAhk9Z5NECbCHkqF3jIHkfgyifDARlubBcNeYBkjzHre3IVyTUi
pG2g+UyExd+F/ti4zb22x2uZ1VxlZ8INbnNp2sI91UZXPxzxYlACRxO1P0MiZBzk
OwAc2gUM20hi2DYL/jO2T3JpTtH8mUPUUNXpap0WdmtrsLn+NyqL5Nwt3QXkgZm8
3g9iiwT46gEEj5Bp02pUhoepjTR/8qQ4H/73JZb+AOxKIHzzBLqCHibvEAuqwhWj
jE5zU3uKeCrMCwecP34PvLItVuyes34Z0IZyGFe1+VVHCYhdTqjB/dPhPLHr3XSx
sqKNnehBCpa6uJ7lIff4X6cWc4a4D6rAZg9ZnyFB15m9NZ55QoGgedZNENE/nd1O
SX/mXFbjj4qUFBsCVEPRz1wThe/5v35ASiC2vKuPMTB3PQovGCgf1ZwOyHR7QhDG
IGZWZhHb+YffNjNZ5a0DLRZu2OUR6PyvR2f8bUWSecTvqbouYrU3KMCHklEv0ain
j9d7LygTM6kCArsvDX0BNyEwFK9aZOFwSObZgGFH1G9BQ9tojlS6S7j0rAFxS6lA
JmDaHUoOQ9ouYSFECOTB+yUSZjI5d3T+AJIg8oMD/zmFpjU7tBOiWD+K/92VOlQJ
EXDkE4XM/ayq3EIz/3UfA91ltVjUnh5TA6cgAZ/13Zp1Pa52qeosV9DADuNHbygA
Vm2ygAHSIslMdIovm5Qxg0irl41KsjmvMUplKMyauSgaWcDjdoD59sfGDS7rNo3a
S0rGjgEVxtg5e9wQ+VmfplW8LQUjQL+Hvr4kJwTI6OL8VuROYcsUjViPgjwvQjf+
BY3SENdnUVrUjwkGVh/xBc5B1EIY+NBTkfuXA+P6rW0PnGXmymBUaYdRGnpQYBEA
5VglrawTd/NRoQ2uTvA0nvjWcSKzqSj3J1hIWBwaxDNxSLECuM9tJSAYZBa2ekcT
6tJwDq/8I+PsAFWXypswLF7MISQcHeaC8Rp+I2JGe5jiZxXtL77Q+LN1z/ipC5vW
x1Jm1X+H7dJUmGrbWfiGYe4EpwojiypMu1/2rvy5G4/KJ6NP3rqLoyG6pSo78m8q
+aJ4tadlvNrTJcGNR5DoMfzPoU4w4a2KAf7eHey22TQVcF5N1dfL8aQcBT2lKg0c
YcnpTC46N6mdqosd5GWyYl+0Anj+28JrH/aXtW4cswUVW46joCB2pb7+VQgHPzit
EuNFthVhwCNZPaJRB6izgGC4jzC0zlUkFeshUKCU5vh/RS9ngqB5yRpD8T/X0J14
x8Xtzxkr65zabkxeEo8St7dkSLaKiLCL6vlS5JEV67jYOJgxd18aOCPNy5FOIYl3
HaBTF/tSNRl+LnfVz0MybSCLrrNTKbTT25Q/N4KmAwMomNLvP2rlP6uNAFI44GuF
IxaD38A0/zjt9xnS0d1IaqwExjPz9cqxZRO2XBv80VqRmV6vHcZFUcQUEshISXhX
RL26FHUfOEOC4EN5+SzBmvTnC+UM5XC9InjRDXRo+46fPuSTkIJNrL/IUKzFyfqE
wciHy9hClxIFWMk+jMthTUKOmIZiwr1UfIkzvveNwC/F9K9w1hwVGMmiypJFBhzM
eJPpF1XWUOH2xeDmL4WQcT37m7l+si0vmgIMmCCxqRVngUf+ctDK55zVkCvkgBD8
8F1eGoJ6o4MER5Yj7+PEdjeyuVRly1XsAACdinrB2+s3HYagjKJ3ROdbC4eBpZPz
OD8SMyiP8nl4eayR8GMGxRKooxuB7Xj1f0avik1aJkDERdqi5IxDFKnoI01HyMBw
GBrloPqr9ELSMSdPsIngBobTpasjyqTrVpvC5rGql3xVGDUiVCo356TQf7uqkbf1
2jAr3RpbHbOX2H3LctVaz05YEH13ducaH/lmW/drEwf6TqXoXeYEOmWsFLNConKn
qfNRubqhc3937mwyVm2+UeQZBNeljjEwGV192al/XtTqMGf2vnLzsqO8SmAm40p2
R+zkb2iXOK3idO9A66PwsinpBuQOwZpmxfPEDzi7mDAuXsSPWB5Fzpupo7uFioqs
WBqnC8VvuYg1cNNZirapIVKUHMoYM1Y12Y3ggKgh2vJ3sEnveKROZte6IAmCcTE7
X3COTOaOLBCDUZhxEO3sA2BA49KK/rmvJ2VRXRRrKPRA4RblGyhp/fGYEn2HjEBv
cl/ckiYgsMdBw5rN6oLmlMCSev9LSbft+GqHSa2ddNxp1xeq1qirgdb5+IVQtRqT
CrMuIdjCjLmId6/XkYNKcL7AhDtxWydHg4vwpBLOadGhoFwp5pVCC/84QZc1Al5n
loKNSSVDevdjurRFeOtEedZwNlXAWL0YwJFJBmASFPpKDh9PJF96z9qZiT5iu7gl
i9iDLTfB6BWhoybgAnn6SRUep1Z4CUD9hSKPhLbeiG8ifAQ6IjRdyEjqu87iNbVo
500s/a6DQRx24P3PdluZy7FSz5IGO9Ue4I6xRUsjgEfQuqlCBvQqxc1iJayt4PlY
/7Kj6F61gOGXKoaEWMOsXe+oC5Xczlm4SucPcINSC/VZsZpMV/ObCJ/O/ibCo9ZA
bw6Zc7q9+oifWqGb/ho21YuTJTroARRH2nMcozjOAYseLFY2x00R4+iw06MOBwHw
URmgqQRd5/2xc9k+2tG9DPsqDdw1DLNJgpIBzYBJE0eo1p8QyfRWPyzYfZQcsmJ0
soRR7vPfG2ujaUaVyM826FW3WZC2h8M0H4Qfpyhza91dzDkjOhQdhdL3zjhxJR0t
Q2GzzzzA50ImRLuyfPBICDhezAt1Id2WTtumehmT/RcewAt4JR2gH1YJM097O+RC
5meCzpDoJOqeNwjZ1ZGoUKGA247X6oxwMshxjAw8Glv0WQvYzP+FRZRwtRI9AdT5
HB8iq2Wlw4uRfyO8gZWdjjs7Qz9SbCBVx7uWOmcO2jpjPcD5pIw2CKkVcCWtv3uH
MRmEkIjfzaT6Ep4JzuUos/Ol6s40rUi3eUdTCAMKAd7+lher3ldDsgBjwyEVPFBG
34uzN6ksjFDIeeKdm88XnJkmPLBAFaEeipxjFxicpPr3KoBimr5K+h7mTzgl/wyo
jJZUvNu8muiP0shsUKPi7N5/mWQiklm5/s5xtPNS0FjE77Nh9pPXKIzXSrLtmo1D
hgPkGxyY8ydT17eZzUa17m4vFlXzg5cHIxCIwlxhP6BY06c78ss5JZPpc/06tcjC
evEBxjUorN+Z5TW6ojLbPt9NdVHQZqmM0iQOk/ZJ78fKmJJ0PrHaTzxMe/hX44ks
EmjK/01TZkqwfLGOiSjS1TO8Bw3t2+bkw/ON3nyjtrQiIoPD+QkF+ekIRqQYyGiO
//EQRelp26lTohwNyHZffmeU4+g2Y4yoBKhLT58rmHNNZSIhC26UudND7OP85hfS
F2d4odBh+70FhKG+Pl3Qta1+eJdMSgDkAk7QJUpbr5kXm/Fdmae1fVUUqHrH9p7F
fDic72T5gyoJJgpZi1/NwYG3CSScJU5CyAI30z8URgMIHeS87BGQkXgdn0SHNhrV
0uDisyVVV2gm0DdcsmLMUXMB1Jac6u4J3JZzYrTKDzjI2xlS4XQUBMbwsidAHG+o
PEQrVneg+mLT/lLhUu+9cC5nPUY5UPaZgEL2yyUUh7SZEdQFP+qcl/GBBAeidzKo
ZFcYTGJinMTObLJqIEnTqDTYkUBcP9SP74P6Zn7gM1Gi9zZTO1jyN4gxUx6p0NXX
kRDrFtMFT/HDdFQKkZ2FJ5i24xEY1Ypeh8k1daGdu4ZfXJOPfGhtagHwvz0nq8z6
VS3QOFNAcky/sdBybriLDrf/IO17PU0cOY4P+ECkbz1kIGaU2y3gIoBZg+p305No
JUS/CRvh+n58l9Aj/1NBQ+teCOrNKM10bkO89sDvXEQmShOJOUxVtW3pxYD71fju
m/p2rQWnAyOLO0yCKjTX7nudsQKTieth+/LKlCANTfZKr15NYmtDU2ooGDLjI10A
PA24bWmWkTs8LVw1o7rPh4O3KFRBlS0/EOrpsVt6g45s7/2iRLAWq1Xf2ZDOT+Uj
vDEo6O3+3Zl+K8XeI8SJyZsBd9xlA7OAFU8lDM3Y+hqKuDvWw/DjkhC+KpRGlScC
gANpANzb/fE6Baia6UUJGTA2MzJ3veKSTSj0sAB+xt+9VyQ40GEWRg/Xsx/+MXFH
t3yOPvMZzcMTPVkUVIMWmJLi8SZbsTKe02Tt9rtuAKQ4E63gb/bEcGLRXRppZPg4
kNB7U27aVQdheVlJbGduohL8NAz/4N9APT5QVCvaoHJ5cAxC3irVGVbPczPjnafo
uuB2lXI0V17GjllcgIlx8ctc/8fT6bd6qGZOFjp+v6PdZElXr2Ht19BI28QyN31X
YY1jGRzJxAqWe8AvfoUC9Fp/o3uWs+sMkLkRy65C9Y0ksUwdIOWC4lXCgWx+mO0O
4+qbdsPG4TOYChHUE4BVUB9PxtSCfxglkeNIn950dkcbMH+UvL6MtIFlEJagFm4I
UbOMxv81yYZww/fxpkN0s1mpwhCVIHYRZLymAotdadFy/fyA/X+ms7QJjRr93f0l
ErpLpePev+ojbszJRDNsggEWy8EnLjS0jPoFlNHotDcwvGi9ZughLT2/tXFuf/yh
XgZ2SUCe8UU9UA+ZBTeXZovIG+VCs+b0p5a5i1taxdhGxJsxMOW+yUoX+T/W3aA+
K+Ldb3GIAQWPMDSJECAMTkm0PE+KvHeAHe/HWopva63qU6oZsxiBu9oLRCL4veXQ
bVGDodw5bhkx91Tchmn4bVkJiPcgT4GKfEd0nLzrPXkkuX8SYR11NxtKwoXUCxqc
mtrKEbp8SApmcFD2ImdI1P5WMYm78vPaQ+b9SsbsFBMvNH3tTHajNvdj3uqKOX2E
tfEFoa+cCCab6FDe/46yRRW9JBL05yI7QeLW+Y/DoADMSQxavWg2HxLft5SFK5QE
vZrpP9DwLb3NV+9KjLsRb9/u6akVZdIsTtpXxsbT/Inw+/gEMtzYoXoac1VI5y98
gj76X1c/jFtGEw0ISLItVoum3wuX13R1gOftE3biV0nCv1hNzSpdz+YIaYqaWa2z
7G2QUiCARPnZs43dIaKw+ftUl8RCDLVqZmpf4Co3F+fnLGNUR6NacPgIcAkp9MFz
xmW+jzqs6s3DH/XGazETPMt/R2QNBe0xdW0AIuLDSF54tSSWQ6G23FjIumgWht3z
RDMFvQRfWPLBtKPxU0BOg1nmHxkKe4JuBcbUoBZKkQratuaj9Hw+23SoOHtoIb5Z
aD1EQS5u+DR5DcSESR6FNR+qPc3zqQftA9LH+GzblMV8OA2H4nbIaLvUj4Z11Pg0
NfHK0d2xVjG2uH2aZSZsQej+ZpTW+bmOOe0yWU5DZimvGplm7hgpaedvspyRNXxF
H0lyn2dmQhppYAfSv6m2M8IDCcBFnFgFXtX+VP1uZGFKUQ0SnM7Kj4ZPaL4XJfnh
eyjQ27wwZlQPlECMRZvhkYnvBtIFlSdzf/i8MahigP4VITKkfwB0O3b8idXPXbZr
EnRRuNv2GJrJSGAZO/rk1YiQh0cwKV783OEyTYpm6614+BZ7IBrmIe+WvawpPhvs
B+fMPZRhIHQqR5TOrIQMwcqNY9x2xqvNUqOq9vJIeYrkQDYcHTCRWdllYpCa4r+W
a7jww0G8Tol5VwQIhFb2+yVJjQfk3hSE/Btbv6l3t9wFPOHVga+wcFmrw5hVd8An
K8e0s/BMkShIcy4njhhLjMtUAvIfeF8zZlew8eo72Us9dOgzu/oYu237hanRCgoW
cVRs2aUqvO7gSZZC8gFvIXyhPsubU1PWpco7MLBKyubUEqHo+AVoFMwZ9ObTvbgp
s7OH16p71fpfOM1ithbS1eUq4PSLn2FKLKyJoeWwgwV7qe412SXjsQ1YiUmfmpFB
oJZrSZwFs6PWXrC8Jgyo+O+GjF/qTXtOOPK8p0EW9Z0HWESDgUNoE0032RjwCw7d
R6xkhqH6eo3cfIyX7sRk9aga+9OE5NfFNcr09qt3gkf9RGSXh56YMEhDUreggibP
z9QaQUVye42VcfqL71TEiUVSRN47Q3zuvgmLKPpaIrG3IcPfN4e6eXHBANqu/nj+
UbCoZjvS7/2/+obVnn751FUQ5mLzLGZlFNmg+nxa3Xw/iyXp5BuW87pivWbW0IaT
D1oBsPBuJM2m2zeOgeZOPTJTALIRLlSjb57wBnAWCwoxvhlRkImpkTzwu8VOLdZ3
0Af+0SLcLWYnrHmT/w5vpIBWKOPGEaDGVxE+N19R2/yOOaI3WeM28RUI2OdCsMj2
iE5nnNc+mFne/JY2KS8hByiCunvGoAMz7aCjz1HgMUrKFNwkPy+eEDSE0cxNqfuJ
dfGrRvw4xQXaBQMleWKn52NB02Oeq82Lfz22oHNN0Pfpm4xsrPnWGsD9NVYm2iis
XVnQJ2UoTcXdDxJ7RTSB4w/YPIOo+sTgfK/8Z9cof8FPWjRFNIlKeC6NoWC1gI7w
sILuIgWnxSGqBwl/ijE8QmAzvh36peEKtHk4KVGZnj+Q/TzG0I6WvTnKr5bd43Wm
o9ujSjgICd6OL/8FPMJSP2ycnb+0filbCKIYNnX8Ioa35PRsP4m1KcbJuD+pcbHL
ccn42ugZrXFYPGxD8CyLqeQHVvWVsswlg1U3kTiBfQxuYxccdK9vYRfc11c3CbZj
ULJ12i//1DalArW0VT43ZeiknF8hvN7SN/0eHJ3J2L+ZVhtR5NlTrv9oVNeIsgoy
0cmeiThcsEFaU+ODqDuxo3nR5+TnraVmdQd7v+1cxx+9g4X6lWwRH7oqYs9ENo9w
MkXLiuwqabmgZI9lck+YVhZCEgp1jfXYxjDGjgMe2gwEP4hVxze4w/o0i35H/zsB
7sae2KHrlCooF3X7GbRBXmYodKcQTHkdy+ykOUVn8VQuamAHcCXiKIMDkCS1Xtvz
e/E2bQtDQTGPEZCRDogkhzrI6tmJd1zts5PudE/+BR9Y9kdhxXHDEGe+Ie1n+ZIQ
Hs41S5+7chafku5XET9ZUdZkMiWJkYkwFuoRaH5GgVCFccHhDIOsxjD6wC2XwEFz
HzEpqLlNLOhZK7TrjDrX2rgGvcfBk2FxJXpAQ9cnQ5m+wfiUa60oURI1yEpJHFFl
Q3+8LH2SPU3twPqs3NedNb6tv6i+tye4eUk9hmJdW4xuD3ncHehOPzZgY23EU44g
kcBLMJBbTHtRyg8brC8A6gycB2gibY5TgBz1CJb1du6ubkd5QK7QTtYj7W6hn1Xg
FZaU+i9ljKnDZ5Fzgg+716gYXMVtPV1b3U6Gp5KpnvM/IMMCkUa3oStiQNVymF3T
OU+gKc5HcMjeW5Sf85itYoEYILcLKtBSBqS97Am7cbXF4nVtL81c+um0ipgDKRg7
Ob+3q8lIxS09xcsV8Yq4mXGl2zzKkHeYDhZIWqQ7/bmv0ngGSdYvQio3wvnlgfuo
fCfRTXDfqzFW/ow/0yec0il6Jp90Bd0gnUj1oYUrSAyrXcbHMrAtb3yQCohkOrf7
Au2HBJRLA0jiccp/2dXJ6LEYnbGLr1xVqWBy6seyd9p7h4LNlQfToZpWBevRCrYR
QODu9fbKqReJ1I/rvrkQUxj1FGOnO2NccJXIqQRvvnUgfG0M3SMg08qJWC1zdfxq
/yBU3iYz6vdFF95QK4nq3HMZpX+bZCtdjKeI04oNycMifgr+XVFY5DvN3SzuAERi
CYZ2+DssfOu1uTztbtvLuHmgAufRqRyIlYUTG+qDThF1yJf4E7nRlM4b93Q62I2J
ZolfONMRJmw7hhymUBBvWZLRdnxCnkpftpOxjVq4F0AEVlrUIk2BlU3RGSPA7xpR
zdVEsZBlXidvuUziL8hEaCIRxjh4DFvw4LLdfG+PNcpXV2ZodnnNovNQbHYcNzBp
dn132qp3TpaytJ3SX0wnPzO47xA7g6JFFyngN5UCv/diH++quccw005JxgixKOlx
l9nvR+6TLe8cMlzyRbS1sRY9IuqIszXa59rl1dgD81IWmgZ/aEgba2VoW40w44l1
+l0hSnaIHE42JbfJGfThgcMJNEhaUoWNDmuhHw6+2h2vC2oERlNs4qaWqjIKplBP
9DCYU1k0wvy1cbzZFK14BYQu96ZGXCQO15Jl2W7jQhJcWZKuAbpceEA/setPgeFP
f/PMlhLPyKnKyyqk57BN9PD0hiPprg5GhE9T4oKWHK6EEMamUguM2hgBTxpT0Yz8
o6PjbKPT0cpLbfZ27LC/wXzwIjlwMlkirNs4lzbV2XQf1yHIr0n6CYOan2Yc95Cd
HT2VdUiiYcJPXh/o6tcP9NhNBlkJoavyntJV4HcvPanTQ7aXymZLFUr97VGWgvo6
OcKJyOuNccgtgWIGUpITy+QTs/8zST7gkMRcaCtDTZAoDN7r1a80ptzINGD+GDeU
T3fB9cPWoztjNBA5soXuJgCpEPwGcUUfVleYnnhio6184T82+9YWR3PkYPDJ6GFC
hpN2T7A/EEOFiHucF0o5FH34gTBHJKlGz5uMbWdKXxiQJ/g45AeDJxk+4rZGqbET
F/g4+pZ5Lz0qDuW9KA0Wod5umbOTRQ4972qSJCi43R+JCTlm8Ovfm51tQuwLU8gR
Kfs5IMhy4g1VlTPDpeELdBEGt4/SwF+USw4OnX+SmvRGuT4y4j6qEYLLwBQpZfq4
XZN7tvJHBZR7P6LENDfn9enDeIeeVUNSTyVDYqtWW+Z+raC3UNglsgVvWsR0D9cX
d0Fegssig9slV5euPcUp+iDkb/zIw2IJqFVTi1TGhzJIBt3cT2055/98gjZby37p
GTC8HTUpokA95zxmHOuepr03RfRsXlIN2BxgZDQvjW1IrQccssxjOyKWbiZgEMhO
mAHOgIyBgdLtBsFM8L0SsSLOZ5dIEW7TOroZKeCvpXggPe8wPg/EaMGBGmMWLx1O
0j5QMDCl3Gqf3bPThJioZKhVDqBd4VEvq/io7rONvfkAWxuCMsPpORiKgsEGyfHM
0X4YVhY3LKu0XB04oMITJs81vA5IkZkehDGZDbSg4CqtQ/84sl1zz/wioWoxGcKC
AKtsvlFU11+54HeL7ST1BSqV/xrr1putm80yNJgHS23SUY2WLsJJWmV84H7Jq/xT
RFJKXvnX46k5RTZN8Dnk+ERoxQW7LPy98Z4CL/h/t0eQbPaT04yVksNUBHZPc5Xd
zgVBRJPGET6Dd1+dlKLeLRBDLJ3YtcQ1B+ZS4nFw5hF8ZqzIL2ILKD50SRWAwUrO
dEO890vnQpOW48DiCZftBfav5zXfcSIJ+8zWJrxAGe7kMz1L+QDJUL/Xya6vjqD0
qbf/VEjhVGBUKqHE23CpoqsAT3kWKncDPD4Lm3klX7W9O1IFhIVcsqLfdaMcMVxs
vEOd4NQ6ckYH/hnoaQq15YyJPMvhR+ALNrwUP0jsrDApHiAvmG2DkDajEPNXyjah
BR7CG9hhoSLY1mSNJwnH9zG2okp6Ioi4IInW/j0YD+arkMK6gws3AX8ZIUkQTSvB
sI/wsQpZ4YLyGtThJO94AN8tqyN126ImnVRgGykMMih9K1P24myDgTgXZ+rN3NRy
D+9Ot62Zlt3WxnKqIKcSCBCDOMkFwff/4IOXcL2ReqU8WRKAjc6alifR4FJfhKND
NKFu/vYQfc9ssDKzjd31yqrJhJ1Cuav3RB6PiLnDrAP02Ma9PeeuIGiAl/4DXx7w
AHK21O7ElEOeObmVvBdj7LHXzil+W+ocNiBUR8KQwhoBvlJ1qpQBR7C0sqTecO08
f0H/DizyvK+DUZOEUgvtA7LNdtETZs3eLndCSRul5x5nok+fe8NPVR8rE8OkSWg/
a+j/hLq9Oe3Wl4KHN1ifPGM+omHuGXb9T2ptDfkq5irbzPJWe/zyjzbNRoUmxO8B
IxeYsrHmaKzvxPd5Cj346LJZJHRMpngJsK3xQ8LTziXssivtpgINagc5xoxzax6C
lnjshTMoBn1tiXVrrRW0dKkdJLcmYu25huHmITL9/Q1tSFfrvIiSwv+/qG/lP3jd
xIDn2KRj0lcemk5rA5zYPCqOBE6gN1uKP72xBhEXK3RWkjP7ezLb5iiT21NhzDEm
x653ZeMW6NbsZeKSNe7uvj+Pv/eGHA8tBGfsFy7NkPqY5XQ8p/G2XvaT5AqyN5W9
BUM19XJ70BXztonh6HLI6Xv1HnOWTOBOUelPGzHSs4heNuGd1dwxqLUIxzo4QVFz
yXNugJ2+gbGdw89xeNHT/7NcPa9CVHY2qRY9Bp/Uu/3Pds2E/bKl6o/Cb2/aKNoy
jWd228+bAecls39gVI0XIzrm9QUHgw2HZvinvgRDJ/ZxWe8d7kFhauRIC7WACfs1
YftYgSUE2eecL1k/Fmh2K3gOyd+vOeRPgP571rrO7bOBSWrJmgCF2Lc2Y32Lyfuf
+ujhyMqoPd8zpUcOQ9tOZGXkIOVevXccF/hXsdXaLXrra+BU9elgBfu3YXLopQg6
hp/SwsZdLGu+HcLjK/szfCh27DZaSy0vkVk1lwK0Y2qh/e7b2HrkmFk9oFvlMRec
DeODWtp/cU2XP/JaDpSYCUMnUMbzTn97ahbRGsHHmpcetSOPOcl8/CCtMuN7SP+X
W5UQ2I45VAVlpesDdI0nvyDVBxlexQ8Z8EeH2DWK7MVW6AX39cdUij3146m/nt3w
n18zNSUyxTuTZYa+Hka++uEcf2jW1F2+sSe+CgBcFJU9U55vj5+mZ8Q1mRwxmGGY
jCanVlLI7mXpoWCS75TU8iaoxg2Dfwdsq3g3lTqnrE35oeIYNrRzUauT2PYimWwQ
0A6l2KOqJqFXzHkzKoqlo4wPKA7/z5IAsrjild7qu4gLXwArpSr8BIOqIPxaNHiT
e6tPOZpcSdcA/H2CRpf97YTjbMmwxTwsKxL9aDYStRrfPCRHmwMUp3OGYwOIGIni
J8gkN1d8doZAae9ibccjx7MXm8CNs3+leC7fOp4/iTBu+kwd9vmYxrb63QgnT73h
viG38bmE05bgfI+G7QOw53mnuFugyewwR6Hyxw5KlODigmDrykeoWDFhutQGEWpF
fqA3ZSwWK9qvXkzMKxarK2JR7H3bBgMQ/YqvG9TyuE9gCwhubJ1E39i7jbqmw2r0
XwJzqYPZwkob7MzTdFvfPxLfv+JnvFXrZIx+Jgt0lhamZ0Fj163vH40D0ZwLVQBi
Gfs6sH+37ZfCgiL9jKXirH312+lWLrvzXwWCSTXvoknuDINUG3H9tlEwkJUiSocn
wxfSOdKeESUsP+G8JATrMZUbm1mrIULlVBM6/ei+x1cIxJVw3GBDDj8LR0sW/9KH
2fqm2uAnwTP59Xi3QSnncz1qMToIdDXQLOF/b8I3owZt9U/G5HcUfGHqwRMeuYWo
dHfLBg0lGLjlUsdAsopKbDLA7MzpoahOMc+EfTe5nZZpLdSCnXnnqDiWjHmtNKxr
WTzS7WmxXRXmwxZxQOn1XdJZesLjgCztXkoajimYHfrgJ0Wj9n9OztZT6THDV/f1
JZAhqSmyr7ar6+kzuKw29lALCPVN7IbhG5WML7PI1ajPzC+jv9YIj0REjitkb9E7
4Q0yCFEbgqdS0BYCBuJ/YyZdeU26TZjEVcvQnXzNMpmk16r4PsXd/yi5dBrQNQLn
w5xpxvEzCz8I8sEuj5gWsPDHB9ZirrUs5xLJUFJhwgfGDj9cvshJehk9DM/mqfLG
SVXtWbN6MeRF2HN4SBVf3YYF4Q5/G4cnjjS/HvT2hgjU14uT0WFzzyJ3+JZpUKlV
Sq349lnAAMD+CvTuK2zEYbTnaWJJK2kfTwCjzcv8D3X+mRVS1AVUj4iHka5SwghP
Bagw0Sy/jMoIsqNIcq00iyZqG8IwX6Qr5HZ7QtQayDXPg8gDkj8trngyRJTyeWH+
9tKpJ1AaA3Q6O89ZXI3LLmNPIR/v9rsweth/mxJ73DgC/1OFLakWUeKwB8hDgSTf
Hr0YMk2MhfTGOGnua9IqrbpHdsbJH+ikvUlGkBMdYSYBfdBwR45EHcigG0VaZQdr
9YGDO7qpbOpmut3Dxdhgu/XxQdiEiNCKiVOJeQlx3VuY6sU0Kk7oZSaIF4JIH7ZW
+f2Lp0b7yuLX2bOIyiDtoiSpH5YN/UOT55z7uj0nxzhrjbOna7bmZzGstksPTJsR
9PaalX/CkH4vWzvbj03OI8whZLWQumClbBzOA0aeD3yxz+PUQx5Eqxs7f+IEdhS5
mzDmLTk3lMl8pXeAF2v9i94y+cOB1XN/dMjSu9TzIXutOPSx4CzTBy1EgmCAyIlM
zuoYfnymTwiC+AWyM9z9f04DMSLdGWOHHupxuYI1EDQ2W74dcG9kUSyutnJhGyeH
OuRj55j8ykQM/LJf69BF27nd+/G/ZJeEQjXtLc0ZClRl9qf4AAn37h9QLZbI0UwV
fhCFZ1uBmNRztLp1LqwvwszJKPwmEfRACmCdGuhYO4q1xRoR2G8Kn5z+E+UIFJ44
VLMSLucSBOMwe35zRBJxgDfsICTgLKJ1RIOyDG/kyJBJH9wZ48YCG8MPL7qm25C+
ldJfepd5MjeHBeZ/aLv3bUt6zH8iaK4L6YWdFV3D6SmrMQFfLDWbsK+cFpfyYzRV
Gr72Q9kyvz5i8BGB+ygF6Py54Y5+mFUmVEFVHVZIYl4c0CiIwjbZGr5JYGinaRaJ
UoRXdU27nx7E7tMYLaoNbmbOTOfTarNDp9J9Zo5ok4QlpMlU/KUfStX2EThE+7Xc
WwFvNY/EKMAUGpIT3SfyFJK9QvnpxLuM0B6VSTWwsnTqbzfauJp45cn6T4tUxzuU
+451wQV0YkdcgneaZ6vvZ8yodwtR69DWFU8/qqoMYHNnt5PFRMgQKCEKhQGZfmn3
3KIbkkMQ5hTjmGtC2CVcVL37HhgI+rsJnC1qdtX3J7lG80Jb4NgHUNUtXdUotmFh
zNWe9PPSFUIGMfwk9QncbQ7wCmE7TZRI+Jv+4hoDJii6cboQZ2j/tJKvltnCBpzf
XI+WdWbimHwPfRYSdTZkd8I/xcN2+C/r6OcgnHrUYeuxtAgaQKc+55aBnxDrTZb6
1YXqOnipXLcwf+PQQ0IxcrKsRFKYYSn5JMbTr6Lj1tJHsv6ziup55deawHhl30TV
fpZodSgV50ZeduyDHrqEzaVXENyF8/OC5TqGBFIgv/KGyPRUMAEdGvsqDh+IHeUD
uvlrQf/Cp7DEm2GZst60tofX6i2MvkrC979a1r5mF2h8eUPLZOoqse0sBurkZdYV
6y5+vR9wArZ3Tsk3inNWwFgwY3F9JqFn53HvXSfNL4XRy1xGE4yXT5ZMFJ/JzRll
z5r68WpOv8hOydCDFKK4iMmNUUc3HFlCebFH8RpNa77cKHw3NsCSbxFfT1s9QTzd
oFbC23bOTX4WlP59ndc7VenK8sB54P7yvGW40i/wSlAFKup8D645HyjozaY2vzCA
BprziIUz3K41YzC2vI2yHLC4G0oFU/BAEVUHQzp//FoKOjOMBzItT71fPImXct7W
8mwVSwUC5xL2uUZNaf00PzjBLwCEj7eV/BSbAQWwtswJGKXna6K08CIU7u7vsJWy
YjsN4Z4YiOQ+AkhfuDFQjf/1DVvwO7JlgmVRyDfttwLCxQQIn2LE547C8LBnjwGX
Kfrc199yXF26HWJ99PUB9mSBIsjfy/1w85c93rdCUwdEKzXMICTDgWzbsGLCiozc
y7dX40KKnTfAslYTaPwNAA+XEEMgT/mgdWWYV9f0uXkvjebAnMTkE+FQkPhIhTlF
NdeOyFmxqm9Li0ZYHuc4YhcB4c0+vcJkmTVYU1rtNB1IQen1ezExnucPshBVgkAi
RGnmti874rDm0IzdK3LJrIl+aXSpRENYsLwsvEH5FWdXJs5xFnZm0sq/45lpYwyW
+qr4qbDMZqc+bOAvaNBst8SE0r02hzihox4yIw02KrIIVJTdNLksdrCGZ+SxYSKr
MirjTuyaIjXRbJHiJpsicqdNzo8F2Xh2z3REhSvedCK2j7hy7Wk5ve4qM0ilUcgF
S3zl+8CrML9gEp58FWNJoEAQQx+KmMnHa08HGj3gL1YftcVAq8ksSssAGotl2of/
Czee0Zs1LJDvjwDc4L3xSfpALdP+WGsfxy4GiTl76KA8ctAkSiQDGY5TrJHTdcVf
89jxp/d1GscJSOHy0+RTQYoxKDqEeI6TrigD3FxqvXhiY9tms6HFDv9DG1nKxdD9
T+T/S/3tcTi7COtLWA2oI2uytEMwK6E7MHiazogsKJTUOWWP3s3CeXXPMk24alL6
SGCUZ4G2kOv3XN1PAAUYhkIimQTBTE6SF1xtsdPCLSwJIpS8soKuwITSPLyPgNiA
0E4xIuMVtrVBFJ8lKQMosPV+ILx2lwnZzr1y8+/IISrl6zyFMYUc8sQ3VE8K39uv
NiOiVfd9GpHNt3S/sXV6plhD2SlqokXvjbh1ReU8xI3E1cMR2Epb/LWeC0LsEiUj
wxC/lKPt2jdHzZta4BNmdfc2PAtQPcvI0TeUbtETQ1oIy3bDfbU3bmVJhd92sWkj
Q/ocm2a5wEszz+d7VfFEljT9r855TKj/bDyzd2kb93JrH+UDxil1wJv92Ko0788C
jf9F+g5XAYWCd7DuVzvnce5rZZ3WwsGSh7sdwfog9Xzf5DABhr36t5BaSn0oHp//
ftbjPG2XELqKTFFOQ3HN7puBeOcrXBWAK2xObJ7Pq4oH4i5mjc/1TkzS7NNBvjqD
wCGEFgPffkkC++kVB5M+7QIApVHNAbklahXdseTJ1Gqqv63Fj3GPaxCueYDfW/XG
BDlAne0Wr5ojPAdzhpG+cG4aPeEq1zvMy8aQyI0DMca2itfLS7Mhhz4E0m/c9XFh
N++D2m7ZgXioiRJd3VKHLaNal4iuku0NZrrB/ZZIdjpGtvODiI/EnLCEVK84+/wf
9PtOJ1eU2WewAK8CNJIIUYNn+czwU7kaR/rHrKMQl/AcJVgvcV5ASzVxmXnPxekH
dn1fJqJoEatu2FfAoJwgiz9ftQBPbSgG0r69ItRk6lMIvf0KUtPYDxKnzQ/aPO9w
X68XqQy6ONOhxh2Yv5KO7mz44ryeQ5lBn2U2BohH+7QvGS6KIZSSnNEAInHUFKeb
RVg74tSstESvHVnUXR/MvnCJO/1/xTCW6kxWmW8G9azUsovgGDi7tusC/E13XPTj
eGhY1mmAE1b0+AHu/5A4UFPMeoIV5DYR/d/jY1j6G0ROti2G4AcD+HWspvDpofO9
eKki2hJyfIXzxtNP23sD9CDB1J/50vt8AtCGFpNAxyofvQFxt2m56sWigEOz6Gm3
RegqJxBvYaFXeAOdyeUn2+8ip9tSytSkkzsu8+8DhNWqv/d7c7BglqYp8pPtKGEQ
`pragma protect end_protected
