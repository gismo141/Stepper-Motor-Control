// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
dMsb2I1kVeTwmNo5ou79RuglEPGok/G8o9hljOolE+pLXzVjbmKGDBT3IWELCMX2QJFqH29S06US
29PqH/cdX7HeXa6jVfOfK5gTCXjsEbCCL2pupqI3hBEsDPLBKopOOl7wtCbou3t/MgTi3e1UOhR8
PGE/vgNRuy9kNXR9yzCsEMIG7PH5GCUUcBS8r0M+ZdoczY21GsOFattREt63cLdCAgKURo1/OLvn
JpL72UZcVA7GOTyeAmKnax+uhY87IY/lz4cZKnaleioX1dxgjAq+ROMY/tsIyJgJAu0cLF0quqkY
dZaixw1qOyqxVn1YAhVWOX4Phg9LgCr1YyhYjQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
5V/i2uCh6zJijS7ZJQYSnBlxFWdCDpZeqW1UjoK9I93TYCwzT/juLFmTpDwVYypQ+ehiHu4/2dVi
sbWn+EXQiS+ppUk+omn9s3Hej6r4fleNgHLfcROroGfB5Hr0AQpjypIkBU6lU9Dxeyz8DVxUpEy5
lclpN7bazKXPq1cqvtZtwdOPJJ2urSlsyFz3xV/XNxT321+YpgH86rbpXqy6DrIJvhxjqFOgQ7Zk
LSahdIZfSNe4GrGMEdXDuJ124+qtt6aYNnk/at5SalbzXslmdMCAfHe/feLE4Y9r+jGH7XqVNtTu
7hx0QtYNbfCr/NFJq4BDaiCIXlbEHf8DxSoy3OHa8bisvBjG2hL08RnxRbg1Zt938ortPS8MmUgF
RfcP7CiZGC75pRQm3qfxMZyg3DlMND8u3vhpCTjksR6mK5Jh9wgIXDi99KtZ9yUt+bUBj3MJL7pV
Dt6l4nSMHrc37Tn5IgYj+4aSU2E2uw6te5yR3C+/v+Vy7EWE7tFF/MZqZP35BQC2k/emBJlVDNZq
jp6PTMm1I/ICH7Fst/3HcA7NpgSFt9exICYxhavWkvmbA0FP078w7laimAtxPTW4o1UVqfvmP89F
HPI8WwI5NIQHQ0KPW7hNKARGsYv2OgN85mOAkCFUF5wn8rZjLAnLUyAZrEMxX0e1fdOxa1Cij3I9
l9ek9f1FuQSicvfDfp6fFMjp2pC5Rr3EawBc9zXm4qMTCa5IJicm9mQWs8mfDOlJqfen+X4kPzJw
lYpaArtHBK/yUYnGXLycl7182ZyyRb7nHO0TcVM194TvaH/c93tPQjqmgICnvHyjuVPJkiSlKJdT
PBXTxdhQA9ie0DZwYu1vjfnZJzfXZ4pns+fzB7xNy120rvOm4DDcbPb04N/vhvVeOp8Sg/i3N/us
Rj8Ds+LZpLySqiMhgFRPfX4o6okAQH6RJaNgfIqqi8dRx24D++XdQkAnpL4j0VuDW5+/Z4L0GN0X
qcp44nxfggfxwq/ngLzjeMMLiGbXsZLuZopR28zr9hn7dDUYQYn2UKi2+g/HcGcMGaEwrI5qslKF
AhZl9MIupHK8MQbxusMYP0qH0yPta9DyxP+8fWGDFGroBgkBXHUY2zFx5LsGSIRH52/lPyH0m+ll
E85P7ttR5w+yY0w3IGYd4H5LiGc9a9urdvP8P7FmVy6zWE3z7XZviu9NpOjZXkRiMeHJcQAV6een
Dw5OtJ/UCr204JdIEzCziU7zNfhpc2pk6WcHL8ohofReUrJzjwDzlA5cL2vvea2AN2Mo1jC7gwa9
cIq9wSWOjLQo2lr98q5zAiLDsE0C3A3YpC13Fwq5CCJlGIo3no0PKT0AOwYafiMMvj7mE9OLq9aD
kTTJ1FCrIVTuBLv2Do554i/ZcCVARA0lZ2WCpfh1GYYIoWrpq569cuJrDpainMSSGxAl4XL+VnXk
gN626Z6iaPVbQksuAEI0dVQ2eV1PYKoV2igNvxYqHAWgrA3YfVnvDRjUJ9MOdS1c7QPHF2+qCCvq
KYQUB2eL5K9z40b8e3vA6nozU9B827lVAnBDn4dvrZ+aJe+ojxxMQsIideWOF8qAHEa6VvJA6hHQ
pL2YULcKLzs0rHv5mdsqwpQL4UEs1dfm6lNvbOP07xBn+ZvFpsH57yl9p3c6TXmHMHbNOfIQLBjs
10qy0qvrptUT35vGn9I1tTLo78l3oaTXWMv2zIbDiNxBODIU+YlAyujln/Bc0I6tXDRX6sDzSw6g
Enrqf5aoAe+E/O05q+cVPfXUCSyXG4OAUBvESyyHdB4+ecQ5fFrDC75biRiiQ/YC+bbWEST50b9q
RyQhzPTB1mKuwPbKxlMrSfTNxcLxzxVWJPAacvme14OPm+7WgXbkega3a1itDx+FToRo8amPpST5
C8cR+TN8YaZXfA2xy5sOfWeXUoOSmrRxjN3OJfF24OL6q1/9PQRWRF7CJsICjwLmqVV2OMb1Jc9a
ECREfByYZguVzvSJ5F9nL1/1IF0vlKbFmy1yTgoqVrDwTLqfYuc/Pe2boG8pEDiw17hz4R/o5kAt
my426+4NqWFMv3kRZJcTk+mj8l7N00zuVtbksZe/QZF55cr/1YcK+ioMiTMIBIkbysRoJZql1kYC
osjv3rYuu5AQ3MU/7PR+M1wxpddtTAaijXT8uVTVmQ86zt7xtYTbfj3aaz0ZP9scGn91Q7tgRaOp
2WQkHMieXImeKnQYGECM9RQvLYtoEJDaWYT27dILAMqmTzrlgm5sZeUk3dg78nYQZSg5VweKDcI7
sCpxA6cdgcY9VAAYW7ClYhQwO+Io9ArlDgZgrs9Hf67q+Z4rWm4qRoChZc7tBuN3s+Sb36lCD3EL
ySetGR9BgwNx5pA6Xlm4ow6VTUbXdV29zgL86RuU6sUln6b6tdfL2oDbwZfkFgfL8KGCtkbl+3ab
NBjaiK8mPtUYlQWf2ZxsNBzmfnAALTCB0WK49gWEKKAcWtfUZcj3Q54E53xV1oz9doQe8/xPoh5Y
2WqlDPvi+y+sN0v8Iestp+op23qe0RG2DWOzLyxCkIXl0DYmrafTPp2JnZ4aAM38PdvwpTQub3GF
O68eyUrd+6PBb0tM4xMTACNcV3BTxE6t0yujQdml0t1Duz0Ah6Rqk19EgFoLskRehoDyj0s1tM0d
Ob3VS5QtW8ENli/kTirHPsFIxZ0fivKUZrHcxUVqZMQUpqRw9lOs0pOQD/y5b0kfp6+kvaDsQKNb
kcSKAb9LweVQLI1i5cylmkURqsWwUQhn5W/X6uzk+WU1KPSBiLey0Vupul/xj/mWENGlWrXBFXlf
wBzyn1UejinDbK1iOKO1lzfzj1QyXhmZwuMI5GiUEV/eWz/wrbCdprx0V2CGD0w0BK8Xrfl7px1C
lP9lqos1b3niSDKj4RRA82qNZw4DgR8v1kQuNZcyB8AkayBbJFXrtz5bvc7me2VEiFVEYzh3uUK+
E5P2Ab6Rtfm9/zw6MeyEGnr9AUg6s5X8gHUJx1A/xVzJ/JMIWkMOW8agj5YhlfQmTuVClQ84otZ3
/OP6xTpk9wmVuX77YwgddaVkXSdD8MyAQnjh88OfIHy33akhbfYJikVR9Wtl7dxMu/c4SuHuJB5C
sTxnbqzjFB2eP3suydQoj0Hosm3HJBab7bRagb8TcBiYt6AMcModDuxFhGILJluqkEBNA0tFbVoK
qQSh4x5U7mqhm47hmG9Rx81TjmuF+GwQ6wCbtPgqgVbbKWMW9akU5JZl7S3dLOBVhLxkdHvrMJ5R
Z8VlB7DswORnjOg1VSdUwCgIQCYRqlnJOZSyIqa5JO8a3QBakdi2AapLt3xjUHjz2BDkJQ+gOW6S
VQdVkg1e8z5wEXOVf6K87Xuk82lvcNWWqRQc3P0A2Ratas0TUhBCTF3u4rf5wd0RIe09R1NDJgEe
HWn+lwkOYBFxnGFJi6EJu0JIRp4bGngyIgvJ7T4QjTTkcQqzA9AucdnMJYvMQYCjWGRo5fQ4nlfb
kysawdlKnsfGRo+ayn89Gp4ImHJgPyTI/Yc7IALy4k3AJ6m0apiu7FtS3MkCYoBE+yFd+mlzWgBb
ANDiqZ49P8ti5vxEnKf5/OJS8FcrKzXYzBCQFfc/4UExzZxSrTQ99SSl8JqpMOgAC+HkjYXjAdi+
vnxscxpGPayr2WFnqmmvZ3be8eyMhggPu7AcLX71CCF5StNPMHyMQbvIpcfu78F2tcbdY6FAZUOU
41V6ldbCsNYJcd7+DVx6f/RWDeCGXXlf4XfL/7cRov4qMxJabuQOig9C0xmhhi3BOuGDhXThbZaD
jZ9rIOYlQVIozdGb6JCE1Zdvp4y2TgNehrg6PFNPhLrVITspfJaGk6XMZaefJ03F6KK3N537/858
chmOi0cphAk5luKDbyJbGPpfxbL3HmwEaekZmFQ0/CTI5Yi3sv44VaNDM0lhTTOSzDZRcDTetjDd
JGDjL1GSL5ruhDzZg6DrkVjwBIdAff0hGalxiCUwA2p4bjcBrC0GHfMwjhJixtMx8PMEHmEXR5bV
E35tzB4KDzofDMZISAn/oko1GMnXrJv74lpNsyLT6Ug6hYbY7iq6JTiq2DJ4fnpPJEcTM1weIfDg
+bgM0z1V9x/CVjEfuVARlMi4wGMWyZCBJDN5ysXqlKtJIHGsalLPc9ZdGWeww956qq+iUmW+UDR0
LSTzMa72qnrNFrwZEVKKR27esoHZBtfI1bej8sH3EeGjLeYT48nPx63dhtKY1FpJudXNPdj14h3m
bxDqQlaJCrFNzJYi7yL72LYiXkFkqc1d3yf2MFfeLufwIfdF3VpEKutJ5X2Yhrt6JNRSWIOpEoXq
xLWSGISiEd9rIWwe8UKQZSZqFywGTPNjTu4rFcBLn82wFBm7NQVYT3u0LG22vJKSozP//kwpK1tM
8rYWXbebtmLMXXA6TDVwwN8DDKIwfc+H5VegKyFguVOu0GYbUWCuOTuV8YSvGkicwLnDT7jKEy6A
7jzVFWlbWs8o6ptoh+6XVdf47Syv71QmwDw5Q4MV3o5xUNM2R2ER51byYioO3EsnvoqqsX1EnKEs
cx5QTSgIdl8Gh1gpS+X11slMf39D3rQnnBj/GgbOhSh4lcHQoyBneG/97RSR2w2Tw9TTq48Gl/O4
GE411psB/8qMCV9C3j7ErsQSMdBupHgaUA3cYYICM4+p9D3JH4lbyBTDM/vILYBwkyj8G+zC2wu9
j/yBKH5wHMAWo4kyxxOs7Slgx+zQhUfcMq1LyU4uB0C2Yin0RQBkOoYLErZliThJqvygvoLGBwrc
R2EAU1goD3iYJZXrlb7/+WLq15CVcf/TwvYhVzuKbAICfjWLessgn51LrJ9mPx7OkK1Ix+OVrKXJ
qZzCrQiA/JsvX3mCpbw2aSc27tViD8av8Fq69SErtC3sglp4eB0OXMXVQ9Q5euSRWFpXvhYg/T4Z
f6GNCDu/P2wsc/1crOcEBtQrRfjftCBsvM4ykNJK0CFIrInkSF0EeJ+qP73OgzbjoU+eZ1fjW/kR
edNukA9om9WzjfIhjSVSt3OcOB4n0TBE+Sk1pqLV9kAEi2uRiSqnxcV24k5Yega7SIEa0VQvKakX
xEAhiqJ0+8KiQorL4Psj+VIcPMP+Bb9NofU2SVE8lAnSb0dVqkRERsRmxQt/xYudCgb4YKaatKQ2
L5aFonPcyMRl4s+Y0RdIXd07ilmA6iWag4G0KUTqe2HUOXPOxZpyoecitItPAgAerY3VoS3sjlEu
9t0cH9rV5iY9Wk3ZEka7zWfI0Gp6hjdCtNJ6gE+UfvaC9lnlx6K8WEuqTgFLlebhGkBPjiv+ZS5W
951lBsoP2VukYAje2QAMDO70PNrQb2dYgu6o5OsYRDZvA3i07Iy5P1BYOGIbyi9mDh9EoCRxm3Vp
D5VFVL3MxiZ5fRbxD0x1JUbbhJ737jWScbr9kkAJIyUMlKH/W1bmErds9lDubg31Utcfw3qhZZQZ
IW/J02NYkyHsf/vpJWy0GRzXGJjS8zJlEHaOctjb49o2dDxjtqhnGBrMV+5LtLOu7NIKIme66A/a
HiC8cKduYQ8BRLoyyJIvNdE8PQw4Oi9ShY8Oe7WeIQEgdfOIkqWAXuia5BDsh/n53ANUAeL2KjOj
lkjPjBZZqK3XcYIImEmmSV2PQ/nrbyFbFuX1eC0NihHJo0ZBXQhvLZpXmnPYefnO/arhvA2UEP+6
EL4/TXVGFsfqpwOGmuCt7UfKJYZr6U5durZVV5Ju3giDTXNLoO5HOTmli5KG2SRELMcueq7egKDn
r5bMdcO67yY73Xs0uA2RvRbdquqeyl9cIxp+33q6Nnka7sKI+WQcFq5NLduRK+bsrkDEzXmSAQ18
7mm6GSi5g3+H6lhD+O+FIeR8Wcs4Jbq+JhbS46dL8WWLA0R+eG1jA/aNYZVR4wIi0OBhGc16JkeK
zj8CY41YvH0bZVBHZ4aBg3dfFMGFFd2drnMGQM2j32FGcxVXCN8pEmEfPCYRAhaotRFYwWSwgiWd
iqaMjoksr0ybMAzQQrietBkLRr0X+WgXMR0j4FlaAMgvxIz5/Vr9NOX2Fh8nEJnW3vD6ydY/jfG6
HoK3DlT/YPsvfiqOa4cwMCroMeuU3ldVv1dQQAto3nI5SU1qbsscduUDvlcwJ6qcpg3Qof3hEKPd
qTZN9Wm86F3JGe/qTQZ613TxRwfdb6Od+LETD2HzGorYwaSczLUFw102gYxvex45Rh22z47a8SHn
TWDIRNAS1MvRu4tR5B73yFwmHufu+XnvpVHUBfnsNoiH8VcFxJ6/W3MGICFZBqqxSz2+5onazWvs
k2ptf7VUQbr8vq/OU+8vh8dvtPhSoOSxP5dduB/jdlYpqqm3gMF4Z3SeEdmxXH2ZFcTlriZBbzmm
ZGSEVHPqT6NEyNC1jtseXSym0MhvxpXzB3k/HyZ9DrmyXXQWwjotrKDR7R/j8mDoNvCIhgXZt3hj
LZCqAH0Baqsl0zTKYj+isHnC+VpknDeVUojlyFyvip5615J/ssAzS+mrNBI0xduI9Lj13XDuER+J
Tcrow797mV4QQxjgLJJzzdP7b/zj2j3xQWGFTbVS6l5GiAZMjoMaYE8RxET7emaUnJLuHf1PZ2TY
nQLHR0M+e4mt7heECBRXc/KOsxsAYVtvPl8pSKzWMwA6C+b2FHVtvbiejYlUZryWrAlNjjmPcccl
8m50zlmxBYO8lG9qo5qc+4QxZA4T5NGLtOc6SDyD/S3Qjbs7keLxU51PLyDLqTZey9I3JIosslE2
m1SYBJ1MgMT0+gOcl9vvnxgTJB8aQ3GOWNAjgEyxZGZ7appPoDh/TdjGIe7f4Wk1reCihDiTOMTq
UZqquI5UNGj4hR7Ivw2705iYye+I9sJjsRW/eFbQ3d6KzD7lH7vG2HiC50Mv74BX2L+b/K74HCrn
ifFkySGe9ywotN0qye8IkpEG3AP9ETxfPDbdTfct/3Spehhd6FwN6VpEXt05Rjuh5IJeInDSJGvh
L8uI4Lpoimls/Gum4a91FQq2jF0MQZ5WHMKL0jR6jBUeRspX1s+KTci7OTR4wfSVnkTtnMnrS53v
BzBKsjN1j7YyVwd1sg7QQhJBWbAPnxfKNQtIwuoYPsBtUbv5pz5odS3ElkUwYE0LLBqtB7E/zRdM
ua7AtHApnIwYbhB+v5vXtav02IDpi3sckoj8yeyHRXqQdPbkP/ozAf6B9hYf2/sDZZ6ggWPSjkNF
C2MIJaYnwgjA5lDxbnHg1jKuqRE53DrqQRpFAJWeIs1YhAisyxmpzNcjbm4/My3iguzYhz43xchl
0/Snm6+yQxiWxdSZAgdBW1Tw7ztBX1M1KggKYHp1A5O/lt7Mnc5V/sFddsY+T5/oY481o5cQ0hlS
YZDwRH1TkbaBZhbc7OOYr1io84824W3D5mLwxtJQiA0+HrahlzE4cQUYQ7p8F4Fp1ccW/zT31Ern
O/mtq+qpuFVrZomLBTenYhfcsSV/Noyw4oNBAbSjaQ1OlXYUEkLKWL/C+APOEY7d3kZwSmJtLSSd
bV+lFYrGQgwiaqdl+gNZh6bmV02Tq9ZTC3iKBOckvxF7J9TB/r0VanDTnPzSmb2wH0scTnyKu1C6
4/C64EsFFIXl019XQ3amIfWVSug5D4DB47MdOyOdIHM3t/zeOzAO7xeUpIIvKa8WrtbTe5BY5IZ2
GysY7bHWcI5z/edYPwloYB0rJzxhOoMI1llRNlLJ2hNLtsobU0ZSxOp7ltnqmBQdA9/NAnB8fRYR
jrJM5/zPb3fK7KMWUa0oMwBgh7QRq9LsKNsQV66T7QdpjMxEWglmyALMoqH/x8zm3x7R3Y0fmQnK
TITd9YC3RVGCx0VMsIYEpSKnSjPK9LAMo+ZidJCAA6cTZRP6CNlpfOZ7nqBkIR/hInWFgwD842BQ
qa+Mn9F/KeQm7Wqu6GK+wXm0dL/ZRcBfiyHycf3hpt/P/ZlZS/68irOuV8uYV+eRoX9xXzKIfNQx
SglDsWqwYjwOmtx8vhzK7iV9hI2sEh7IhQclXA+AvAN+/BjWMs5VQnuwGwBWTg6HkGJuMkr8z7tO
v++LyOiPWbv2+YNJoKldpCsFODaMUp7nyANvu/9PQ/VG7Es452THmxx/0XMUvhGtKk7vxhacDmrN
k/R7axnvWoE9DTGnjYTxI+PB9sZDpqdSXVd7C2WK+T2Zx+ZQ/yqMjru9t+rLlmJAfGaroGGtD6fv
qbaqjkmFzwTrQ/6BZyuSNgU9I24ERkh2Udn1uwTQmfykMsrLbiR7Z9W/KrYFkAvjjZJu9ujfPbfE
uhO2HpBX6vhV5UvXpGQU4fZMv1d4rZ6uxWCZ/Y3GhGSEfN6jlkRFsC5SI5EsguUA8SkLsmOCnzSZ
aml4inIfkfBfvZKH/0VnBU4AiZ00wzqYG/Q5yb+TPXPrNB0sYK3J2obBoDX6/t/wb/l6MLql2v4K
5P1HPCcHXseynIRt2x5CXWyV6IbcM8UKCPkq+HEWyEeYNiVKB20mzV6b8NK5JphfamMKswArTJNt
hG6GGtS10nqRsz37ocYW0aNELfh6OgxChB4AhaNr1Qrk/awamBOtjikd9DF1kgbvrDzwDG16vAsk
WreqzNo79uouQmjMpPK30QcadJFAlb0mnf3rqMz5bw4MyxyxuSzHGGfKB/B5OQkvMbsllJOTIAxw
zMrxgxoFcuqPjN/2AbFK5Z5xea4rGgkXAg27VZ6C7Sz91Ve6TaxGrkot7iPQUn657n1ODauqJcpl
zMx4lp+lpO2pCDmDe2hiUUwM3B76Jc+13mQbeEz8E4OKhdeBRA1WhAbpca5fXGaTI73sc1OOJEVQ
wSfWGr2QwtbJViQ/Ynxf87qLR2iDX7SxEGm2qR273WKTxkB7N/NsiUC6u7JfJmkeYhcDlS12dVh4
gb4oSbW1TwJAvAF73gQE97J/DDlmPepPrxjt1JSUgMq0HVC9bBuEOnGqEiDMwXT/nz8g5zN+fnZk
iS4rMFZxozQsMtsZhK/cRXTk71RTMp1JqlK7lWknTMp9o1eY69wgud7n16P6wBhV4BW5s6xbkc51
lG2Ko2/w309m8V7LMLPLCOO9wocmZFYziVQARG/bMnQ4OGYGrbCiPk8lcsi3n7V/41Jnbog79YBP
ta65rhFEMgPY6wSshBoXs55XhQB/vhi9+ZUO0TMdMpO3r2YptuThI+dHNN5pZpN7N4oOFTucvYI2
hRUJVV6v9bgnqPJPFlgiQsn/rMjvItPib73hFFXPpKkdtQtG6zrXYbO7pyHJ+roevcz3AvMTTGYm
jtsO6H/iYQkr59iYt2mqNsfEQXc2TVV0H1UEgkekINrvn+CBZrKEBx0E18K9qbKaQfviEFeZZgoE
iH4RLm0bwoItVMtoyUCv3D5w2zsw0lDZpDeU8jNUaWLNgxvM+8+f7wVCJq7BrCS+7DXRumpNtfzu
UjHIMtDN33ERJQDx9M8VgATF3U4K9ThuHb8uHXQqsA/XprG9BmoymoKC1r6BdmGAK+oJMVSu/sGB
mioftmouzYFKRB2Cns41OTUmgxSFDI1293rzged3DJqfrJeSOKiAwUzhcoLsaiNNIvmxCtmQyC6Y
A30yxC/gsEhsMI0eCkedRmbTFBZP2GwT8ebrm6uxcUPj6jS2+mkrJLIasZ665otHgEWXiwZqrXFD
8GnlxMtLnXV9K+lDtPN/yz0hi0j0yzyPJkl7NzzbO2JTu/iEnh+/7cowuvqvO6PCIPLiEoOz+eHn
p6uIICoVJK1A7jls4r1kFTarw8lbGf649OwVBAPtWXQ98XFaua1Uo9PQEgIF4/rMEInEbpiBS6TC
Ti/k0KaAfihhjx3jepUzKZpcIVJjLojIQbKmezxkPAJUXGFpIu6T7rmAn6ZR9vttHlsDzTthinC0
mZSS4doO+kYNcvXWFTRsuZ6hMjN3oWkOzIQH46BIYmOP19ytRNsUAXQs/ddpUjQNLtw6wIpup/mS
uRy7z+4XyQ5ouoBdgsSpB6KN4XmdYdzsJ9pTFjkkrqPSnj2MMjhhC7ThhOWJ9EnhcjcZ2HqU33Fx
q4rxe0z2T2nLYQhvl0MV77wsNxZleBMArEulqi6sP0ZGamUEClW4qcLuOpz8C1jcJVyTRc+9d5OA
9U42KoyuhaAn2Pj+XHWtfKt8DgB6114okmhqJhCQ6y20Qsw0syJS+xqad3mktJv2Pu0CFjsfcxvN
bFAi7qBZLVNpNq3XtCZjQv53a459GO1x9Q9JiX/MojuH/YP9OI/ypjsS0ehYWgRMJD7PtawuDdwz
7WrI3ydT1aWbx5iBVydNyh9lw026F6e8OvRVifldiugKJy/78GKDFedl9/5ii4es66fZlN06ZN8R
XN10y9I+nt9huQbb+LptolzfmL6p6g9pTIZrA92uhVEB96890eS1O/S20kWMasADF6Ahb5ZCX7nz
s3xJOOSnAzofDwMldciexRn/6PtpTgw00VCdo0P0kTBrP9IKtRcAW0WHuq1O8fwnhk0x6/tZFnme
YeNjJ8jkVr3LopPBjVYw/EfO7JJZNvQzP0Lap3MEt0gsFDsedJoUv27jTdfx7hgpyq9yipqxF9Bc
dUuGqYmC8fIaVhcuNxCdm2eL5KumXP9nTRTSXXq/dRNMaY2DZjbkY+6HHKt3mNReTRlOpwpOb5F9
H6NVpBk1Wu/ASv84SmBuHNC0kVUCDkLUg3Ujb4uVUYQEfQtzWqrPY/4I8DsSJg6d3QvYXbZra6Ep
2dUiZCwU662Z3wXlebg6sjnNpa4xsIwoorXqvUgAjjEWmJuzrM+Zd4blqcdkCYhI3Udb5G1ovEgP
SB/czIbJc1qdbo2yTc7UoS3CBfO3R0E+7c9Y/cPPCLTwLm73v3SpqlJymwiaALNuKZUNNTDq0qgV
7MOsyykmxQ4fWj6Q6ppvNE+qwADUqdid3LPykD6toCYt0YapRXcqVEocGgbZExEJflegRx8sH87L
QB2uwdpaDnMeF/X0qcB8a7TZvPXmBYDOKTxuPLOaQUMtm5XSZMwUwd4vuN5yMSsh3MAuAZ+ppL7g
Ikt41iTWKBPSfZ40wL5DvdKgzAUKJZpVWaySQyhXW1tgCb5ULPGrhO2jxVSXciYwhVWnbaz/646j
RoUtmpKcbd3xOC3V8N+tr3PKcMzN6MfNpWzSU2RTqMzyp5Uugx68qtqdHAlhyrBR495TJj2ryeEd
C7JLpFkMhDVhNXy+iIKedJGl2KCnxaDEbB/h/KlAIf8B+Q4LnqOo0Yt58hp/fQvkd8tamSbmJCcj
y5mo3ccoYG7Ck+iW/XgoqBkUbdSJIdluSo5eR1gsJZLGlA0ZZaLZ5BoVAU4NBujBx1+ude4YeNFH
+yFSQOBnYIrggcS9WeXOkckXPsCRnaNmFFG1tV8nnJ5z+aAuuOMugRZ7L73utgoSFN03ajd5vPVN
gbx4JhmyAIrd9etGfvOgEvDm/WAEgQdnSLAAppjmiKrEPQlAmh9A19UKs3z7WmUvxdfJQ/djwusf
7oTX9NfAFd77PBrWaMTqwL4BVbUBstZPRkMjHq6s0KW0H+YIqCfzyy/uAxctgKXWGXkuemsN/6Yh
YkvgehEUDpmjuIY86FDlcfw+POfeBYNfTf9e62uTlkBAwCTrNXnpMiJF/GEy5DhuSZM9j5gwDdWG
M19Eq9lnX+Zy5aa0MJo5u+zOxbquL6C5o6BgxO3VOI2wN7fQZCS74eBxkoExkPKQGezQ8tzS12pg
K0Eq0dscnU7Wf128cULT5Jm9NZSOO1X1kjutPe9mde5f6/cAUtOKNBpmC6VJbTcEptuyB1QJ/jOw
4AIuwJBZNA1ef8jGkg9jLxyCJX+uv9XA8TbVskp+73hcnMbS+n1cidcAY4LRxwer6k8gbwJn0UC5
5irwsOf5/BPuAPy4KyiZfGEbcpBxIMvb3vUtxx0Dn8G13FJxjEROxiLXfxxHDaAzThYMoSjDctJE
ymCqYrthbp4QobLEq++fMx+/ClXh6e3sgEuiaw12hXhCyFIlpJ8GniFozXeAfW9oVaYFu40QECB/
HjfKf25k8HUysI+41vzGhxqxX1z2j89G/bD6JsPvkbX//hjmjLYcVPPrork7YxqCCHUTaxvqizVn
cc+38Gjm73cYQCx5sM5074ekD6CyQoe/13Tr5WIOlMqp0DRjZUYRuqYrfEkWQmL9PQEgskghZWWm
9+MUMuuczZVI5un7YRu91BCsTohQneWLZ/fbEk4QcmPE41TUQf/zFhkKbuWV5RhNCuvI8Srswt2e
/gkr5A8FV+a9fX+RHVf+A/+fMjN0HmW4Zg2bz8q+y85hmRS5vWl4axbQmpBVkleH3Lf6QLlieyRp
Kas13ZXORglCFuwBprQoTatMHcuQSsoaOYq/4YUYtEGJ/Lgrdoxhs06PX3Ug/NfOyVQY+qO9Tb6W
1en6P5Y4GT9gS/wdYgyUlt9FHsY2MNzXNAommjZsMMb4CHvzEyr/AkrRw9VqWqghk1qbTvWA2SOh
/BnDq+DhxZgotWgF8Odk0VtYa/0hJIGoDIBNc4kZ5HXnt8uH26gWPuw/k8AJlg0YE7o5AD4Sz0iW
5M4M3E7Vzw4sMROgExlDlJmX+G98GtlUvMiAfEhQvkEjqUdAjM7m4TW0IKy2CjCB4bws9IDlsoTm
K/ivge+DEXEIPsrWwmlaHZJMbS9bpqqruCdzyCSwsY58+T1tob/Jgd/77A0Uz6BY+5PiTdR6W8oW
UjdEHouD6kgz2u65aQCp1vHmwHbjQHtIdC+glLifTUM4TJgFpATI5+lo1fIr0FyOazJiiKYGHdKh
0KwVbqVR7XM2B5CwNVb8cqbcrZnhsa9+KR/Ux9mk3gzYcPMAbXUx1i1rTBEco8efIJIa2F7Sql/J
d6vjq2R+f9gHq3xXgdcngh7LmxrSZfGLgR7L5zEcpCMVTRRmDW0evjWbnRg9Lm0h/1dJtSQ1KuGJ
U2ikVTyFrjzVRqXkRHRB1KOsA16K9V6IOWMQSXAIM5eG/jbsfboqKxskygvjR6BvhAUlxebRDvL9
HxMuMqh0NNLUKcmVakERi6hK/h6dMgLVmmFE4hJPADK7kysjY3Wam1d0oowVeMSPyMkFGFekM5nK
Ed6yhujLBekmLqTxUdXWDIHiiTJkDbdOJ4FL0MJD7CHLAYhBV93e+wnsRry3v+yQgLotYVGuCWK6
Xc9Cc2dmmbRjcDIpZQPMztDskD09REB2mkCGhYeBx4WtcNIjNYfC5QOvxQ72CRXtBG+9mznjt3/E
BmIYZS41z9IvhRePIpqjXAr8GWKUbOTrYp+kyccEjg3N+2tXq1uEnE263mwavmpAcbu8KwtaENqu
U5ssMT2rqhy2VMe1ezUzLK/zvniJIR4qHyQl5E6s4Rq4K8cxVhWKR1F46UB0ZahLyWimRfPDeHUl
OWVRZX/NX4Ec5xLVoCRDnZwaRQd8GU1sgjaLUO+3sz4vH7zZ+EELZhqXzzuxjQArJXGDzMBT9zk5
oeFj4m3ETRJkXZTHS8SUsSyaj9ArCzdVt9jN0f0w1xT7a11KoFArygnlIQs8X0ez+FBMbdaWQft4
s7UXIwJKW7NsQvGe+1g/Exg4f/atZjCcGDcTiskHsr8XNUPq//njB04ozQPLCSAtLjbqOhn3ua52
fh0iSFNl50TeRaeifzOyI9wPHKP1lJ9DEupjOz/SObAo5jOJEC7GfTdLCcUx1kY5lvhMhecic+7k
OolCHe6mSwAB+81LmkNs+OBqIT9LL5pddRDrouxRkeH66BQifjzWJDGGv2TaydaKaPV01cvuEjbq
ZjUCdo60v1lBgT/pGFhIc+RbnBzq4WGCUQAOFqPZuCxVur7huMEqRdCDFufBTTskBJQMCIpehbK1
5JBgiwSCQ0AO03ocSNirL6EzKCI6Mm0qlYygX3zSHL5bDUjiDZLoSC/1SanV4vvxz3mzT2DoWMJu
/jpkqo27VzswISAM3Dia/OUXNDHvmOCYjoGRzTqbOMkQd6R5qQ8g2YZAyN2dvXfh4HYQbGWXa4UC
3JhLjdcW9fKDCS9XVGYCK4cNJ8l1xsM3vvDFjCW9gPpyvZXdn9tEMQOIk0+FWkw4JiHD/vIZssjX
Xv94xEz0tE6gEKfrO9wRVFWyhb2pY2L73tJzcRHYY2jsoDC7Z0cRQqOwMkb4kL1Vl9IDvlxhG884
if9I3LLjYYsSNvhsJlJ8LYY2JR2rc3FsaPmlIG26ws9HkFKYnuzH75Bcz6TpLbRWLDc0PzE+HDsu
1TTJ9fPzpJrFQdma1jBDMRDpYWynJ0lMssT0UQqQ2y0i4zL5jMbERAR/F4RkgYyLqvGr1hcaG9w+
bnz4Z/rAzOAmEgW3fqpy2595H6qAdsyzxH4f2I9e/dCXTjMdaiPzC8xy/LIpjXv+axqf2EpHjTe6
k6Ls5aZpMHxGOsIXL6CRHv3/jj798dPlRF5UoOqEhKhQUj+Yd+kgFSf791xeqo8C5Dedsso1Xeed
rr68N91K2bmtUqpAbhzSWas4sqXTpayIqe6hWoIioZAV10JJ+PpSBsrXlR6dqO+Rws6FVHyV4H1h
8+TPvT14RIUFhDxZAeXOyk02Ublhh5gzJHoX1MwaihfoxpJP1WXxbz91AdfyfohK7IqLHcnp8zxQ
23hWTXTznIvfmD8dYCzjMF+kbmlKNv/srIdg9US30e9cdgUpgsImCt8Zml8qODk6d68tXTPfYm2K
asitstjuVcIfrFvifDSLioqDv46+Pld8IS9xnaDGLgOhrjwkfLQj5kYV676z1EXX1kVIHALhzDzW
KwHl0EvlpoNME7oQJCi5F5nuIlvc8ANVknQcxGvzvcaDujlslbUmK46RlxRwV8LEjvmUflQBeqgC
sPvo1dSgjtGI2OonqMzlsPlvfmA7pPcqQC5Ddpt9KV6dcZzjNHqAxrtQBkxynV8KuX2J/CUj+xp9
iliex1mxi+y9GsfzLn0kV9IvjXmn2xD/7C4Vo3BjUhkLjh6eCuIhuhIijXZcIpKBt8J/LUR1TEoM
ZXM+pqRpFBaPcks7PuiJYBlUrg7gmyGyv4a3ToevAtnCRzvkKgluVkwzzflmZieTCJeSMw82d0TM
A/VszNC8EBZjzy4UFjQbT5DzNs6XUcTcR5LSRu+Ky/mp4s2mvyyJZsmc2oO2FCIUjoQAsd1HhdsC
nKlJASar8B6FBxRatWyvAT4mm1F6pHSqIysRSbSYZz9hGj5W3H5LFH1TfCJyMoMQBp6aUVpwSWRK
dpgIxtvEhDZ7phkv+zdI+/HHG5T/s3nsYI+UQiEoJivtTpr3jc1udw6D77I9JF0wKQfyggYK1Sl8
8pxa8Y94uXMYE7+MFdOsMXzyEuzJEb+YuT2I2H6pdxxObFUrDZOdLKnSJ+asmsoM1twlZtb4K29P
fjFFYMsxVeUbYMVeflJqMHC/n3Bwm5HNvXea1iH6vShJ5BTz0O4BEkr4z9d0QOq6IqXUPQdUICue
Dpr45eKvRZz3fYM8fcCGUj0eFkvt1rZ7g/iBk9Ihju3HbBW69i/c3qOA/CzJksE3Sjvegfl/IJrw
oDsTuG70xCZr1IunoTAE8IvPlYifdU6OryHKg7KVdyi1kpjZPgJ8IsTJX2Dud1s6NoZ0Fk6Npxm4
6ILSaSBGLkThVTR4FhC3WC4VYV5qoEZVsw2dqUnmZEe+FhvN1jHE8/iqVlkvqgYCWx/qpcmFiWfX
PEai4nD3XrZiFWm2+MZROX2nXkG0dcoUgMRCDbNNDgQFpDG4ofwFUxTOUaNGr4g0QmqT2YpZ3wnM
J+JdG7FUcaxODlxl+hGfoJom+4lR9YgJYDGL191qmhiIG5oO/j6eTcLCVTaBPPb13UUWiUuSYOAi
`pragma protect end_protected
