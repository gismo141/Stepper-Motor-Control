// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ha7HtMch3G2Sn9jlfyvhrW/cZBqO132L0m1pOcTDJIaY/4Kw2OWipTSFIYHJ7ZcpiY1Vk5v7Ngdm
WAlWvOAGOryTTH2DeL7Ubu886Ad4CH7Hsnmsggb/Lq54RFzpI7rd6vt7JGFn2gdn7lK4vRu8YaaX
PoiGqoL+FXVi5Kqs7+923KR4Sp5HkSQczeIlQHZkkv0mZtY4RTx0KM7YlSDg6Gxh8QvR1nQHHfT0
GPKgPXvtRJqmUF7mCeyPCeOPY6vcxaZUq+IGOoEI4wQtkQRrcrorvtFl46OP6E5ZyCgFzAvo0ciZ
SV0JXzcmjvxysygu4Blspm0hA/I3JU0CLvWXVg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
HUBdyazvkpZ79spxP5fn6A/onqicfvU4Ka/r8mCjsdXY8XhncRzKZTdH5d2MOYy+R5MPSVcz6Ww3
z5wAZB4Li8tIHMdDc2o4I5bd28yX/iLemRYxYwIa6BiU0wVTYay5fUUwtTkXkgWdgGHYIv9NkdKc
a0ALNBnGapCtX88oQ0mwpafHbtDph5yehhAb2oJDz0N9c9dzWUX1DLur0JnROnK7j/6zXA4HGfd2
EWx6f6eirZd+npalIowINFPGjTHG70wWKdnV0jpTIRKcoMhdtiqQq/9Cdo2IwAcC9hkOXm0ElHHw
C6ZDutShl22E9MN3FqUXLz1fle0W8d/HRvBoci/pojiEFFS1EQo2gsaw1pjjOD+pwnLTL5Gmj2Dq
KnxNmQfckxQndsVAfD78wwl64mcBNmtIpygSv1REyI09+/qOrGLNqaJ/qyuxtCtUd9alCIrBz4L6
B5uDAn8NoG/VhPd8JW2gFNPLO+PyZISWd7hcrBJ66bHbhWxzKVp/hlHazh0sSK7PYdPKHOzMN3Oc
i/HPsWktBjtRYigri7PMt2yWBRS3gQHov/Qk9YDeBQqtWdldAPpYBjiI4m4/YivsQ/qZ8PJxNayp
PXcqfIlAidOR1Bs370tt4/CfOm/sulVAqWqJVTvXO/RbPsCSsSV4mILE9vQaZ0cdO404xdosyYdq
O8YVSWG88EbCp33UPaLuHMkg/9qyuUAWGMdz8OafdFIIqchbsmCjVgLIHKl+yq+9kMMxnb9Av5Tl
dderxllNHj8DVkdGBnUBmLyidOHpUqK8VkgcTReMhDY2LVNEh+VAC8Cl1hxHb9Kros4FRJMqirb4
YS0+LeP71IjkPjnot6gH50HoCqq/kfR+/a2g9CjEStk0TyM6FNooF3T+jZZq/S7dVpJ13daaAdMK
koqyEsCwJrLzmh1wc5PVB45GINBmY3EIa7OQ78qvjXkd7hIGvZLKAN41AkrRoCa7gsCAaro3EGKT
UzBEdwvHSqchJ2Q1YBWk5W1+b6hTNP5y4M75vNMHVS0LgLTyw631NZddXpLt8YtXmVNAS8iWw87K
1XVTdio4gVup+lcZP0i1fXqCYBLtTykTVDnju7EjQvTQVprRhVFRRksQ87lPJZ1TLfKMS4aQTztr
982X+k+7rl3RP7SnW5izGtXz2XfPaJreH5AERdjXu8tCvxEUbLC4ynOOqDPcxRtka0T7ngB7x9nD
tw5RoPTnqvNGNpgSYTjqXMfHJzNNeIsY+vRBEkwDa4he2ZcxqvNRdvUhGwXQwC3R0RpWYVqLK3Mt
DW/QOICAIPQFy+nyX9xcGPnod5s+1ZDMWsQqUKF8F11+0RPIUrBJ6fOGJY3DrhrMI8ACmS8NR0kL
P1WHiY8R0M1KRsfKPQDanEjOLMiz45kAZ3MmiUm/QW2biHOeeRFhAq8DAVFu+8cH0Vo0S96yKBws
L5vD8Z96ftYMry5egrR7jjxcRFamJ2wIVNWsKn6DuBNgp/4GdnhWM1xjvANTg9gdPz4jtJ3SyHor
sUUgjqOjGq+lA3RfTU/V5M1hiN2pEf3aHb372k+6XmMpWIZfYsJBoZzoxgln6kc9LgvxZKBvIv4J
oHRXAEn5qFCAjnqA1E/tx/ZejaXt7mwVXl2N2xSM2zGst3SB9ucnIF687WdbJUunqkf3THizb7WN
DL9dgLAc9uEbOus8MOEyIwfzWJ94pKy/bFnMJYxzq7fxX0xxuctHWf6VNVkveSbKdyJp3IUJoRjA
TIXCiehiouynlE7ipeDBTB+HEBVwrJpe5JuwT/SuCg9PukwutaBivmNEjUyCWMdmA1H32PdVJa3A
Agf766f7DJIXtIsiJoI5QkKP8CeUHKGhT9AJLPNm6Tg3V3oDXwenb3+BKHUYACL+nGJd58NF++B4
7W1tP6jN3F5P/UnmJ3VT1dTxyrfCpYFztRSN3BOSTT9N/c9il1faUoUSHD1BRrUfX+VSYFojlhoj
6dc3MgahujH6/Sk+Z4bsn5Kf1LSzhHc3qt/7yHFpsZUQMHkDzUwxwW66MvxMwFdk1w4eVVCwhFcQ
agCtIMfPW3g6k+1yrbFPdz0UwmWa28Cz35sWh8HBE94MbLafAgkrppxIrCh9j8natcTDwSAEoBUi
4eEob3g9QTdftGBpdmym4JJApl1pjAG/psYgr8LXhbFxIBIu546f8uOd0K9NJZeMbjmRGmTLkr4j
/7sj+g/VtDGtJ7qIqWlYizpmQFLMYd3gernhrMnPzWVESXUQtdbTUTCIbCiRE60/zkMh/0Co9n4R
hFLBvTc4pG8LREg1qI7dM2DGwgPpF3DYyKWOejaBmseFLKEKpf+6Z3dFbX9Ek0VR4MY2MQTviwOU
genMGsrBXzEHsj7i8uto5XMhb8LvfrEazt7tXuYBN5llIkGLdVHQeT40INJNMI4bmapDbTtXH571
YrO32VWYVvw4xVrabcX+e0Dbu48Unw1cnc0DNKXsm0TlnbwHq4HclHH8zWvEmPNB9iNeE+Q1h7Fr
qttOFLDH1C2ou0kDqB6C1uy75XjTM+Jr5HDhFhWkc4ltj+cEa7Vb7kID+TgNWdc4DsqvSbQ3AZI0
tR7XXAsLWAQDDInrK/i/wid1DB++oezOuXV2DN+WnmSlaqnW14vst7ZXrgIQ86gWaZbA7apa6+eC
7rXUQphKDrtIT6cNOSnG6YmdMuv8ooHMf1KD8PHlVedN5n420dZ5VenXHgcKYwqi9kwJW601F4my
EYW4pbJFvQc/8AtHVi+khpT8VZh7Klr56EaasVxuTYdNSVUVNbRmNdIbMAtc323rfSL4Qldc9OKy
l9N8Ps3PkH+QIfhfj+CUkC09ySLLtNl6vQiFlVyzqf6m+xa23UpoEyDYn89KHuTByfHPxr6vLz+f
90ysTYji52PVWA2BOjOxehpHFNbVtcaxzDS1SXGbwMW+2Ggr3+MbSY/2zetjohfEFsLxW/PByTW5
NJWgfYOM6ZZKeRZ7p5z6+Kbbw30jQGMNwMM1ShWPO17Gkg29f3Q9Vv1TsCJtwUBH2OazwV+/DL65
nILnjV9lfpchQt/F7wSGRcvi3f5fYbh2vv+Gkzy9C0VzQ4aw5O5gaVRMbdufD63cED8fYVK+rgbF
Lm9yYnwhuBLEaE0B3dR7tk0ZVeGf5abdX2aHRlNguyiLmepmX0XzN4duA8M6R+fRaOOK5Haup4rv
iXjAn/q+qOW0ASJWw3/GXiYFf+xqaMjm4Jj9oJp5FKTQwWkS5GgoVeBdeHz/Z3zaaRlKj2rz0ZW6
acHLTS4V7ePyUHi1PZbRTGxhlBArjaQJeMcC9tBHVXleNL4cgpo350QvHT5EorgnBe18K5YB+pko
UvTIZCSR/HmSxTsvNiLZdJhrTXmSVQDelTYoIrUo3nek9fPS15deWyvT5DmZOYsSfsKswAiRK1BK
mDI1aYFHnwGO58L4GOInYiZymeCWU4UJTqgCy66X39X/PeP5AdPNc17/1kjyF4i6D2Jj6yBqD7PX
47x9V4RsPNuLOuzssoMdFTB4QrT9+dMEQyv5XB6UaoXYTVfU3DQkOqKEDTVItVQqAlhs924Mzyt/
YzRc6PG+GznijQd2OAlNVIWOEU8AmRnXKqs/Dfh2PSTRB64VMp3WTqHYbp3LXPYjOLB4kZBBfMLn
43s9d/4HMSw/ZuBXm78BslJeL76wg8sOgQLq6DSOJpm2/axZWV5IuLwIXrs7l1Oa3CjISyxt3Wbt
ixAFLIcRY06Bv0MaVanrlUgnTG1Wupz8bblZyF0XhP1tv8X1hDUMX3IY0V6BqJ+FaNimxfeL0dXI
BTwaZ+azVKyubcZulZGK4TRcrgAVcV2J1Aj9jhL/94qWEo6mjAPyzQ77sNuQJpuhzbsleAQH5A59
J9YSvdH1JklIaB7TBCSZCSdaqcOm0EMhyAffsXScgmcGe8/k+y92CXKOAOiXTc7M2Yvm7prXWT6/
Pl1lan/IDI5d/O1mI6AHd83okWa4p+L5Tmcga5yhiReT1RTiBhjPvaW/C26ushJKh485iQ7TJuzj
AaR086OjRChzB3/hdY3C8WG29dMJIJchsdjsuq1+9pk/7dkUNhIv0XoaxuDr0qWHda/0zwOpOGMd
V3MUzbsQIpXLj7A9vx5kcfJiLEvvFpLn2I2uAMUmbeGfL1xDcWW9nvGHMp/dcWr7e+Uh7lie48Ut
JpBAUS2IFfTMG/0LS9DUwGUt2ar/tWVi2SS6yAjJKxG+fDKDqxTQEUwTfL8FrL5pEi5oMjtLZxZ9
yxHbelk0a30i6uZvuXhN3gd4gNV4kEY+glVVvgDclIFWfYuKP2D44bV/YjsvK3LTZiku7FY/sMPl
3vpPfH1Ebu63yHjDT+9VEGl3cISi8JYmaPaxDkt4ac3F9YrLHfzieWo87sztjQqeuHKPdYXp9zYN
tnFVOi4ZlddepXVT9c5tw0byvgz6Ru0rLdmwqJew4Z1rsBaQQ32arhfi2tIQBsjHDIkBKTsutsx7
3ofymFkb/oxK3AXX7Pnhwfo0AWC71wAC8Gt+XpTvhZ9ZHvWRJM6LuZDJXWg0owwDKr45TeOA+T2P
ItgOgDVCS8QjjYZ2+Tja+BeWqtT83OJNMY4q3QJINt5hlWrG1x+HXBA8wdvyc5R55bNfNlmuVkj1
0MIv85Xk5c5+V5+ljw2IhJLhX/12PQtsja0ac1Roc7Xmu6YKup997QZ7YmrHEUdL+/gdzZA9/izY
m8cJQr8RvxSJvxO1H8InCeFhGUZlZSL+CzgTDj74gXxz1d3vs6njKf18KtqksW+81ebYflAfdVOv
dEVmoHipB9AmPYlfH+dbnXBI8Ps+nS+fHC0ZIG6jhx+mC7wLdbPu1Uljrkxjy/SkOyR/aosLsFKo
FyIyljseMKIao3nJ3c4ijyfnRLqzAFRP1CsXbAZ2Lag3vWW7XeH1FWzq1UGF9ELowmFeY4SVI4yH
bp9xEjxQ++vZAlgZqBVgVYPdDmReu4xnVKvXjV2tHG3eNcHbfte+AhxOg5Q//BZ1PJANa/d/Nr00
IA919Bfqvs4qVIZUCagF34CmBGBsqK96sCIxR5fZH67T2khnayC7iipsDwjl4T4fY0tJnz+1bi8X
LZ9qoTIAfSQKYyvAFs8QQ8Qo26c5XJTBMiolbWrUanGrvpow3+efsM4zd0L4wFlaoMNUF4sWrVi2
veD1UtxtBSmLcuyWFqz9FbUbCsZY/4OUVAo+LR46F9krqJEmX/l9bU5ajTiOvXpurwoSqaZcjslc
9UmDedVZnF1WwqiRI8UTmApf/VfsxTfwRX1i81rt7FQD2TLIF/FOSXpuJySUJQ3RQY/i2F504c1V
m8vN1uMOD/OZ8uS4uSnXHlZNR5TsU5LmUCfpRpqT9fkSrL42CYwkO4lYHJw27xZHqGdNFdK+p9YX
X5ctAff2hT6zf0uYyL3x3rQnAHp7Sr9TwIoD2NVXYDAlcE2zMk9ShQvVjhmtNDM7GSZijLipFzPo
bm7XSW2dc0wtEZDu51QfauthceQI8Jl48c61+vx8FXeBNsh1G06bAbhdwbCAltu1wAy1I0MtKmlY
4m3EEpgkOo/uNmHxhOL1N+IYp8u+xAaCK0ON1RXHpbtii/LT7wC5JDc0s298rBU8d5iK3y4O3DQg
CEr2d//kur6nTxGujbAvr0Z3U3tYQ6CNJomLVbi5bP+dDlODHhg4WZeAJaTDuo6K6fXrvwoeKpYv
swQSoQTk6PUGWVYPEPMrNegCLT7iP04fIAHU5SzKNodGG3ari1RVDw2YHX0QBLhxRdX5+k/NG0BI
hFHWXE3KvqFPvKALOJNmw8GCE/B1E/W7Ba3l56duSmdoFYc2G++lItKXi2iAfvvsT8FAlnO4QlB5
I00kw4B3uv7STrMk9dMLtZds8tT4ueeNeoZnYn/pxVqAVE+vmE2BQW9fd3cxQRobkcxqhIY3IAWD
73pc7phQDNKhxWm7Ze1b9zYFrIL0LJTmZVezznVpBkr9PQGJ4QrZHCzCw7yw2SpzCpSt3F7NF/AD
gPf74YYpTN0fjTdpv9+rCuHaHucoh5Xb8Nc438F8gYul8wMdM8pQLhrySrv1hQ88xQPsJJuH4Bzp
C4X4wWGtQy/LSvQljW0kP2pv6/RpgvWKu2Jw6/U78kOvakJfvIe6gUZJ83jATbfSVsl9k8LYtocu
sPnzxexfvLQzgOmN1fQfFPebQNE6gRCiZOJdRzUKGlqcHlIzbQoZlElVIvlx96zft3n3ngisipZ1
+JT9/3l1WPVAA2r0KM0pkojl6ctT3iSPJfkERwC5aY/J4llrueVaclWeXDnyTFH/LxBJhm9QX/V+
iOl/bCcGmUoPIWNGlwSllzR4ilQbyfl5LzHVn7P7ohfITFMiX/uHuep7oVmoVGLBNDvH2M3g+w6D
wv9sVP6ilGyW9DxzXyRIpVQW/H8RiqdpsPHtDMHJ/RFNZRrs2rlpBlJ5YKeGtG+bkx1e8LsYHj7q
JnChnLx1XHr5j/+OJbl0WeFBVYPESekNo0I7VK2FkmeAWlh/Nm7i674BGvXckO5a+54jrvWE3k2T
ZVPGoA0YSwL37ZBpSuypfxmUWgDxDXSjjgEQpXrtlNdWI+uwx79PiV92TVPH1A/tiyK5XEAFDZDU
QvMpv4zk6Ck7YWaC+JnqVQk2t2RSesHvTA3hauXAEDj42emiGW91RY/gvXmnFmdGOwyec0Iqs8OU
I7BdTuumrPxahp2vRR9nA/1pULOeaHOfu1JcNqFig3qmECNeQR80anYX/N5CugWVUzJjiJDQN9Sj
29h8a8FdbvLajUhkxNigfVzvU6MXHAJvzQfT/v5gmZAQsw14ceLSacuIkBi+PZiosIKoH8ox+avO
zjLj5BtSh8/U+/qVm+uV7psjrp11RG+2wW3ppgc+FYVhAznZAcr6cYxgyrhecTSAose48HBleDug
KBAM+g5GJOYb1+bT23fk6KfPAWIf8dNSOcB1O3o9h5HmhqzLFolleoEmqT6ED08IdC/QNTN1BOCN
lOl7FAI1vwjQ1HdoHKuztierFfOy8tVoMR32/eogsof2qdOM8jj3OVFP+GB9kWMI7qBwlDWM/L6E
k0wuIfGdkEaL+oGUQKywXaJhICzKzHBGYzZf2zdEJQ+nmdZfezv6H//RYz5QPM59AhGccn/VIsVq
Uvhvv+X0Gb46Cw2aAIk+Edw2hPxH9tnn8OIMByeHeF8VtSZCGdYfbEO+Q5WXjDY2zI9RcQoit1ou
C7J73h29OVL8iGGAHvh476JKGu9C7MxP7HraOejiLUfbrYq/oL6s0aQ1GfISdod6wURn4RNyOkgZ
avZJsIpiJjoRKFY2QqiO1YjPzLJJo8/zt/fZBdcUhmQG1JVByFAv2/8sJH57tBx93mIJnCby3cpK
igK8OYyNN4oxwRZfkPhvexmm8YDGQzWrDpJOVJFTqSI06eJeZzmU8nelWZJmGsiy4m+LoMdbKlvD
nT0sdnL2rHWJZ4TPBO7Xs2YGymnfS/Q4Tr4Vc8LSEPq8ozpablOL868ArZh/fy+UBS7Ewyk7cZtr
wgDIblvqC0vPy8/I7F1dFvzfpMxz19UxQT8Jv7gLXzY/qqg6MompXUwn6MeOJXwIZGQY6Hz2u1Ji
mJjMwORaWR3cW6ndHM/J2V/RvUV2bMAPI9ybdxoZbvpWR78VUExtlKGJw9sYHJ4dJRz9mscVDqH3
E1ZMNZRPocqu4zF3zgq4PshQzjKG68KRefnqM51v0lLqQZJYsEw+7cSgOHlyEjXbJrvidaY1HHdG
fiaDnpyXz+tz53Sbq9o8Bn3+a553SH9hF2KvykS+H+U/8G9GO6FgUIR6aQu80bOaf++VcU3RqLtS
K50PIEnD8QLOsY/QMVwIo5EjOlXFfByXW7ty5PyqxOLHmp2l4LUB7jCeuNPoXIqfTfInbPp0SzDk
h68y+B+2V1Fx1WVmbItXodGtFE4WyavKRITE0XOfMlianhIkd/1KmV+0I67RldmO120/OVT+3nFU
BVgNp1Tzky5m2ToyO152tx7M8k0KCvx7Lh6kxV0S5+RI6lHoFTFWaMsAdrB0C4ieZ/UAymjEbNVb
OHOBX8KXsRlOTrKJLlULYxv3MNQ7rgfcVUh1HgOcPbn7MtSX1T+z28ADUTCcrjWzBwaewN+MhktV
U9hZbSxqs5hQqVvQrPoEqrMCq6Z6lRRiO+UOgr4v6mVqP9vV8g/NVlq15fMnhQHneLkVP9G7x7ke
pYVjMEF8kalxTI5OzEBB6+13NFNKtvzyPjWTsIM2j4tyOndPA/Y74tqMXKkSCav6xcJWi8iDEpHQ
FSb+hjbsAZW2mvA/l8znR8quQKz679LuR49Ar1DNCNR/BLbhgCf/xC0eknY+G59RUVLIdkF+hDZ2
YVnyJCQLQORc0QP8K8q93UAe//gO6qrQWswEVp+OLqh85Y1qfiTIFhGylqrtR655fXqxVWJGl3dM
8hseSB3gCMDgY4gRMfp4XbNtH38CnLE02s8TuTQoAxzXqc07HaegdyTNXQ3bNnjMuo2oh3u/w93Q
/zkgCC91a0onjuv3NRHYWI4Sy0GaT4k0V96GALKG0/nQDPXnfo19/KUIgKf/w056X1mLicPWMwfO
I1AG/UDVBu/cFTDqhVDKJObzYwHDck53jN079oTHhj/b+Q4CTCy5NckXqHTtj0o9eVK2wUfbRqru
4BuOdG8USJQmA20q06QDWUsBU4KkzjaiZZAyKwFmjk7x713VNXRYzU1SzeLTo0oxZAEREDQ7I2Ps
DT31r9JBFmYK3h2stLBF1HjH/CRe8m77i8DNbQQiXCb/Bw2JMNHQlq9IqszF0hjpnM7lF+btAO65
Hueq4tVVK2XAj8H4yh9d5seArpXUUl9EU4ssLWsTfxtYS0YfUvaUB3YdPsDA/xbTbPhAi68Tep/P
KADgw7mMEihfAt/BU3crgvAHOghDtB8Q7Dwo1kO9ealrQ1nVjU5zXBJ86S7yxySQDgBtJB9nVPqq
UiJSvC9khFvLpkLm5t+fEdhwuMkSTDbZAD+MtppKQffw0SEH5dx4AUf5vYNKL5mjht2YjbLjoBVQ
4F+rz+uLw9Yxf4QRMqtVvFSTpwH4n5g4jnfID6Zt6K2p39m6TXpavYT1Lv2+UMHoNP3WsxRo9oDk
wWDo68khSs7VAo5GdpnTAZOqTS4lLj4iz8sgtUSZCyMdcRGpRO8SbL8CyP9TGPjhovbi9Nto5SpI
47vzzJ1WOvcSSa6x2Tl2TOZXch7exnOew+xkhkxlhp+a1p6nfDE5Pft62Ko4osjM9+YI8vqX6woO
ECJFlQCsI/Ej4BjFDSl+j1vt8BFI2tekXH9iKhqBALN4gKG5EoqbBaZSF+h/75RHkxnsJnmipOEw
kVq5qkJEel4O9TeJyNO94HfawX2LMjd38mEmCnMlc9+Ot1QF7+LVbsHwNMG3SMPzg+rkzT5H417X
uSl1TacRTotEIigM/qMxV/1Gh8oJJrXan7Zmx3UHQO77DnggXwBerQx6VRZl+YK38Ade4VVUWTQv
p2X0Auqw5Wru+8nlg4nNOn7xP5xCr+cWR4QZft7Yu65Rv2UV7eTaUZToE91u+Tk4UyKGTvcqVrL3
0a3BAk++2ayYXiAlEsLJqruRMpEwIJRYKjBxa4KXyn5VLBKlii8Lg8oHLGOQVI54lymGlerhPHiC
ZLIg+5MixY/ByseSwVIRoJmt0Iz0jwitboShH3T+lhwhnLk2kLCd9QFBSGfuVSxXzD5BGUFaOVyg
gkRSw++JDUzcN2oCxCxDrN4M+2KGWgAyFeNYZ/0f61IZeAupkYqowExdARw7NfQmBywgqlq5F+K/
yAFLkjcWNNw5vCgc/Ze+/p/KJKt+8+Z85xmF/9D6LGYBOv7OAJvxdrjmnaHzusoyOtFgOsXX53N+
NFxweSK69a5YGUStYH9W11QagNbLH5GdvuPyIJaqJ0mx744pOQGmxtATapsmU/Hh943TBScz2CI0
aTh7FOl+Kqmnkq1KDfNErXGVKUP4PdfeWuIcEIcZUlrbiXNioQo+31Bi5U3Ltha+7klpc2q8jJeR
fs020UUA39bK2Ml0/4cam8XTyv7xlXiK83VM3BxfWSH5dtpqrC1PodN7dVVlbYvDTVz8FyxXFfqg
/L4qayWik6+uSnoz2tlAaBhCNR43NcoJQ80jej8BqpWIbYyMKxmQ2grs/k3BK1FRq5iYH1ftcm/d
jzY599zO39GGjuxrJKZI+hOGJKG60rya3H1JIkBxK963GCXCJDQu5dxHUgg4DCqmKhm10IHuuosW
kpvHJbEFNNzzEhma7cqv1UFPC3LNENQRREG40VVQR2Z3FMtsDbuXjc1G9DK+d1G0PhkmzGFQSVsZ
p5ircQHJHxvxaWaBpVgAwsc/g96j+jKn3hfgBuRiZu3px+v0Xiff35+UU3JoGwjzAWMdHMsW/dUA
Q1L9qVOwinCKf4GjcPQ8jhseaNC7evdXdhdlkBGweQ1W/F0D6lVDFxW84u4TqNcxcfZZ8UWCYKA4
vQS/yiWdqVB20UmODJyZmI6Qpqatu5r6fZd1HPgY6CDR+muzFEL4yegfPmRj/ZvbMIYPIIE8B0gR
Zzl5KoBY3ryOaS3LdTUedJJLcn0ntNw+tr8idFuVLvx6z2yUrSbv8n0j8jAhQrFNF7a2peaeQic8
/lLT36KNeKmijxB+b9pXZkqWjdD2eCj7f0CuE2LskTvSJKR0
`pragma protect end_protected
