// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:02 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZR3ik0g6fp3Aq8oeZZbEFk6eb41BsF4AO0s22sli4VGJ5FCA8bV24/mMXtCn3uM/
FkrfVSUCSUnYY8LFTPxiznUYwSJfH3SIE0Mn2Qf8EywgQENSGDmdjOsA6cw1b+wM
2Iu+J6Mjs49Ei9B+krWRxWVGy44bmOsCCyLLL8kl3uY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
ft/Ze+SMBKhzoBOpRKDGfZv0HZthrDbvc83+cwxSETY1ipyvUAHIn7HISeSO2AJk
9dg5TK9bnTwJJA2rOFYQEm5hihbgpcMUmoSXT9pgylXygSfWGAydBcTuukJM49MY
svhgl0xZ+L6Sxo7ADYQViPm+BudWilpZWthhZvkNzObclgIk87uG1hRyGW8vntef
yPTTOuMu97V7OfttHD9BfkyBzYIp3wHwt1YbO/cKRdY43s6UVzA+dYviGLDLuZuk
jMcDWy5JNhgph9/mIazV8b0UROzx0Z5E6oB/Nj/8+5tENro+UwRIAX6an//QGngc
W7zpycWqzmfZ7jSXP7RKQE6i20E2EUN8pbJC+DTaMnQPfqicwe0xK5miXfATxjXB
uvcE0taJJcfYnGWRQFsoOMuxS98D/P+O+bebQsjVu+C53c1hbMDSVC6V+jA+NL7C
t+yUsxwTPYOxguPtv+T2Jlj47UJp5i47suKBmTI042nQgKED6mnyZBmfWh070WME
iLUSHL8vXFk0AKRO19PfL3A5qDFusGDYi1qz5qCEp7D9knrKLNkSP1iTV7WsEyOf
DHMNwSv+GUF6dDQMa/ITgQx5wSq5VbBr77evUq0AEZT/zHcFMqgA/7nvJNwVRlT3
oJ7qtcO/WwAr2u6fg4rM9kk5knwz4JXDI7IolMk7JEB8geBwqtvqUx+4vbW7bIXJ
f6HeFQmrz6JwFHDIaKK0e/lbQ4T/Qpkk3/+g2FfWkiBgQjHMMlOvYQvA58RFm7E/
APcXkH8nMhCKiW63ftGYuNFJBUsZEPGINUmO67ue++UA7/9MOXt22rvz4jfkLE/M
ARW8OjA2pDqygK6Q4ekHGRSYKE7C20uwc+6HDlpsl7tU4GtX+dCofpCEq5shQMQz
fyUCKT08dXjEldPQC1nfRje+3NZdu2uBhom6FPGc/Xc0ZpnQjGOoC7QP8MViRLA0
WF8Z8Gu1uECmL9nkRMBOMItunYwpYD0GF6UDEoB9opCv4Lg6Wfs/zrCfnWLMAQad
1BppCn5bG4IKDB1koQbBBfdfnLXGsCIAVQdIMh9DPm6Beu5PsdE6J/owBEgu73Bq
UH9x0HEyyvKdSZWu81v4oea2MIOcTqCJ07EJOg0HhnqFw9TIC0yw3A0G0p2xK+/D
C0ipvekeXWRG18AG2Ryi6FOEoSDwtg+0V6G0dmruJamVATA0rgVlnlmaZSPcpNlm
b8NE7anWlUFala7N8LaAo9lgUxDcf9FXaDffrmy+TBXLlipBQUXA5xEXbyYJGm9V
TL4kcMN8D16NE3Bw13i+a9AtGF9kHGwOS8RS5F1bKpaBvOpTMwlEAdd6NxqymfPG
Rlmn2YxUcXaU8KgUOgBvTUwaNWet4VEs4k7DbeeprF9X8kfH25oofHNc0JgII3Zd
25wIOh63njO3LJXQi0KigkG7wou/pTVybPki6h9CakFnl/y2Kg5lGZvrQBBguNM5
YCi6u8lHnaimq67un8t2lVNhVbTat78coMUQPkXN2XLMLJRBWUdU2w6lIv2UC5U2
uYHYfaDri0h5ejoP1MdAv2zPuMhiErS4wLCMDed+TO8+VsKsJeLYuU8FHGutGE8J
D3xZmmzPsTWbvfSgS2QuE5pGgzvRKXIp+CCIx6fKhzSZix1I/tuTSn9l9A7nqhOk
dST4pH+iFojuelkppIvszkyy+kSS7jy5oPfu+hmYy5bqPM9sW919PbmCuqotrxP1
gG17b1+Bz6J6/aw1pY9N2/kg/r62OhAyHvdw9FsmG7F/Lhw9TCpm1fZiUZxCiQaa
PdSCgbw3h5CMeH8+E9gjj7rDvT8sByD2fi41Evtl3rMkBuIB3j5RGUwSizH0C9S8
7rnINLV7HDo8URlRbmgGAEYw8BuTppl3TMZVSWaGwZI1hDkHMPDT5mG8X4pzDSBp
SUc/7hs6z06MiGHqBl4TZ/qvvRZWVOdq/VI+TUSrhpzKNdUxawyvD4rXyR8koEe9
mK+YvagmuK/+HKDtcs9DVZRvWEhn87rX+nHYSfoJQgL+otjFr5pyX46M5PkP+qJT
l+189O/9jrn4X3G1OWUwRgsgOTx458ZlpUiohAC8q4wJ6v+f6dYF7iHcD5rcYLXY
XVtd6Z2NscMmkGSp7UWtmx7CpHNxYV6nJ3JVqd1KtKYFy0RvX14Avgiu/kLfsezF
EuZcgCk7yniKa7hrO0Q8bAkLDcyx8T2/1wFW1VpIO8C8m7SmqZ9Cy2QGkAJ0Zp/J
eUctFfIspu0r7Vq9XGgA+WFj91hd85QYnux0wQ1BmmB5v+oKnBemBrDFxGACqpeh
7QEMZhY+o7Sq4R4KXQAn1+oww4qtJ8leybUaVyvDIoeZGqF8VgAzp7K3F+BGO04J
ri+bksllUkdf7zoPwMRnEB1N1YGtzDR8qWb/+N9mp2uPgGiaQiOEBg//9do4IlxQ
3UiS1Jn31xQ9lLCJ6KXahXTSJpJbvj5PsgG5oYoI07LInmVg2liVTK+Xb9fpVMRD
MLWYpwbHO66hQLsA+XCCQnPWonPLP9irVLi2UfMbNbnsJWNuPMKtouRbFHo4L3ML
WCZjjcQ2uRVszEM/z58AXvR4QMrzCmQPuVyFMBU26mJj670DSBh2Ach7nbheFL8g
btbYF8TK4LBqCuK5qRQijQ/pJmHydykY6gMeM++BSwMmXZiRKGeMPbLSQ+ipfSWu
5ozJGuGx8XVhNW0ec1Zm4oEW0y8+jDFzO+1lB2HiI7CxiFkkxE1u8R/swfyy7A0u
1cmKMY7XuYIGx9B3r2Hg8DUrOv67QrLYngeXGWELwa4xsk8uGHTVyQly+zJ0SgLH
OC4cu7IKNeJHtIn2S+WPxJcPrpyqlMO77RYPt8c3pKtMM5WE5CN4M9gRqRoaIs7u
B/5BfLD2K6sjF1Bs2IrO7P/VuEeqWxwRBZu/AyWdF9354s2V0tPfIuQXZvJUaDB2
DDB+2Nd7kqi0bDnY7X2yWlkSUKHlWiv/Pv9SfSJqsUtqyfgxHG+Bvvv1K4KqZufl
aGbYxPrqGTQXIntxrdaD1pHAn0+Q55b2VdAgfeFBYF6tDelBW8AnMLhXTxbOKWFF
SjCSbWtwdwM8lfPGTG5G5b0c2mi7Ipb31MgdQJmAryQ9MvquLutTSJ3ZuCr7chHh
dV9rmiNPMhkjPAnZd6hA2dG8AiI0JW+5cpgSXC9hpQO7gfPdiIV+0byakPA2LRX+
eu+4oEtMD6eAS0RUV+xbo53q6pIZuvz7fjFEzWpQkqIEvZJhtpXf1BDqFOYk9MAp
LFBPAvZ3oZxkEzyc8f+FsiuqIk1qm66f4fBbwCXbV7vRQbwYE3LAcdlLr7srRA1d
wcoz3p8CkXvVxrUJY8MujdKAWeFv0PvPOSOXmikH8ZULhBQUwCRbXaFl2Dl6a4et
nZVegEP553nradY6XMuv4Yp8Rqg4VIlaksr1U9HPgFPwJdzrbGjafM4PLzieictb
NH+UDTwDrhd//f076r6uLrDEh8sPQhxHr6qP/ebHbiyOgH57+giQ2Fbk2FpUpR9V
ZA3zqG1AAbGJfR4pb6jRsDmA4addPRHkh3ZCfl2YHp+rGUQmCzF07qXDNua1KKOs
D9XryXGvvBiJrEbTPfSv+53tzqt/zEGUs0xREMAdD+S2ZKnQi6/AlszztepqCTb3
HzlAF3WG6t7BgaHB4aDgzsAnx21dd4dANO26NrEtUe16xQej694n5V/95Kb2DsqN
LgEMmnOz9HX9c1JxIn1il6VFgutb4YJEWNYN1bLILR3qGJyahPDzLO+NsZ/rIaT5
etXxB6IPV1BZQfGhRjbMkQTJ3nH4L99P4naI09cRjYan9hXmT/eWqhkyEWvRx7dv
OAbU8BT4iY6t4G512j+swD6reAmVKfZq5L1z3GU2Ua8ZIMz+kZhY2vcb0Fw7qE5k
EbJSxTLz7YWC0UiMhM8WXRH2E2SYvQovsr4xTnLqC2HlgLX+g4ym6pGydJG+0Dli
fmfBHzmFgxU1sJFLXkk1zWfwuiBRpx6xfTUrXHxZkHNWVU0bkqlWD3YmVapND+TJ
aKLBvd88VLP3m3RcbxwrPGoLqaGvgfTU+oqV70JmU6mmtKFBn+cD/WwxmTjy4xhV
lX/dgrTHx/6woP/1n6ljujxZa5gKNQ+2+Xk2S/kvY2VNs2dVUXwGSv2iHrmwU8Qb
Zpm31bfJSjG7B5fkurpBPBfF+TImUTfymMbBkzAIqqc/TEIKc7N4HCuu9iUjTVMN
4Obsy/tpY6eNM+1HrPfs2bQA/hQDa2ed/hThw21KL+czEtFKutb2kxvEFQfuFywf
dv3HQjgW9CKuEUulcKamqtJtVzSTy49l/kbyO6sBIspz2SKmMgG/mD8TfJmYldOl
3cARxZEMWx1HkSGNq/jEhpKJ39Ys44Y7p89YJRgfcb04Fgu0YErleR5fFGvccIYc
LUTjxdTgnb2QRcbzUHjdmdvYlAX2Gyv4rI/D9kakkRnbjWBq5ut8375VXLOPQZHb
hpM2VQxi/FYIQQ26ZtyBzVITlDuTjx+VrTXg40CKpExVcPYzRA0OtE896jqhkd31
Cmq9yjy8BAASa1lJlUZafjwGK4cfeJxBAbLRNABfxFvaXpJYFQn3IvkyAz5x3xHk
1FEJm/Lmc+W4c8i/rJoUiyEWlUY71vsl7ni5+9L7HQruuzMHehzRk/IlExqv2aE3
oDZi3Ruzyz9fHAA3JTBhkoaqcrYf95NnWy2rQ7Gp9ilVMg0IbFr/tWnjwkJioEbV
XZtgbimyLZY2mCKkFGUr5Y1TkYfGCOa3xyG01w/WRrwuVYfHzSm/YEWi8ddJkpov
+5ptmUZFJjrfO6qQJXZZaAYC5mMOh/rpkt/7q8zEv5eAwm6I0GrehgJcVUwf3RqR
FIb+IOvjiXbUFtgSKULXBoAwG2Dm44Y4PXV8Q562DrF2p8YQEcyZDSQ0TikMGEQX
7V7kF+gLbewMbpPvB/AxUUtVdCyL5844UYVuRiQ3Gm8eqE3ZVJfFMNrGU3ZTTS7P
A3Jr+kHN9+ZHHZckzLKL2ReOI9+x5NpOhbWIJbs9jGKaJd/YBsKTj1IxVWurQLeP
xfy8XY0rijGlxx69mCggZ/qlvaedkpWs64dWh8OtvzMlybqD4ebEMqv15PGSykpY
Z9jvjtlFuUpMLRirUdEddd1fmwEttvSsvbuusLOBK+1yXE8naGVFABiLrCW8R/xf
hadi0oGRsWaEF6ZmTIQPupLlrtyWcj6266GPZmsoXGhgz+WhgWP2Wk6Xfzi7bZ+k
bXW4A/Sis1k/j8aG24bLRqCB6KcBBcCndb735Rr/3PUyNb/qzaoMLs3lPacfXo/D
5h8TCFB8wvByg2BDuIlbIytVqkVWJrUjauj9nITk7qNTxh6hKGj25s6Na7eN/sli
u00luNd93Nixucx+bdimOe+nda6O99nyZ016//cWm6OQAaxmFa5+juAQUdQBzNHn
J/s8fz+NA8OYXaX68BTOgiYdeUThkNgdQxCT5OxKdYTp7Y9L+XwuW3PnHEh2X1wT
H9tFZdenqaiJc8Mhx3ADQ1XKO036NempebZsCv0yctri1VkBFNnIleAqkpOdLYN/
66oaZ5znuPAUD++BkR8y1w1xP1J5l5XcRFWqDejOmOPxxHvX4NY8aKuPXvwACAd7
5R0E6QoLVPKiuByYnU1uS0h/oxEdC51d5nT1If5eFnTLGsiUSx/c07E+PBs5qpui
x1OP1OjCm7+teYzvJZHPlELU2YOxS2E6AckWszhob1krHER5/SFT1Sv8vdngy/xF
A09fpFkJndwca4NJq9P4KaYK/Ngq7bniFlbt+Xr75zHrr+0BRhs1VcEutIBgCHB3
bSnawYIIT5UC5MfHPQjNiOUba0OCxtvSOao11FOD1npp2i9vcbO7PAquk23U7JwT
r7OzrKnmfSmh06drkBzd7V5qJx8iMjExVYqyezmU6PqIPIbIF3F+UDA5AKcNSARp
gphgzSNjvAHMMOvr63WLwGqPGf5H5uhElDhoKkn5dkrQ70cu/YpmB+IOao71RNWQ
6I33VXAkc1ylog95T6ncgne3ZV+4J5PTwQefD7kupE58EbKHzEQB2z7KZj3yIkL3
LuMaWSMf/LvUSRYvInzT6/d9ZYx5F7copXDD+FXxYPlryRotGhBs+57QsDyX1lvf
6UL1e7mNGH58tvaEWFSZivBSRRNtFdWd0Ib2J9oEiks1vWSVKlPkyDReeZBN277w
z67EFyNHyceOfnz3pYQOm6jxvxtDV0I0Aof9MjJ/x4+asoPjI0/cPMCEBRDbZ7b6
dEOGneSus+K4oTk0HC52blXikEwtTXv3/KGN1qHUqCeR24+YwIAoSCAxQZkp61+T
j46swvyidV2nEQW3kos/OoS3q35q9582WzoZn0oc3ovoHGjJ10kp/rPYNv6IcXqX
pRTbXvpGk4HDlIUdRKDBQGvwhvjViv1s8cmK3eDpG+82ojLEWJBgGDB8TPE2lMH2
bMTamhwvCZB/DjP8wIkgiQNMiriDdOdNKUk2jSLkN0AhLyeBZmb8AlpRzWF7qYcA
hVpaRZFwoBHAlahQH+5mNoYXJhDrt7nvHEiZ61WShD3k3H0YCDNDgSCP4Y22cfdC
L0eL1sTS9bcnVRpOl4nrFLTirioEgnla9YwOigJkOHSd+6pPQ82ZqjZhCY2oe1BA
EKNfHBBwwWzV4EJn/u85rwZo+b1sfGLtR2akl1+VhiYq2IMTaXhlImm/8YQcB3A7
/CIKtOrxHPU94cQPWBQ98agFiVJ54BUtMaXfqOpYiO64TK+XqjIWYcOJg6RrtAMW
fK6urhGdX781hnQuLxh7AChaP5VvmXbSrxN4+2jzGLyiuVHoRl04foGOap8Q9D/7
qRM/10GS2ODyykjarbKcGXISL7u2zb0zVVCE4Nmm3KqqWUazYUHRSV3CU8YfCLK/
kjcZ8dy7C6tAp2+IgMwDeS/9/BIRrUuPhUJ7GNDFhlgDJs0wXfhw6X7lp5ff6MgR
ZrVgRMLXtFBtn+Nx3odVrYXbsb6wP5KvV0vFtS3ng1fnHZa8OK0S8/lq6EtuZaYS
wcXrQcsbEuDVig4FVRqytYIoFJm/oEokZXSQ5hXrIo+y1mAhRA3iVQBJ11jbWlR+
gSNC4PRP9tb+syUGkoh9KPKBMWUImXSncpcwzvmP+vMpJBx2tWc4ZNZyvn4OOSGH
luyZEXTXPujSkjJY9vVIxkBwG5rBbjuEC+fe40EjI9UgUHQ0lr01HFDlC5+OeCRy
5VIgjHCTHsBkH8i+W/8SiCKa2DB0skC4ATPifA0VQDLQ2SfijyeBbRpNrzgyJI5p
agDmjkq+gZNZbrkt6tOuTqmpEyl4RfnxFOwqMwLQ1voXzAP3AykHgKo/0uZ0+/Pw
ssAxVux/0anuebAnncdQorEOMgqH+v3h7WUBaYALNm9FPJqXIdXkv5kO6fJBW62M
weXek+mc+SVVHHaCLCnET1J/B0FMtJA+vyEqKy4HhPCLB2307oEXbTZmxXmGjLiu
l8YhZY6O6/vKOwRBH/IwYU9qfrFnVE4lILwLaYmEFp0vW9OjPC4G4+MYPPw+ag5s
CQANo6dCgysa/CkWpDsV2TQCRZ0D39HPy9ft06/YdEI=
`pragma protect end_protected
