-- StepperMotorControl.vhd

-- Generated using ACDS version 14.0 200 at 2014.10.27.23:20:06

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity StepperMotorControl is
	port (
		reset_reset_n  : in    std_logic                     := '0';             -- reset.reset_n
		clk_clk        : in    std_logic                     := '0';             --   clk.clk
		SRAM_OE_N 		: out   std_logic_vector(0 downto 0);                     --  sram.SRAM_OE_N
		SRAM_CE_N 		: out   std_logic_vector(0 downto 0);                     --      .SRAM_CE_N
		SRAM_BE_N 		: out   std_logic_vector(1 downto 0);                     --      .SRAM_BE_N
		SRAM_D    		: inout std_logic_vector(15 downto 0) := (others => '0'); --      .SRAM_D
		SRAM_A    		: out   std_logic_vector(17 downto 0);                    --      .SRAM_A
		SRAM_WE_N 		: out   std_logic_vector(0 downto 0);                     --      .SRAM_WE_N
		SW      			: in    std_logic_vector(8 downto 0)  := (others => '0'); --    sw.export
		LCD_RS         : out   std_logic;                                        --   lcd.RS
		LCD_RW         : out   std_logic;                                        --      .RW
		LCD_DQ         : inout std_logic_vector(7 downto 0)  := (others => '0'); --      .data
		LCD_E          : out   std_logic;                                        --      .E
		KEY     : in    std_logic_vector(2 downto 0)  := (others => '0'); --   key.export
		HEX0    : out   std_logic_vector(6 downto 0);                     --  hex0.export
		HEX1    : out   std_logic_vector(6 downto 0);                     --  hex1.export
		HEX2    : out   std_logic_vector(6 downto 0);                     --  hex2.export
		HEX3    : out   std_logic_vector(6 downto 0);                     --  hex3.export
		LED9    : out   std_logic                                         --  led9.export
	);
end entity StepperMotorControl;

architecture rtl of StepperMotorControl is
	component StepperMotorControl_CPU is
		port (
			clk                                   : in  std_logic                     := 'X';             -- clk
			reset_n                               : in  std_logic                     := 'X';             -- reset_n
			reset_req                             : in  std_logic                     := 'X';             -- reset_req
			d_address                             : out std_logic_vector(20 downto 0);                    -- address
			d_byteenable                          : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                                : out std_logic;                                        -- read
			d_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_write                               : out std_logic;                                        -- write
			d_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_debug_module_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                             : out std_logic_vector(20 downto 0);                    -- address
			i_read                                : out std_logic;                                        -- read
			i_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                         : in  std_logic                     := 'X';             -- waitrequest
			d_irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			jtag_debug_module_resetrequest        : out std_logic;                                        -- reset
			jtag_debug_module_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			jtag_debug_module_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			jtag_debug_module_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			jtag_debug_module_read                : in  std_logic                     := 'X';             -- read
			jtag_debug_module_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			jtag_debug_module_waitrequest         : out std_logic;                                        -- waitrequest
			jtag_debug_module_write               : in  std_logic                     := 'X';             -- write
			jtag_debug_module_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			no_ci_readra                          : out std_logic                                         -- readra
		);
	end component StepperMotorControl_CPU;

	component StepperMotorControl_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component StepperMotorControl_sysid_qsys_0;

	component StepperMotorControl_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component StepperMotorControl_jtag_uart;

	component StepperMotorControl_RTX_Timer is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component StepperMotorControl_RTX_Timer;

	component StepperMotorControl_SRAM_CVGX is
		generic (
			TCM_ADDRESS_W                  : integer := 30;
			TCM_DATA_W                     : integer := 32;
			TCM_BYTEENABLE_W               : integer := 4;
			TCM_READ_WAIT                  : integer := 1;
			TCM_WRITE_WAIT                 : integer := 0;
			TCM_SETUP_WAIT                 : integer := 0;
			TCM_DATA_HOLD                  : integer := 0;
			TCM_TURNAROUND_TIME            : integer := 2;
			TCM_TIMING_UNITS               : integer := 1;
			TCM_READLATENCY                : integer := 2;
			TCM_SYMBOLS_PER_WORD           : integer := 4;
			USE_READDATA                   : integer := 1;
			USE_WRITEDATA                  : integer := 1;
			USE_READ                       : integer := 1;
			USE_WRITE                      : integer := 1;
			USE_BYTEENABLE                 : integer := 1;
			USE_CHIPSELECT                 : integer := 0;
			USE_LOCK                       : integer := 0;
			USE_ADDRESS                    : integer := 1;
			USE_WAITREQUEST                : integer := 0;
			USE_WRITEBYTEENABLE            : integer := 0;
			USE_OUTPUTENABLE               : integer := 0;
			USE_RESETREQUEST               : integer := 0;
			USE_IRQ                        : integer := 0;
			USE_RESET_OUTPUT               : integer := 0;
			ACTIVE_LOW_READ                : integer := 0;
			ACTIVE_LOW_LOCK                : integer := 0;
			ACTIVE_LOW_WRITE               : integer := 0;
			ACTIVE_LOW_CHIPSELECT          : integer := 0;
			ACTIVE_LOW_BYTEENABLE          : integer := 0;
			ACTIVE_LOW_OUTPUTENABLE        : integer := 0;
			ACTIVE_LOW_WRITEBYTEENABLE     : integer := 0;
			ACTIVE_LOW_WAITREQUEST         : integer := 0;
			ACTIVE_LOW_BEGINTRANSFER       : integer := 0;
			CHIPSELECT_THROUGH_READLATENCY : integer := 0
		);
		port (
			clk_clk                : in  std_logic                     := 'X';             -- clk
			reset_reset            : in  std_logic                     := 'X';             -- reset
			uas_address            : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address
			uas_burstcount         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- burstcount
			uas_read               : in  std_logic                     := 'X';             -- read
			uas_write              : in  std_logic                     := 'X';             -- write
			uas_waitrequest        : out std_logic;                                        -- waitrequest
			uas_readdatavalid      : out std_logic;                                        -- readdatavalid
			uas_byteenable         : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable
			uas_readdata           : out std_logic_vector(15 downto 0);                    -- readdata
			uas_writedata          : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			uas_lock               : in  std_logic                     := 'X';             -- lock
			uas_debugaccess        : in  std_logic                     := 'X';             -- debugaccess
			tcm_write_n_out        : out std_logic;                                        -- write_n_out
			tcm_chipselect_n_out   : out std_logic;                                        -- chipselect_n_out
			tcm_outputenable_n_out : out std_logic;                                        -- outputenable_n_out
			tcm_request            : out std_logic;                                        -- request
			tcm_grant              : in  std_logic                     := 'X';             -- grant
			tcm_address_out        : out std_logic_vector(18 downto 0);                    -- address_out
			tcm_byteenable_n_out   : out std_logic_vector(1 downto 0);                     -- byteenable_n_out
			tcm_data_out           : out std_logic_vector(15 downto 0);                    -- data_out
			tcm_data_outen         : out std_logic;                                        -- data_outen
			tcm_data_in            : in  std_logic_vector(15 downto 0) := (others => 'X')  -- data_in
		);
	end component StepperMotorControl_SRAM_CVGX;

	component StepperMotorControl_SRAM_Conduit is
		port (
			clk              : in    std_logic                     := 'X';             -- clk
			reset            : in    std_logic                     := 'X';             -- reset
			request          : in    std_logic                     := 'X';             -- request
			grant            : out   std_logic;                                        -- grant
			tcs_SRAM_OE_N    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- SRAM_OE_N_out
			tcs_SRAM_CE_N    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- SRAM_CE_N_out
			tcs_SRAM_BE_N    : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- SRAM_BE_N_out
			tcs_SRAM_D       : in    std_logic_vector(15 downto 0) := (others => 'X'); -- SRAM_D_out
			tcs_SRAM_D_outen : in    std_logic                     := 'X';             -- SRAM_D_outen
			tcs_SRAM_D_in    : out   std_logic_vector(15 downto 0);                    -- SRAM_D_in
			tcs_SRAM_A       : in    std_logic_vector(17 downto 0) := (others => 'X'); -- SRAM_A_out
			tcs_SRAM_WE_N    : in    std_logic_vector(0 downto 0)  := (others => 'X'); -- SRAM_WE_N_out
			SRAM_OE_N        : out   std_logic_vector(0 downto 0);                     -- SRAM_OE_N
			SRAM_CE_N        : out   std_logic_vector(0 downto 0);                     -- SRAM_CE_N
			SRAM_BE_N        : out   std_logic_vector(1 downto 0);                     -- SRAM_BE_N
			SRAM_D           : inout std_logic_vector(15 downto 0) := (others => 'X'); -- SRAM_D
			SRAM_A           : out   std_logic_vector(17 downto 0);                    -- SRAM_A
			SRAM_WE_N        : out   std_logic_vector(0 downto 0)                      -- SRAM_WE_N
		);
	end component StepperMotorControl_SRAM_Conduit;

	component StepperMotorControl_pll_100MHz is
		port (
			refclk   : in  std_logic := 'X'; -- clk
			rst      : in  std_logic := 'X'; -- reset
			outclk_0 : out std_logic;        -- clk
			locked   : out std_logic         -- export
		);
	end component StepperMotorControl_pll_100MHz;

	component StepperMotorControl_SRAM_PinSharer is
		port (
			clk_clk                 : in  std_logic                     := 'X';             -- clk
			reset_reset             : in  std_logic                     := 'X';             -- reset
			request                 : out std_logic;                                        -- request
			grant                   : in  std_logic                     := 'X';             -- grant
			SRAM_A                  : out std_logic_vector(17 downto 0);                    -- SRAM_A_out
			SRAM_OE_N               : out std_logic_vector(0 downto 0);                     -- SRAM_OE_N_out
			SRAM_BE_N               : out std_logic_vector(1 downto 0);                     -- SRAM_BE_N_out
			SRAM_WE_N               : out std_logic_vector(0 downto 0);                     -- SRAM_WE_N_out
			SRAM_D                  : out std_logic_vector(15 downto 0);                    -- SRAM_D_out
			SRAM_D_in               : in  std_logic_vector(15 downto 0) := (others => 'X'); -- SRAM_D_in
			SRAM_D_outen            : out std_logic;                                        -- SRAM_D_outen
			SRAM_CE_N               : out std_logic_vector(0 downto 0);                     -- SRAM_CE_N_out
			tcs0_request            : in  std_logic                     := 'X';             -- request
			tcs0_grant              : out std_logic;                                        -- grant
			tcs0_address_out        : in  std_logic_vector(18 downto 0) := (others => 'X'); -- address_out
			tcs0_outputenable_n_out : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- outputenable_n_out
			tcs0_byteenable_n_out   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n_out
			tcs0_write_n_out        : in  std_logic_vector(0 downto 0)  := (others => 'X'); -- write_n_out
			tcs0_data_out           : in  std_logic_vector(15 downto 0) := (others => 'X'); -- data_out
			tcs0_data_in            : out std_logic_vector(15 downto 0);                    -- data_in
			tcs0_data_outen         : in  std_logic                     := 'X';             -- data_outen
			tcs0_chipselect_n_out   : in  std_logic_vector(0 downto 0)  := (others => 'X')  -- chipselect_n_out
		);
	end component StepperMotorControl_SRAM_PinSharer;

	component StepperMotorControl_lcd is
		port (
			reset_n       : in    std_logic                    := 'X';             -- reset_n
			clk           : in    std_logic                    := 'X';             -- clk
			begintransfer : in    std_logic                    := 'X';             -- begintransfer
			read          : in    std_logic                    := 'X';             -- read
			write         : in    std_logic                    := 'X';             -- write
			readdata      : out   std_logic_vector(7 downto 0);                    -- readdata
			writedata     : in    std_logic_vector(7 downto 0) := (others => 'X'); -- writedata
			address       : in    std_logic_vector(1 downto 0) := (others => 'X'); -- address
			LCD_RS        : out   std_logic;                                       -- export
			LCD_RW        : out   std_logic;                                       -- export
			lcd_data      : inout std_logic_vector(7 downto 0) := (others => 'X'); -- export
			LCD_E         : out   std_logic                                        -- export
		);
	end component StepperMotorControl_lcd;

	component StepperMotorControl_pio_sw is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component StepperMotorControl_pio_sw;

	component StepperMotorControl_pio_key is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			in_port    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			irq        : out std_logic                                         -- irq
		);
	end component StepperMotorControl_pio_key;

	component StepperMotorControl_pio_hex0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(6 downto 0)                      -- export
		);
	end component StepperMotorControl_pio_hex0;

	component StepperMotorControl_pio_led9 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component StepperMotorControl_pio_led9;

	component StepperMotorControl_mm_interconnect_0 is
		port (
			pll_100MHz_outclk0_clk                  : in  std_logic                     := 'X';             -- clk
			CPU_reset_n_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			CPU_data_master_address                 : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			CPU_data_master_waitrequest             : out std_logic;                                        -- waitrequest
			CPU_data_master_byteenable              : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			CPU_data_master_read                    : in  std_logic                     := 'X';             -- read
			CPU_data_master_readdata                : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_data_master_write                   : in  std_logic                     := 'X';             -- write
			CPU_data_master_writedata               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			CPU_data_master_debugaccess             : in  std_logic                     := 'X';             -- debugaccess
			CPU_instruction_master_address          : in  std_logic_vector(20 downto 0) := (others => 'X'); -- address
			CPU_instruction_master_waitrequest      : out std_logic;                                        -- waitrequest
			CPU_instruction_master_read             : in  std_logic                     := 'X';             -- read
			CPU_instruction_master_readdata         : out std_logic_vector(31 downto 0);                    -- readdata
			CPU_jtag_debug_module_address           : out std_logic_vector(8 downto 0);                     -- address
			CPU_jtag_debug_module_write             : out std_logic;                                        -- write
			CPU_jtag_debug_module_read              : out std_logic;                                        -- read
			CPU_jtag_debug_module_readdata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			CPU_jtag_debug_module_writedata         : out std_logic_vector(31 downto 0);                    -- writedata
			CPU_jtag_debug_module_byteenable        : out std_logic_vector(3 downto 0);                     -- byteenable
			CPU_jtag_debug_module_waitrequest       : in  std_logic                     := 'X';             -- waitrequest
			CPU_jtag_debug_module_debugaccess       : out std_logic;                                        -- debugaccess
			jtag_uart_avalon_jtag_slave_address     : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write       : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read        : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata   : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  : out std_logic;                                        -- chipselect
			lcd_control_slave_address               : out std_logic_vector(1 downto 0);                     -- address
			lcd_control_slave_write                 : out std_logic;                                        -- write
			lcd_control_slave_read                  : out std_logic;                                        -- read
			lcd_control_slave_readdata              : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- readdata
			lcd_control_slave_writedata             : out std_logic_vector(7 downto 0);                     -- writedata
			lcd_control_slave_begintransfer         : out std_logic;                                        -- begintransfer
			pio_hex0_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			pio_hex0_s1_write                       : out std_logic;                                        -- write
			pio_hex0_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_hex0_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_hex0_s1_chipselect                  : out std_logic;                                        -- chipselect
			pio_hex1_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			pio_hex1_s1_write                       : out std_logic;                                        -- write
			pio_hex1_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_hex1_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_hex1_s1_chipselect                  : out std_logic;                                        -- chipselect
			pio_hex2_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			pio_hex2_s1_write                       : out std_logic;                                        -- write
			pio_hex2_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_hex2_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_hex2_s1_chipselect                  : out std_logic;                                        -- chipselect
			pio_hex3_s1_address                     : out std_logic_vector(2 downto 0);                     -- address
			pio_hex3_s1_write                       : out std_logic;                                        -- write
			pio_hex3_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_hex3_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_hex3_s1_chipselect                  : out std_logic;                                        -- chipselect
			pio_key_s1_address                      : out std_logic_vector(1 downto 0);                     -- address
			pio_key_s1_write                        : out std_logic;                                        -- write
			pio_key_s1_readdata                     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_key_s1_writedata                    : out std_logic_vector(31 downto 0);                    -- writedata
			pio_key_s1_chipselect                   : out std_logic;                                        -- chipselect
			pio_led9_s1_address                     : out std_logic_vector(1 downto 0);                     -- address
			pio_led9_s1_write                       : out std_logic;                                        -- write
			pio_led9_s1_readdata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_led9_s1_writedata                   : out std_logic_vector(31 downto 0);                    -- writedata
			pio_led9_s1_chipselect                  : out std_logic;                                        -- chipselect
			pio_sw_s1_address                       : out std_logic_vector(2 downto 0);                     -- address
			pio_sw_s1_write                         : out std_logic;                                        -- write
			pio_sw_s1_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_sw_s1_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			pio_sw_s1_chipselect                    : out std_logic;                                        -- chipselect
			RTX_Timer_s1_address                    : out std_logic_vector(2 downto 0);                     -- address
			RTX_Timer_s1_write                      : out std_logic;                                        -- write
			RTX_Timer_s1_readdata                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			RTX_Timer_s1_writedata                  : out std_logic_vector(15 downto 0);                    -- writedata
			RTX_Timer_s1_chipselect                 : out std_logic;                                        -- chipselect
			SRAM_CVGX_uas_address                   : out std_logic_vector(18 downto 0);                    -- address
			SRAM_CVGX_uas_write                     : out std_logic;                                        -- write
			SRAM_CVGX_uas_read                      : out std_logic;                                        -- read
			SRAM_CVGX_uas_readdata                  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			SRAM_CVGX_uas_writedata                 : out std_logic_vector(15 downto 0);                    -- writedata
			SRAM_CVGX_uas_burstcount                : out std_logic_vector(1 downto 0);                     -- burstcount
			SRAM_CVGX_uas_byteenable                : out std_logic_vector(1 downto 0);                     -- byteenable
			SRAM_CVGX_uas_readdatavalid             : in  std_logic                     := 'X';             -- readdatavalid
			SRAM_CVGX_uas_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			SRAM_CVGX_uas_lock                      : out std_logic;                                        -- lock
			SRAM_CVGX_uas_debugaccess               : out std_logic;                                        -- debugaccess
			sysid_qsys_0_control_slave_address      : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata     : in  std_logic_vector(31 downto 0) := (others => 'X')  -- readdata
		);
	end component StepperMotorControl_mm_interconnect_0;

	component StepperMotorControl_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			receiver3_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component StepperMotorControl_irq_mapper;

	component steppermotorcontrol_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component steppermotorcontrol_rst_controller;

	component steppermotorcontrol_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset
			reset_in1      : in  std_logic := 'X'; -- reset
			clk            : in  std_logic := 'X'; -- clk
			reset_out      : out std_logic;        -- reset
			reset_req      : out std_logic;        -- reset_req
			reset_req_in0  : in  std_logic := 'X'; -- reset_req
			reset_req_in1  : in  std_logic := 'X'; -- reset_req
			reset_in2      : in  std_logic := 'X'; -- reset
			reset_req_in2  : in  std_logic := 'X'; -- reset_req
			reset_in3      : in  std_logic := 'X'; -- reset
			reset_req_in3  : in  std_logic := 'X'; -- reset_req
			reset_in4      : in  std_logic := 'X'; -- reset
			reset_req_in4  : in  std_logic := 'X'; -- reset_req
			reset_in5      : in  std_logic := 'X'; -- reset
			reset_req_in5  : in  std_logic := 'X'; -- reset_req
			reset_in6      : in  std_logic := 'X'; -- reset
			reset_req_in6  : in  std_logic := 'X'; -- reset_req
			reset_in7      : in  std_logic := 'X'; -- reset
			reset_req_in7  : in  std_logic := 'X'; -- reset_req
			reset_in8      : in  std_logic := 'X'; -- reset
			reset_req_in8  : in  std_logic := 'X'; -- reset_req
			reset_in9      : in  std_logic := 'X'; -- reset
			reset_req_in9  : in  std_logic := 'X'; -- reset_req
			reset_in10     : in  std_logic := 'X'; -- reset
			reset_req_in10 : in  std_logic := 'X'; -- reset_req
			reset_in11     : in  std_logic := 'X'; -- reset
			reset_req_in11 : in  std_logic := 'X'; -- reset_req
			reset_in12     : in  std_logic := 'X'; -- reset
			reset_req_in12 : in  std_logic := 'X'; -- reset_req
			reset_in13     : in  std_logic := 'X'; -- reset
			reset_req_in13 : in  std_logic := 'X'; -- reset_req
			reset_in14     : in  std_logic := 'X'; -- reset
			reset_req_in14 : in  std_logic := 'X'; -- reset_req
			reset_in15     : in  std_logic := 'X'; -- reset
			reset_req_in15 : in  std_logic := 'X'  -- reset_req
		);
	end component steppermotorcontrol_rst_controller_001;

	signal sram_cvgx_tcm_chipselect_n_out                                : std_logic;                     -- SRAM_CVGX:tcm_chipselect_n_out -> SRAM_PinSharer:tcs0_chipselect_n_out
	signal sram_cvgx_tcm_grant                                           : std_logic;                     -- SRAM_PinSharer:tcs0_grant -> SRAM_CVGX:tcm_grant
	signal sram_cvgx_tcm_data_outen                                      : std_logic;                     -- SRAM_CVGX:tcm_data_outen -> SRAM_PinSharer:tcs0_data_outen
	signal sram_cvgx_tcm_outputenable_n_out                              : std_logic;                     -- SRAM_CVGX:tcm_outputenable_n_out -> SRAM_PinSharer:tcs0_outputenable_n_out
	signal sram_cvgx_tcm_request                                         : std_logic;                     -- SRAM_CVGX:tcm_request -> SRAM_PinSharer:tcs0_request
	signal sram_cvgx_tcm_data_out                                        : std_logic_vector(15 downto 0); -- SRAM_CVGX:tcm_data_out -> SRAM_PinSharer:tcs0_data_out
	signal sram_cvgx_tcm_write_n_out                                     : std_logic;                     -- SRAM_CVGX:tcm_write_n_out -> SRAM_PinSharer:tcs0_write_n_out
	signal sram_cvgx_tcm_address_out                                     : std_logic_vector(18 downto 0); -- SRAM_CVGX:tcm_address_out -> SRAM_PinSharer:tcs0_address_out
	signal sram_cvgx_tcm_data_in                                         : std_logic_vector(15 downto 0); -- SRAM_PinSharer:tcs0_data_in -> SRAM_CVGX:tcm_data_in
	signal sram_cvgx_tcm_byteenable_n_out                                : std_logic_vector(1 downto 0);  -- SRAM_CVGX:tcm_byteenable_n_out -> SRAM_PinSharer:tcs0_byteenable_n_out
	signal sram_pinsharer_tcm_sram_be_n_out                              : std_logic_vector(1 downto 0);  -- SRAM_PinSharer:SRAM_BE_N -> SRAM_Conduit:tcs_SRAM_BE_N
	signal sram_pinsharer_tcm_grant                                      : std_logic;                     -- SRAM_Conduit:grant -> SRAM_PinSharer:grant
	signal sram_pinsharer_tcm_request                                    : std_logic;                     -- SRAM_PinSharer:request -> SRAM_Conduit:request
	signal sram_pinsharer_tcm_sram_d_outen                               : std_logic;                     -- SRAM_PinSharer:SRAM_D_outen -> SRAM_Conduit:tcs_SRAM_D_outen
	signal sram_pinsharer_tcm_sram_ce_n_out                              : std_logic_vector(0 downto 0);  -- SRAM_PinSharer:SRAM_CE_N -> SRAM_Conduit:tcs_SRAM_CE_N
	signal sram_pinsharer_tcm_sram_d_in                                  : std_logic_vector(15 downto 0); -- SRAM_Conduit:tcs_SRAM_D_in -> SRAM_PinSharer:SRAM_D_in
	signal sram_pinsharer_tcm_sram_d_out                                 : std_logic_vector(15 downto 0); -- SRAM_PinSharer:SRAM_D -> SRAM_Conduit:tcs_SRAM_D
	signal sram_pinsharer_tcm_sram_a_out                                 : std_logic_vector(17 downto 0); -- SRAM_PinSharer:SRAM_A -> SRAM_Conduit:tcs_SRAM_A
	signal sram_pinsharer_tcm_sram_we_n_out                              : std_logic_vector(0 downto 0);  -- SRAM_PinSharer:SRAM_WE_N -> SRAM_Conduit:tcs_SRAM_WE_N
	signal sram_pinsharer_tcm_sram_oe_n_out                              : std_logic_vector(0 downto 0);  -- SRAM_PinSharer:SRAM_OE_N -> SRAM_Conduit:tcs_SRAM_OE_N
	signal pll_100mhz_outclk0_clk                                        : std_logic;                     -- pll_100MHz:outclk_0 -> [CPU:clk, RTX_Timer:clk, SRAM_CVGX:clk_clk, SRAM_Conduit:clk, SRAM_PinSharer:clk_clk, irq_mapper:clk, jtag_uart:clk, lcd:clk, mm_interconnect_0:pll_100MHz_outclk0_clk, pio_hex0:clk, pio_hex1:clk, pio_hex2:clk, pio_hex3:clk, pio_key:clk, pio_led9:clk, pio_sw:clk, rst_controller:clk, sysid_qsys_0:clock]
	signal cpu_instruction_master_waitrequest                            : std_logic;                     -- mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	signal cpu_instruction_master_address                                : std_logic_vector(20 downto 0); -- CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	signal cpu_instruction_master_read                                   : std_logic;                     -- CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	signal cpu_instruction_master_readdata                               : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	signal cpu_data_master_waitrequest                                   : std_logic;                     -- mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	signal cpu_data_master_writedata                                     : std_logic_vector(31 downto 0); -- CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	signal cpu_data_master_address                                       : std_logic_vector(20 downto 0); -- CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	signal cpu_data_master_write                                         : std_logic;                     -- CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	signal cpu_data_master_read                                          : std_logic;                     -- CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	signal cpu_data_master_readdata                                      : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	signal cpu_data_master_debugaccess                                   : std_logic;                     -- CPU:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	signal cpu_data_master_byteenable                                    : std_logic_vector(3 downto 0);  -- CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	signal mm_interconnect_0_cpu_jtag_debug_module_waitrequest           : std_logic;                     -- CPU:jtag_debug_module_waitrequest -> mm_interconnect_0:CPU_jtag_debug_module_waitrequest
	signal mm_interconnect_0_cpu_jtag_debug_module_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:CPU_jtag_debug_module_writedata -> CPU:jtag_debug_module_writedata
	signal mm_interconnect_0_cpu_jtag_debug_module_address               : std_logic_vector(8 downto 0);  -- mm_interconnect_0:CPU_jtag_debug_module_address -> CPU:jtag_debug_module_address
	signal mm_interconnect_0_cpu_jtag_debug_module_write                 : std_logic;                     -- mm_interconnect_0:CPU_jtag_debug_module_write -> CPU:jtag_debug_module_write
	signal mm_interconnect_0_cpu_jtag_debug_module_read                  : std_logic;                     -- mm_interconnect_0:CPU_jtag_debug_module_read -> CPU:jtag_debug_module_read
	signal mm_interconnect_0_cpu_jtag_debug_module_readdata              : std_logic_vector(31 downto 0); -- CPU:jtag_debug_module_readdata -> mm_interconnect_0:CPU_jtag_debug_module_readdata
	signal mm_interconnect_0_cpu_jtag_debug_module_debugaccess           : std_logic;                     -- mm_interconnect_0:CPU_jtag_debug_module_debugaccess -> CPU:jtag_debug_module_debugaccess
	signal mm_interconnect_0_cpu_jtag_debug_module_byteenable            : std_logic_vector(3 downto 0);  -- mm_interconnect_0:CPU_jtag_debug_module_byteenable -> CPU:jtag_debug_module_byteenable
	signal mm_interconnect_0_sram_cvgx_uas_waitrequest                   : std_logic;                     -- SRAM_CVGX:uas_waitrequest -> mm_interconnect_0:SRAM_CVGX_uas_waitrequest
	signal mm_interconnect_0_sram_cvgx_uas_burstcount                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SRAM_CVGX_uas_burstcount -> SRAM_CVGX:uas_burstcount
	signal mm_interconnect_0_sram_cvgx_uas_writedata                     : std_logic_vector(15 downto 0); -- mm_interconnect_0:SRAM_CVGX_uas_writedata -> SRAM_CVGX:uas_writedata
	signal mm_interconnect_0_sram_cvgx_uas_address                       : std_logic_vector(18 downto 0); -- mm_interconnect_0:SRAM_CVGX_uas_address -> SRAM_CVGX:uas_address
	signal mm_interconnect_0_sram_cvgx_uas_lock                          : std_logic;                     -- mm_interconnect_0:SRAM_CVGX_uas_lock -> SRAM_CVGX:uas_lock
	signal mm_interconnect_0_sram_cvgx_uas_write                         : std_logic;                     -- mm_interconnect_0:SRAM_CVGX_uas_write -> SRAM_CVGX:uas_write
	signal mm_interconnect_0_sram_cvgx_uas_read                          : std_logic;                     -- mm_interconnect_0:SRAM_CVGX_uas_read -> SRAM_CVGX:uas_read
	signal mm_interconnect_0_sram_cvgx_uas_readdata                      : std_logic_vector(15 downto 0); -- SRAM_CVGX:uas_readdata -> mm_interconnect_0:SRAM_CVGX_uas_readdata
	signal mm_interconnect_0_sram_cvgx_uas_debugaccess                   : std_logic;                     -- mm_interconnect_0:SRAM_CVGX_uas_debugaccess -> SRAM_CVGX:uas_debugaccess
	signal mm_interconnect_0_sram_cvgx_uas_readdatavalid                 : std_logic;                     -- SRAM_CVGX:uas_readdatavalid -> mm_interconnect_0:SRAM_CVGX_uas_readdatavalid
	signal mm_interconnect_0_sram_cvgx_uas_byteenable                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:SRAM_CVGX_uas_byteenable -> SRAM_CVGX:uas_byteenable
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest     : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata       : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address         : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect      : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write           : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata        : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_rtx_timer_s1_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:RTX_Timer_s1_writedata -> RTX_Timer:writedata
	signal mm_interconnect_0_rtx_timer_s1_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:RTX_Timer_s1_address -> RTX_Timer:address
	signal mm_interconnect_0_rtx_timer_s1_chipselect                     : std_logic;                     -- mm_interconnect_0:RTX_Timer_s1_chipselect -> RTX_Timer:chipselect
	signal mm_interconnect_0_rtx_timer_s1_write                          : std_logic;                     -- mm_interconnect_0:RTX_Timer_s1_write -> mm_interconnect_0_rtx_timer_s1_write:in
	signal mm_interconnect_0_rtx_timer_s1_readdata                       : std_logic_vector(15 downto 0); -- RTX_Timer:readdata -> mm_interconnect_0:RTX_Timer_s1_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address          : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata         : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_lcd_control_slave_writedata                 : std_logic_vector(7 downto 0);  -- mm_interconnect_0:lcd_control_slave_writedata -> lcd:writedata
	signal mm_interconnect_0_lcd_control_slave_address                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:lcd_control_slave_address -> lcd:address
	signal mm_interconnect_0_lcd_control_slave_write                     : std_logic;                     -- mm_interconnect_0:lcd_control_slave_write -> lcd:write
	signal mm_interconnect_0_lcd_control_slave_read                      : std_logic;                     -- mm_interconnect_0:lcd_control_slave_read -> lcd:read
	signal mm_interconnect_0_lcd_control_slave_readdata                  : std_logic_vector(7 downto 0);  -- lcd:readdata -> mm_interconnect_0:lcd_control_slave_readdata
	signal mm_interconnect_0_lcd_control_slave_begintransfer             : std_logic;                     -- mm_interconnect_0:lcd_control_slave_begintransfer -> lcd:begintransfer
	signal mm_interconnect_0_pio_sw_s1_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_sw_s1_writedata -> pio_sw:writedata
	signal mm_interconnect_0_pio_sw_s1_address                           : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_sw_s1_address -> pio_sw:address
	signal mm_interconnect_0_pio_sw_s1_chipselect                        : std_logic;                     -- mm_interconnect_0:pio_sw_s1_chipselect -> pio_sw:chipselect
	signal mm_interconnect_0_pio_sw_s1_write                             : std_logic;                     -- mm_interconnect_0:pio_sw_s1_write -> mm_interconnect_0_pio_sw_s1_write:in
	signal mm_interconnect_0_pio_sw_s1_readdata                          : std_logic_vector(31 downto 0); -- pio_sw:readdata -> mm_interconnect_0:pio_sw_s1_readdata
	signal mm_interconnect_0_pio_key_s1_writedata                        : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_key_s1_writedata -> pio_key:writedata
	signal mm_interconnect_0_pio_key_s1_address                          : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_key_s1_address -> pio_key:address
	signal mm_interconnect_0_pio_key_s1_chipselect                       : std_logic;                     -- mm_interconnect_0:pio_key_s1_chipselect -> pio_key:chipselect
	signal mm_interconnect_0_pio_key_s1_write                            : std_logic;                     -- mm_interconnect_0:pio_key_s1_write -> mm_interconnect_0_pio_key_s1_write:in
	signal mm_interconnect_0_pio_key_s1_readdata                         : std_logic_vector(31 downto 0); -- pio_key:readdata -> mm_interconnect_0:pio_key_s1_readdata
	signal mm_interconnect_0_pio_hex0_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_hex0_s1_writedata -> pio_hex0:writedata
	signal mm_interconnect_0_pio_hex0_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_hex0_s1_address -> pio_hex0:address
	signal mm_interconnect_0_pio_hex0_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pio_hex0_s1_chipselect -> pio_hex0:chipselect
	signal mm_interconnect_0_pio_hex0_s1_write                           : std_logic;                     -- mm_interconnect_0:pio_hex0_s1_write -> mm_interconnect_0_pio_hex0_s1_write:in
	signal mm_interconnect_0_pio_hex0_s1_readdata                        : std_logic_vector(31 downto 0); -- pio_hex0:readdata -> mm_interconnect_0:pio_hex0_s1_readdata
	signal mm_interconnect_0_pio_hex1_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_hex1_s1_writedata -> pio_hex1:writedata
	signal mm_interconnect_0_pio_hex1_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_hex1_s1_address -> pio_hex1:address
	signal mm_interconnect_0_pio_hex1_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pio_hex1_s1_chipselect -> pio_hex1:chipselect
	signal mm_interconnect_0_pio_hex1_s1_write                           : std_logic;                     -- mm_interconnect_0:pio_hex1_s1_write -> mm_interconnect_0_pio_hex1_s1_write:in
	signal mm_interconnect_0_pio_hex1_s1_readdata                        : std_logic_vector(31 downto 0); -- pio_hex1:readdata -> mm_interconnect_0:pio_hex1_s1_readdata
	signal mm_interconnect_0_pio_hex2_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_hex2_s1_writedata -> pio_hex2:writedata
	signal mm_interconnect_0_pio_hex2_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_hex2_s1_address -> pio_hex2:address
	signal mm_interconnect_0_pio_hex2_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pio_hex2_s1_chipselect -> pio_hex2:chipselect
	signal mm_interconnect_0_pio_hex2_s1_write                           : std_logic;                     -- mm_interconnect_0:pio_hex2_s1_write -> mm_interconnect_0_pio_hex2_s1_write:in
	signal mm_interconnect_0_pio_hex2_s1_readdata                        : std_logic_vector(31 downto 0); -- pio_hex2:readdata -> mm_interconnect_0:pio_hex2_s1_readdata
	signal mm_interconnect_0_pio_hex3_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_hex3_s1_writedata -> pio_hex3:writedata
	signal mm_interconnect_0_pio_hex3_s1_address                         : std_logic_vector(2 downto 0);  -- mm_interconnect_0:pio_hex3_s1_address -> pio_hex3:address
	signal mm_interconnect_0_pio_hex3_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pio_hex3_s1_chipselect -> pio_hex3:chipselect
	signal mm_interconnect_0_pio_hex3_s1_write                           : std_logic;                     -- mm_interconnect_0:pio_hex3_s1_write -> mm_interconnect_0_pio_hex3_s1_write:in
	signal mm_interconnect_0_pio_hex3_s1_readdata                        : std_logic_vector(31 downto 0); -- pio_hex3:readdata -> mm_interconnect_0:pio_hex3_s1_readdata
	signal mm_interconnect_0_pio_led9_s1_writedata                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_led9_s1_writedata -> pio_led9:writedata
	signal mm_interconnect_0_pio_led9_s1_address                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_led9_s1_address -> pio_led9:address
	signal mm_interconnect_0_pio_led9_s1_chipselect                      : std_logic;                     -- mm_interconnect_0:pio_led9_s1_chipselect -> pio_led9:chipselect
	signal mm_interconnect_0_pio_led9_s1_write                           : std_logic;                     -- mm_interconnect_0:pio_led9_s1_write -> mm_interconnect_0_pio_led9_s1_write:in
	signal mm_interconnect_0_pio_led9_s1_readdata                        : std_logic_vector(31 downto 0); -- pio_led9:readdata -> mm_interconnect_0:pio_led9_s1_readdata
	signal irq_mapper_receiver0_irq                                      : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                      : std_logic;                     -- RTX_Timer:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                      : std_logic;                     -- pio_sw:irq -> irq_mapper:receiver2_irq
	signal irq_mapper_receiver3_irq                                      : std_logic;                     -- pio_key:irq -> irq_mapper:receiver3_irq
	signal cpu_d_irq_irq                                                 : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> CPU:d_irq
	signal rst_controller_reset_out_reset                                : std_logic;                     -- rst_controller:reset_out -> [SRAM_CVGX:reset_reset, SRAM_Conduit:reset, SRAM_PinSharer:reset_reset, irq_mapper:reset, mm_interconnect_0:CPU_reset_n_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                            : std_logic;                     -- rst_controller:reset_req -> [CPU:reset_req, rst_translator:reset_req_in]
	signal cpu_jtag_debug_module_reset_reset                             : std_logic;                     -- CPU:jtag_debug_module_resetrequest -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                            : std_logic;                     -- rst_controller_001:reset_out -> pll_100MHz:rst
	signal reset_reset_n_ports_inv                                       : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv  : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_rtx_timer_s1_write_ports_inv                : std_logic;                     -- mm_interconnect_0_rtx_timer_s1_write:inv -> RTX_Timer:write_n
	signal mm_interconnect_0_pio_sw_s1_write_ports_inv                   : std_logic;                     -- mm_interconnect_0_pio_sw_s1_write:inv -> pio_sw:write_n
	signal mm_interconnect_0_pio_key_s1_write_ports_inv                  : std_logic;                     -- mm_interconnect_0_pio_key_s1_write:inv -> pio_key:write_n
	signal mm_interconnect_0_pio_hex0_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_hex0_s1_write:inv -> pio_hex0:write_n
	signal mm_interconnect_0_pio_hex1_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_hex1_s1_write:inv -> pio_hex1:write_n
	signal mm_interconnect_0_pio_hex2_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_hex2_s1_write:inv -> pio_hex2:write_n
	signal mm_interconnect_0_pio_hex3_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_hex3_s1_write:inv -> pio_hex3:write_n
	signal mm_interconnect_0_pio_led9_s1_write_ports_inv                 : std_logic;                     -- mm_interconnect_0_pio_led9_s1_write:inv -> pio_led9:write_n
	signal rst_controller_reset_out_reset_ports_inv                      : std_logic;                     -- rst_controller_reset_out_reset:inv -> [CPU:reset_n, RTX_Timer:reset_n, jtag_uart:rst_n, lcd:reset_n, pio_hex0:reset_n, pio_hex1:reset_n, pio_hex2:reset_n, pio_hex3:reset_n, pio_key:reset_n, pio_led9:reset_n, pio_sw:reset_n, sysid_qsys_0:reset_n]

begin

	cpu : component StepperMotorControl_CPU
		port map (
			clk                                   => pll_100mhz_outclk0_clk,                              --                       clk.clk
			reset_n                               => rst_controller_reset_out_reset_ports_inv,            --                   reset_n.reset_n
			reset_req                             => rst_controller_reset_out_reset_req,                  --                          .reset_req
			d_address                             => cpu_data_master_address,                             --               data_master.address
			d_byteenable                          => cpu_data_master_byteenable,                          --                          .byteenable
			d_read                                => cpu_data_master_read,                                --                          .read
			d_readdata                            => cpu_data_master_readdata,                            --                          .readdata
			d_waitrequest                         => cpu_data_master_waitrequest,                         --                          .waitrequest
			d_write                               => cpu_data_master_write,                               --                          .write
			d_writedata                           => cpu_data_master_writedata,                           --                          .writedata
			jtag_debug_module_debugaccess_to_roms => cpu_data_master_debugaccess,                         --                          .debugaccess
			i_address                             => cpu_instruction_master_address,                      --        instruction_master.address
			i_read                                => cpu_instruction_master_read,                         --                          .read
			i_readdata                            => cpu_instruction_master_readdata,                     --                          .readdata
			i_waitrequest                         => cpu_instruction_master_waitrequest,                  --                          .waitrequest
			d_irq                                 => cpu_d_irq_irq,                                       --                     d_irq.irq
			jtag_debug_module_resetrequest        => cpu_jtag_debug_module_reset_reset,                   --   jtag_debug_module_reset.reset
			jtag_debug_module_address             => mm_interconnect_0_cpu_jtag_debug_module_address,     --         jtag_debug_module.address
			jtag_debug_module_byteenable          => mm_interconnect_0_cpu_jtag_debug_module_byteenable,  --                          .byteenable
			jtag_debug_module_debugaccess         => mm_interconnect_0_cpu_jtag_debug_module_debugaccess, --                          .debugaccess
			jtag_debug_module_read                => mm_interconnect_0_cpu_jtag_debug_module_read,        --                          .read
			jtag_debug_module_readdata            => mm_interconnect_0_cpu_jtag_debug_module_readdata,    --                          .readdata
			jtag_debug_module_waitrequest         => mm_interconnect_0_cpu_jtag_debug_module_waitrequest, --                          .waitrequest
			jtag_debug_module_write               => mm_interconnect_0_cpu_jtag_debug_module_write,       --                          .write
			jtag_debug_module_writedata           => mm_interconnect_0_cpu_jtag_debug_module_writedata,   --                          .writedata
			no_ci_readra                          => open                                                 -- custom_instruction_master.readra
		);

	sysid_qsys_0 : component StepperMotorControl_sysid_qsys_0
		port map (
			clock    => pll_100mhz_outclk0_clk,                                  --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	jtag_uart : component StepperMotorControl_jtag_uart
		port map (
			clk            => pll_100mhz_outclk0_clk,                                        --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                       --               irq.irq
		);

	rtx_timer : component StepperMotorControl_RTX_Timer
		port map (
			clk        => pll_100mhz_outclk0_clk,                         --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,       -- reset.reset_n
			address    => mm_interconnect_0_rtx_timer_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_rtx_timer_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_rtx_timer_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_rtx_timer_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_rtx_timer_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                        --   irq.irq
		);

	sram_cvgx : component StepperMotorControl_SRAM_CVGX
		generic map (
			TCM_ADDRESS_W                  => 19,
			TCM_DATA_W                     => 16,
			TCM_BYTEENABLE_W               => 2,
			TCM_READ_WAIT                  => 10,
			TCM_WRITE_WAIT                 => 10,
			TCM_SETUP_WAIT                 => 10,
			TCM_DATA_HOLD                  => 10,
			TCM_TURNAROUND_TIME            => 2,
			TCM_TIMING_UNITS               => 0,
			TCM_READLATENCY                => 2,
			TCM_SYMBOLS_PER_WORD           => 2,
			USE_READDATA                   => 1,
			USE_WRITEDATA                  => 1,
			USE_READ                       => 0,
			USE_WRITE                      => 1,
			USE_BYTEENABLE                 => 1,
			USE_CHIPSELECT                 => 1,
			USE_LOCK                       => 0,
			USE_ADDRESS                    => 1,
			USE_WAITREQUEST                => 0,
			USE_WRITEBYTEENABLE            => 0,
			USE_OUTPUTENABLE               => 1,
			USE_RESETREQUEST               => 0,
			USE_IRQ                        => 0,
			USE_RESET_OUTPUT               => 0,
			ACTIVE_LOW_READ                => 0,
			ACTIVE_LOW_LOCK                => 0,
			ACTIVE_LOW_WRITE               => 1,
			ACTIVE_LOW_CHIPSELECT          => 1,
			ACTIVE_LOW_BYTEENABLE          => 1,
			ACTIVE_LOW_OUTPUTENABLE        => 1,
			ACTIVE_LOW_WRITEBYTEENABLE     => 0,
			ACTIVE_LOW_WAITREQUEST         => 0,
			ACTIVE_LOW_BEGINTRANSFER       => 0,
			CHIPSELECT_THROUGH_READLATENCY => 0
		)
		port map (
			clk_clk                => pll_100mhz_outclk0_clk,                        --   clk.clk
			reset_reset            => rst_controller_reset_out_reset,                -- reset.reset
			uas_address            => mm_interconnect_0_sram_cvgx_uas_address,       --   uas.address
			uas_burstcount         => mm_interconnect_0_sram_cvgx_uas_burstcount,    --      .burstcount
			uas_read               => mm_interconnect_0_sram_cvgx_uas_read,          --      .read
			uas_write              => mm_interconnect_0_sram_cvgx_uas_write,         --      .write
			uas_waitrequest        => mm_interconnect_0_sram_cvgx_uas_waitrequest,   --      .waitrequest
			uas_readdatavalid      => mm_interconnect_0_sram_cvgx_uas_readdatavalid, --      .readdatavalid
			uas_byteenable         => mm_interconnect_0_sram_cvgx_uas_byteenable,    --      .byteenable
			uas_readdata           => mm_interconnect_0_sram_cvgx_uas_readdata,      --      .readdata
			uas_writedata          => mm_interconnect_0_sram_cvgx_uas_writedata,     --      .writedata
			uas_lock               => mm_interconnect_0_sram_cvgx_uas_lock,          --      .lock
			uas_debugaccess        => mm_interconnect_0_sram_cvgx_uas_debugaccess,   --      .debugaccess
			tcm_write_n_out        => sram_cvgx_tcm_write_n_out,                     --   tcm.write_n_out
			tcm_chipselect_n_out   => sram_cvgx_tcm_chipselect_n_out,                --      .chipselect_n_out
			tcm_outputenable_n_out => sram_cvgx_tcm_outputenable_n_out,              --      .outputenable_n_out
			tcm_request            => sram_cvgx_tcm_request,                         --      .request
			tcm_grant              => sram_cvgx_tcm_grant,                           --      .grant
			tcm_address_out        => sram_cvgx_tcm_address_out,                     --      .address_out
			tcm_byteenable_n_out   => sram_cvgx_tcm_byteenable_n_out,                --      .byteenable_n_out
			tcm_data_out           => sram_cvgx_tcm_data_out,                        --      .data_out
			tcm_data_outen         => sram_cvgx_tcm_data_outen,                      --      .data_outen
			tcm_data_in            => sram_cvgx_tcm_data_in                          --      .data_in
		);

	sram_conduit : component StepperMotorControl_SRAM_Conduit
		port map (
			clk              => pll_100mhz_outclk0_clk,           --   clk.clk
			reset            => rst_controller_reset_out_reset,   -- reset.reset
			request          => sram_pinsharer_tcm_request,       --   tcs.request
			grant            => sram_pinsharer_tcm_grant,         --      .grant
			tcs_SRAM_OE_N    => sram_pinsharer_tcm_sram_oe_n_out, --      .SRAM_OE_N_out
			tcs_SRAM_CE_N    => sram_pinsharer_tcm_sram_ce_n_out, --      .SRAM_CE_N_out
			tcs_SRAM_BE_N    => sram_pinsharer_tcm_sram_be_n_out, --      .SRAM_BE_N_out
			tcs_SRAM_D       => sram_pinsharer_tcm_sram_d_out,    --      .SRAM_D_out
			tcs_SRAM_D_outen => sram_pinsharer_tcm_sram_d_outen,  --      .SRAM_D_outen
			tcs_SRAM_D_in    => sram_pinsharer_tcm_sram_d_in,     --      .SRAM_D_in
			tcs_SRAM_A       => sram_pinsharer_tcm_sram_a_out,    --      .SRAM_A_out
			tcs_SRAM_WE_N    => sram_pinsharer_tcm_sram_we_n_out, --      .SRAM_WE_N_out
			SRAM_OE_N        => SRAM_OE_N,                   --   out.SRAM_OE_N
			SRAM_CE_N        => SRAM_CE_N,                   --      .SRAM_CE_N
			SRAM_BE_N        => SRAM_BE_N,                   --      .SRAM_BE_N
			SRAM_D           => SRAM_D,                      --      .SRAM_D
			SRAM_A           => SRAM_A,                      --      .SRAM_A
			SRAM_WE_N        => SRAM_WE_N                    --      .SRAM_WE_N
		);

	pll_100mhz : component StepperMotorControl_pll_100MHz
		port map (
			refclk   => clk_clk,                            --  refclk.clk
			rst      => rst_controller_001_reset_out_reset, --   reset.reset
			outclk_0 => pll_100mhz_outclk0_clk,             -- outclk0.clk
			locked   => open                                -- (terminated)
		);

	sram_pinsharer : component StepperMotorControl_SRAM_PinSharer
		port map (
			clk_clk                    => pll_100mhz_outclk0_clk,           --   clk.clk
			reset_reset                => rst_controller_reset_out_reset,   -- reset.reset
			request                    => sram_pinsharer_tcm_request,       --   tcm.request
			grant                      => sram_pinsharer_tcm_grant,         --      .grant
			SRAM_A                     => sram_pinsharer_tcm_sram_a_out,    --      .SRAM_A_out
			SRAM_OE_N                  => sram_pinsharer_tcm_sram_oe_n_out, --      .SRAM_OE_N_out
			SRAM_BE_N                  => sram_pinsharer_tcm_sram_be_n_out, --      .SRAM_BE_N_out
			SRAM_WE_N                  => sram_pinsharer_tcm_sram_we_n_out, --      .SRAM_WE_N_out
			SRAM_D                     => sram_pinsharer_tcm_sram_d_out,    --      .SRAM_D_out
			SRAM_D_in                  => sram_pinsharer_tcm_sram_d_in,     --      .SRAM_D_in
			SRAM_D_outen               => sram_pinsharer_tcm_sram_d_outen,  --      .SRAM_D_outen
			SRAM_CE_N                  => sram_pinsharer_tcm_sram_ce_n_out, --      .SRAM_CE_N_out
			tcs0_request               => sram_cvgx_tcm_request,            --  tcs0.request
			tcs0_grant                 => sram_cvgx_tcm_grant,              --      .grant
			tcs0_address_out           => sram_cvgx_tcm_address_out,        --      .address_out
			tcs0_outputenable_n_out(0) => sram_cvgx_tcm_outputenable_n_out, --      .outputenable_n_out
			tcs0_byteenable_n_out      => sram_cvgx_tcm_byteenable_n_out,   --      .byteenable_n_out
			tcs0_write_n_out(0)        => sram_cvgx_tcm_write_n_out,        --      .write_n_out
			tcs0_data_out              => sram_cvgx_tcm_data_out,           --      .data_out
			tcs0_data_in               => sram_cvgx_tcm_data_in,            --      .data_in
			tcs0_data_outen            => sram_cvgx_tcm_data_outen,         --      .data_outen
			tcs0_chipselect_n_out(0)   => sram_cvgx_tcm_chipselect_n_out    --      .chipselect_n_out
		);

	lcd : component StepperMotorControl_lcd
		port map (
			reset_n       => rst_controller_reset_out_reset_ports_inv,          --         reset.reset_n
			clk           => pll_100mhz_outclk0_clk,                            --           clk.clk
			begintransfer => mm_interconnect_0_lcd_control_slave_begintransfer, -- control_slave.begintransfer
			read          => mm_interconnect_0_lcd_control_slave_read,          --              .read
			write         => mm_interconnect_0_lcd_control_slave_write,         --              .write
			readdata      => mm_interconnect_0_lcd_control_slave_readdata,      --              .readdata
			writedata     => mm_interconnect_0_lcd_control_slave_writedata,     --              .writedata
			address       => mm_interconnect_0_lcd_control_slave_address,       --              .address
			LCD_RS        => LCD_RS,                                            --      external.export
			LCD_RW        => LCD_RW,                                            --              .export
			lcd_data        => LCD_DQ,                                          --              .export
			LCD_E         => LCD_E                                              --              .export
		);

	pio_sw : component StepperMotorControl_pio_sw
		port map (
			clk        => pll_100mhz_outclk0_clk,                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,    --               reset.reset_n
			address    => mm_interconnect_0_pio_sw_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_sw_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_sw_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_sw_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_sw_s1_readdata,        --                    .readdata
			in_port    => SW,                                   -- external_connection.export
			irq        => irq_mapper_receiver2_irq                     --                 irq.irq
		);

	pio_key : component StepperMotorControl_pio_key
		port map (
			clk        => pll_100mhz_outclk0_clk,                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_pio_key_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_key_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_key_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_key_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_key_s1_readdata,        --                    .readdata
			in_port    => KEY,                                   -- external_connection.export
			irq        => irq_mapper_receiver3_irq                      --                 irq.irq
		);

	pio_hex0 : component StepperMotorControl_pio_hex0
		port map (
			clk        => pll_100mhz_outclk0_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_hex0_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_hex0_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_hex0_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_hex0_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_hex0_s1_readdata,        --                    .readdata
			out_port   => HEX0                                    -- external_connection.export
		);

	pio_hex1 : component StepperMotorControl_pio_hex0
		port map (
			clk        => pll_100mhz_outclk0_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_hex1_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_hex1_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_hex1_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_hex1_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_hex1_s1_readdata,        --                    .readdata
			out_port   => HEX1                                    -- external_connection.export
		);

	pio_hex2 : component StepperMotorControl_pio_hex0
		port map (
			clk        => pll_100mhz_outclk0_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_hex2_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_hex2_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_hex2_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_hex2_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_hex2_s1_readdata,        --                    .readdata
			out_port   => HEX2                                    -- external_connection.export
		);

	pio_hex3 : component StepperMotorControl_pio_hex0
		port map (
			clk        => pll_100mhz_outclk0_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_hex3_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_hex3_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_hex3_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_hex3_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_hex3_s1_readdata,        --                    .readdata
			out_port   => HEX3                                    -- external_connection.export
		);

	pio_led9 : component StepperMotorControl_pio_led9
		port map (
			clk        => pll_100mhz_outclk0_clk,                        --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_pio_led9_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_led9_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_led9_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_led9_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_led9_s1_readdata,        --                    .readdata
			out_port   => LED9                                    -- external_connection.export
		);

	mm_interconnect_0 : component StepperMotorControl_mm_interconnect_0
		port map (
			pll_100MHz_outclk0_clk                  => pll_100mhz_outclk0_clk,                                    --                pll_100MHz_outclk0.clk
			CPU_reset_n_reset_bridge_in_reset_reset => rst_controller_reset_out_reset,                            -- CPU_reset_n_reset_bridge_in_reset.reset
			CPU_data_master_address                 => cpu_data_master_address,                                   --                   CPU_data_master.address
			CPU_data_master_waitrequest             => cpu_data_master_waitrequest,                               --                                  .waitrequest
			CPU_data_master_byteenable              => cpu_data_master_byteenable,                                --                                  .byteenable
			CPU_data_master_read                    => cpu_data_master_read,                                      --                                  .read
			CPU_data_master_readdata                => cpu_data_master_readdata,                                  --                                  .readdata
			CPU_data_master_write                   => cpu_data_master_write,                                     --                                  .write
			CPU_data_master_writedata               => cpu_data_master_writedata,                                 --                                  .writedata
			CPU_data_master_debugaccess             => cpu_data_master_debugaccess,                               --                                  .debugaccess
			CPU_instruction_master_address          => cpu_instruction_master_address,                            --            CPU_instruction_master.address
			CPU_instruction_master_waitrequest      => cpu_instruction_master_waitrequest,                        --                                  .waitrequest
			CPU_instruction_master_read             => cpu_instruction_master_read,                               --                                  .read
			CPU_instruction_master_readdata         => cpu_instruction_master_readdata,                           --                                  .readdata
			CPU_jtag_debug_module_address           => mm_interconnect_0_cpu_jtag_debug_module_address,           --             CPU_jtag_debug_module.address
			CPU_jtag_debug_module_write             => mm_interconnect_0_cpu_jtag_debug_module_write,             --                                  .write
			CPU_jtag_debug_module_read              => mm_interconnect_0_cpu_jtag_debug_module_read,              --                                  .read
			CPU_jtag_debug_module_readdata          => mm_interconnect_0_cpu_jtag_debug_module_readdata,          --                                  .readdata
			CPU_jtag_debug_module_writedata         => mm_interconnect_0_cpu_jtag_debug_module_writedata,         --                                  .writedata
			CPU_jtag_debug_module_byteenable        => mm_interconnect_0_cpu_jtag_debug_module_byteenable,        --                                  .byteenable
			CPU_jtag_debug_module_waitrequest       => mm_interconnect_0_cpu_jtag_debug_module_waitrequest,       --                                  .waitrequest
			CPU_jtag_debug_module_debugaccess       => mm_interconnect_0_cpu_jtag_debug_module_debugaccess,       --                                  .debugaccess
			jtag_uart_avalon_jtag_slave_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --       jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write       => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                  .write
			jtag_uart_avalon_jtag_slave_read        => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                  .read
			jtag_uart_avalon_jtag_slave_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                  .readdata
			jtag_uart_avalon_jtag_slave_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                  .writedata
			jtag_uart_avalon_jtag_slave_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                  .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                  .chipselect
			lcd_control_slave_address               => mm_interconnect_0_lcd_control_slave_address,               --                 lcd_control_slave.address
			lcd_control_slave_write                 => mm_interconnect_0_lcd_control_slave_write,                 --                                  .write
			lcd_control_slave_read                  => mm_interconnect_0_lcd_control_slave_read,                  --                                  .read
			lcd_control_slave_readdata              => mm_interconnect_0_lcd_control_slave_readdata,              --                                  .readdata
			lcd_control_slave_writedata             => mm_interconnect_0_lcd_control_slave_writedata,             --                                  .writedata
			lcd_control_slave_begintransfer         => mm_interconnect_0_lcd_control_slave_begintransfer,         --                                  .begintransfer
			pio_hex0_s1_address                     => mm_interconnect_0_pio_hex0_s1_address,                     --                       pio_hex0_s1.address
			pio_hex0_s1_write                       => mm_interconnect_0_pio_hex0_s1_write,                       --                                  .write
			pio_hex0_s1_readdata                    => mm_interconnect_0_pio_hex0_s1_readdata,                    --                                  .readdata
			pio_hex0_s1_writedata                   => mm_interconnect_0_pio_hex0_s1_writedata,                   --                                  .writedata
			pio_hex0_s1_chipselect                  => mm_interconnect_0_pio_hex0_s1_chipselect,                  --                                  .chipselect
			pio_hex1_s1_address                     => mm_interconnect_0_pio_hex1_s1_address,                     --                       pio_hex1_s1.address
			pio_hex1_s1_write                       => mm_interconnect_0_pio_hex1_s1_write,                       --                                  .write
			pio_hex1_s1_readdata                    => mm_interconnect_0_pio_hex1_s1_readdata,                    --                                  .readdata
			pio_hex1_s1_writedata                   => mm_interconnect_0_pio_hex1_s1_writedata,                   --                                  .writedata
			pio_hex1_s1_chipselect                  => mm_interconnect_0_pio_hex1_s1_chipselect,                  --                                  .chipselect
			pio_hex2_s1_address                     => mm_interconnect_0_pio_hex2_s1_address,                     --                       pio_hex2_s1.address
			pio_hex2_s1_write                       => mm_interconnect_0_pio_hex2_s1_write,                       --                                  .write
			pio_hex2_s1_readdata                    => mm_interconnect_0_pio_hex2_s1_readdata,                    --                                  .readdata
			pio_hex2_s1_writedata                   => mm_interconnect_0_pio_hex2_s1_writedata,                   --                                  .writedata
			pio_hex2_s1_chipselect                  => mm_interconnect_0_pio_hex2_s1_chipselect,                  --                                  .chipselect
			pio_hex3_s1_address                     => mm_interconnect_0_pio_hex3_s1_address,                     --                       pio_hex3_s1.address
			pio_hex3_s1_write                       => mm_interconnect_0_pio_hex3_s1_write,                       --                                  .write
			pio_hex3_s1_readdata                    => mm_interconnect_0_pio_hex3_s1_readdata,                    --                                  .readdata
			pio_hex3_s1_writedata                   => mm_interconnect_0_pio_hex3_s1_writedata,                   --                                  .writedata
			pio_hex3_s1_chipselect                  => mm_interconnect_0_pio_hex3_s1_chipselect,                  --                                  .chipselect
			pio_key_s1_address                      => mm_interconnect_0_pio_key_s1_address,                      --                        pio_key_s1.address
			pio_key_s1_write                        => mm_interconnect_0_pio_key_s1_write,                        --                                  .write
			pio_key_s1_readdata                     => mm_interconnect_0_pio_key_s1_readdata,                     --                                  .readdata
			pio_key_s1_writedata                    => mm_interconnect_0_pio_key_s1_writedata,                    --                                  .writedata
			pio_key_s1_chipselect                   => mm_interconnect_0_pio_key_s1_chipselect,                   --                                  .chipselect
			pio_led9_s1_address                     => mm_interconnect_0_pio_led9_s1_address,                     --                       pio_led9_s1.address
			pio_led9_s1_write                       => mm_interconnect_0_pio_led9_s1_write,                       --                                  .write
			pio_led9_s1_readdata                    => mm_interconnect_0_pio_led9_s1_readdata,                    --                                  .readdata
			pio_led9_s1_writedata                   => mm_interconnect_0_pio_led9_s1_writedata,                   --                                  .writedata
			pio_led9_s1_chipselect                  => mm_interconnect_0_pio_led9_s1_chipselect,                  --                                  .chipselect
			pio_sw_s1_address                       => mm_interconnect_0_pio_sw_s1_address,                       --                         pio_sw_s1.address
			pio_sw_s1_write                         => mm_interconnect_0_pio_sw_s1_write,                         --                                  .write
			pio_sw_s1_readdata                      => mm_interconnect_0_pio_sw_s1_readdata,                      --                                  .readdata
			pio_sw_s1_writedata                     => mm_interconnect_0_pio_sw_s1_writedata,                     --                                  .writedata
			pio_sw_s1_chipselect                    => mm_interconnect_0_pio_sw_s1_chipselect,                    --                                  .chipselect
			RTX_Timer_s1_address                    => mm_interconnect_0_rtx_timer_s1_address,                    --                      RTX_Timer_s1.address
			RTX_Timer_s1_write                      => mm_interconnect_0_rtx_timer_s1_write,                      --                                  .write
			RTX_Timer_s1_readdata                   => mm_interconnect_0_rtx_timer_s1_readdata,                   --                                  .readdata
			RTX_Timer_s1_writedata                  => mm_interconnect_0_rtx_timer_s1_writedata,                  --                                  .writedata
			RTX_Timer_s1_chipselect                 => mm_interconnect_0_rtx_timer_s1_chipselect,                 --                                  .chipselect
			SRAM_CVGX_uas_address                   => mm_interconnect_0_sram_cvgx_uas_address,                   --                     SRAM_CVGX_uas.address
			SRAM_CVGX_uas_write                     => mm_interconnect_0_sram_cvgx_uas_write,                     --                                  .write
			SRAM_CVGX_uas_read                      => mm_interconnect_0_sram_cvgx_uas_read,                      --                                  .read
			SRAM_CVGX_uas_readdata                  => mm_interconnect_0_sram_cvgx_uas_readdata,                  --                                  .readdata
			SRAM_CVGX_uas_writedata                 => mm_interconnect_0_sram_cvgx_uas_writedata,                 --                                  .writedata
			SRAM_CVGX_uas_burstcount                => mm_interconnect_0_sram_cvgx_uas_burstcount,                --                                  .burstcount
			SRAM_CVGX_uas_byteenable                => mm_interconnect_0_sram_cvgx_uas_byteenable,                --                                  .byteenable
			SRAM_CVGX_uas_readdatavalid             => mm_interconnect_0_sram_cvgx_uas_readdatavalid,             --                                  .readdatavalid
			SRAM_CVGX_uas_waitrequest               => mm_interconnect_0_sram_cvgx_uas_waitrequest,               --                                  .waitrequest
			SRAM_CVGX_uas_lock                      => mm_interconnect_0_sram_cvgx_uas_lock,                      --                                  .lock
			SRAM_CVGX_uas_debugaccess               => mm_interconnect_0_sram_cvgx_uas_debugaccess,               --                                  .debugaccess
			sysid_qsys_0_control_slave_address      => mm_interconnect_0_sysid_qsys_0_control_slave_address,      --        sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata     => mm_interconnect_0_sysid_qsys_0_control_slave_readdata      --                                  .readdata
		);

	irq_mapper : component StepperMotorControl_irq_mapper
		port map (
			clk           => pll_100mhz_outclk0_clk,         --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			receiver3_irq => irq_mapper_receiver3_irq,       -- receiver3.irq
			sender_irq    => cpu_d_irq_irq                   --    sender.irq
		);

	rst_controller : component steppermotorcontrol_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_jtag_debug_module_reset_reset,  -- reset_in1.reset
			clk            => pll_100mhz_outclk0_clk,             --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component steppermotorcontrol_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_jtag_debug_module_reset_reset,  -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_rtx_timer_s1_write_ports_inv <= not mm_interconnect_0_rtx_timer_s1_write;

	mm_interconnect_0_pio_sw_s1_write_ports_inv <= not mm_interconnect_0_pio_sw_s1_write;

	mm_interconnect_0_pio_key_s1_write_ports_inv <= not mm_interconnect_0_pio_key_s1_write;

	mm_interconnect_0_pio_hex0_s1_write_ports_inv <= not mm_interconnect_0_pio_hex0_s1_write;

	mm_interconnect_0_pio_hex1_s1_write_ports_inv <= not mm_interconnect_0_pio_hex1_s1_write;

	mm_interconnect_0_pio_hex2_s1_write_ports_inv <= not mm_interconnect_0_pio_hex2_s1_write;

	mm_interconnect_0_pio_hex3_s1_write_ports_inv <= not mm_interconnect_0_pio_hex3_s1_write;

	mm_interconnect_0_pio_led9_s1_write_ports_inv <= not mm_interconnect_0_pio_led9_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of StepperMotorControl
