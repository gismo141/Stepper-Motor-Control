// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
d2FdIVohCEa8lkkq9c3Dzv64vGOi4bfd/Usjc8BjzkUtaX2fEndXB+BlO5akqFyoYbQiAErmw8dC
x2LBGDy9oINya2K9RvyYd035tM2GDbB2rIETJsXF+mITQSYoUFa7oa3vN8ha1zGRAOL8hRIXK5To
Xbi1PvU+EsJc9VjJnKL+bgbAYjbxOSyqnds3rDsMHs6ViREj9XS2XT3a7DfDbLMWH876WFR0Q7uo
CwKQmA+plfcbmDOB2+HV81UV9pAniwf1Q4bZTTWAdOGRI9qyI1tnQ7QgoyhcIdb8ijoROAponOya
9Fq6Ls+KmQb3mnEfctmNXnImQtZE9pY4flH/4g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
XwFT2DAhKhPVmbLPd2pDqf8MdjKKHcTc6yRZgVRLkRzlk9ko+VJdKcMNhRLGcKbhzlPusHT65Yxk
U0DdeuAAiRaOR78AAkTnEYk1ZFS5xLhClsxP8a+aBAWAZtLDvUd7Vs/k7Z++nhLcYUjx/eUdRyP0
UuoeGdQwqjZkkfxk4sgO2eCBiCM9h10VhMVsEe7nJZOdvf1gsINObPvGOIg7K7VbhW/SRHWhLEG8
ePo8d78A6DeXhomSUr2NHbWuV65tF3SJN5+FA0sN7oYyUbkRYMGlgeWLqARyoiitwVWbVcME0Upg
pRJDpLNZOsjTDJyM9lVEJfqzjqAkFPlFCI9ZcNE0FiPUPqKeacZOAdK8vRoj+iota0VSs0R5tw73
xHUnRaTJu++pb8mkgXPEdcaHOBZusq6NvKp50ZMIUbo8N7Bjpt41hxhD9m3JHxRf5dYrVeZLgJBe
ssz73nclELwFI5MthPaWiPb95L3YHlWborw4P/hiYG4Y1KYuJBljzYXq9iPSKqKfqSJy3WuI3jBu
O1mgVyAgijlkmhOJzoQtwZ5YTDp4CDqWbIeVSHAmyJsYzILC1ozO49ijwU77oahdzQA4f95WE7ny
gvYA2hvT2p1NsMA8d5eFLgVKONMYFvCU8eRLeo0NVjijV54ggsNlZIufTLRLVXq6QyL5F5ph/wLm
hZdHSRczq4a3nJBx/tS1/eLFrLTOI2r5DgmUxLJQj1VOFkKojevV1+j+L/atANaXe9RaFxGh6NSi
wtgL0Bp+XWaruItvNbD0ySc9ca28rbTczAu47PTVuX1czdZISLzj2R5GsedGxl1uWAAoPwqiy7Bi
mD+56RfJFXxTeoTAYuV0ScLqDt8eVvW4dP+JqAHXriCX9ppkRunkCpcIlv+VrLDAIwOBr8lB3brX
R1X4RVfRnQnyPy7Cl3YNihCqq77d5MGK2ldHF6ldzq9f1da+86qJaMyqQG5lbluT0VSYYf/Je0r8
q8llf3mxrIb3qQWJLVLZHT1B/bRirnJ0Bo//pcQmCQPpq3uWRJ+BMCW57+KQ1RrKmLx1z9autxRb
f66fK5EjWtM45xM3HYViEIC7Ol29xqX0EmJhRvPksfm4uroDh23KiGO5rZ9ETBlpMFINWQr2qYNC
fUSFc+GKq6oHIXWjn6ga5rInpDYQTHeIPyzScTNDed8hdit5u/Z2cnYoaqOfOx+sNn+to1nFxBS9
ueFv4d5419K97mRdvkLl9+ECnE+952lcV0inhfIJa/EWFIEbd5lQo3vJtTC7pcaCWCSqyfB3nKqE
xUoKaJfDD0OJ4vQFgdcm0cQy9iTE9dYdgysIML3+PvPRhFAMkkvpwm1dFTwNYJG1n+FB0dG33NG6
cJIoK6+4/nd/PPmhxCp8063o4di2MVZIC+4TDE/J+WAmaYY7VCO9EsBcNV0Ta9sEBWlk2cNPS5UP
XIqvsUWWyvRA9cj2p6feP1uzS/TYaMFgwrx6gBgKwwBiBEmVtZna43ncNWbj8MkaUJtFSjZYiacA
Pt43hjiIV1T+/we+wXM5X4GZUlzq1KUQjRn57AuOwwviMv3L35S9Zv1bBCOihX8FQOtmyKrsa71x
GTeY5LrP6WqgAL6NPXyUHpCav9UQu3lh/NiqoX3wK4yOvv1un1/O+adwVmeHyF8ZQGxAIZBBdq0z
bXVTwojzQr6IoHDbsZ0+e+LPEW7sMdJgZtZhefsOsn6JrsIDFjGpJ1vsfdcvtPgN82XevbN/yyeB
Sbn1IIpzaY0aALVjIPMzbl3e+OzMlv5ikpGaPdidHEAevusj1neAr0wYJSRnSpJa6Y8r3YOA1KdV
DzZzmIVIRoc3vwBeIATKgnYKPUs3/p3S0U8bGc6Mi28uvwHJ82Hzv1Km3PSc+EVlJRxhOVTZIXQ4
tyNSx+OZztfOpnSvZJwfOZ0/SMTOqy8/z4gV4gCtbB+lbusy/LtYudEM+JaefS7ujjl5NoQlLq9t
QIH7CaAHyrDFDld9vHOx0zZSP9mjcq9dI1JE2kh5/H0o74K2jwkGHy5huVsRM8/gbs6U8QJjuiZ3
yaY7bJgSDM0re/KCC+r4w6K46dsVtNHs2OD6GkQjYjX2Kz0TZxPB4Kv+gr85DdoZwvx6P4Ydfjpp
JEf/ib9U6NvrgBVn2GH3ZHzy+0H3N+BfxABsfM00T77hK+Ebl55qwkWFCIb33SOO37dn8d2bOUqi
xIwsZFr2cHXnlGj8G9AXBDaPWlHeY3ryFRmyqQNbyvBrfWz19x6OSHXkXurpRIBF9miMpQjbUS5V
/cnc07+hJtXSnZ9IfuYqWXrdItfcaTv+/lMTMyV6jOBgpa20ODM18UgPDbfAw1Dyjc2MuyO5uz3+
AFcLtSZX4CjKv8SvOI45imAdjy+qZHkcyYaaCE6zFp/h7T9YKYTg6DPcrWWbaQDuDJiKhS8mpOJ2
HbbGOEtuwZfgedW8OI/nwxNDjT+AL4U5bJ9v9U+Tz0joeHYosCdjv+42de3pRcKbXPiDzZl/Kyzk
r1G24z8RjZ6UfZYOTF9W5wpaFw8UWaSM+/+Qq/KEP2E4K7juVSfJ3edySOTlTSVvmeY0k6QDzRBi
+H3ddyy3BtNBSuptolJGC/DDoM4oPDnULzsGlihqvSj91RF5gqnKg5tlYrp91Mrig+zbS1+2/Sdi
DBtL6+1oqTiZnJZnk22mMvRpO9NIiMGCvrPCGTZX7oRNePrjp/v1oO3boU/Dm3YJRsGurgceZ68A
VTRPRcHYjK8jYSiqLbZmIHf3CSoeAVLCtH8mMWKeB5UncaMrlIksTUN7wuUB5k+EXUvTkAzZ23Px
7ol9FbZifb9+ABOklxye9zFeEcqVCbDmS2xaDeQziiqKSJQB2lTB80cLpHZnVmaV2NaMlJCCgyUq
vb9MsAArZK7t1MN1v6XNMidaAcaNUCmC8evoRyN4YdYtD8PYWY6fYe/pL9j79kZoWjK9Z7MhhQl6
7eNR//NAz93747z7L1vdzuYb1GgUnYpPvEb5rePeLrtjHVMgF7DJClUfUHGKYDUPYMnH60zFU3ds
H/9Mh5etroMIsBwkadC5elCS6/WQ0HkxIa28AfDwtRXt4wni+ZyC6zGvkkNopBL7/kkHdx+z9zbt
GYSX1IGx2o9cfHPDN8fOePXXvrJjSR0je+1cICCzjTEYILVq6n+EAxX/83blcPJ4q5WEKSK/Cdgi
nw24fXk0JGTp/vpFJZmbWSOBbGKZ9osRxlppbzC+kclfmTgjq0knlzWgimduyforEjLv1QY5zIvG
31DsqBM7YXWHtTIKLx323C7FeEtHMAHOzLGPjsapUxn1dzHz8Xd5PBTK4/q2Sp6Cra3IWBFADKh4
twDAqHsEqqhm8C6JXEqSAs8w9jHMt2ptGBlG+ni2CgadQoU42nAHBZGHmnNTNfCm1TlzHyB9Ojdg
DhBdXvdSD0b+nxJ1fUM5Ic8odDoBXuHG86Q9fhjSuOCRfu/UkKQ7oxRLQBV/VSoqdpepnOT66BFe
Y3iDPQxA0nchw6+Ajn2C5IrMc9qsA6EUSxu85lfuCfhnPrWaxhZXB0PaDBJ5CXr2nvZL2nJa+1Y3
GdtI70TANsaG/QsxoMLf9XUe5GZ2UuUexJJzaLJWaUlT/lcjWvpdujIwyYnuA28uUw82ZR1sYXiH
Jj9qrWJTZMw1SPo6xIVVK3pLA0L/VyJBn45dR+5mVdu86qK3osQk12ewxioUARmFrS9HVfl5QqUw
majUP4/lhSkDCgcTmHOTStGfGldF6Btn8oED6zUvq7e+8iOZs/8a54OD0OBbaCdEkHYBR8GEVq3h
uVyRBYrOh4CUzlOD7+64+4UhHOlXyELQIJexBOgllGPP0ixalz/RzvVeXK5zdC6tx2ek5XzOn6VH
UTFius4JCosj+vGr4LyfumEf9w+pReT175TI6CexdzPlZ5tp6u+/RwnNMA94RpJPD3TcvknHG5bo
5MSLYI4zE6AiUIvlxNAFGPKixhXxdn/FMS7ptYWJkiU03OMh4iUtbKO+Rc57C4IfvG6zk/GsftTD
woCKPG3BdZrUIQL/Dq2F7ttquAhf/TrcLplbzoE8KDP2oDEd6jKRtGzy/EbnsGpObOz//0jWBO62
ebu0v8U3JK5sBG5ZroUyNqpyxM+xmC+dv4g2XzVNcwuodYK1mPf7QC8oOwoQ+QeuLmx+lk8lgZXu
K9lEXQ0R3517IS+WHjhneGhH/0I/uxojU7XPGXnaNkdgvNE0n8yR727syXTtOahGTYqGaIkRiYDX
ygkEjR8FO//PzMi2Ow1euDnMy9X9ccip0F6PzkD/XPO56RJgyLqH4e63L+8WSHFAUKjvXtSlPVho
oqTPRDpkXUGlTbLjk3B6dyQE1fe56xg9V03pZAywtwM23RZ+1zQ+Ss1hr+tQKyxv101GZ9nBcjo/
fY4K6r3yoFynAVf+y3l2usscHpCe1TmLBIAT5JwtN9IkRF54PfsK8kSrdqX58PMpJrXisvLoxmM2
4kSRKvAn0y18Rv66bajdx7sBsCPhfzXWk3CmC3Z0n7RGTZK9PlkFUp8ct7RtK6ur8kwE+aQ95EDx
F0fJsEfBRl3dBq6aHjSnuDG+6ZDMGuSxnN93f+cNDMOtX8j24uAkY4TFeo3jmxM33gtq6n1keiJE
cZdQzkHP76DT4S2FBv46A1F9z94hrdMfJSiqHoZJGl71PqZvBS3zly/oRzhSLpxxb15JO0Ux5J2k
vnJ8BuzcHjzE5GDCZSHhMCh+Zwj0dCRKHxmFAXh5KltfeTi54pLmTcWFfwljcwh8K0poNEmrQolh
mi5QQcnRb4vKlTc4LSFSUYSP1zC1k7xfrfYhrBtAxA1Z2KP6pps64JDuA9o5+ZR0e83p6E43Xskz
i9FZO4KFibqpNs3m9NcMlBkDL3ZwM41N0F15PUh2cgc3u+Ju19c3viU44aUtMUXXX9K0tCiC4/m1
dPSfCMBmRl7LfrrIqNr46CE7CMeDCZkIYhWCaVIyPlJMl4wAEYMWcaVs8tHA/s64yOfBGkHNiYH5
CJox6cgT/UTCR37puE37GFsr7v5P3lzbfWWdQgd3+iofgMwqx2GnzfUXtJblRhaPRuP8BP9Ad4uA
HJ68mIM/40OHkwvenxajnmJxpo9OfVNG8muixl00nldmvVW/4XnbfVOXjgk3e+jNe8yrUn6sHS3r
XGRjhZBBdaLFFTFI+K56VCJdgh0rRWs6tuTT1yQq+Lozy/rSmr5dY0esaQYge7IO3jC7n6DRZt+r
3OSE6Q7vDfrJt8N9BTSNoZJqcUPqjJmxDM98IuWcyHx6k1qPAIswF89Tv8WYeh3YHoE3KFzcsYZF
z7q7/+/VbgEPwSGs3h6NZdovBVfEXemFU6+vySfAS2gsNSdZyJdyBeCY71UwCpdyedMlA8D5wgPD
LvpiF9UDEBzV18tdX3SyP/mAAEMiY06JQk26DOIVAbRrVNgru1tQpPQ4q3P6Fe/+BDuWQ7Npi2FN
/FH33FlHpmAHy9/6SRBazwUf3blK7TYgheLIi32pIlOgmCN5PpbV/TLxcSTlW/1OOoDtZoKlVpdC
rOLmvY7qqk8eSceEnEKPnVFX8rUDFTpyorKSQGlcpc50lMdsz+SYNz/ZKsuy2TGCBs14EwDkg85m
pCa5l4Vk+7o4xVscFopnKCmCgy93pioj4p0kGZeMEvanWthuRvPw7mCQn3lFNK776I+Q6d97MOjM
5E1ujBlCMrfk3xYRBKX2kES9uKBG6epZ+ZdwIHPOxkfZ9bO/20qhNEaEx5HX8T8LaflyQ78RJVMs
Zyz+VPxnJt9YJOE0u4LpH0JURWJedqii58T8+FRftjIijaDR48PFcQN4UzMYaxgDO7pteAqnb8SH
Rlr+RhEaHaiWiAIAAu4G4+ldFudMYUbqyE3ZLujbQFd7UMY49biAm93KKRJvGAivtVoY9JG5og6A
5WjCgyN138iL2rOMjZjMBwTuS9/PI1ASFRVOJ/Htq87Fg3Bd8fBoFFEktCMqFjTwn+LoNbYSZ+xe
83CwKIZK3W/U1urOdr2e5OVT2Q8oCJ6tTVHz6/Yg3wUFAwv5oqhHooWPD/KGUr4RuE5ywS1jm58B
hKWlfxo1s2WRnKXv3aThN6zd/hOIEZGMVCV7vfdy6VfpOJZ8BMVnaQkCtO9HiJhhRPALtVJka+yx
eQ5DIBmoyPhfJ8XXLNwVnlmcG/qHlHVyJ+RbgTS+FwXRIuD+gbycuA4x7jvlXu3Cxkrf7FQ78vpt
s0jvTe9/1NV3DGc5a/lPk6IpqqFMUvQbPBnvgYqhJ0oS3ano9s2MaLBpIcBpdN6ngZw3JXMDTfot
NDX01L4JdWysYqUaYKcWFvGlBUSHBmhiY0dgynk2NA02qLw4yEaxPmTDOlNhGLgr1xFbxwzHbD/O
8dRlmmfNTfg3vQMGAzDRnPRjhx3HU68zp6QKyHItlQ2JA7dpnmK4IBIxCWB0ML76gTBcO8EU7fWr
qFoKnGd01eaVu43cx82p2aXDWhS13Df6pbNU+1wKRmRFbPGA4HFVM3jfchj5F07KGsuxL0PCVpnB
IVqs+Ld3qtcQK5seIF5bzY/JH7hsBt28oZ9nypW4cd75M/sJAAIBP/u4+uq4+7YyXKAH/2Ee2xCP
wDYthusoSfMyyT1zy3up1/B7WPc6JDSTIG1Zv4odpCTraFRj/FuETwTggIcAN7sGfm9A3sRBR31z
o/JE5DFkEUN6cDIUR0F3rzJOf4cvkW1jiQhWxwXI+ijBzW9xrjGMw3X12Kzuhn8x+Sy1wpheEU9h
FvtVGvs4Klou/c6EnJXQx7jbCw7JjHwJMbwxI9tdQesDewDekmmHX06mghsBoa/jHfQ6XJ5bUpRi
yfGqIO1tiLvabiK4u3g0Gy8f+J18+YIm21q8F+9+83xX42qiSHON5tBG238kAI2HdFczYlr9TqA/
OmUgpWtDU7UEFHsNs19jdN8xIly+7exIjl75P3kB5iIHfqRA/SgwwdsfLSGDR3p5tPlIyjeWt3HT
gst16FY4ZXd7tsYwdDLQM1VuT43EM7EOolXWG/nIK7s1KjSrG97LGDO6d6PZT9jAYYnyoraHQpOn
OsqmBgTj8DESsua5rJV8A3+Yd/iA74eHmMWmVHEFMK8NNif8Gptss6tciFbyCncO91mT9eF9j6k4
TUBM6BSEJSA3BM+q1OhpYMeLppN3/BFoiWZYW2s1vIeizOWfnNW0USAlfhvXUG3dvxtUTCZo0iLb
E06fuPMyC8G4vIOoepu3HY1rHNhdN5/Zp6Bbr0npUi8OienK7zbP4Subl1MYeYXmTjOgYX39PLcX
P76xYRRFN2SEt12C/Jkl8u/a+DRU99JLPztQKdT1pwpcLKeAj07O2ro7vIW7ZEsFiA9avchCDAJ0
Ibrhm6qbepAdY9eksQqrgKp+vptiVdZugWt9s6HKJKbrgVhS+yheE+ADShGCSMboiFPQ6IjAclsV
St/8u10ZoqR1JJYc9N/SgKKdKi5FIvJc0cWhnvZcvR7ob/oBMCYiAu/60EV0hPjZro+bxpLb1hQ6
1jG7tHkepH62/hwubdjXHwFjhvm7E/i3ZLTbFRTViRrqS42nuV/ylDmUgBTkI2V27d+/HqZnbDKF
QQxhQVfLO6yJQBfVKIqmJxJigSvJlqXS3PmpdQH7hsQl/c5BOJqGKMqK8Pp+9AASlatmI3nqZJ1B
B3wqsJcY6nNWU5Eej4FVSXIEVJ33W4vHHHnRluVhhSebuoULc2utq4WtIV1mZ0YyT3ifARxg76ob
E2E33UiaH98SP/7N1GUXvf8FgrUxfoU98JX5XH8pr//hKpOiT0L6Y9RYocHG62HB8wnanc+k4L/L
+pUxF5t47KCZ9ufmM3K9bsMl3v9+lRH8yqVmod3cwPAuYboqVbFEbbxe7tfdLJEyObLl9DGlGD4b
yhY2mookV/PU/TI7l3mN5WVr7qeb62ZSocjouC1Jqit4+LwIK5gypkMe1OYXE6YMJWhBbYc2GMwJ
qs2a8jz6r1hXG9TKq6oL/kWx3edpFBvHm9EXz17MAzif0meenMqHc0NFg4Rh8LFxPRzTdIlYU6fS
oH5lEP9CnnMWz12vLVy1ujTUW+BP9g6qAv/iLIwNUcPEjz6QNdiB4IXHQ9KxXmvybT2nG3l9oU69
cZ+XQnBBwRB9mGzuBiL8NsLwsGrUJYqOhsHKB8Sd4zvqKHou5Um4RCVF08x19MnmY+Va30JVyxyQ
Br1tP/x6uaGBw2vSK7w89li5JHLQeyr3yl7/1IjRvnSlAH6GBgBY7V/EFM83sjVCFpnuwVvKpMeQ
OoyPUmjU/ljf0YWeB/FMgbrPHfZzr6gP8bIjoYG3CQy6H97Jld/MeXphk0rl9g+YpRoE7eeuE87T
IwG89qY0OGnQSjXhLye6nKQLBRg+L5LxAG0IApUUrA7N33l6R16+whziQFKwsIAZTKzPBFAHpKgX
As3n+9NLdTvSN8NO0DrnW84DsXg4HMd69p4xZXUVhv4x+6VOl68Vmwgz9eLyvW76iiFg2idp8XkD
BT6P0uUD7dGyWIGIA3V6ve2j0on8CV53jwiZxhrdsSJjKfVNYxDOCAFNygo3AVoPw1oIeIVc5hdK
yWjLoJwVihoc80CwCBIF4ASJGyTEXwVHVxrRYO2/iWUFbzro+LXukJVH8VgeL5AlOHgFgbI+xcbJ
aOJ++YZKauv//HOJyc3tl9dLt0O0CxAfZQRwrPbh7NHnsCZBFLOzgjRkUrejIE22fNdW5mMFLa1C
hN9DszYtTcVhLsvxlHUolmqWUi+uS8XMmJg+H9obdVuxg7kXL2xcyaxBwFAmYSSgkJ7leqd+T5aN
gx8XwqkilugChBBUBD4PHvQ4uUiQLg9be+BXg8K7HroGws8ebNtQ24j5JFBb8usvUkuGtRBsumAm
hsvsmoFOgONDdhi2VVL/v92wVMF2LFfXm7/0xXP3tidVsbugW1+SLuYxQIBVvMDZZqWTtgLqu40U
51Qhl5OpeOzjjb5/quloRyH3KDZ2QUh9u3Se7eXlLgrV6dBb9WM1vuv7DJ05iLU/vCwHuxLegkGM
5zkmgNPdtxmDUFgwSQGTdw2jGxI8f+ZW7b/AmHGl7KwuZS33PGFAm/lB4pT4d1RK/Gje/fwJWDPd
tyz2ne3PNmYDpKxXp8nQtAkm4GDgjCI0b2pXj3+pUmPCfKCmNH7/R1bweim98NtaRjIn/Efy7hHo
AL6A1nJ9vrljx4h+worYcc+ELUZYiroNbrq5A45kDGa2s2AZX0T+O980F51mqX0ZAMg+DZQhZcn9
Wl5D6Hrt7Q4TW5j8UYFYN0V2qVyIGwDJTIGsXNQ/bJECQ50owwXaKH8Gxx91To1l51yFYhrBDX3J
smSObwlXCD6tl13SthnAz+7kYxvTLT39OzC+0317S/V8LCd3UHIzggIRp0grwod2Hv+qJls9o3Zg
aRWUBv+/BPJyAiRHO6O09fczFSh+RZPYJ1ZYekLLRBFkzl9RfLQzcay7KTm9eAbcQYn3vtuYGyM3
XrfhYS18CykcA8DPCqvozRfRLLxGM8qBQXxP1o5lZr/RiHOaoN6k9qbEVIseYFnDL/QjKVW1NMS4
DX4XxcMYburOeCsn7K3LzYd2Tnb1LRm5eExB13Umu0cEV/uk2OcQBKNKO0uO6bF0qYRUE8bn2Zt3
xE7kxEKOu1yYBPGxOtOgKNAqIknesTD2txdCVoOmD4SEwwDmaovrqemq1olQUVmpH9GJyPHrCtnJ
EExkS0YSr25UrEa0iF6XrpHk5NSdsigiJ09HT2wKXta56M/27Jo7Ech62x88bTZxQE5i7VZfYl8c
QZWE5Fs+tfSafHtlMwxXeHnlOUdtbF+eAyBRASrJjgWMEa3UH6z5BwOv//JVKFr1aw31nTszAv4f
j44cNAVNSSr3gZxPMj/i7A+QnS85e6Ml8XG7g2YYrc1HJfIk9qONKSeTGxmRCIoozpXqF2CJQN+X
lm5MQ00/Luw96iRQ6lM6BsRZQeCVqCIwT6eY4N5WxZzzKHtpIgzwZT62xhkVvyoJFhFi3D9mE2Ot
mtCOhb+6ZGKoYaVGRtUaYY9K0vvH70bZrc3m9fTAAt3oB/ZUbabQswTRhVS/AR7WihUKATEHMw7d
T3F8BH88O++gRn5zfQDAqXOeIe+Zd6kuAX1gmw9bsmh9Jj6cfvVHpTZZcXcTqig9i2UJB2Sj2WWl
mMDch5f1Ml/l/BgHedz9nanuwa2H5AFYP9fSspBokdD8o5IgfvOP5625QkF14CmmHUPwZKy9hzcs
BRCe0fF3wWXeOUAERVGuYSZikBWa87hbL2nRdn+Db0lhCO70Wlv2Q6VVoYYyzi/goyF+Z5dVY0Cr
kOxwKAgk1rczHy1Ez1siFJtG4pJ3XBLFWgHOqCB5bUBRbjw9+2seVzjcLM2QsZjIQm+xzHgpJYWr
Za3C+dK4n0o0MI0qK0zQbbUp3hYYcKiy72Cn0zCfrhsHmvNxMgWTCvfTNwDMdtfnFPFt3E5+qjXI
2kmUG7+MFUnjlSxA7lQsPG1Rs4jTML5l4jlj/5f9k9PzmEbWNmNphETCC/RF/xwaV0na7Dhy0wMF
hoh3CGWojoW8t+Hjyyd0JYq8WbBzcitRaiHmb9dFS6pDpwr7UcIc0Npsl9eByJMtMtbY/LlhHUqi
8genAYx/P+paa3lvxPn4kgFsZurp3qjc70sz4wC53nwROcWHkTmdCsQiBX7wjOV57WLrunULqrFG
R4h7a8A+plYZk+bFyAf/lbEjGvP/VgT/wXvQ2D6iJfMFPHaF8frjI/LBzHq8f6nt2WrwwdwFrK2U
370Q5CzhrcUfI4DoUROXYewsJxZPWcAzwD7eGMMaGUV7+Rq4vKfrAE8HIUjaanUQrEIBAJQDh4cG
bMKDADjAreqW9LjVRp04C1IA3azx2VWa4nJm7ovCWpE9UhoBte4+tEJIESTvGOLZ43njJXtV9tI8
EAC/QCLbBX6NY+5vPhPuBuZGIKRd3NQDjwm99JA38pGVVSU457UPd/VoCiKmsU/64A0vqvTzenQA
MJd1xUg2gk3q9ZLzVLT/aOmmNG2gp+shPAWe9w6oOjdx9rsUXeqav9xV7JtxGyhYU6Uv4+i3T6V8
CLaPGBJx/ysVDUwdHqJbbIJCZEd0FHVYSTFSpVtslSfD24byfk9D2RHeGwLJrJz3WMcsrV/Q2jaC
NVFD52TBNpwMTKtanrJwd0TY6YFwrYhjHmVpJXciiR42oFsb1bwQw9JwfkhHOmuGRfimHqr+93yV
Bf6wtWvJMs7lLUuUMXG69QWkfojqm/uMUvYeuoryIk/wa1RZZJCxFcojNz3e2fZynBAX3GGEf9kp
ootcLJowgc6Oppxk3F0Aw+HVTZHf0w4cOOSdXm6k+vL2ePtjO+nX2i5JrWlP92Ca0+HuOTWkPMjU
RvppVzFZJPcXxN1i8BHtS3m7frrRWP3ZOoEGwPKwKNYYMz/tJt7iiyEB8d6xvSUnYrMI1q0GMlLU
W9P40LChzz4/OtYxrcv2wR0AbcjbRot9TdK7L68s14apYs0W3H2q3TlDI+dLHr9zUEAgavvPicbn
15Eowm7vInBAKT1nEpSD5hrmcP0pgwjfiLwUYcbI2iJtSdvM/8H9i7mb46qr5hksGpN8emRNslBN
poYCl0dFbEsyZquQCvGyeuWVqIjSLOSvfRYVtNLPHw22d0Ucfw0vaw4aTvJtxz7K1u8ftugNSRWY
/A8j6KRPJ96KYHIbccGrr74AEgnEqXcAiL4OzpOZK75k/21QECWCOuI7hDW5iSeCkcNzuOd4Gmnm
tzlk7eVQUXsaC98EDVNbDD+HGRBR93YA2sDeFzkC/4su0hL3kNKpNywdteSTq9VXEsidB4uSfH3+
2+feAdBLTgSUmEWJjWecvT/6HZWBcieIO4XT/a2wAZYAhrSsng3cYy0c1z5rAWMrm9kCeIFeOisI
dfYTj1ZzOJmh28GDBBF6NKTgWMTEHW8b2gGSwhaMEIw2gw24IxxFmWUE2ywX9u2HvSOtij4LwMF3
jAPthRt0W5WVmr2TXRJlXPxNUJ03mVyRJxTlg1h7I30ErJGVZAdHxIaueZUkV5RuCD2aRorpvb/a
LlQLtPzyRkl/uegxtPQfbfY4kk5xZXnJ28nHA/dtD9jmt1G/qMKhMkCn9PDdmOHp9aW7NgmJxDty
hMGDcY2nYl+3ycZjZVRSSR+M+x2GqOnV9zlQFUv1S0UxHK7W0E5br+q+0J9B7JCrGOIks38++O6k
p7OavwSkpNiON5d58rwMkgMM3QajlsRPJ1p2bAmSiN/tNdFsR7BMb8g1bLaHTYujI0NdVeMILS6A
bXUUkUFcUnEGR5j6ulFbzXPHqWYlyULviOIFMPK8eQe1sNyejhjfVWVZBo0A3LfHMHOzSoGclRMW
pKOrbdN33gOB0gySzMJT1k2MugJ7hLJ1vtADXDzJ4qu2NgUhi4fcTC04eM5jOJhYHdoSrq/SDA/J
+FhjOGZp+ltepdIxeBHi/JxgflNkRNV4W1cFescf586LREdpXMaaLVuREcvTBu9BpAU9wNUkFdOm
noFsjLTv0WzuBMic4iyPgHm0opywWSJ/71VonEzwQB4DNurq5hwijs+VIlKQq5/BONRpEksiHSXa
EemOhhoZfDM0M+cTFJYzOAm4m65ViquJaZnUA8oQoA0Lr8fMGzQ8Bevp3wsBSxiyt0pjc8pSeTWj
X22+sQ3G3Q6BPgRBnwRZXXIsi3hCT0OrD/HxjxBWdkGo2iqOyBxiWMN4invjzrq/I7MmQULka/YN
SWJCf+jOnOX/+AAltEopfZhGZoyTYRsuXshYaRJE6U7g66zAOp4pd9yMDaeDp3ZwmD4+CTX0oyY/
Bn0fWggaTxUQKOJSywNCt7ApL8z19xp2dKzEbCbKbFq3LrPx6eOpndrK9v+tODj9xhqvPt4SUFXx
UpV2IYZuj2y63W2oP/mX6Dz2JgivA0xEsLWMDqc6yscKTfOz3Grap38Tp/yhlZbk0Q6INvq4T5wr
FAk3GEtWQehmLivMqffgZfTfHS7pIhQepB/UJLZ6x0YjzaiDaaR44w/eHwdsdXD6wo3GIKwwKxjB
YR7P/FcGop82V4jziyqA6TaOg4Rhf4lMzV1DMJmWC+xFmHmJ09Qpc4Rh6KTj2XeJMlqE7iy6xZG6
uLeFPk9sQiCnAC2s/+Q+ebK5lVzbi/wt/hdEEp6fNINqrOh/Aj/K78NFwr9QmgDEebGm5taI2W6r
YpHfzSapGRObYytJPLJ3AW2uOrRz911VDIzSLg9j8mGvGbigY9no14BEcyjLOmR1oGNkRJqQaGKN
bQRo6jSf3AV4amhQmWs9z9vefsjaX4AE58SfeHdzPKr1ZLBxvSZjtHvbf3j8p0PpKumxscw6alw4
mkNuS1dHxrvcnPRMcL8Irk+MJTfXSBbPZPY7+VrUOkJNDQwXlTjffJRuuykeQgMGiBiOJJnwkZJE
WJBxh5yRcnVutPzuGRVJjkP+zXOaSwD8FBcBCOQ3qPCmobOZf3/l2SIsbrFIk29YzRXLn/gzAW2Z
b973NXmY5ngdArEbon7dilRspqYjAJjvXaChhJBPyxJ9qGDb3pF1BRl4C17UrNEMRc7u2EP6AblG
9HE7+917TIxs1sn+gjDkbzzDS4Irby7lgT8uL2ajkh7rOGopEkbekWqjqY/i/ffgL+FHq/tkhcu2
9NZVQG0t+U/eq5TIs7xr/I09QG8llMuNI6zxtkZbSDHBCeDS2g2KsFNXnSdmxw906sqQJJe8xYB2
n2fWbEIaoskKK0VAVHCRsut+lEaqtiVPy6BdeVmMpwI2tmy5UARpX41V4r00upYrXWF+cCJuXLdO
ySHn4HDlQrxqLzuHEiaCytAabWopzI3xX1XXQrL3FceRrClfZYFsw9Bah3IKCGbh/k4/GoOb/zgj
sEjVEYyt6gFYwACp5a/scRCv2b1nbxpoZL+uP/DBnuZQo3iw4FlrxY96gx+mdTQbZyaAvvtcMlej
kQMp0CaIScfsY3b8FiaAgT+Oz6PxdSoG3cTkGkQmi+uC646vClRof3Z1FwgVVNI5ZZ5wU/I8TzNH
tCyzI0O0Jc4sk/Zn6Ncyp7EYuWzLskxJSHM9dLbe9gZsvdFscKHQlS3xqsUd4wTjjkZdUKXzCi0Z
lWVA/PNrbKB7rI8+uPO+sIwfDjyytXJ/L4rqMBBw0KJm04t+WahuMCqjzEgMTnr8V6ZVocHKXy9k
VLCwvEHuJR0sAb0vO1/aDAdu/nSvgwLFrZ94mCsf5FazYkNEt+eE5cuLQXq/PrRPZaV1Gy2a7Ig0
Ch04OaZe5lrloBGkPLpFw4rwLyorVgKIMq8RyKu2bqGuFz/6F5EzYV29bPr9w1XG+S7x21zsw7YB
gl9K3NbgG2puQ5l+X1HylusxllzkaYjPoQNbQoIjInFSbNudhLkk0CVguAKV2Z7Bq923fFPvPpU5
omTVfg2RPMhxZ3DIE42dDrIt7l9DFskMNUC0KwFPFMMheqm7lMJP7kgCDzBS+gEXfZ8akx3tOn+w
HFcTuz6n29uZMB/i1k5W8NgOiRvsgmgsuflMrSaRAg88zU+f28v6DN8pKzCeXA6nzlXucfg/HKkX
Hr0LWU6GAZ3Ve1c5pNYje4cSRUMKSt4biGOnBD/ns1YnU4KB8HeY97Qjqz7RQIFziwRUi8AgHDjY
EH1ATmPaKqOavVKS2LyBWyzKDIjPygHwe95OXcf1cbq9zJCDFLmQAjbhbnw2DpoZ68uxRmlRLXHn
JVoooJqWuErKmUfty1E/5cmP1AWRR9/Q473jjkJ+hoIXfCzqYJDA4tI7ysO4HiXoEJ4iIt8Pk75T
RWbyZg4/3viXIPIwy0JoPnKGKGLVHaLMzT0tXXQ5B1KA0GPwe1UlFmvoaMhju6citUHs41PCVcP0
W/Zu1DtIHNH589Z3xf73eDuxPGPk7Yk1cH+NAiJ/ysEICIDpp4VwaVMcDHhKCFrw9Bj4AVtNBjAv
9CMjfnTp0pI1Ig9LKczA6VNeTNKHL+22ClC7LdT/zpvcGVR51QyJ9JhEVg7QZEzkz4NtNRu2jBrn
2MmZrH5Tinmw51UKYxYzOOfIajIsQuTh4zSpM+ph0ofaJNp2LnITsamwXej4OCCzMzfva1bfEPwt
0TffvZPFDhD0OsThDuHJMo7UOhgAmsRrVC7xQWEYdDOquVIojxFnEvlUSe0hNMryLfHIHdwG5nrA
qKjA96NtkbcoHqgKtRVFGviovAd/2id5IrD9MOkkjraA08qVfEazvAhZH7op9XlPeeT4MeF9GMCv
gCODTna2OE6xbGCGuKAVv/VT14VS5POyXknktZcn2vWU4KkgvYYcLcLvfjdQkA9bSbuS60n3sMZ1
Fv+bEw7XzPiT9QrZ5xGHuWYRqjmNcRMlFjoUZd2tTaXZ+XZmNS92b4p2wV6/nXuTj/8UG9ls2nE5
TVMCF9l2A1csj3FRDqKu+2Lp3zCMGg7BAKySaHcIaWbFnxvXq4LpJXudzvdqNr76XhBvMNJ8TW0s
Z/HKmpZa4m1QzhHPRh9sHCQTSFVZSdxarZEmJGYIXM9KLtZqJ0yPcALjUzJ9OZo1KnTPU/YMKzMY
0CurOtAP5optYA+1x0/7CDKkdkeAcnIsYItILdpOiz5QXaaRIaQCiROKCam0LQsjOiueWF7GEMyP
uyCHccfnV1cDn8shV8V1Wp7HxObLQDd1NYW03IlNNKwBBm8ZVaJgMKwU0kr+sWg3Aui4kbUZGYRz
d/3ytOT47oWvYRFRXd54umEuwHy6LC6N17xy71TMFgNmDFjhzzDEAVtfgcPbqY5Ng3DiyltLxBb1
9dNV1pRtFnP13zJ1bOmBad6elCfbzixIjMH9HlGgSfUj/lth/dSr0F5AqkGSY/exsjmzBTLIG7vt
eSrVe/mfVaF1MfpEbj5tmc6EITR+BLtp+4uuGt1EmtT4BaBkDneVUEjM35NmC3yoMjCmafR28zYU
9PSONipJKsgMX2GZ9dMVnNqwPC0mDFtXhq4pLj+12jeu3kllBfJytK2Jpstl4gH4alWMpq7zQjGB
+v0VoGbhtX38BTz40a7qO9qGrI2XBuRZkvjFCXfbPuVuJ1oxENUfZ7mNg22NqOY1oHH9NEYiXIT7
Kr6wVxVDVMHM6XDyT/3V5qWxqIKHzm8SrUr6qcizh+4xHddATXw2rjSBV5ODgvVBAyxbZYvzeGRN
YxiiJn2lNXVxyF3DeaYJ9eNVAfBr6+xyiZEEB2WUZaHaVLcI1Ef+WvCjo2qwZuM40Nl8vrk/M6jo
4PAY9Hu/UY9XJSmoAcI3AFctw8M7ZzrDS8LW01sWdzVoWSfw4pgjGYvRs0skfDV7BuiqpabsXtVr
3d/0r4KWUU1autXMv8NQfYRbFExnOzbLy5Wqw9hva7Pr2obP3O5qb9mDWQv5tqaM6tV1pYO9W/Xr
OCq6lo282//g6oWEqAMcDYaNtt+UO+h11hwIonYVt03MTfH9lVVPI3/bMtXuc+Ey/I1XW82flsSn
BkaGuKTXp6sdNx36tObYLKwxZ17EYsFPhbZTqpIHDX5YoLvvrdDZl44IHyy34cScP4CwLzUBQHur
hlLjNMIc+6nRuUFEzbF1zvD5SRPmGCvC5faYj+vyE7XWW7tTmipPJ9c4mWoREbY/wNO4iCzA4R0Y
rKds7pLvXYE/35m+zRZS88NLpwTH6ovQfaFKJKvtG+ZK00UFTuiN97vIZut2YJ3FMg56Pdc+nAwG
pnIqTSdehK7Et7WjMemE/steDQg4nKzpaZDVipTqawEgwneuH/CMBv9T8b8Na3641uJbBdF7YxIl
6d57e4qy+IlX+xJSGhfgKvWxrSeymSwzdzz1AE06Xi1q5GDH11qbjt0Bfyjecwb+higgOXmJQkZn
otUQyL8/VMvT8b7uOXuRYWikTQfkATpNyTv4EMWbZkJBHoFD0mPHW0+T2GiIQpKd6EgwQY+fNXMB
bzb1t1FYisRoNMVO5R37NlUQcj8LAh0aHZZ4huiw15yURNWU0ktmJYdZyZprcHAvFRa4NUyKC1ez
laCTM2wztiaJQZawvb3+7SCecxMTnEk5Qn5P0Dzc546205Nt6DOO6ll3YcN+s1sDSnE2m/g+KpOd
u8ettOqGAuVKa9AwtleayW09EzVTU9Zyc30s5WktBPdOXQnuQdqrPJObDj2Kwhy1WKwMUuwebMOA
eWbHX8li1VQherZ0qahbw0Jza6dGoiXG/oi48vHbcDN7N9SLbWDihkEy4MsusTCX5xZRZBoSqSeZ
GuAfS3sewjOlfKxVh6tFuRXYZOfSsk5wv+RXefB1P8UXq4EC9Rb0rXj++ypbgwH9mL6oizGdNr1y
OPI1amxM6wCiRCK+oZhs0J6erbax35L+aDzDcMBzusRRlBHmz7DF85hQCpUn8LTw6c7TKeOipEm2
A9R3h7krZGrhGuqXBOYy18sEaBRuc9P8C295fVBvlBUYNGJAoYQe+0ZlpjYJlwVwl13uKHWf+NgN
RzenkCPOGZ9ShsKcq7+8f5rNxTGmREIgtUgwqjgMW7QXH9yTRQL36YyKKGw52Un5FREXR7lsviuV
WOCqW3UUqNgXkj/WU4+KSFMt3XRLcPa0wtNK/IDDtkO0r1jMRmXxf5Fopj+pkwmLvILPBzXQbF2W
+qk0TfOgQklKerSXqkempvarnR0qEq00p+NQamh6txNRqxSehYYjZ6OY7UD6X5odSIRyA4qSeoyX
MpI0CpYR/dHn6ocds2qGKrDXpz11WzS4DWyKWgvD7EjAuhy789QUDqnlhqKF1yPcYldy0/3sc6/j
HIIlDlEu4WyO6I+ZOBuNMYYSpTDpPXzDRBYE5mIggacxsK0uGSl81zzV2nOF8SO8D6NaDWzRpE4C
LqqGxGw0DaWV0DqD+ai/hPPisMVrwoZfGEdZqpS8zpV3RbJogdEs+jp7OR9JGEyVo+7hnjEVYTPw
rDFSnFIfG/nj//VDySa1vKwfseNP/0s3seeS0xhQV2GX4Mnm3GAKFYMCZwSdkX4h/UXZn6/Sl+3Y
I1MDdNDwdagA2iJ0jKYU9OxL/xeR377IxMvuqRhL6Ms1HiPR6Y2WXa4ihMyyLi/zCkVOWpDF+j6K
HDCTJuMgudf2hkZeAMCcZS1KKeUGYycipfXKqf3lQ3wlb9RUtd40vJ2S8wvZzc/dYKnr6bId4LRw
3kVS7YgK8W1v2m7zxbVHfK+oq8AQYUkLPzDiwZludn5oUakqPgCh5jtdNo5O03p29non68kZ1Wpt
qoV7Ob1RAqAwtLwWe48tRDpRwp233Nfi4aTJ81BmZBl3D/9x9oY8z3qkkW9Odba/i6ycchioh8WT
es9TJBYEWyMUdtlfFZd5NHNNJHlrQFwrKU+xz86/IPfucteqMSOSxMAxl3Uk0qOeL1i2HivE20pZ
ki2NHPoElgjxcOb8Dq8SiAoast2QNOW/GhSUwWjBNmGHo7Q0ko/odl2vU1KD3O2VzgTc/XMGTE4d
zz7SMx6FpfCwn4WmeVX6tIY8PCJD6VNVJ/zaTxbhF5PMDVjwNVycab5fu68dryTQVCdiFgNjMg9I
0LU4Fsq0mFsbyfSFSzKkmslRp18awnCop9UKfSm87rfoRTkU/JwO0qeJP49IrMYZBkuLEsnIHb5I
/lprqFAOgSt5/cgNvdnN30HFQJE4YVGPgZEsnKOUvgMIV9QOkW6husReK8InPb04jtZpx6cFIDaj
98eJF1fPxBjfAw+1thlaUXPIqoAoX08w0VYdM4pB8SOj6kmuXOZdG9aGpYxixnvsMVSXY0+HaqSF
SKl5Tb6nwCrq9K8NJeGqGAKkVHLKThc2jBTAXHZahQkl74HDH66quG8tb8P7gsDhjC02t3rHWEm+
a20gOTFkWmq13j4ZWSDUoZEfMGTfPClhLXB345AagwSh6pvsu8mrx9OJG9TrdF7XpLig6kvIDbHT
D9YB+egVyLUsPOm58NmGkcsEP/FRSw6EDl97mkR4mWoV4xDvKb51WvUGJiy9o1U9XM21P40OpM2+
ukzcjLIE9yMCl4zPcU0xnCPP1/2Ey5kIXJLelbO/a4QLIrBgtqz1udgKFZukduW0lHvMkPz+8AbK
PVF0C9KDZUpYWm8GFE0InkYulwnOFgZloTMTSZjy7czX4hc1DQiWGmU8EwHY5Dh20g59l6SMguA9
OS4P6p1t02uctBNpShJTpm95gdRDe7+/pfOXaacaTv4ffHOIQPXN3sM1vmHeEpBXhTeXQ6BtZIBm
bbSi3WP7NhrQM2cYMgwyw4tYeE9nfDiLhmcG8kLSmIoCnC9V2yx1zqrNhMdC/ldNYzO+4vKE/uoa
dD5E45MRB9QjCb+XnHnoVsSRVVyh5Tvima9URRZUdoxUBYiSPv1a7N/a29UJCLJs/KBZUj0aQvks
I0A8veIUSlur/P76/+QNbL9ifevwogYB4UtUgNEz4Fo7IzI+LF8tyoq7dD5kIdFDZKqDanzFRT73
35F1ST6EO88lJdm8/i9egwhfeaZkCg8Y91O6s0nQfViDuuz8UpOgUiGP6mlotwcvQ8q6ewtK0G5Q
Xkhxs9lT0G+e93VobBJ7XhrqWwXtYwYsSVViFEGco1k/Ku5DpDMfp6iprN8Tyttl5RWxElYVDcNy
vNxC4yHjH5j5QCiYOlMU4ATPdwVGrt3rRZ5w4hyfiQf0N6eJ2LCy1suYNpiXkPIh1LnUvKPrC+MB
/babY58Ut+RDWyaLVvjcBMMtsp6hpilrNwUo3w2YozkBGTJu4A5QuRGa/5WsslO/MfDl09jop5zM
XwRimo8uz4Sm0Cxi4UazLMwRi+B6Pi0sa4qRS7WitD9Ds6vTNc+ftr+HD/7LZRtC0FElJd7rNARx
R1i/mP4mGjtpdiv7KyiuwmZxqLiqKLvBYd1BjLql7FFQKY+p1SGesxkLDudvsZq9A8QDCjPhDjth
gCPMIUx8DENdNbtXN/LVCgshUgHrSaCxUIEUkWe/4IznHo2Qwpt9FzKiirt84QhPd6R4TvcMX9K0
ZkKhlH1iAQhLDZD65tURhNA3vZhmsSOMB+Krr0HGOU0poIWM/7WB/MoJm23m/ZpVmE8yXiDixOB3
6FJPkT3xJmeocT2cj+d6PqxpunQaWf71/4ulIPvIVGwUF7nVsvcsjf0nTQaK8O5jMmimnXZI3a/X
QI7Khe5++0pE6FYofrVjVwxp2EY4oq4whDOMUxHIb0GVxZtqNq/xVy9pb281qQ8LRxXzz9W7WqeT
h5CeiiZ1miOX+UBMgpSF32/PbRnNc+NECbx0wkEyDEykw5kQzWH4PkmWN/19KvptCxh6Xob42jQq
JrHPTnm72P/EdYRHE6aVxF0K8SNGF0gGlNE7CRcIjwX/jISmwKMc2MLCoznMKLtcIv45lMFdeuvz
oDLrS0LGgEuxdY3JwZX/+6zT2UniF7RwT54ZTtFSx9nnbQGU9HHakuVrO/A+yrt4tbIOENouwLqz
3mLAOkBNkx76l3JLCuhqFWWfB1N97uZ5rMWVyfHdTDtKpqtnb/Yj1LeMHQQ5MWWzIP/4iuWM1wYv
b/n9uBhnOEFox+2jOyt13gFCM2e0qy22ra+ujw0W0paJfYhPjNjiz6zDa4LNua2mtdr8/YblQHGy
rGNJhOTvZ4qICpLTYh+OOgOkCEWZ5T7jQQ74zLGE0ZNkC7I3pbb78ftbkC7JEvO3q7oDUw9vlFJ5
a+Zm0RH99oiClcTuFzICdTO1KBPt9g9kIF/JLvBbn4aM9kv3IHSDK0NJCnsl5OdEF3oyiAo5pBlQ
Z+vvNWgisaxXj9QtLHcZc268okYaoasgDH+XI+THtwsJltGqXCHGkL5i6+iopmfJ2tha+Rm1t2kK
PGKg1i72bq2gqpbM0R//ayEIA8HW49qgj6XJUS6c6pn6JXcItFZd+u3IPpaohzi6fLeCvHrs5OMl
7DfvGMIIaqKVpWiecaSzbgzbrmzr4KSa3huCHJdOjkIBsVgnrLk2KpaT2/a89gzYa3pkcLBglCof
eCxZtpoi93sIzxHGKZrWqmIfv8lgrvzowJHLXdBQ7MYC9BkK3ghQpOsi2pXdIO1C7XRozsFPzxTy
WWVvN2vWTfYzaO0O2fnnoGrEPNkTVMRCOCVZMDQXF+uJ9Qregz5T167n6JDMwtbUYJIhXtkboraI
RyA/7fhmJ3Z9KfDrCjy0bANqlZy05ng2/vtTjuxGxLp6ak0b82HlyvihvDVK+H8WXkoXDBWCOfRb
hHBZ4jcbsbsuNYMbU84HLiqMoJYFB3bHLZ8dZv0k9PGILMF2Dy+v5ivyg9bSZeniSGTbC2kZ9P+2
jzo112K9mAwXbjcXe8yZgjv4NzAgrqjplZe6RmRgAyfU+XWQILYURiUKaM59gJTamO9BTDLfkoM6
jxDdgHIqXplYVesz/3WPbLIuINxeb5PkmQ5ivnF+pvDvHIUwGb57kpmfCaCcAdKk/rUfoJlUg8ZS
C9EMzX1nv0HuUQxDXCjGWM+BwSjK/7PwKrk4U4fYSj/wWpM8IcrZdV8x8rE8jSHHiAcw5RjYwOBd
qLk7MpSkyCPja6gNvW5+aKJ5OtDTg0Cug5MCdkoot6IfBozdUgIdsbWJbdu1QTPLCeSKN0lGCQAR
hoVdbgQ+JFcuzAbgDTZvNZmI15Z2KoLa7J/tJ4UJDdT/H+MnWjT7a6S6cHcRSsPyOPtIEi26vO7U
m9CAjlFr30a6wWwoMtCVEtQcmH4ifvUVGdPkWJQHSyvSwT+LhIHH+kTkCfcEUQ/SUrOfx0f8c+nM
e1G4VXqQrqX+WYvI43tRdpOrMkAJqG49YBq6Z+Lt1l1Y5NRXp7RGxoZ/GH46gV0ql4nJj7100Zhr
91oT0c7XlXLFgMA9jp+g+vDTwo0e1ONCu3jLjywo2Hyz4rjVaP/X0HU3IDNq3lrKTQaXAYsPPq19
Ap1i/TbPaYjZX0aYjeuf2WbBlYwe0WEtzAAlKLlCJY+Vcx4utu6aPX/LsTUMDBfgiOh3yzdnHGwS
x7uSgfe3JWn2PtHzTPMfIPgOHqGlSaWc0bcC6PPL+XsIddVZCKHWbwDBc1aVKi2A0HPtlj/5ZCLJ
ajEH13sw3t9tV6Iy/rn81GMLprO/h0TkgIEeyBXVbxPqRk1M3lCv2TXbVio05L5w8ZoUkgbdXRDn
JkQIakCrmSmPzLwcpdpUgaV0VRlOUg8hUCXDpOW/fhq9fHjzOzxe13rYkYaRByhxq+Sp5R36eksu
82iYHtzlPpnDgPwMCTXipxqNf1a1iAWKprg/1sJ2raEYof0CSBlCTaR3/hoO+qwQYc9BNIdDNSpg
NsMETIG5G9tNhK+a1zeAXnW8Fit6eUZfGu8P8zbTqYW9jL0XZ2kbkm4VmCuAEMnAi7oEaZIcXGOa
lW/dzJQ7G16750MKjFFnVuDAuSgt43n1sW3QKzyK309jauQiqu9Z/j8DHI53Tk/ldqtvZpOIhIeS
vcp6qw6ZCX7o9U0WrC0m9MD9KK+Ryk5oxMwPKetiduMZSzHgbVXJJ8Z6hfmUk6HjpI/p+GEFB0gJ
4hF6rIvNq4gB5ZRyxevBmyZ9A4EEMWLU+65Qxjg6T+fyiEThhcnSy34GyLxgbgKTQ1WZTtvuxjUZ
ce1xZDKkFZsSJlRVpKce/HA5PgXaXcAihVRWueyteaUBBVFGgqsZcr2oGwknmlx81rHnOANesVaW
3eWhPdFF6d1E3IiduW2wqjMQjalMRi29YSKzjqpCzRTasZqNjWBgwa1T8x/BXaAyyNi9kusfqaHV
LeW8RHO/WEKja001SgIHhIoP2EEYknDz70cD52Y25ggMk/CJfw9U0jl0wfOnVh562WCvovlYytj7
5SDZGQk3Kbb/M1Q2rhG65W6yisLuU9rAZeCjGZck47VJREfBcBsI0XpTCRHA/yJ6JLt8u1ZtUnjC
mmbnBjWtC/ucKKI5s+iCKUdII5yi1+hj4h9XD9y7wt/TvSTkpGUQKAHR0nZ2a4SM9NF5EeUo+jN2
bok=
`pragma protect end_protected
