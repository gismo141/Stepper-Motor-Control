// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
THeV3ijsCsW/X3roQaRSCcINdPaaiY2tIEseRqL9PRP18plWyUwUyL4AkqvfQDKL
MS7Fjo/Q/gmdCQb31zz9s9XT5xLHDBKfx75mHj/F7zMU9nFIct4V/hM0cbNfAh4K
eBDcU7rVLskQacMh9PMQRuhYe6HM+xe+GRDTrTDYR4Y=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17440)
71C/1pdE3bwBmP33Pt6+7ykwJ0VLQ8Sf461BtsX+z1H1VdfWMmZioKFF0AnJSjBV
g4w3KiyZa/HJeHnWiGVar3cHTjrgsw1+YsUGg+wF9idOo7Rc+cRCeuRWBpBppR98
/rF5Yl5ZmmKs3rMclrgBKF8yfbzEDS0kWKibQ0DViBf1tnJQWgJTjw24L+YENwyf
DnEAIQMEXH56ttxYMtMn3cRoITBhQzDIn3SZcZqL6Bw+R3XyCq5XMDkujb9MdQyW
pFNmFXHeXs/XpKmV4DEBQ5t8vgibTE8s18BTLbuqD/fbel7dEbWwNmMUHhnvzUBd
dBjrytX0wclIvvowicHzZyByjR6PbY0GO5B6UDLLtRhYcalgLoTHYp148891tVdh
JXSFEcezr1JlXwDil4Sfimhga07VD7MBdDkhdyR5Ocympqp0p2NDFYueuTwW90Kt
IOlY6E/Fub1Gz6PHyhY5zPtLPzwlUh5YIDIHey51qtjZbsMaFwmf+oLrzVQZAXp/
i8c0T+WPtH89RZJsfILOKVEm+VUdKz8QZzbvB0qBHCQo1AIoOJBFypL3TmPQEGw+
xW8pwWlMvFAHsU0lToo3rCvTBirk8k92ERKyrCiNHaNvZ0YGhvlmWP5JVSrf0i5q
Hmw59Rx/jAT4ep2m6Ed+yLNxDozCDFginKB1U5hj8l+qLi0uAqIlgAK3TldSCFTk
x5KroYg0rkNTZdBwRSGR9gGEFSNY2ifXbw3MajU7bKwYDNvQ9eSwOktD3BOvuQiB
sL3mQ6VAjIOue1mRxxAZOMnqPGUei3DbV3j1vsMZJ0Qi6Y7+8XXnUHFL1NhexAvm
NajTarH0Sr+ZIt1HcM+Mss7wUz2ZJS6aOPssLyAaM7iv7w7PCga9H5n5HPp65pTA
EYZap4ZF8t4OZs2Xu4iDRA6wZ1aNVEUpilTQOqIJjmmssLO6KY06vGx/WmSG5mZc
JhNxtnoS6WU2AqgjOFU7Y7D1sghXghZIvL+8uXjLN/iKwaAhBFDtFk5JRJcUJK1t
IRjEquppu9OTZ873rbmgLwLiKKKbGYPQW90U8WG4Z0dvgqhmtgBWBUzhFo6H/XPc
1qHDGAbgnpvtBs/xK+XHoIFuDYepy0w/ju/zLK3syumqXFWeMujQqhCNiZB92IPQ
sDO1HioeFGzBpYO6dy8IYVqpemJZ2i+vbFoREIoPuXQeZi+AWOBwrFis0e4mnfUC
BbQZOw5kcbNuzIMEsfUMBh5XQzFFNEu8fPcsOCr0cO+S4BGc3bsLQweBnjDyfLLU
3f6NeDD/Bfly/KiajzahrW4a8Pm7VMAKavjmWQ3mQyGphpaxSGsrkl2ittrvKpkZ
DwGnRZ1VK8TnhXMQHF0+6PyvOormXgBpLXYODlaHtINU5gDuy2DiKbinNxpp6QFg
3YNhdOYyv4w031Ns10S+0+xXx1Tu7rpWI7wicx+gzGCCPhjuLQpHXuJuvr6fJWqU
ONyFypxPCkST/JjAFsEF49H+e+3bTi4uOvrZ1I9GEdLw4xXOR0A2k+Yhub+wm013
m0U2TjCSNRneTScUhZwiQWAxXI5NjI53bPQbbYTqV7N5eGoZ93XPw4/YuboEY5VN
zdnuIaRuc0iGdBUN2XHdfonEZugV4n6MkMHJsRwl5Mx90Pd2onFNBKHE6R0L6fb8
Tr1ioqapEWemKi1YZejNSclg1GMD0VeoL3Z0lEKGswmdir37CAr9fOrhVKkZpYwv
PKyCVa1kEpgKn9QIc9k0eXZsEH+DQnQZb1SY1TQ7Aza/Nn8AtPYgu82FJyED11pU
NbfE7w3NV30DLx6/VCbDTG1PW9Lx9QFSXHDZm9DRaxKgyhzbgRqT++GFibg4cnhj
dKEbNbx499MzItuj4a7VzqcaMmD3Z0rqY12T/LuZ1VEXEi7FZVSgCw0p4rDGjePP
LhMSAuJW0Ud5o4CQMnjT+EluRWtslf3Nm6jFhK5DxyMCyAjg8KwH9JOvCQGw0Q7C
ZCBFzmsugtpOPsXkLtR49EGzEDrNr+HNBWv2VebmTBhaRgKd6yZHNY7oAgcQ4IVy
77Y6tds1aE5oPrOxEzvwKv+Sss8qtSes+FDq0vnh3FssHBS3V7oIzvmkb81P2ofh
hJiVAaQaKporxMIqDNNkVhoaF3n8FW8bm2i+DqQOqKLYmL5dfK38b4aIoa5Urw38
l6A9r52z+A2w7N30V6dPbplJtATjESwu80YHuNgT63JTqOseFju/Tj8bDyBBS80A
n5D9yb8QeilzNmel69dF2mELuy5pRxK3MRJRXFsemyPnkneS4TCq6LaxLReEOtvs
BqQUiYaAGsrts8Bo3aX8QBkxy+peBXt0HwWkfqdWMWWFC7GVzpEpqFeUEpjwmQGV
7zEpTQX62FhO2syLtrrjEg8UzVs83sSLSoV3FWgQTTXO3f8DfUiaLwdXfkSNMZB4
fIC2TyrTdydHJ2GZsWPqGtjdDOxvX88U0fv4e6+bnd2bnnHJUmsM7Pur6UcKWlHE
6tfainYaMsEfFC9p53lS24Gwve0OHkp4R8Crfv2WnYpzlAugNyG1ZrP33XSbPLnK
GmSHz6EBLk/ShcEM9NNOgKt9kw/1mb3IuEJbmrL7dOT8qfCcYBCq2membVfT8QZ6
RdH2AV5shYuuzE2WB6Ka4R/Q9nt+8y9tQJLg6Pf0sxdk0wbC97VDVOrDejD/RLs9
IAwCYotn5WFpsWcZtomYAROHa3hkz6SCH6CxNK9jPSw1WtmFcUmtoF41jQOfsj4J
9CJFSb4L9KXKfRnjuwApKAsT6lyjEIvLm3kmvBfECqeTBMlRHjyNA97i3FKYUqdQ
btiXv7Fsk6HKSeBcfl2hIsn405oISQW+efyFsPTHPgjXqyVwLt656WSLU0s7gx4p
ig6DyVTmngmzVpsxQP0TpMPgrX7zKfmJ/AbwHA9qGKQq1jQRvbIbNi6ik39kYz3Y
w2pZh6ZDhQemUMuiV6ZZD+mqmUf6CvEjbSlICpXNiUkc83jyv4Bbua8V1OY29zus
X9jxCmjqAJdHQqaAja8FKq5k3K5eIPWP7AoRFKFGm2AODdaWLHkJmFVm8S9gyzZI
dDgHdBzG1HWWBc0FDd0zL9bAGddSO1gT6m8zxI+qh/v8ZpX1Hxnz4K71CVDXPXwl
yk/J0cbsVhYM+Ow18mEnQ47py6+sguJusdbUgotmBJ4lT+sMTOkjgGkWklX0cPrc
c0NYrYV/xSV6DcdXW0LcWOlbgt5f7qVtBKYKQqOjXfLbQvUHfeUEcdvNEONKjdHQ
wAa5mIz2FSq8LroNcfF8kS4zJKsQe1qWrbsvgl6wUMHdQrwxqR492MfQjJgsykvd
FRHB7gC7eksoI6cU+cyat/HU3oIHBB1QY+GfyhyQTHWBJAgXlQRgMWTML2qFo3MV
PXogXcirCocia/61LWdvuH0VXm9Up221KRDCHPOnO1Axm5BBjfJzORCoIarSk9V0
yNhQKgQf8kbKDp3poHqEff/6duZNwxxs+nsVQqe1uB5UcZZfCw49srVqrmLYFzIB
90vGVFmpq3oyPA/rZ2X7fQc8bnXnAPBiG9IQ81+Bi6rxH2G675sU308MPUYDfwiZ
Q/+SVvhIo5kJymwDf/o2phkAPI135omQwyx5/LIdYhN2Y7x02GS52WD1I4tRgsiX
vcZvXUkj6LGqOpU6hPAQN+eTLVMQtRUR1tdHHWEmThxDxriilxYSL0O3jWzDp44n
47AuecxQwCbk9aLmFuhUkqWWjsz/pmsotoq9IMGZwM6lwyFnFqrMHzS8GZtBqUiO
vLHmCTI4NchXhvn4zNPHoNFK1BkFEf/0Nh0T/Tk7o5xigKzYVFdlMx3Oj83o6UwD
FQMxbq5KlVYMjJUGhc8izER4FyFSI/4UYc31AHQuc+gTZtWfCjQKTd2ywS1OO5Xk
9B4olNdp4uddrkiOEvJILcZB7pzfM+vq1TwOjDVSgMkzYcfSG4WWMF38JuTzM3M1
07rNww3kab/WeQqjD/TO2mpjPnRJtnc8D3ar6XjHs401P+GdS9a4EPzPFVl7wJ0S
D2r0Y5Ddh8qZLHL7A5FLKHNWbbPPjwlIENPgDFj/tpVXcQs3XvnJPCLz/N+I8fq1
UUgYZM9j6nNLYGA+D/DK58w/8eFB4TkG4jFwJvPUkXIb529bJq+XUjdrf7VaQ6rz
1ilG2RY/XvUjhnOS5aEOnfEizbBtCq4aDQQ5dD+FUDMesDONfocDiLozGd0iw60b
z62wBM7IOMa1IWnjjuuo5M1uZOPPTxblAU8ham4WShoJNS59H+dgdsccCOvt6YKT
xedYerTvFBMtIYe+8j8YxUMvYgfzR5cwG+N4HlxW5DEXxSk3dXJZr/YJzKE7OZHl
pfZCwrawRILqBYtMxvvh7WjbVpQn/Q0eyK25oCT+/owOiFhU+ZkkoTmEqeIAFcdz
0Eq6JSar6bXjDIqEwc71UJCZov2hi5VXTh0EVVe0uf4FroduyMslsQXiep+oUjmP
7Gt8CUL4KmlHOB4KLNimIZca8gb10aqWmYgmNJZTyM1a5/bp8h9znJvZ63Yoojnz
0/b11j/7u4HHtTJ/O1FPafKz/FcWhQHO+6/ObFM4fDrOo4WfamgwjGCYaVRFFJWh
FzZnBokP6lMWUgBGY3G3tXZN4gH77ZJUrWA01kdTyu6Q6nGcckv7Rziz7eo8POaV
zpaMCq8XfWYhPw/VSvH7IGoGbjLNSgiQRjiNU6bsW851mPCOaukbAnXcjGwgelqx
KmN1+uZSKnsAzVOj+Z0oU7IL3ZZ/31A3WWM3EzblSTAcUSVqOG6e5LtNs8IYCaM9
jKamXosKFb+xd28fHOxQkd9HTYndIDn/kJkwyb3vwUSO9CqoS8Q1WegcQIDWH7q1
UbbxGRvKdsEQWy6580aTOQH4PuXHvozS8CYy02ZWDjpmGvVdFR/qO0Ut0xHJMMxm
LHatIL6UmtQOZ1wlfwLzF/ZFIzPOkxl3ixA5b5cXsibp3w+mJerNv3Vg0/Fbl4Ld
+XwupcqhHhf86uWH64r0XaREX5XrPVoubXLsQk0N8f1LeZs++B8Un1c31vj+ugua
zNBD1IKLYy24j8F25dl63gMUM0XQ0ammo9tqa7igtxRd4afWYpFBWARWtHzfX8SK
fB73gugDuyPAfFo0ZxjmtfIswbXmgT4BYbtQjaDq6OTSu735iZMfleoHqW4Mo9U9
vVVJdf3c9aE7MAPTV+MhK6alN37lWI0rsU4qAPF+S33CoYd9CYST+pw5vh42hO8B
6M9rjDhiY9JZUViwa1nrrosSvcdpiM3MaVACSXGfA8euF38B+bvRFNgN06PwIxVr
5cie9DN+LiLyNsMtgvMxXXl/2wnQGlu90YqG3+fp5fOs9IuBf8kIVVRBs1gbFwnx
kEOaWebw638XinVUnwLIjBLSGODU2RQvBLSFSX2FcYkh5JHqbwkTlYi0JaJ6iFXK
N8Pr1HTD/Ba3Fo99tR/KmBgQoGsXBdnJL/mjyJrXbHaQxObJJwu6S3SjbG38cPeH
mj3vQmp6InfBghfzvmNbCpvMi9+yE3JiMPQEO9B3RydsuOViK9KkcbQddddOtsl7
4KNqIXiXtNoXw9WgUeDVE88u0NKuk0hNrdkzjuFuSAIbF8/4YZXhtZJd2qILowuV
1jffrbmFIqmtLcKGJUQn4zc2VriITzcbvBg9oUtJCpMD1jZMEOn7yfHPToO4K+Ru
VtVXRcv2hIpYLLdXG7q/mT3Htlby2AuqDvkb4GSpGBq5BwMbgdtC+e+iavpkZmb3
wYp/CJH/A78/WniqY6DNBjKYF9TNRXJQfmzwDLKFtYHOMQ9ZeUAjkMpmttF/IqTh
RLN3r2yAx6ArLCV6Jce29iUJWglwXeTDtd0CuwtfQ9WmCXTlisMDWTgnXu19Udpp
Kyju8tSaxmEkkl1tlMkGlYjycCRTlS/PSqG9ee2f+OZQhZV+4OdeZrV4O02eCO7D
PLFsyfEPome+LvF6FVgLO8yL9AtBt1/Lfs3kdOWwpp4co4Zj11YZRiATHuEZm1Jx
RGTnVsr7wsmYKCd2wZyCoHEk5nJStjmppKLZGN61rq1/nbcu6FBT4XjrWQvHP3ll
MlzlYSRcB/Kgux47caws3+u9A+71Y0TwzuUeFu7rKg6W5pfDwXePyIjSsSKwl3oi
O6Aivk/mX907GC6Nw0+ctJKfbpOtqoCoVbD+l4VrE956yfjCyLz+tv6E3b3lSpwv
1B+h8Btawz4pEe2KohflNC2Ta2pYeS7ObbW1mjHEIPvMv2Ijz0N0WbVHUr9Jz5Af
ey0LmMBcz9UnQaq+fYKP505vlaXgdtjEsIw0IwKLa03MDJa3SBZQXAkK6OIO+0rK
5gF9jy0xGqMQnNaRG9BczEpx6a7JqoR0bp6Lvaz/Nf6rQHv9FI61yOKREJKChqK3
iUpV5SRZ+qTyTpa1uc790Q1+8Hb1W5/9tuBRY7P6a9EgmClxQjEVKfeVw6lz8yZ7
Hl4Zq5za/S/ZH2yqrVKydBdYJz3QRlfV48aCA0wWjpKCItda6Cd+DgKycEGcHfGK
MTB9s/5/cPEwkc4jVcUOoeSA5M7rWPCwUv6AAwkx0ku39YQ7ac5sKihGtP8BWu7u
B+hva3uOz/2s88Gns0lHNs1s9Wxn0w1zpeiIWj0le1afa/+dJ3a8MXoUU6ly/w5n
THXHHQVzGIoBgQg/YU06tKAe7IFibfjM+nFHUrYiG2CsLNroggPT0Yv8B5JHE9RZ
gbT7U+2LKM4acNSx0K3YiBnDCEySDJ1RQO3drQZBVJJRqpcMelRDDW1IuTj8Iy3+
sx+X8gOkDahP3vX2HrPq6U4FfJjusoLUrAQsmzLAVG96iYFGlXxJyOarlisb4Cio
RNZqVDqdHQMMH66AXSzmy0Pt4eUyUljP6zdFYXR9hsYDZMNpILGqZD61S/FFrTUA
6XmH4Tmoted0WgVauaI7SdB2l9jb2zLSk6DLt4L9Y/n2kwvapDfyIZwV2SN0ytc3
cFeLPHDplB7d3kw/bCtis5DxpBm4K+kU+NMwwlYKybKUoUoQEiTQQ+5bqGE0HRBe
MdhCwqOzIcDnfY2ykS/PM6fGmE1FQRTk/fEFDvGjsHZvcuZB3Cav3Vc7Ka/kyfJV
MLwHZ54yFU3qCIge4zQjqbOK4fvDZoCOLOjOOMH+9W7AgNxg3s7M1mM/wt0ku3Wl
WGAesLpw8vsW9p4YYRhzDix7db/HB/QzBKPamHEcajZX0tWNSZNxoDeU1eju0TgY
a8b0tOPJdB8bxdjSeshj212hLDWSYahVTmMNIsBo97uBf8vWJ5BrQrWhI/0IGjXC
qikBGdRFeGDfkPSUz3/DGrVP3g09WDohNaF4IVglPAUepF65ZgovQ8ijSu/JFmJ9
2Xnqlw1EiMxhvywMkFTsK/vuupMi4bLhpJYXWuzExqr2dHkJ1ffW6yL719pSLVwM
RWC90KPZg4EF/clG320vqa2aN9YHW17vOT/Muea6w8zwyyBay0pdCu7iK+wL2Eqp
myRNn17r3PfKcZ3nsrUw1NSWrSF+okEftBRRDKf/9dosUTBzS67xZhjhq4gW/63M
171+TT0P/La3sqUYyFTSEit6znm84G4xfVVP3Z7QMb3vPk2hYXOy/fP30IMxF0mB
ujb8PLoXnSOCPMBSh6uC9UT10879jdv+H4SuWB86LKoxPIqET3V/HdqtuXdns5Z9
aNnE1Lp6CaK2VGews+iuddvGbm2K0+zs9/LIMI1sN5oFQS7rk9OGsgaf5iZYwsbH
uAjQyEl/EFVjWX4bw9pYnXbhuc2yPiwhP+iHs57MflbVucS1gB/yMJH4rQ9aCwJM
zPMROpZdIVP8ZU4cakFLZSuVbeaXH2y1jqUh2TeIsvv8NZ2KqVDGdBpHh/XCe4fi
j183iPXHAxnnii0gfMu0qE1LKCpEsKt1fY+KJayudPvugn1++YuOCPe4c6QUcRHl
9E8zEelEsSegHyyFdRDvyrG5Mg3mXzLxaU8CX+RTrzoVdON3OvPSUp+IPdpQQ9xx
BE3QrwGPqtt0iRAR3QiQq0WgOJcayye8gN0dHoF9yO8e/uqQJEt0yGcBbNDUVhdD
UlrYlvOHvNWLAgDFYIcwlvpr+0sKQhtkwkGTZN12BytnsaDy4xisDXVRBgBnPeRI
eVWaCQ1Yhz0Xl6Fx4nbvTzHJDwYaBqoeaeYq61Cb4YMZFGZWGqDkTJqLQuA5EVaQ
g0fT320FBxwiu8Aq4iTQiAXA6XoiPA+pDs5/LZmcO0ichKYqgflMfkrirNCaychA
FiNTuVFo48S5/V1AVOLjj2+8rZoKElBuf//ZC1uVF4d1d/lpFzGjTw/Vr9XassQ6
/9IMGjYOGFdMcL5evEiJ/OMcG5C/4Ozmf1swHn64gAhWAkU6dNzQXHl2wyHVVhbs
zJgKtfwCrh42105lPOjld3zHCYSdx+YAgildrrA1s8WNhX/HeLpgR33oQ+0gTcl9
ga6jklGqRKN26tiVIEk0lpLOZZAX++RAb2sS6tjibjcNMwT6iSxOXFTqJinpb/Yc
pevVyheRjTq5Q1jNQsKztyGrs0HsDKkMLP+mWr3a7Kw2mH3/L0LVDiOZ4mqDn3dM
v6hQ1QjeoyIhd2T1fJ6J5LF9dlK77uYYvJveXQrUCR2P4/oOhGkhtFwGMptXNC5F
0ti+sP1lf3Ynl7A4Yq5FU/JhZefCmI63e1v8MBtEYsGRP8a/n4k9I7H9ae3Fcr6n
NBYbqSjnWM7gRWDFRQlF5WR7Oi2ToeAL4qsMIGHs1Q2GF+b9siAj/BO4PSKyJz5E
hBgE8ErmJNhECTlL1AzQeNyutP1BuuPM2k+fLcl2wMMV+GV0QiVkVZuF5+od1Ffk
Dk4gqY4CTFY97PlJZWZ4UcNEc+HJefVqfNK7cwqrkHxSmJcDD1tVQfnqLVCEpLFg
OvE+FEtDw9tLQSXrXpxQJeKeDucr3hRiZRhpoO/wha5aX3ipGnrKHrnOtxfvbrgB
CuBG1v0S95yS2WlBHXe4wcj7WTCf8ha0HE9smMWqA61fcbdCZJUr0DyIRrjZfGtt
+VeGrJ7NXTSA6eYsR/lP6z++Aa3qqTob6jI70igYZ/GX5P1Pj5JqEBFB+aB+ltwp
pXEd7FPH7q2xIDlU9jjhF1clfBKQZJxroPAN/n8nf+kX9FOkbBdcGFY1fLgRLCFo
gCfmMsBwRWjAd4k8TiwK7itGR9tES7RkQMBQFHnhfSy8Zjd8WE3s+YlKsUQZcWbd
ep5C9HO/PAjyN3S7itrsaraM81dDdTgIzm+s+RtyY0o1wunGBrfI021J29jhJSAH
ubYgu2J9JkkEUvD8gZQDdCM1saEA8SBShkLgBF/J35Uj29QCnwicBVxwCfPh31Gm
0O8TkfFw4FuxOAPp4pw03w2D7h3wOPSZqPIxviW5b3hRYbYit2LoMSIZKuQSO6wR
Wl8MGljoKFDkIlUvkksFP6r3Fr0uaJxW0mu45/MV3qxVOgMXWo8ZvPi9k8rV8ReD
BElFrrRISx25uqfmqbKkGbxrxod52JgerU/NMDp2y0ZYLpMOjRjjJUtwhENHyllJ
ua1eoVmVPrTQmdIQg995ym3YNEGTc8QTRNfZ//IYCWIhNr7ialWFWQlcTkQ6N/zD
CFYVKuhuAlMqY/wAE657wcBDGo2uAPaVTL26sBOB7e8aRu5br/3qEJifZwcYfINY
9XHAq/yOSCsJLRdQpEZIgD5pIH7Pdds1ucWVfQml8HnzCor0S5OjfjdgeVtGhzjz
Inc6DzCmgxzLWxokZQll4XUU+1eo4RZccJqHZTRiOQG4Qbafz6QNTSW81eZwj0Ew
J1evbXc/YY+dw304ZHayEfVdlky2jbrPvan8zbUHW/kpoB+WPPzvVgjcK/dVfkha
oFbi6lQlxyUNEm47+oeFWV8BA4OhdsGweJekb94kMq/JprqQ00oOkOhNgSjxuxEj
q5GLVKeGmB56l+M0gfi/1Q7bxRF1JtueBpRAunCvm7E2QGY6ZLZWqPHTJs/VX20S
290CTsby74EfMZBB0iqef0LP/dh6inVch3hFVAkw9dEoB/dyaqMax9cOQJurLstG
EFc1vG4NaFQHmuMaFqc2Oukn/DFT5N1GC9KYDijUre8Pbdx1t4og81ogm4K15wCa
fyTO1dT0KIgCBVP/MAYLYdPdN29rp9UIYh4UKD51ABmMFcF7dWN/Ag7Yh+2kFY9R
i9wjLGG1BdMQdyFK9wtkHN1LusRz2KimfLy+ssxiXBgjgBHxYgURlQd8dL9F5y2Z
O8N2SflPcehZAwuNkEgOFlqKbMW8sTktuFqvHY1VGR/7ZekVq4f8n8SDyqWdB9Ga
Twi/zVFCE0voHq0uMJ9sNFmTptWC5EAe0j8Ujy5YWYwl+SB6TETvLOSQl5Kg7uvA
/XFt0ZcsYaiwwybEH4CO6I2bwGIchA8o3YLXv0RKuMw1VwQoCh9UyP6K2XXEqOC/
2h2el2myp/4WDCBUZ6m+qAHKUqxLVPnxemQKQWtOrXjVfRMo/iS4tO1foBEOXU/f
GlksxOdaL3fMwhwsW/Aa26+z72UTpp5K/aQ4P9SzT5CFIawbZ+D49kP5yYSHQ4/Q
9zz22+/wPlE+6NbIkH3JA85cV7zH3RC2vls16mNuct+vsYJF/fCvpqdQTlmH7HIN
Yq5jUrUusFm8SqyBr6QArz1zfJE856cYtrdUzHj6J4Qv4cbQdXzPisU2WDU+CDee
79mej8Wmqz9bVJLAnW88tg8TkSubrzaQBJNuxWcn1gQsRnIV7RAxqe27sKJ5n0qn
L73CPG6D2EKVdcyBg+eN2ZcEr2iZ81bCoBdtrzGreGz74t9BG8+SFspMkPLAFtZ8
twbN8I3IB6g4lW6GpYT7YCaFvITItmn2mf06QvR0RqamUc8keXK1DYW9G7odQSFt
+lld4yOu6R72Qfvi5BKSjuUxuj42j3WSYOb+RbB7MrwadHDQ5yN2lgBPVnu6wAA9
v5C/ld0VauDWfY5wp8kinUIq9VA0hwQPAoo6xkcpES0Gv7/rQWbfe0PVPGjrccUg
Qx4miwoiE99qxJ+4+QYnB843xZHxsn397yTc+c4z1jnEENVqAM9EheKYROJDW4RR
CFc8FfAOqMYeaP/a0xG0QeiZpUdAsaxf1IDmHkjSnVs+Vcd3VzsHaVYUrZB41qKU
JVuRUzI8gKN817F9e3SQWxetCi0Ozm1ApO6u7pndf8/hfozJZv8K+ud5NJkcd5qd
d97U88xp76rDYYxJrxgxI1TyJrzjdY2nLFvT7uvVcToIU5uhqzHSj8l+QGSCI+tC
Po/f4t69QsqqUbRJPAL/Rij5/9xQlRh6tj3ftfi13wPvcnSklvwJCDfBOOcUgSDb
4Sa8epTf4ptZ3mx9q7VZP8hQKQmQNchYvdUuMh/x0EnExvV+Z142RP8m2buwl1/C
g08NRuKpiN12/H+oNqljWFBM02PVQeAd+DeyS+zCdNaz7GxqNp4TLtxPDYIUQfaj
7Z0X+wQ56ZzpjzUqdk36AVyBr0YdQky1L/9FILKyHd3CqBxHwMGZimqQzeY1+2U4
aleD0CyKsMReeunq1liWp8vDvDzp2u1P68Lbrt8LOMmJ6LxUBJDvF4gWnwJf+f6G
6L+nOEz+6LTFRZX0UbtTpaPJyMGvXcoXEqyyiLH1dC39JOdMe7GO5qug4/FkWIka
J/VmMoVnDXUE1dKOEj8Xg46x43okisYwoJJRuJVbGkXQg3OoQau2CJCPa9VOY+Hj
kdIx0OgmcxzOE0hkdTSnetr2iI2kuU5SbwVe6bhvt69lfMzoZW+twTkMuqnkIXUE
ReDCpsZQkvbPqJuIQHazvzbMy2IpluPTYwDlTtq1mntjzfIfVYiczoWL2IY7DK7i
pQBWWw3r1P4Lf7t82V1FXN77AlJasWnl4OaDNeiopiM2yQ2eQMj/JgsalD9bR8Me
oDq3DJOk6wBXrDG6eF7w39pCRei80xFvIEWOdWZNUdOstkFOQK1OpdbsGCnuFASQ
L5l6zsbo8NYNSFjgsOrS2c1t4ICmMdVxG3476KV8lsXEN43C5cEkSFXLaNRVlmbx
xHCj9eiAj+RXujS/8++p6HYFUZPsTZiplaeTOitv1D6l0gfYeb3hF90GM2+GA9uC
fcunV+wqPgPXoJIGAkYjgJU8Gm71/FGeVykNYxUTO1zsM36puX4191G65pK3QKQW
cZ3E3w/r+w7oYC/PHwvD31g77QrgTzfhmVeQvBTiWFVJzw4y4xq4mXWtteiAesIT
+QECJI9WpVTNrYL1grQAJzsoZIu0ZvbbCvceqtsoIP/u7kiLUN/jmmNT/g56s4xx
CHt4Yq3aBMbb1dZ7hupKECgoAoOiHC1VKFaz0+1WOCShSZ9pp9dRo8eALcj1Zp0H
2AROJe0qfWml3Fof71nlF7GDawtYkwk1R79WDFxe6rhS9KpS647Vx8OvQwsBSqYL
JabmjghKMg+ETb9J7ey4po+5YGUT3v1NE1lHQlLq6sQA1b1l8YjC2anBrgf1HcHQ
i2WJjYwmWi/mqYiu5A/XZ6o2JvGCDGovAdkSuuLtqGr6lcqUb56AzT6midZKhBQS
3/pczWyUYfkhebtJ91KeftsPRxXKufIgB0oNS40g6hVpWs6HTuR5K2JfVWX9e16d
XFxnajIrhPrAuFtspBqYDrV2H2fkaxhxo94Rg7FggTilnGNMhu4bDgZ0yFg2fMst
KHFL1NscTW3xrwYz400KLpgNwZhWhqZxS60z1XU9vu5f4lE6uthb3xbytxpTm03q
LKnUhioZcdpGyMVVHHLX/O+dMNpE2qmzH43pkAc1x4IISxQeQlkYRAU6VO+gsZrQ
YMqQlpgNlJBXHOVyBMiuAgGyjyuRKVkhZbFuawpHq/u/WcJqO0uxPkcQ8ppdnoEf
lvI8C6fgmQ35/wRxBYBwcyNLwHD0p/TOCofw6RzEsI41voDXjtqHqdVFSVab1sZx
6FjELQaqpWvgjCybAlw1azylMt1Uu7AqSRsTdAIt5u8qCYLQRRBTP9ofOqRZN29U
0CrYsmxpVXQMhXGVYcM5vgPo8paxXi8raEMq3aM51eSes8qFqxeVOFIItvR1u9H3
wp47JcLmk8n4XYUfrfUkOyCuYd9bzdt21i9MBSzvABBkgnfu5p/qtjS51ejaMmvg
eKbNoIWDyN4LxV/a/kIg5A6xNHl56EtsKLYZnrlCDIn2BLoJuUC/qWTb+TqJveHg
arnaDz2WESaGNmrpJ4BDwy3wGJkQvPkPZWj24G5nMWi2Gv7TrGA8cyEKo9Csha1p
vOPutPpMHkNcAj9+q5hu580ocSmpsb4rl1d/CODA+Lzk3FecQwtcXrmmRfLXkBrT
AOEmAvGi+BoRP+ecK0z8JI0j4YWePPhRl9sThXBx+JCdG4Q9t9HUFHwEfLSWmM87
BL9pom0ujzIhNmvtnZcr61iaul7ei4xdsFQyJCfsOUZmxkcT8jajtczDplM/ha16
5fzXtyxuOQOeGnAxyX1pPJJ5c5OzJgOGZuY6OY7Z2+wv12DRMbjHfbU65fqC80D1
b8Ksewhad3X9C6oGnvVUZ9nIkfH3VlyLtRBb/7rF7lswENYmawn2X2rZRMNMgK+8
brU6bf4/dewQ1UnJ01dyONSqu54BeN9Gwq3BRiXpNZgomJOF8QjenVYgU8yqfp/w
n9Kx6jwYex7uddPNnqCLSmvlYjKegl34LoOFE76jwKY1rw9F5UlwHcBZXqoLZtPm
WOq31zWQJdIvC1dXBEf6tr6N4v+fjq8QKlpOHXNmi5skj5Ff3Ki0sHzoGKlsqUTk
g1UBscYpsDVYGQPeHqPwzua2Ut4jDWp8Su3UggBBoT0cBYvvNfCPVAIj5f47BnjX
LMX9kbUfgqGHuPSYs5sLzPxq/tphzbI2IFS04lFogmISLcHZbhqYNZjtBJgnqoBz
so2nYJr0DTn8ctf1dDZnE48sBHycjvTvIf9m1kMix2IviYJ9JFtF1VHE73wU7Im4
U0d7BkuCnUzACllHTJgW/l7+Z/Wow/XhrmAUFDWSFk5mkLtPUWtyyqoTlvxLG3r1
Fu4ng6ro18+B09DPiOl9EgTehwtzzOC/jppsjTw2YjZFpwRzoEfAd5tVhn7ez7c6
qzMTsup1xVLm86ElKXQMobkf5N/yXPV+F7DJIU3mVCfwBAgtqALE8h+snstbQ1t5
PQijfC/ihJj6Le7QTm5H06NQOVqmOuYUcBoz3sDP0glAAtRIadplCTIsfaQRjvwF
vlKaflQXhFCUs5GDgBLth6VOXxXD/jDsJIyLcm++npAdWKzD2pl4K+Yu0lZVwYTY
c3dw6BPBx6WPeqL5FkK72XBmDqSxxLqlQRh4sxqJStYXDwFvtxMfkRQxPUttccLI
aUzAKQG+Ty1R+hijPlHAVtXFK4d5T1oKUIZsOPCtH09gzGvhQalORxKAhrkI9Cb5
Y35SdoUygVit04oQ3zerrdlY0a6Bb4jZDT917a3Cz9Y8CzW19uJJ2gmVHDkuGsnp
kPyxDJHuYdo1q3kqtfJQQ6dkCLJZokANtfB3D/8CnXyzQFr6ZVdpeLgnea3Ld60Z
iGiOdW8ET/tZ2gZ22BgttWHIyRKdXR3/GMXF3A89krdJtmZBbHaMkW4OPVYIbCQ5
OtR4ATrOmHWgNZO32qid6YFiNRcvnnyNEjgC+04xPniQc16r+g3L+1rtghfMnKn5
Rdh4s1S9C+AiMfrlAsa53aLvgJcwgw3VnL619tgeY8IOt45kSEqTRa2t1XF2ANTL
pFWAAHjKGkFbaUZmLz8KZi+vHI5kPmUY+sKXolQz/63VE0VSJ3QFx62Ur0QBM+xI
dUyBo47ZP7ZUmj0H9vjpbMinUlLsZv5Y6xqUP2w/HJ5pLsr4KAaZh30TEB5FHT1L
H3Rmfa5C9V6w0Mg56kwvqx8uYee+8EvWJiwg4x0cNVt2zJLF3PU8RoNMTh0qf7+v
NowxNzb4oW10Jpw3T8UFYGgk30xLyQTEAjrZsS2TlmNVoP4riL5GUTeLvQ5P7Fwf
5TWXCHKjCViR/8eY4QddtGkNMYhR9QDn7izYJ3oOF7PvS2qf+lCZChXZcBHNOaOt
DO/FaFaYR+6tSMihT4n84LbdX8QGFyU8cmI85nthS6X6/pUd1OL41ldJwqTQhYVO
CGNfs0Xd7emqMq2ccfuyssWn/G36atmo7AkX+/X/KWohCQJzijIeqjYOPq+bLcM6
9DYalhWFvbBwsYzA3h6wTmuqSmqla94HGXkbkg5IKfNFQEFshA2mtJRfGJQs4ITz
4bjhVAx0s52PUWdYea5BeGmo6zSQqtGGn2XsfynGcEnQx/1qvYkM2bB/MgaYl499
JcqyEhXaISfJYHkhZ0q4Xc2nBl/zz1CKzdO1wFSmd2LuFnwqVHs3ah6EbLSJAdQr
vhMlvUq+CiTMSlTZhHUy5Yh3ROaoGfmlHmn2r9Xvf3N5hQ4fwQOzlnZOF8twr9Sy
GDvn7Yp/xBbnbGtWefW+bXeZ6gBNmMA/gWE96JG7zEJHc3NbB6TyWRrCIdE7ajeb
S14Eh2EKBXNuVsOCLInoHRLwejRb+N+3Ce4MCujooQQb9bgzJ8XV7m5c9Duy/fKY
gjLQfieRF5xWvtX9KOHQZf6OYY6aVXEoOCb72QBKA2nnt229nt44Yfc2pzEQ2vnh
oG8HBLOAiz4awCgoTS3FcPnLxpspzu6ogpQ6v2KLguGdeuu6/NNmiEJ7T6Jezo4A
YMV1r/6p5dHzUoOCtJqk6DKWi15fyz9AmzWfjaMUyZUmioFk93vZSrCbbgugHv+H
wWrrqiexZBVhLu6xtKWWd6BBgk1cv8xmfIXKaIquixyR8b3nCnQOy1t5zm9706Xd
lLjWWwl+Ol2eByZkEP0Q7IwItoiiATKnsZV//S5y7tfw6QMQoSzUUFeX+IFNMS9r
aWfXbroyDVMIXcq73nC5cea9/65rKS2/Cte6auVobIDZJuiWbqx9nhdm6WqzgFqZ
mmrmPlk9Rhs5uMeZAwlQGlc14wVL1c/rjPuB/X9tBLy/ZHc9DvsIGnhDGHloPreF
+yprDAM2LrtI3QiPZJMsFG1FfwJZSlAVDIB8IXB2r/hffawa+HD66318fGQcf0sK
w5/HmFkMSE7wwOpDOKyyVpv2qCuRu9BShjovOED4CfsPTIxLmOUDUXUbD7zmkMhM
FfrKJ6V8HFaPtNxDp0e06tzpw6L5yvioOa0OOsUqqKmG08aaDad0NoJnNgzBRtaN
I+3yX6/NOdIDG15R1rtYVK8Gz6MPc6qUGgGEWOiTmJ+k6FxsNXPak0gPx2Hv3xbD
7lX7ua25/CKRcbeW8gqjyS5a3Ny39LTB24WdEyOv9HDcukW7WT9gmL4KEXPL9X+X
C46BAGCdd8g3Ss9uVfptAYi+dbynfTwOTLXhEZ2iHuP+l+15sMxjiMyVhDFwuiQt
h5S9k+MdyFfal3oZWEiyDHLwElkpqJ8XQPX9M6wVJGuKpJ4QRyr9B6ZfKuUgFsQc
3ewXY38eGVJx1RTstEKd+UiBtRv8RulteGNTpfyRkiJQCQjxQQG28FMgwTScIhFi
hy5I4zf5ryykCzMRxyfvYP7EI7Vh3zSU0czCHm3zjbPqNI1S6kxd6PioE+xQEdN9
PAyc41StDIeB+nXk34/bFFZCCW3WFpf0spsCzOi3E+cPlbxC4uzJQoCZcQmgfwGe
7WOlR3WhhLcP/MhAEfXWi37jzH/k9IF4rjFcVAIrNNZE5ty6klA83sw+eWvAxmTt
JPMtkJC6yuKHbP2lFVIzzsuFN0NQRu0RfLcCwpus84bTAwhSPTQl8L4fVqcdtHQQ
ZZROqLL1H6oh+0jMrD20yHVXiZytb8L+vpqfXHnJbztYGnuvKgB5mUiusKXH97CW
Eek7kjWGyCSasLG+4skQZ81g30h/vT2pftcbgs3Rtcr2hnoIM1aODZ/Q3eFKCPTv
fM410LVdCLLkbmh9CLJW7dka7FQR3G9ke37CGQKj9q7+SG+U8MBt5JYCtl7Jwqud
WtUVoyujSQcn/w9U/WK/kiY7Olm9pdRm7Abi+QApjVYEOD2RKEc6jEiaHnCXr0DG
XNvsoX3D2ctecQK26JIW78YcwG+ZpGz9CancRiTzCwD9nIKyvw7sGP4ZhLYEmAJS
6RrdyaFT+9IoVPfW9swJ56D9nxB5ZVXrjLzzO9vRqZwdWf/vb6pGvon1zssUJ5vK
2fB7VZEbRnHszUzHlAYK7730oUKBL0cMTI0ChmnNiD/NPzP+Arhwmfex/H+hpd0V
Gt3NsbE+IxLy/DHGkRkbaaMshvX/Q1EyFDxr4Oa1rDjei/NWabAhsxLFn7XbnhxQ
gPjO+K1j/Y7yxuUSvwqVyWRUw0EWry2J5ko9oqgWlJ+CXarISnbhlT6MVTuI36UG
Pk0bjNHlB3N7H5iHBtvyOlTVK1MTXUFkVJXP5ENaXeln+q0AngSZIW2YS+3fBcY6
kXyZiZtCz1If0br3nnk9It6Qxvu/M4oIFDmZJHPTJHjWxFL/AGJb6F+UDNFXUoJi
QDkQ/gpKmeAmGGX63sBGLwdkgIIkYdX3a7tGs/Gommtn1L6p5SdkOroo8pz3swFr
/NiCSiIeqrdwmbE5S2oAIfzgvF1KV23jRmcel2KZlXwCHpknhL1+K+aCbLv67tq+
Rq38SWkRJNbtQEImumLqSJjGMCnBneTOqSdFERUf+HWr2iWzgduvxSJPy0Ak0Ba0
Py749Hfv8dMJOnz0HPjolybLzyAgId1nX4zeCiMfWDURZgpiNls9/hgLBTw1UvS9
ItiD7f0zX2hk1yR//jXBZsvoteO2eY6qfsdYU2GwJ8POa1CxIbYrwMUyK3e65Kk4
YIJzWAnUYtx/+lrLt8L3Sm7OZe/xBIYcwHaqxVFaffye9OH+qgv6ulwM6F/ADiTe
9OowH1KW9OiqLS/ORXFBPwfbEe+nfdWqFpsHK5dog34FMJkzvRfJ3wZQqXf/a3R5
vuyypgG+rEQGU+0Ffh4smr00v6Vi8bWz4pDeRmG4k++9+A+0rSHTU6DTCiZ6tQcD
FarbiHvh4HilJTligGU+9N/rZuiWjvrcS2ekTTo9StBNfPUyOuw7k1/M3xD4Qik6
N8P6ZPZwDnu8ply4PMZ/kTvHuZ4eqSVMKqtedkyYSCZ8vowyI0zoEWXsQsqWdExr
woDJUJaW10PfmXhoyxdsgJNyJr2epeJcGlQ1zv9U0fGR1gO1V87tGdNItmIpo1m7
EsIqO+1uxXP9l6VtFA1lZBX7x/HkKE9o2pfKE99+UoTXqV8e4OLUIN4yzAWCLhd5
iEvdQ9HQOhg6DwImBlzVeV9mxdBP4Lmlz3y+z3NC8wYQCv+Cv2E2F0jCKHkUlFmp
0hbfeLAPgalwrTTp84avWjzaEZZpQGBWTv2EuDnsBDkaHf/v4eyeDlcQdvtuFJMH
ab/4DVmTK8pymnl69K6OEbh1PRwQBST63QAqBXH/BzGrWynkCsGhm84WEPdcMSxB
AxKZB21z/6unwq0CuFalk6/SiXHfcblrb4SLJPuXchK8w0Ie1c+Pdz+b4pU8GcxB
WhjpT0r8bFs8W5/dtrTJFx8r+psMbZdg3307SJIA9pU4I0aO+iEaTqioNnSCzeml
2uT2xUu6iHPxkirUlLLbcjmoowQzlN+DWgKABQxBV1Db8cVHldScRqWeEfuMhiM8
FmMD+OTqpn5wMAnmuDqNypo572UKxMNSZ1OfUO/Ny0dAxdLL136GPdeTnHZNgT16
J1ZWUc2kvoGaOQfAW45FuD6193t0LayabxrSnMGPAWpL2nmTBPLKePqTb1Kt0IPI
r9CzVKhsqomxeFYHi+mRAyZ/oF9pvFdqtBOe5ETFXirfL8xS/RRxz9u0vLIMru9y
yK+pj8142v6zI6n6NOiufxa5fHjU3xnluYjVfoq6q1nIS8K9CYBouq2OluL5w+sT
1SG/I/TbJono7k8YOeMwxOBHzGo5cgxv5Ka6pF/CMF3Ws4v6c3CjhZ2SojepS50p
8zMXsCrFlB75EyN0C3SqXh6f6ocNuIPwUR89pUl/fkq1bwmiR8D41Eqm0ExtjtOH
rk9D5+EmFi8G3Sfdt7GYpuzn9FP/DbCj2CoHk58k+Z6kqJpv694KR0GeTIhTGEwF
/Msv9Sq3ZXUCBWdCzUHYtmTY9r7R9YdyLQPQwkXbJiKWVnz/HUe78pHz6wmXCcVQ
mlppYK8ARyhOiSgMkCasatADctwUwm7ql+1hHSEK4FHUweg2xXbT3vHHOocw1P/5
HSryrQLYaut474+hQ7P3pxH+/t7ixKhpU4KRMWFTcOSkLeA50hx2xxQuWNdUkW1v
Hek5kXVrarqkzhA2nEEbkI8p/BoP7n42lz/BKEIVUDVm5vh5t2OKDvaUb3btn1dg
KKMwe+Nuoi20G/liJk16HashbpMDcgUdWqJZoP8NDtW/LgCBAemAn6VozmaGeSu3
4cus4RzyoXc6JUX55QkjUb+FU8Uvh2k18EiXfWrV5Kf5Vq/Z6NBuVh9c8XkZgo4F
ipjYquJSGvtPWA2AuleYavtxDO3MwoQHRhhDjEnC03dXKQGQyZHKW+5VZAx43vrs
l3+czt892Jr3++LuW/YcNtME9MSG/eZEgV4lsH8icO1FmFWDhB15n9c241QZulMH
/SLdb7aGZl+3xOcSsbV83ZwASqHT5RR3/tjQ/KheuZBp+v+vp889GZtblA5bL+4J
g9Q91mlAM3Pf4Joi3FYKWXq90Ltxu7dVOHdAWEOXDp6SXAjSsftjmBqX1QvkjnBx
iRpzHaefx6w+xBhoRGcUVyamzj9pgiQX6m+Vc5kXTFCh+khO3R+PnwZDP4acwThC
cGwI1VV5sazw5MDW9ZtMbD7b/N9GCX/7oLTVtNuBHDDMuZHwzGvyU5JjEU+lNi0v
gMEURNO7kLQJX0OS9JnOE0K6CepYx0Vze9DOAr5RG79AefxDzSUD10oEMkaHI0tI
c604Q5Wzl3z2FOIjkzsTka+zNbaICObk7f4vZXgJaEg8VNizyPBYTyr8VG37n3eW
pRZagpknuQ3TJW5Z1aHZRUJ0HKwsP/yitULnJYVWbrWKoF7b5uNzS10FCvOCFqi7
pAnQOmvkjz6xdtDR/TC8mtY6tOa+8BN++Qrqb+tvCq0VO+8TYP2vr7FULyhbiQQ1
eFkRmTM78xv0NwW0PCzUUzz7Y87xrEueoehiXbXd4MSOxdRmsWakrjgMN1Et1Tqr
NFvVB/wu85Ax29pihEt8dRKWoDbXOWd7x2MCsUpRRYH2A3FQ2+kvPTwyDfMXz/o8
7JEZ+BovEfXA/2PAF37WbPk37e3zQTxxleTvZRybgvuNNCrbrtDlD6azc4ylgLvY
p2OebdyhjEglXElmCFrWrihmrV3cnyqEcnINmr92sWykP/cKvEsigd+2iuF/3P/c
uASXPkieAshENt9py+D+VkVl0QbySXtRHgXKbgckSeMH2aDt7RqLC219xOG5x4kn
te6BiEDMWElQgDmgrmFzXyZIRWkrP8zyBsIDKMqPRdq1tK22M7jQVywC9cxKnI/4
enxWgcub+hnozY9wnHY9hRZfjLFNT/a7u8fgJRIMHZbzXFCzyqDShcMzugDOYhAX
tYhwvtEtCFoNiFgbT2ehXEAsf49cU7D51YWOmjVJ0UGuHLas0R0xn2LEUSCf+YyC
udrCTDs+o/YRCP4LtmvueL2mOu9hcgAo1RZzzWuMxYxUnHHDli18IdJjvhse/xTM
rN6mRYSrKJMhjSPiEdX1Qg9u/4bs2DC+oasn3GrdSWPySYbHVkpTC4Nv9hYvfBHk
ngVYPjTYtdhMSa1FRYZgu+Lc8obEfujiy5XFIFoi+A0EeIQIJ2GrLP5ZazdtRMd7
rJHlA4Pn8gKJIBOYq1fVF3dejnAEqgZyL+e0nga5H8YzYsu8LB/8sc/LyMEQrhgC
/gs9/U2/fSe9fZz5CNsLOudVOTGx8hMjMCn5GG+VN27LsNWNaxgRBog7xkAPNWXq
odPQFRPCgWZWwfps0yjRw6c0DiHXkaYXJOORsyop54S2uJ8OCr5TV/JaJEPAAAgx
kmfPb0Mr7vJrq2qDN5VAPBFupCYO2oo8z2lOWD440zrlhNBqgygGq+MR+oTP6DVN
w7Z9b2dLaMweevqylfbaiInd8+aEdiPRqy11ilsz9Ow9GK5gwX0HLpNgWPfmSIg8
W5rjMpGQD1fjfW+Kl1Pp+3QryGrIbSXf6NCrv0dwczIoQ8OeWpTJq6R5R3zhaSSl
sNkJGVYcs3FjcvXW9IiqW8dvYX2i3RUh4jPTpNMp0O/sfw+3oXPPerl9ojVTLV6+
yoiiFCJ7HaSctLwbroCsmwLId6o9LwehkBL0nU7EMIj8eqsetTejFpiw3qSBOfBf
9pppDhBEcoxl10OQFOcOucuo6yB8apiOM9KTJunyxCpqoWGyyXiPY3+rgpi+dVJs
c1lZGq3ZeTpAOCpuendApPTyoK9PxVxNBgkWYwcegFCc9H+XojdE/nQ3exXidiOf
AiDiDkRTCRvlDKZMpFEgT+oIHWN/4KYNNmV+7bf09b0OZfynk9eNm7BDGIdQ2hCa
J3zvoj4zGexwnDCB4/ELLqrdCLblR2d+GwJNjMmFKyHCKmHL7YEuz/+c7Y9pzQwe
wXPujAt2n9yAxhbfEkwNJAtUbHkaUYaA7pynZmXjP1RKqkLPp5YgwquRjOR4pJ6d
H4j5KepwKVSgpZEYSKhO5zCHnQomXtbKwQrLt2Moco0sR+unM0RtD9H7YlejOnoM
qTSLyCUgBh+ROQQf8S0ROos4D4Ggg7SvJHs9pSHVHI9arWyqFbd6iflqzEQAM8A5
OoaKQuNui5eSZPhWyFn510NirkKmRTCDwwycs7TK2p4oHIgdCaj704coKhYLEfkz
+jj8EXCinWDqdnCfNIcastuX1yaDXxksN6n6+/MN0mbHfvoHkHIf+ORSA6ZLwwqF
k4Ksx/MB3wp+hIWoqMpdYn8pPnxxCqNF/p8JbtnUmJsBK7L/+ie7HcAbbb1VjtXp
apvbgk2z8Xs9lZm0NtATSAcztcKJdRKOrCkBUVa2q3cClVI5cSBr4kN8B63YMwXV
vtz5bonk2YTH/pZbLSSNavjXOHHpZT32DEcQPzzEjrRSuAxy5PB0ImgWxCc/rkmG
INoIfGqBEkLqdIeB03Tz0HOyQe1e5iLxPbpqZ+aUH36nhm0+Maser5OuJj5U6KDu
yTyAgm2vIjR2whoBFQZK4C3kwkkV9MlkIDLXP/WK6Bw5X5WiwJYcCcf1ZT/wEDRS
wJj8+g9d/lItBjf7hZrUJjB3I1KM7t4s4ctygkR3T/ndYp7KeCzLWh+JDjMAXrbW
Y9qOB0X/d5OICK+5nCMzLgFRytNQ1CrBlUYf79odOHqaIhtWhThcphZFnfIjNxgt
/ExrERHkDx6pRvI0p2crH134szpKWmxvUEzf7ZhI1ZG2BfuMWbQ7Ue1HCoOUEso9
fEinHT5+Bx7MYmd9TCCqYzEf181wcGhMwkptyKVHyCkYc+6P6YpfewiMAi/eVy8E
kOwJZYdIXWxvWR13cJhyl8LUgLni+nUKdz3zXffkCBkYFWILG0CcltZFuhkRosAj
p/XWrkbZdrkfILF3a56vCVTR7hD19R5B8YvQFKAUD9AMxQVk45zQyB82SJ0efUPy
853FUKPQ1HWhBKaQKN5iNRkCYdTKcmqzYYX+vFxj7cgHgTxIo57o6ZuZzkM3G5i6
98UzJvFG247psuctjzi0L6qwLOZ+USXBI1ykZ4V9zQEObuoBYRLseSzQGF89rjIb
CnrZsqqUTsZPv3RESCcoVr/x3P4WIXcBRAtkqOUaJCW8aoX+xlxfPPwGmV9q9cCE
kL/M1CoNMkW3UMWM2dKPgYc58fRXjJC7KX4G+i3hT/gAaYZYclNm9qHMuWJjo5TC
FVNeWmvHkSf+2UoZelDkqK/rEfHjToz1npvxg8Mpcxsar76qberKmM7OAUhJVNHk
qZyqss5Ft/l2+O7b5g3OX/U42/4y1cOu4E1MMaFdbkDTOziR5/oh8i2jOpWvGtdh
1N8QsJUDs1xtKWV3EwFXspOt7pSeUrR1SwcEeFSMF0P9blIZL+OEGyhUJO+aHtNc
Z30yth9qocq5RqoHRp5bid07gMJi5FbBHJ3j7qBMMZbY3LIGWfFMCw9+BdNK15vi
mQS9uVzciTHfJIjyiFgOmHH2gr1SLbiiCz9AUNGe70FTHUd8jD8O7jsi2IrpzuLK
4O4ZYxoj7Xl5ooBSa/6YQfiQ2dzwtVyYgMgSyAAUu1V5xlQL6/xICCJIcrPs35+m
8Q1n5BDijcdHFMOXvdNwKA==
`pragma protect end_protected
