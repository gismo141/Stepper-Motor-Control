// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NT5KiYp1FguUlB26s6pypL0KY+mWm39+EFyK18IbMITKWtfQedDCsHdZIr+42bK+pOgaV1E/+7hM
NjrrnyyUGybI8YYhHmVPS26e1xudqmQq4UXcFNKjGb3fInWM3Fobz3Sep7fq+6nksTwCSvSE3V+B
hXEFpk26fPaD7hEvatUivlijMA7dhG9qszttDNMDSiB/yBT1K5JnM0nIJFpXGSkHmB+EhMFGG5V7
yWJfvoTyr5ZJ4g8+C0y9uXPqcx1vqFUelds/KA7l8InI4kBdMArNUXocRnyOLn0wTYXt3rPzLNuh
shsAY070wcWOo3O9wux2HcdjNF63+Qdw/zBKDg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
5hcHUhPXyPpkmQ2BLVJ1Dggujc5SLvl3oGMgFrh8wieqFzEe++eNtdrMQHgZJRBT4dr/iNjDmMF6
5udfnT1HL8qXsI/8hBNHo/+ZbCJZUOKeKtUw/Wp/Q3eObD4d1NVPImiaK6EuFfnGGJdwKys8I3ir
VZO+l5ayEH+5FWu1F2x+h/j24hAUyh/Afa6FG376CAkxOt9y/Obzfm5ZtDGU1VIxv5iYc4pv6zOa
ysZVN1wBMMxeMs7hrsiz7XgkQ3VuIWivPOdExtt2lTvFgaLzOoHt38m0ndgXgjBELFl1Hi2HJxqM
0T5yCwg+KMtu+XWN/+fuBSwNYLev5lksB4s+sNgk38CThWaEfdERDlXfm8hipQk7muFNFjZ47no8
4wh/uEgntWxQmRhvRl6FdHd7KdjLepxjzL9ecf6lajEM8ArwOOhyHGss77HWU5F2hUDDNBfPSidg
mIoHdpo0nHG3jnuBIcV8OiT3o/t13fYIV65LcqBzaBWJxH06zGmFHaAVWPhoZHWxseb1D2/HVjKi
4sCxZYr/ovE8B2TxX6Ct2T5/oMblo6FSks12hG1zgafVvak7VDoN5T3/nVmjEqhlVOEnGNlLIFTm
ewqKodb/UuSTT5Q4XOu67oc4i2RsofoDXylbBavirUU6TdMaBC1MrdHvUhHJFJ5bSJAlZzlGccOG
5biUz5UocHlyMv4pngrVnpjzGgkhFFKK4dSAYfNcjiTPA5q6kcYtlK41cQrDE8rVXcCEP1PQN5FK
z9d2FZjrri5hUuQqt4wcbSqy9RUPVoTQy8JibQn7ySFTftppDgsfXnH/eXH5Abyl6y4H6RKJI/l5
IqvvU2kJgxF4oQBJkO4FkMxTuNo8nkDmGAA6r3RKTry+cfgAfbTatfebZvzcILlYb11tO7GRKhtj
O52AKWocS2akTaL1ueK8lzI1cwB8Wpg0RK8JjLAKCwL6RKqTJxsWVuT/y7eKEeJE8DB48zg5HYnJ
Z9vdYMBuu316xqRU/JPU0RjjuHyh59WWdNYa60xnxMXmum77gDSo1GuTHQUcW3QyUmOmHU9H1B9q
3rVSXGA8Z3HFz4xDlBAPZDQ7vRHsD5ln7+8usas2vW61hD53KnmYikRmoCnnauBN+cqeiUo4BzVh
MH2wkEHpmdx19cF77K9lrkAXyePMzfl/b9D/j6Oac258qGCFxdn+0lW/VFGuYp8csaUNyajRKppg
/HpKPn911Kyf3BzUGWGCxu5/5KSYwbSxWBqJQO27v/b9Z2ffNZC3BvsdbSk833FGE+jmiex4hrSh
6Hb5epy1Wjy3H3UHrHJrg/6bDbLldjAshizwRJuGn/TYRMZLNq1SxNLznQ29cfxTCUYlXlcBMCha
JpbVHdN8/FSqo5Z5GdPTAQSNomMKZBS5Oer+TC84c5kIvMUU8gXULEU4UJ7vr/YK6XjwRqPzL/Kh
uF57TNlnWE6m3+O9Mp1rokUeW0TlIyFgRqTdpx93Pt8RDz7gm5s2dvAmglz8NdkfsnMq+Iw54X3C
gQq8QR0y4ypVUsf6lGksVUb5wkPPlzwObViUzmWIs2N3x/mKEfU1uQbhrn2KPMdMkiH8egDSyFrj
rTXeyXflzRaii7CWwvhrD8K7I/d2k4SIU4yCKeY7oZP1RlHYUesT/1hkmCAVMrcSTR1gA5fUMwil
ikAVusG798boqhu0kzxtA9arM4Ip22p81d95X2M9BEQtLC/LYUfUO9iEaHvdYZfTLDqiIybrBzmR
Lh9wwlsttgAZVU89wa+SySnzm/OLKVJfAuSHjOoZ001A8eScCX7MuWWdHg2QVz/oGeQMuPLpt7Ak
Ywtf2IjVxABQrWKairsj/1r809DJ1q86nmgVF7o+7groTCLrTbaI4kWyMANrsm3o7Wn2kNaT7btt
zEoKu9d/D9/6EYdYPFETrVWuhMYV5RsU/BdILGfbun6YxJRehQ/KnkkMnA0NqRfRJMmOQYCksTEf
aw29Xf0XQDigUXvjF6QtfvB8ttUpoAy235FmKkDrTiyEinRkzxtIkCEj8LJu/R4NlGbcMRF6Azqa
S90yd3PtBs/VbUyfcKeLJLef4dqCQC/fEiHFrW7nV99zDuBg5g1wYmAngIOt5FxobKZjchPms14b
ebAYphDSmy+fIqeVIJ2a0bplKAOPwEk6TrQbe1q/lhzUBsysJfBsDDYGvr+PWYbtxciYyRkF8S1W
P063j9qwmr+Ol+6MoIcTWOedfZt8pgBRyqNoG6EfpsI4/LLUJ2BY1QUhqBuZANFMwb7kaS/toKxF
4IFjsAYFwNt9Sch/OB586285Au6xU376lqn6kFLpIbbWCwiBtEFc6+1p7VUT9+BKNCvRa0w1zj0N
aSweKaqGHwRyV8+TfdAHGiMIWvI5gMm7Rg7ScEWOdPu5dBrC9yP1nlS7MCWm852HdEiidZ7k+u4U
m+kQ1u4eWEB/thjxbnZfJf26BsPBqzAS2b+7bSU7jmqtkyJEQNXg4SRUFNpxD7KyTNbZr1v6lSLY
rr1ETqa1rNBA4HzIkwK74TVI2KN18yHr6YgXWbXYM7gTCkPhsncuXW4SlWVYfDQ6kco0foORYX8d
jDWftLLxNAwTVxcEJcNjD1GvWTe6vM8+GrarbrQS8r6s5dix+eh1k9OaWy4khQzzKTMZytausmH0
aH2dhaDo/B1BoLZ3p66U96Fbj1siGAWY9PYAfkQWaQ3oetXOpoy/YfuDWuaA2sR3pfYKlaLDAgqg
iUBCNSi9v88erikGmubfkGUI8ESPKtTqab5puGEszzdbCzBF98VLA8QHfoBowIF4/h+xvVby7+V7
QafSeY6HBfJBj1aF7EXg5Kjvh/rz2rIthMbjQ56sMVKDu1maGkGBxnXcrfTXKVbYjk6v8AP+y88T
HulK8a9CBI8lrzfDFwsnGRaCuZbSDA+vNk0fF8J45jp6oBJOYvg1QVPtEX+yZTIZv7UkrGli2nVS
bw8ycPlJcAdwi0/jFTH4uUnQVFGuvjwsjxfWT1c4vydtNjq6+wIyrXct7ZNhq9Ek9iV5LB87hUtR
rPbpiwo2KEtqTTGJk0Bg0uApX22OhFbQg+LbZlhduucr7lAnUmcyPXAOb+VcWu5z5UumeR5pwYR8
9Szk/hPZ5q8BKPM4lbencjXG4b+xOHEoEn921cCZc7SPQwXn28msUp1RCLYN07zHkZuRyz6Vl4Aa
MOEBR5vzp9oN7o46iLOP6un6M3YVekl4sXcBKF6xL/BPiAZGScmkGs+a7DBIoo5VNHXM82AtQaZU
WPE/dKjdg+bVY+3lrfV1S2OckaXvKl0IPzpEAH+qqNlZdp2Bk0oEIhwunpDjyQJxTZVB1p8xrNj4
3xXhoHjBBt+kzRRhw94sGbWHQJBuTxQRq/U2iwsBO5FgdV46jX1GS2CBcndiTNpMND5NNjVGaAWE
IQGwDMBkmlmx37Ms6XoN9cY5ZeB2djJxSVfdkEhwcji3OCbfkVqpUYAL+y27woH6OE+0TGjsn9KE
XuJrD47K4P8vNfaXRdKFF4zxaKN6WV28PsgWmmNwL1rOSx3srqjW+iWMWBVVcvzxIhjf/cXWWbs3
f5Y8eKpvgwyquDI8vWRFYnhLMi+HT5niXEH0K9WCS4yEIOGokiHYntFKmsnvOkwoRy8ed0cjtaOD
Ofnlit5CfSrjp+HAz4ca4fXLK5LTHMC66Q1e4M97c/p1fiJYPoezkGwsNMuVw+Am51g3xev1qnmd
VQnlUZoRsRK42BYQ6bYUb26/y0bj2FsT2cHv+IfcgBn6I7KtoqAVEv8p6c8XnRbMBB4WIR5liCGj
TZoSTJ3YjqGki+NDvX/ZFJAaAbLNpR6qZV1+qlDJNd0/WE8wlO/OMS3mMoOJpM/H4HBtmxmE3O2a
JSFcAKx+NVbwt2/23m+gKbDkI9yE4nbtyxGASodjFRf9qO1TQ0uYQrR0am1zY8KpoP3k58thFC8G
vpW1ghqbgqCMjaIGrHZ29M8R42j4c7SSoX14YXDazay2GvAHHrWLCTSk0bYf5JdLDtDMgTqKIoqQ
uw5fvcHCCzI0ejuo4w067Cl0RdvZwykUL8lUxaus0XbEq7cI4F6x5hKIR4V9o4yAYJEFpgg8g0ww
pbYElhQMEEOM7WkoOEm8Pdu4QlCyF2XGLxgt6Vy/3i1do0Wnpfb05vVQGxpNKs2m8LYXbQYu5dhp
mI4ZRQ5Rd2WnFV4qD5/s7SUMXXYE7ZOXilW6Fr5FtqhkGoi1dhcur4S02xo7ZeX++gpYrNUtnDVp
Eb2OrNUTr9wr+lPsMf06tSGw8szEh34EDriHA8d8wPJX0BGXoUWNhrdKbmsRS2CMZK7B+bYubZbt
8UNk/9OY5qnUznfaCQv0MbWx3IdYZzbM+zaCgz9w/gLvej+N3TqZamzY8rKOPgoeY/tA5Np7HVIq
f/h6oXht7vRv59qIqUgm0z8Nl4Zw5zqP7UnPW5jstczeJkrcLJMkTY7qsZWADKqLlJMQYTKacjN0
Uny3RQ40sTEMGNR9aSd+R4SeDDfodJuVR1bwohS+v0i9wi3gao1EtiG9ZEs0zWfllgPW6yyx1hYa
oSlyilLCOyl6ZXIt0DV2zRizzwYugfFkBjeus449Wi9VzOOfP91LceD1VsHB7lAruMS/TfEAT29W
EnEW+YbWY9yzQ154vzPvOvDWQnLlh1ViP5OuIgvgXXnQ3sPAgQ8oUwMWffqsYmR0vYRxyIu27i9P
NY+TPXL2/NZv6mBZAa9J/dtf4e8iCziI5oFkhUSah0QmBPhfodfAaouUa40wd6qyWOG7URes/zy3
YL/UZC/Z3qpRyraFjEZkQ2+iswlAnnHzB9tT6aATZceVz/J71wpotRflI3OUfdDtXtwMERjzUpMQ
w23CKGYx/P5qXXodbfaFqZbIQ6GDbOvl0Btehs37hJeRPI5lWA1FM/bv/Zfd31+YY1vFQ6xUFKDM
YijIUtcVDlD4gS4sUd7byNNNSGNznG5qNS5AzHVOXMVNrwXAw1KgLkvxDCQzGnycIWhiOmmJ2V7k
gsQWA7KnBmoiHwNPE9bVV6I8StvpRRltjFb3eHZZE3B3P5FYu81ajdrgpEh02fmXJ3NBFPplyXH0
gq4EJwq2qYjLtN2WiabYi78k4QHGWcnZT80P0t/yMN6kQzxiUkL1Fdsd/WWHwh14qI2JFSpF7a+8
wzxPH/h2Fa76T7oTkIy/7epT++BVT9FHr1s5p4ur4ZeE/M5ijfDzpeauIkI/fnO6ETSQr0O0WbCs
3t1cOX86hdhDarntRB6+oHyNFOZDOsXcsCGQodIW1Xj9wXSjQ89Y5diF7RmmRnBX9AQVe3rPhiVL
1+RbSMAQQSOYvobW3bD1zLmTxNtLJXQlYTeAPSiQHpZRQB/CKk06hnAtmscVnmCZO1MguRFumgHn
pkE+FXIR4h5AoxqagYI8Vc6V+Bps8Ym4LVvVtibGT7ZJoyy8YyWHV9wXe4LS/MiZUwK7c/699eq7
PwiG4gt0tsODAXr69XcwwSzaY20GS7Mi78FS4ULNePLgSezczSyrseMMqftSnoGyvy7I2zORYh61
s6UR1dEPnMMXhJAmYvhvYHCWg4lDCKjJZ4UeisSW3R441fCjiQogaHgIcRaYv8ccAww3bCVijdl9
ujlAyEGG/C5AsG0oGfPdv6NLNv9n0Acxd562hlpSAbEHquf2OJKNY79nuoIAcPetw/FUnziut1mf
GN5dHOSZEegn+REzyRUmAlOyos32smTMOrRoi1pGV9RumJnAdnwA4zBqEbkTXGaYWXnppYKqv5jO
Rik6uVwsaDM/SseB8MRTPO+ExshRD3uPGSOe8GCPLgM+rgReUMjhSiSoQLvVkxaUK8t72tgWKDlX
j6edTEq77YRR211dwdCJcl1FUhOIHn4yd8HJT6BA01OPJOOZXpGB9d7H1ypaO1I9qHb4XfelLgeF
7M5Fhu5kRHyMNs77jp1Y+SO2XtaIWUNUyObmeS7TW+5Wvyye4ukdlsuBUOZVNFUAhOMi42vLByVi
mlwVSK5woi8DVNCJ/yuy1WmsfL84Q7ZSNmbLcD2qYu79D/inHbQl+DxNKqklJJEyoqZQ44lo0Twy
lZOBVpFpQemZdKu+fuLhaZONDKi9FMXI3Py9hcgXXWA3XyyrzRbqOdwmSnJBOf+hRqIBkKzVhjZR
VYEdJyzoNyGw285RWboykA+MM26w79TmDpNpk/SyB9BB7tLLF6qLIiNN+C+q3v0YmqoAVrEWddI4
3AnkbTznRuH4GdqXC4qAOWG9ZMJR+oxJfQnLwm84uKiHDaW8HsAqxAUEzQNRzYmXm5qZqSyS7tg+
Lard8c9xxTtYZ9YZxMbjCNlHNCaZXTvTb/K8b82dHmOLoCFcKwqVhlOt3c10GjB93fXjVosNHaL+
4zNjax/V9V3x0sdNoCLn+VOIqZU5CoFLhDTNN6+AckG9CTDil2VMMdO/Or2scNeKUDGd/2j1UbN3
d7p80Tg/aA++YN8alYMSR3H8lY32CcC6xlMxRfVSzhf0RP4JZiUyToru73ospo5vHtuwNdhatS92
GVodQWAmNpAw/qruplwYQnMRzEvH7LjiiRwFV5YEBZempPZc7LcMm5OLzfXch/yy6idlADjHtlRK
4Vu6Cb/xlwFpQWHoA8TmNLB0EF9DNauPIujH/ebLkvghWkDPtcJgNiJ061UMDkKBSXsGQpBESxMg
cl2gKkt/m/xblaH/gn0WUHlaxfrFaipn9MXu2fglEfCLmpRtiaiE7YBKKMy6CVeW5Q772LB3WmfI
3bUKsl79eazvLHKydJDT225Txx8WaN0Fr3L0y7Y9tCHUq3ThFOrDnNRlffIdU3spTp4D1/j/skYb
3/ZNz//O3JeirpzMCHK5R1BRJjoPV5upxyp1erfD3qjkrv/eM6LQk5vjyVijHUTDckYOWtv0rWJv
n1NObFApNKsLLDgfLi+BWrEedJJ2FxQXraNtvUgJY2xZOIGiTzdOnzQsw4W+uKKm0F5geqq8nlnB
Qt5axKdS6wCR5V6bZsOajnTDf5Fmi0k/hHZHNoPumw3uBu8qVsONrPDbXBWyl3w9gLZH7JzIEv5H
giNJr7Y5wqO0iD3sauoo6q/6Mey+ri8ciBLOgT9ehCQMX8inElpPdK22+0Me37cgIZH+wshlc/Gp
Hu/cRZaid+L5sA7QgiDUjdoePTpDVev2JTxWNgM5OlD1YU4Jx8G7XAgxOoICZGBQ7qJwmuwsuidd
706uHJhoA/xlhkJj05Mlxj2+ivzyCH17c10fYOhSMgWqxYf4mHD3bYdd4XQN+wgq1THIkqTloJQP
f/YEc8JRKQWgfcmGeNA6UdnV0Ou15hjqRCUzNqSFqiPwt78FkvYl2eyzB3V3dddlCx1FheaEl9kg
gXkoD2Qdr2VXhclwQX7O85cgnXP2RhUc4MPHFZ/R2bgMN9gwrNS59TL9Mkq4X3fGESi+GJ/4hxj/
UxLDyKd4ie87ULjHlqHFlmIGWPOQPoU3+etBoMiSc34i9qVSakP1U2islcp+E8WlhMon2Nh1qKnt
H5yLvhwY0Dr3lLrioLkMKTHUaj9mWpnH11OMrKDfrs4aqxGaytsHOR4MbWWcR1drnHSUdm544OA5
NPkHyiVF7ftaPlf+0gyMurwUjKuatNC/epLgMheZU2JuxSrdYaVwJIZZ5tTN4tUauAtXUPC/fOMD
9BhPHrSkBMOFWL/25V27DyX2hxstJK/GMKDfXZVVH6zVTJROIoJQsciUS2GRjRDCsfaucT1VqsHZ
23JSdYwVvAPSGZ4SpTg5nHfdXWN9mb9bz8v6CipkpsNxf45QLC90FZpkiTzWHDV+EZB3WZ0f+nT+
Mi3ypgHuXMuNSorvWWiAk20nKFoVSGcjUg3UIo4wyW/xjjsGTXQlPaYBivttYyhq/Qw024jP1GHR
fXMbUO/IkiBEPlqDpf+w+zJBpEquV8x2BjdfZ/B1ubo/6kQ6PrBWcYe03xebgaqNauEHOkEW7xgP
PifSldgr9k/Fd1kOB3JMLGVlsxlPH/UnbXZMOhaukvi52rS8xGr7j+QWldHMCO5mPvGXGdxucXdv
p/uscgdiBBZlOod70oXEV5OamaA7QpaLaMCBEXRenQfYYHzSmVerP9RxyjdD4WOGUWxuedWmLIBp
NK5ddbV5AraWLuRlpELzFUuyN2OyyvucBJvueZN1VBhXruzw9728KMUclB/a2/lzzZnR848W/f2F
dxFBs1C+l31RI2ird1nS8o0BsPIKB7RRV7HiwHk7n0i4aTQopZpnx2zgJ9rAwye8A27vCyFQwjfq
1HP+m6m90upB836urMuW/K1RFwHbP7/2ilnlU0YllAx7izQHGCHddiCt0w7OOKKwUG7/pZTrP/aW
6eMFl/ursQ3ZVMU2/lVl4FFxHgudItprDTyZmABQrngPThn3GstO4aGIjxRiB7DrjNlnA6O0D0Wi
5S9t+Dc/q2p0yksKI1DrlBBj51sUXsxcVgwBrXwmsGXoZpAP17wi0GY4Sx6Vvrg/Rg5tLL1HlAuT
1v11tVaYqq8TLNtYDX0/k8XYN++v+qqLDE4LtXSpKSulTCLGh5u+VTOxAV/aXvPJTf8631Swia/W
Y2lT6zOOW92pUD3G7Mqt/QwNLMudw+aYgTjE5Blqd4uksWVahDyrLQDGiKB4EnoGApW0BoC66BWn
Kxf85CRR1qCrBLBSYayrE+xOayMSeLf+Hq584qguj+dlDfAx+MwxjtMCOz25Bns1bd6a2DvXF0wQ
uP4pRR+rukR/pvC0D6Kmh2P6B3jmLL/3d+kw1aQgA0NFpzC3U173NnajSnSXDrDOX9eLbArhEbcX
cOnZmCQGOIV0KZS6JDbiXyc6a0Wu+NOfxRJqit2BFEAIcZWnmbPd7ueGRZ2xoV7gPJ8hYy5JtJ/c
yhc6tmFMMPYpvTtHDcaB+QB4U5do1b1scP4Z9B3Fd090yhEEqGQTVmNy2RTMTcvhRQYMz6tnQmBo
KYvtjBZvYxlTdj4fuXcPdSFz6EX/BwiGcR7wceGpq3BPEVdDTs/VNDSrVEdw/4t9p2/ERXQ6eptn
qqPxqlqSKDyVwbzoxwtyVVNpJIX8WM0LpS05cPNppeLCyS7qdUhBQP4t2GyTDLSkBmbmZelptgVM
NYiA1mlxVbOgDYndXU6IxentbUlkfNf6HlozcmdOUV86bhyTrd5pMT82RYKb+D7IaaQMGMD2R7BD
nZW9Ks7UhHWyAocZmXIPX7kV/vZMRUUQ9I7CWfJXCkYH3phi9abAT+vkBL3Lx/598D/ptDHUpbFi
FiLbDWE/QbccjKaRTIKHLrtIRL6AGmytq9aZ6JA/U+sTX0VIKGfBakCS+tMfDqNH9xaFEC8XqPhy
FxRTPJutsDII4RFoKw9748rE62d9juymhvKqA92S8KIcXIFaef6zMvwArfM3GjmtBAZ+lWLgC6BK
3WtDvjHADXqj3WwUcMtXsFr7PMNXBIDHtyfV5h/Z5vaxbu/tiA2Bt9qjRZAy+5jLjNvMvKHj+Rmq
wy+ZhJa/gRp0p9ZIszOqc1GYBygeAmLvT0c+VsTpDBtcXVR34+hwo2weDqKe6jqPQglIgPEPs/5V
3J3eRW7MjkC4HQAMwbJBWsAaEBWTj+kVeHztHZrfsGFyMezYG62hhAHOYD3C2tLwZYXKVxkHWPw6
Oyv9ddkPuAJC8dUY39/4GGeBb5qVlfoC550dwMl3UXFqY50eXhTBntO4OqxbM++8ObN3FZapcnmj
yrA6PW6IIbTFdfFNO3PBUm6OOSALhzSqG6nFdgbLFztnqT+L8NHKnFU666b0p9k+wRQ7WBLpyatd
tG9ehalMwriNQ+V+P9lXWCoUxez2v7ybFvE9fhHrkkspHWE1hH5YaKWZo174EgwN7cAuna7zTfJZ
HJ+BKsGb9fg9cIeB7W5hXNLfO1BI8ASe87Xj/7Hi3u4+NU82eYFYC/xFsCmDdNzzdKaiFpw9H8P1
MwBlmc5F+Po9/SpIfx7BZwqMckZBNpwrDDOP0OItcJGvKiUWVtMYu4KiwWHXQz+4GSgjF6odWVgK
sAq/UJyDJsamyW4eWHxldHrEvueAitaGPoYtJLWfqyYMUhbcTjKSo0qEXCDNe/FMnxpK2MEbNn5N
IG4t5x9eGODt88OomxVlUlPrFcItCa18us3lQy8fy7W+vpCiZeFpTXg4n5E2LKZLu3xAckxE7IKt
iI7eWivlC/xmZfb7lVNoUcSjDrpG1ODAFTQPNpQllpR01mqgGxmCbvU0xOuQzrw+EYlAmsvRIWHl
hnumSzydISBENmq5FvSBl+NlWvwVk5wTrjtHcBsOuYhi89YHxTKz9AG9BFYo6PI2LWaWFMsnT6pW
X/FmCEAosH4p19VHFFX2Bu8Mzuekrnrq7zXnT1LachuR+SyHd8vXmRX2M1FP8IQnpUfHBjPAzYRW
05L4CCsCUk4Bae6JbWxl6ljtD/ljmi8jydW+4e4hr6HnUKskhBLSV3xXd3nFK/rW8+YkusuAUq+j
LbS33xc/bc/S7FoXOrrgxX2iPcxkG+2eSS3tjJaJBNJzVfRVaL590UlBt13tRvle7Wpup9iNTqIG
NzTfqYtYmeyeIzvoOnni1bGA3aLzSXJLy6MQW31ulrEQQzw0mnfyYfVHq1wt8+9vayFDK8nlPr85
nrOtxwXwvl0rpOd7BmWsmo3y7izzI9ZutvSP3TQoWo+Qjo0u80tzHjAukJ8Eo5fX+uQiCLmiYQMl
PzAV0Dh8n7+0Auobkmbz7S9As9rk3W/Y3pbj4qVCVCNGsc37DlHUrqfej9qW2vaVuxcJuDJTzQU2
CTfgqyfqjZxtYFg5rjOdtuugE3sSe30+kSgN6nuNu9O5/hL6u65VGK57lZbFqsn0rGhcRo3IPzi6
WDndKrT7dMUkr++rGzC+2DgLXmzZzJeFOzsRjBeXZAKdJCojd6sbrJSbNH5XIAfWs3w2kJHFxEWX
HjN82wNhp8ERQ4uh739qykB4WiizFTNGik+HOxbcGbbmIJAFEfDYvgkJxw4hDer218ZjF9XbkvCP
nGIZKY9+lIAMYjBNZhNjF0kD7WPcIUh3Ior1Y9qJsnHI06NFqST1EqMSCn/q+t/5YWhmQX4LceMT
Nae1wOSkoOqudhHNQQKn1NrItCFs4UaZ8Als05oiJpgnRNrCBtAXE2Boi1LQjwNAC58UZ8HZMl/l
DUslyT9AR+os9/2O9TmeWvIXh6QBnMIk8F6O2vsqs9PG6vHuxq/TW7wYIVxLSIn+1F6WWD721CJ7
Suy7C4Dms9ivqDeVokrum2G9Wd7AqL6FRV6PVMH0FNXpn/F8qbo0C6wiKeEQ9D4z4N6O/ZV0k7xP
dWQ6Zs7EvqjFDoaRCFum2V2s0gGepb3Z/RWezpp7O0+Bbl0enqo7jPrwTMNWSJvAAYLP2jdDIvuh
0EKmVc3je0g5+5PAPWUCCr2niNcyV5TDHxSKFkxUXvqc10qogM66r6bx1O5L1R79oOELOabSvz5G
99qb0tkL2EVEdD1wsGpfrvusvAg1aH3HkUsbzz92tn73+ZOvZ3oxP3plqZsJGgMm/mp/ERFr87E+
NBRLjdO5aA8J4Qh4WP3Dg/th2Mwdu5Qfg89v3ijlXwi16/NeYZEZ3cPggY7d59+XPfWx2DZxeNMe
1GiUD2gw7VQwRrIBEjJ/TWbg6bFgdCkWKQZxT5KyeTF5RnUW7m4V3EYuWE2kGmuYAF9fQUjykXqY
Pth9ExZohsEiPKd5uDD/G09FjPOsRptTZy/vXxDpliWDrp96AdMOiCGEBjpdnFv+N/I5fPZ6vyMn
40GjhejvugLyYqR2Ycg7uDi1WlKDAR883c9XGx0fPZK2jr7j6VpR4a+sMWNNFNDQ55jTNRnk6+2B
uDNTpVG2EVqaHsWqJo2+m32iyA7Z4ue7AMRFujDZ5IyeoqH6CkOg1w75rmULXb/ha0rQ6L5z6I37
8jgzE/z0Y1ch/7SwVuU9uyCB+0mLgjFRhQVsPa4PB0+dKFtc5eCdJGEHxB6wyKH1t/0rBjzuXMsc
hViW1OptVCULTmEXj/9q4CD9+5veBJQop37gxV6O91bVmkYOjQhEwwtv+x1hXKTy/uRY2C6VQ+AL
xvtqe9z/daie6M7CStdCH75W7nKmk/9WYUGMPHuDd2xDIs/GsjqZAfaOumP9k/fNRNJarx7xSHWV
ljTkIqU6uzlXgD/P5+uizhiZ5xXuEXCzntpim3p81PZ49rXkauJ01IgbjnqI1EC/b4wGcrbO+/oe
xfsf8rEowFnLXAgal6BLIfJHUYPicnlA8T4lJIPjO7KuN9Ppvq3DUUJa15JsGINb1S90xBA4XBfb
d5945hIavzY5DkU71CwBV1bANRwVYPNSLX9spATv39p2GnjqT70UAhvmoPOvR8vl8h9Z+/0q5Nxc
cOVNzrMsYlrCIv6ocqD/o0/F6+d1sCzrJowNpQsw2KdFpF6W/6rfyu67+jpcRR7j0JMNasxwwUB/
CvMrtBMoxJjiJJ8OVhXZu8u8f5luoJTTwupEls3Dyl6YR7rSCA8P6LWkNjwOhfusvqSetRnGAhaw
ReJTzV6coSRpHoEC/l4YgBW1/EvMOb/0MVja9iWFwXvDhIKy4ZSG5lMOB9EelaGZ9fhjewet0ZUt
wdFIa2VjUyyq1L5Ezx8ZZEWcr6v9CCik20VzKg3/bnOmOso2Zbr8jxDx0uNb3gRpHCxNOCw1jZ36
TkTYIp4qIOg5ConBB6NaeLtfp7srg9rs/O6W0/RRY6Z/K/JntpgW+CsXieslNAGhpUc14zl/SyEg
5fBMVqb0c0RQFhov7vV2QoxjrFBMplJBmfHZbA0QzeKBw0U5wNIB0beM3TX0VW4v8LBoh24QQhsS
LVs2+errxKwgg9AWhuKzhd1JpnM+Rxc6MV5Lk6wDpNE0Eq+6Fuo/Qiya5lGmUQfHtcrcJtCN2O/1
HD4+tN2w3OnPdNfn6NwN8EvjOHtV0ml2M+3C9874so5BWIUgadDc5GYnZ9p2qw0WaUWxUNgZkX94
WxumTNa+B5FhZe1/+t6owuGB1oaYpWnK3gbrNPwbv6jSx5eUCx2uAiQlR+C3Ik7pf8GouIdHfjBB
vH5OEBiuoRpL9Te6SF2M24xOi1nQR73d3USofFXv4H3WPAXpg4nO2w8mHEoFGHWPfysGCfQt4vRK
npcFNTT7WJJKcntyw+B9CacjgMvGmKvOynCy6aUxBd8FjN4vKov9GXe8GL3Qa//dQgDiagQOAWPI
aPXuOpm8laBEBncHeTNXoYkKjtNpeTBozkHn6bd1Iw60I1NtzP9YGFEXXzLqbTY531ja5iphPOfU
XfAoWy0UnaTaEZQBNqCbpRvzdRyy8yg+78JXScLfWBjkTaxvK41enPRFRd5iiFBrNrEXf1R3KNru
FvxqKGZSyTC6fJcxcZ18zh+w/w0wrGXj+fIOlqWvvVPZgQqSmUC949IPIatViU+qHxsAOptuNWWq
XJ0hxtQjbhGyiA0ZhXe1afpF4Ajv5ZvaBHqhz2p8M6y/wRsJtAxdM/tZF75wEj40bKwp+vtg/0SG
rjp0iBo7abIgMJ4Wg9Ylfizxs84Iz203z2Q5nnZF790j9r0BqnN9RSb1hGi1tCp7ofFhVx54kmZu
0ZJTXfLcggspNuQ+WHsJn5aVazeq6ia4oTLSnOiNpMNpo3HEPyFlWkfe2z+vPtGWfsHxxon63YUm
hfJ9jGnD2zMD6XZ51BAhmtrr/t97cqt5rPzcKbU+jUI9gBclxzAdYE/vyZeEasSKiBFiwQeOlwX5
HoVeZedVHcKbT/x8e55ohaHAbB2aU79/DqEC8ROfMNnRl7tH//6c7loEFWTTPALpVg3JTOPzFn07
kfW1ruV8iQ4YlaYPaWAbuXXsRUlGb8E4AL46Kdzh9LxOimypFBjSO4DQrnYknpoOOcl1q7J1vCf1
cEtRNJuh/smoQvLrIoZd9IjelDCXLaqEbSva0uIFHEmwx+YgFBqoKtoJeIx6xEy6LL+jIR+2swYk
JNQH14j9yh13XFdMEy3nD90iqNmiBH6YloFHzmOSlevTArFsMa9EZ1fRjOrn+7kiE+ORzip5QLx6
/XOMFb+pOOZkuOvzWFhIS/uDYol54TFzGKpvm/M0kRsnOkbVx9mAAB6cfCLVLrGdyUhjrgCshxCm
Cf3oH/qqtvz2H4ISA25vQsfTUrFg55lM5FO0WMiGYBhmjZwNopYZNn1yx/BBH8MA7xXYVDyVguiS
3Mvcy2fnlNvc1OwAb91DYvCJXl1YeKdkI9W+jjKw3n3StcstAB4RMbdh0sU+mOOpiRZjEUt+nwnu
VNV6D+Ftou/cbEkZ5mSJc9ZaTzHhexHtU765ZURvhoEbFVQEhORVnqJZ0iDKgLv5MRuArMQhtvZq
OW7gk5Z2RcGBfFf8ruFzCTpTRsoC36JhVXJOrdHEohQpOudhr/z4N4lFjkmXrVB2sOt0atJje1cy
BZg4fSIls4IDFspV9D743PzdaBL1lnyr5WqXmTq7bJNEIEpykq5u2vXSLwSnMLX2RmWZVPhuPlgb
YmiWmJbysqzllsRglbprMtHxGvMyaw9e8xJmtQz9xOTm0Y8FRxzQK+zy0nRVDkvmKRJgw9B+yUvJ
qsVKkR+fXScq5DEkEUbiWW7x+U6hhKoCrnauEuzrzc7XvpCsvTlIJxwlWiyXM7xJ/5u4UaI2/n+S
lL7YFNiLHj1KibvbnVtt8atuFPNDANbRNYUDn9ofcwyTPKrlY/iBsiG8D7HDz2+UPiyptFrON7tA
DYF/Xfu421iy86NStIZnY9ybTPF9w20QGFBtIJGaY7ARyCjbW8RbFXZZdlCYgab/P3eKreALAvbD
+WQwGRlv9tW74Qtqz2TwSCFSyIKnk8zUuXwU3TU7V+AuKDbr01oT5UOcpkSoVoHbQ9AjYMDFYRiw
jUNRRrWbBxfDYkf3DWcHfkZhkE4ZC6B1I6FSdvA9UBtmoccdvqGDAsoXcI1kxsT74UcwznqK4rFQ
6WEW581Fi7qFk9xJfklq7mipFlv/2BnKbG7+mDKewSIPsLmHNXT+daweNgLGaToPgKssAt3zH6tz
pL3G92X7o3uPB8rYXEFTDkcYwAojSnYEDCJTSljIYuMJ8NiPbfRIdzUinbb1cXKoi0DFoCl797g5
QuhhIIog/yevj/SoWYCBItiGwWxIpMHCJWjTCliRAOnZRpsyXQXzm1BoO18JSlNCtq0imQZ4AmCI
9PJjLwr+UK9xNYWMHRYXW8M/lXq139ax9Bdn1ddVi/puaOZaT7YQ6VEA0jANnNoQ6oMOJWKhtBvR
7K39Jwxh+FMf+3AQNipIXHyrcoCI3ED1jPH4ACGSSWojXDRHNn4qVVMwYwDOSTHclcSvyankaYOB
HtpEpM4Q0MOHCOuDTp4Wzi8/5kprOXt4RM0kamrve+P5v/h43EVQrF6UTVH2HIUmjcbQ5qxdquiv
DhFF45stFInwS7FJo5cBTIkXRgazFFBj6MtrUkUR9rxLg/ByvZO4LdNhYnUYJim+ynEKEsPcsYIl
shCE5Q==
`pragma protect end_protected
