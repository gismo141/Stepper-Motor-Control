// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
I//GZe4YalrzLA+54J2WzVN43BeWZJzAfV78RiadjYfua82+94ajtReR+EYc9QfuaLzK3vSfJIUo
TNtAV6x29CGWo8ypqjHZR5g8LtY6nY8IQGbjNfaX01ldjfN3auLKqjLNAl8HYe5nAefeL6Hy1cUs
Ruv/CfOwHOqYCYfeU+yPuoLvScDNAmkIfWJaHX9HHj29tYh3y+TNGYI3kHRMuANOjI7QlazFIBbj
I9mfjO+IdTpZLC8Zc3ARDBpJER0eiq9Umu3w8lIJKJCAL0Gc7EDcM13ZD0qj71IwDqp651cx3+ec
8B5WsIxZIqplTZEOEsCIIfOwxo+AAAUEuY9Gkg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
63x+8XJIWaRTX6YtZjfRtKEGa7ZxP2Fg3VMcIdpbs/4Z138+iCFi6We0Tzpg90CizVIGthU/KR1r
okcvtSBFyTJ5yX+IEgs4ZyxnstIU3OIAA25Haj9YpKRdHgD/gETFhyB/8g6lWN2MnrQcF/kuXvaS
Qd2PXHbYozrjml3TpFWjITWmdPNWxx1eAkAAtufdxxVL1G6IA0dKP4DoggiT7aPCE6yq/NyzKKXX
y90JJexBNzwnu4t399mqc2tJx8Ew4AGbysVx7YajAOE9dlv2XCVbvln5kOZFy94x6I0jRxKKB2cm
ebLOMv2u0YTAOKJAhxiHCl1KEUseujcxH1dJJMEq6QIsxgEqGmFFtZBhIj4ACrs+EVANzffQyOKv
heFs5SO29wOb0zgFAyZpTpWXAXCTWwHqKqZNKI8+oPoslouhnq+LE3ezMcO3Vfl9zrGzpSBXmLSa
PwarRWT0Q91bigdNICr0849MAZYUF7SUiEgLSt7dro0ti+/ro97SSUZBs+oq6q4P2qmBHr8iAejr
AblvcBy5W6Rejemj4wbZiLAB5DlBlnStJ8jTLeqEbs7WAqKY0vkdA0DuIq7+wSC7QcFpS6VRbrvX
V/u/w/L2pvBi7bl4ngmMrqZMzT7gt7clkpmgJCMjI3K2ehJl55VE1/HcMcd38Dge4lUvrjde1csc
T+lYXXdz3VTmQJDklxUTZTs59HtEKnKvcHVyi6oYhySk5avzEGvZydL0U4BN2gWJoG9q7UeykHa+
TRIAmZXVd3mCgUdpxqB0XTzvf2Gr5bNb0I0Xxbcw1kwOdc4fc0C2+ZYUxWcLso1rPOzalKOO1929
rlPQLKCucvWW1uyLIRrjqp7DVJxZF2PnoRAysagBDy8mtE2S8ZSsi/Z0lIJ7IZ4WIIUn64MbqUq9
st+o0w0p0iqIuqzh5OJkJ8Nd+bKFQGcTcWt9jHhkm40pFwtOqX+7u+joIem5ZzfH5gYmVZVlpq0o
/tSODBx+sEfQBUG3ZYna0MJ2NfjvTuo9dFwGm8yRxnDYeaf+qZgL5O0xLr/XxBsmNx47xm9N/NEq
pTO7CB3o2RxvbYS/k1T9z3R0L2YRAgxP7+dwpobO13RUiaxI+z8mVbN7oamQIBO2ZPp4SNQWL6jZ
RKaoBIiWnZRkjsp9OGRpk0dqe4TRaVw27QgowJFz4yAI0OuZ3LmrAPQEZXIKtQAHM9WrhVsAq5Qx
RppnfIpQTP8qdLkzfOCfqKxntLaDjA0vZYAF8GxvvzAYsE9K7UMz7jmvSPqnedB+kXNLzKPUr8jp
w6Z59/WbvP8x1cZMyo/3UZ+4EwAc0jmVkIFhSeBUYb8bIIGhPjOG2b84zHsvzSkibBwuG3Pv0b5F
+2WjprHLbGjLyktHaAdFwAOj3qDh+bIOlys6ru6hlH/5dX3opLG02c7N27KQs6A0VUss2X9Kk3oU
NlFUqnm+kw+TN8DkMA7c38EM14vZ3MW64iBWk18JoMUipik9uK+GfBNtANGSJAVtCNoIDiP0lLnP
VeWK71MxExdniYBX0sxm3JpDlegp+QDcEqlhOtyHwar8dZXonWg171HSRe2lGYXCpQgFTaFKDxNB
ZDkbZpAE4BSO+kLkO0WiPN42wg1IKQ9BoVwl7j5qdv5RdyHyVRCAgHDbyImLgTRHSfHXvrLrhJ3F
/odJIUJ6WSss7to6WrK1HFlvLvWUv+JR/c7IraSthVTQYlozLryZpDOdr0tlsDRTpA6fsFOkA9kB
fACcnPpVvIZliSJ2TfqdYRTHZoPgdOa1HDonKtSDRHixfWj69Ia/nTU8c3aYzE/Jb2Kfe2yo/e3W
yj+e1kqoM1cyh5o4/fbHoUdB0Iuy2VSDfCjjV3WVy2xe/e3yi8foP4YkWS4A0iqoCaRgORIMvbHB
wyVJE30sqpo4qnHrroYjf0U3R+iPd/9xUquqEGcjG2C30Z0QXDuQ4dN6Q1n47NmLkaEb7XuByCky
AAJUU3j+qE1YAWo5g+KVozNsZffMuXlC9C9L6X8e49i/LMZTh+3ulnXkSV+n3gneqU1BV4whZgx+
6QTsD13Dnuk+1npJPQhHFqls/EscKU8t1JaCw2aR8rhu1IxTmK671DIQqFF5d/1wnBMjWT680lP+
5YBP/djIOVXkrEinWs3qgDi5q8DI7F59UHQyLTD4pqcQxjKDE9xjre81kGwKCvw1Yoo5wb0OZHVQ
P1oTgxkGKoBkg9kA/SVNQMB0LgVLqMync7BiEcrLtMd/MqLGrz6cHZjvbdvImisVh+GO8WUEVaq/
K7wiEHOV0YUVOJDQt1KtYMBeMZ8nYgRdPUThzjm2cM/9jhUZAFwQa2K2V6s/5akScbUlKB13+fP3
fo+9wAAnxs1ZXX82IKsOl9GFHDASIjxB6pTPXu4NE8eD4rMOLvoceEfSvCTWvATCF/0s8tIpHlIH
+/VRcR30f4QzRi7YlXdHhpDm4tguFyCWYDzIVXRPAFR+hRjGyLvsgxbQu5xAeesUUvqqmf1YmZAG
+UXS35EatRvPAximoGBoGHEulPlwsrRMYEPh/2KMEY5AGD32oio9k14bgxX/9sYHp68ObrICHqai
VKHgO9lHGKf781JFGEFKVAd6pvwDAuBVWqyiypis+bwUmuzyljulGg25LPLJ4Dyl+b+RpKo7sMde
sT7jqJAGTDTIXV5J1A82H1J1l79PWoZzJ/Zlr4z8BQV2qVTD9mtF9HJ8ZKt5FyG1Ehn3wnvd3CTx
M0yOzF2ut6Cf1lIdDtlHUkyVARaz4n5WkNjHv3jMS1MNSGiRHRX4YdUtklcdLoWI2cty+l48DMSO
+Zpg9uoNOspplS8XLPdGvqTFp4XzNrBy3qYzOuBdcRAdOec1NDmt2Am8NCJIkCQJcL0/84a4pT5+
ZKYn+1KZjDlKSNxMG61jUu788V/tgngRCdBkih7KmeeaNFB87EoFyN6Rs6uBr92Y/pBaiIUeOorJ
pfBmpHAlf1zzPkL8D6aI28l4cBJIoXIMhPXDGkWXmECbViD8rsUbJWriyg/uGKa2JSSllcIJKWKV
wrcKmOcUbKHJzmKu+KzDr7giv6nM5tf9YmvXq+XGqv0Rc3suEGK2X0mjdj6kahH5g4ZxQeuxPyy9
26sJ2BnmM9hJFt+cS35OigFnCE9+lPHM7FsSmtctVlZ19Kua7V2ogPj9gFDvoow+c5G0PaVsYYyg
JJpVuS9fSVVaT+3/2jvFgJRyM19djAmfjEgPZtALMJPmnjcjzdZf4rz2vSqzgWxByHZz6lktSDac
4EmdWIlPMmzEQCA3IzvSY1Kr5K8qCfjyQGM6TZwe6XnjDj1pYexJevR73PKIQ6VXRtYDCbiz1QNn
S5yjIKaCj+rCBh51Z6GaI2wC7Vl16DiegYl/6XcDGooDFVm1T61b9sPK943xPavI6okqrO/h3d4g
fuDWXmSC3oGqCmBGl/ZhVuDGgoFsDB4FCkexTXU5qXhJoAbOeDTN0Y1qwjrYo624fqT5aWxw/1ZV
h9YjA7t/de4UcuByx28y5xZB38k74dZZk+So0632LjGVfNUkAgfW1eTUvKN/DkG3zye4xwij+cO7
XlukOjjhLVghN5LcEPwfVtC6RbbkPJcL+zNtrIT/DCvUQWrSgjqK9ovUa8Pg6oAMuJv7Nj95UDue
g1F5wtO8ty6Agg31xRuTmh2Vp6IIuXZRWrT3h+WdNvB6KxdhjfSAjTupx355eT5/1/muAH93mhez
wx76VeV6pTJYFpAPrp18FhDiOPbW1TRvhhrM3xljpZMKOoBYfF0TcapiszoIKT8sNLgOtv6oE3oH
cCIAgTGNKOH+DjdxTx7mViFS9WYhLi9T4e5VOl+C+d3u8OEY81SGe9Rx7jSLjnmk6WmBufomC2pF
ZDjXzepxHoDCtrv3Vn6ng/qbFAaEG9pMCT2ObdIcK9xIOSWJUb/E3Q/v4dHELQtVGs1CDOZcwtLN
WFDynmBGURv0P3c3R3D7RRXxQC67JqgoVV7/d/ZiuOQOJKJ8Y3xHdrCPG3f/FSChnBRdeQRnYzMP
u4iar/QRQYDTJKqgxWc2wHr8yC0anzL3r+jaPoIJHBUJIPukVP3ekqZTg5H9p1+vQ9dOM32F+veu
iaBvPGg3aiPfyP8d//C3ny/KyOP+cX2XXd7+HpLdmKfC/8D+AWJpvfJhWFwtcnVKocl7AuguHjCu
exes/D9rJwkYCayZ32LtI5SNcgH/BWpVlpsG26eAqyKsm99hME8uvLiEZLBqUb/YJ6o1X1tJ4NnG
Z12sPOkcrmqBuDTNTU7fLo0F/kp2adMHIeBIwVQe4g1phIQrbgJYvAiXrpUr+qwO4Wq9CNhsSF2l
i2RNwCASXntfivXmKW6f1F8Dxc4neN8P/LK8bdzOYc2mSMO3Yx8Y2P9MLZrxCmVMZppA2NxBVyJk
juuqKLkPTmSrMShVvQX9nOrO8jjLb7eir7buMdODg9Jem9z92uhe83Ko8uyyUSBnUO+ITvL3974B
DkqOxYZ9eEeKGd+TyGk10No167RUcKY1DZ9sL79eYHsCcnT8/rYRrdTJwGbZchKVpYvfmyHPTmS5
2IfMEMIkpyvLI5ZHxXb24/FEBWcGCLV3KVXXwBPJx45Lr3KuGl9Q7BRqfVpxEK43UCqsUWaamgsx
8JcAxx0XiDlAPzQbT2F1C6LytnG1fwjP1H2WCOiFc+2GjMII7u114q2xU/K9TlAOKAcgDFAgZ/UG
jDR6YDbzGtgnNYBJnSr5D6AZpOfc/xWLE/gWpmZk6hNJ/OKHZDBDOad5snSGJrZWOec2wBpHguFO
ACFwUB5aWpLw1U4Cw/b91Yj/QRPhhbjvWbiluudJtYJeP0hfvmNy8dywlvQ2wEHdz2mI//kpydmz
6xINYQRfsE6NfslpUYyr8hyKHYzlBYv4bO8U4dwvjB1Qjz8qOBsHYh7skb/TvcLTzZ+kHmnGwILn
oxRXPYvRYyayUWRjhAC56VfO6PthsdDLJVlRFgFqHfRQzgW0oTCShDFDjFB+m9J5QHo+a/sHy0hi
w+O0DKKYec+99hq2NJHWLdb7Lxkdr3/tKLNIB27DCddkfSm6JCpgT/zQxHMTiv2lmViNWy7Iri62
rdFivsTZqU0IuexKnzFanek4z/8/v7ciPUiOS5Zv1kpPn8UrRGqmJOjqsB3HrxwJWAYXXRSLyCwE
yOv1Ba5dieUZ0bDBSOB6ArWqFjs/5Yz3TJyfkyGqVESuqlqk3+/OwhzTF0j+IlAt2aPlhl59cfJP
tF023xr/C76YYqp/JI2S3jokYhkgOqXvExcvY7OAvhsWe+AWK3tI8XGREKntc/PtIoOaB1jPSZiW
Mlx3J1d5cXzW4htHwz3aVrIvNot7w4g8KpANzcHXwWaqdG7YIMJBh553sEOvYVrba6ernRmuskFI
RU57gZXeVNZhGckat8KsM8rEo1deU/lvHRTcM/VKyteXsbyu04qL7C6WFzk+2WFbxVCGW5qcPoNG
rHsFTGB2/H6QPM6wRvofPcJ6tKHSD1KmnsUgf6briCxlD8m+AYitk2CJllkEKZOd+i9qWxvbuQoT
QPudQgZs+g2QPGkQEOs4202Hfi1ADkThImhjZu+RhDrlMJpv5mi50Q4iprRaAvgtYAUIGK+zFY0e
F8OF+OAnBTvvq9OSXtz0xpJZ9FETPKbrX4YroMEcChj6jQSm+W8N4Q7y3aIzkhIrayAhPbAG+R70
Tgfr3ma1OSafiB0HpAlLxUzZJDlx+cI45PY2A/423zKpRWGu9XieYN4Kz+nGcK3+bAedWHIZAvo3
NeqbfY2/4K+96wtzzF/vEzFSBQZhJUjECnHAcQ1HiV6/LOsk4QLhNNEV6pMeL7JEwnfGE7AQgwOL
0La9/9pWp/0VsJsDM3qKLqviNXvpX1mydWO2XNRb2GVrJCSMVh9+leLGwWDs3rXnAHnKZN8YbltT
wt7iuAExrRXpsBF4BXXgDzfRW7U0CEBD657s0BIT+9yfXscamdEsy+rhbYrgO8I6C/OfxVoEgBuo
cDo8y2AxvQtqT2eONTFgn3fFElfoKoh4OLzr3Ic4qG1dZHxAv1fHyZRRa+SGrlBA2qERCCGqvgfa
TV1bv3abIus6alva6yUIWTBTUdh7nsp9cRyu6IjZ5hv7gxm80KjNcLYrMKOWRV3ofQ9zxu3qt64b
xXzpYtBEd6ts10iNcmKGfJ497oqsREwjNp4eJIUmBAFzHFRxMmsBU7O1jqhCHxkbbltMQtqwwdQI
b5RCKDV/smHB1j91kHusv34lGzba4lrhb6XKvvszPe5LQjVDBCs7teG5gDAeu9YX+4qzVEBbvW0B
KS+xILYNTpl8KQBTbdI8i08o2LkUo8qBZSRwTTCxrefsXokex8ehd0dtVp0uM8nKojy3AHynjWEB
weCMtgLroH5GFiFjBNZZoUPc2KR8fLG70bj9sWpOlTM1v/DXNz2V5ksGAISjhwRrh6cvh3tOP33U
UY8z5VP7Bo7q1GJEC1ZYB1ENpNJbHBOE+qY/JQzfj+iymueYc5kqpC7gKKveRS37U8bCkkw3ntky
D11L99BEUkml+7aMl/I4Qv/10YeRALgUL6Bl0vX8gBrjJ1taELCb5JrPSX/cMhedIGG4DC69RRju
FC3fF1yTsOMyuh1NZJRwHTIg9GUWo11mkzAMgZPopk/90ivc5HW3mm63tA9o50XCCK3USmdnyh9c
TdnIxR00PAb9N52z26HWuhkJkVzKhBsnWMkJEvj519iBRU7NUk/te+HxeHP6j8JZy7Zoi5U3D1tN
nYazHNtBiLiJCpLDsdRVTR14tcL99yQJE/AqiOyGdabG0sCfv6T0IB4pXobUMi/q+x0kAjL98Wyk
E8KL8puDRG0Etr5jull3Im7w0W8i/HkBJrvKcZQdFz/UON64Sqaxj4Qw/hIgHgGBrwcKAQL2Wnrh
YD6GOkf6mAc7GGhvEc8V6i8/CBIsEcRxfYmmjWVRF3UugDibpJSdkT368e74CuLQoLF+5HAiXSB9
xNUHBoO5HWV+URuuwtZaiVQBPL5i31vuW78OBP6zOzLrotOlz5yeHLPVhdWxrgBmQjQCj8pArq2E
yBacT/4YfRr0E6VBATwMmT3qb+5K+PPgKOfUss1L1tLW5UYVS4yLUoLvr6OaDYhhKI9Q7q4tvn42
5mUf+tmatb/PpeZUCkKAE13XP00nlaFodo+qnGKCgWUglZ7dbc+bigZ4FJJtaoNAtIIbgrYhuA0J
VWjI1MOuuH0Iq8UXCQYbmvKbnAI9qqTjUZx1hqpbStiq/c7a97ZGOUFPwxOjP6y6wzKzIBzdEr3a
esKjanKtp/fLbponYfWav5vZ8nWm1VPPZxLuN+wt+dChpC8kRgKKBxgvcFyGlLhRoWhTZXTRdl2L
ji7SRaSvdD04ETYC4MQaUsiZhtY+d7EzjBv7KfyvMX42vMQNSyldNoT74WfgkwhT6AC4NPc49oDP
MnbIs/T9OsIc0omugVkjKi7H7KjGRrWjRZfVxESVYFfCYqBGjkGT3XUWxP5esLelJpVXvd8QviEl
puPYCgetLgyzEGO1S4c4uNmeqjr+Hbpe6FFJeqbRlIbjjDkStm9SsSI2EkhTMfQbi6380uRdFdr3
PuBC0FDjo58wozjyP28KbKw1fE7QQTXn19uSdQ9XqnwK3eqtDUk2shCaLEL88TPiR+wZKWCEVgUJ
TDubm7nLFljIX3QWcFQm1PSDDy3xC0f3IrFLuLRwQPpchnyl3SdF5m84bIm7NgSzKjEqjixp54hl
lPVgGMQUOEwwHGR6vVpaom6yTcSK8ZoY90Tz+22anNnCje7Fiz79g1cWq966m07XJ06JE+Y+Wypp
NcdFRmW/n95KVD9WyQ3rRINnNQoWb6YYs+RrhCo7XpIowH1cYpmLr+nJAsp5Ie3Yoe5nksNv87fs
MWdovtqyTJNgxFCUkBDDiq46okDQskjVeN0OTdE5jcfgW6CO1qSkyUFES+a5korMqhwD3a5ZSPbG
PtoofpnIjxgozj5vUuQhfkHsOL7WANSkVB9H/NgGsWfQANe2s46cs9kk3pFZKlgXlU1RIn8LVRZu
tDbiKgCgy3Uqn2M8jH3CH7IAMhktRg62FJi8Pci37T3HKiY9kVa/kJMITGvB9W4zU0ewnIvrhloa
0KdU0mUVLlsidVVgCGklQKBvowZBSVb5rAyDANV3mmVrkv/WJ6qYTxSB17K4KVyCLC/4+oUG+Ayd
eI/+MFHTpznZpjClFW+1KXkWsezLjZyyG+7013uMXJCrkgQnbOdOmI3qS6muQ1vanaOAKFGJWkzr
T7tN4Au2EY0xkEBVZg7um2uFooyxDZfFJyhYeiNuqD1cUco4DQCzvC6DSdGoEarqS9NEf2krDW00
1BU++B/7uFqAgQXNkH73flS1cBg/msZHI7MeVgbJN84nNuBZ1Do6qvrcGiu0oqzwA1EuXwUVndIN
Oodpmbev5GfF1AzwN7gPCgoohYQbew5MkxuBdNW5Hjq2miTf/lQinFB6gVu0w08GOGIWHo7YwXjy
cguDDzPXj28Q0EDW7KsFSMzIgVd0lKJNpt6Q052m+pD5rydMYdrnTkQLveBUSl5RIj1d9837IwPK
3Z2OyXt5EQjAXQYRncAI3W5e2n99TTCD4yN5dsYLflcE487WvaZ2P18KuU/FiyG7wM3TB/Lnvwt5
zxUITeQ79nl+x2hbzPoajg68zM8tvy9+AGpN0cAxw/KjHiN9WlLlUqwwWyto3aJRk8I8OV4JnjH9
1LikEvEU9GkXAWL0+rZu0ebnbKkB4pK9mtV83O3seujvPeG+JwGGd3ew4t9btKNXVJz+2NWN5W/K
RGQFFTiU/Ggds5rOrJwKXF3tiOHpxdP2yJnbZzp+wkUSGwOQkX9LDNw+Smm+pxF5SgzUb/4jSo3M
nLcTnC/9HPthV7g7yXPZayyfRzbXq9VXNcNVWBmTkbdRZrEFsHd49H5B/TsSzWDHY/SLyy8GiJzn
G2RsawJiC4SIJhZkOrN4OEfyk4i+9GAHwzB9UoxKgaANVm60Mln3smy4z3HO5sG99EbEkqkSrM4y
LLLIuVt/onS6NAq25icxRKx9IVX2RfQ8yFgBZMBXh/Ae310SvokJ1a5av90FRwjhb7Uf3OMhdEzT
SDU3y4cXtu3xzFALfZyIVmbS13E6nuaiEP0OXdTwWMvA4JtjOdAyHo74Tse4STOn6uN8zKTlwVlj
SQiVv5GzM+Ih3ST3wlXQ3FYV7HQeuPVGzq8E/MjtVXzGTr0KqQXQXEiEvQzv0UkvOkzisOMsCPaY
MWa69ZVTHs8clSwaMTlEbImoTdKw5EF4kUReEAVSbmM0S99N+SxHegTHTSpqFAiu7GR80sESAOlC
FbgjCzxfyjMabpRxQRBUGxXNiCYq9OvABMaGGzQpOBgLGcK17R5pd6tUplGdv4yziyU7yDDSSmj8
zi22G7EwINw/n3PAFksHZ1e1esxCmRiwohUEHGzEK7D2HNioZxXoTAPPHStYiXLMyBLJ5UkIC1/4
TP1sfxuBD+AXRskP4eahGHHL/sptc6sQ/OCQXdAFQ2/xqr0efTArerZ7tGkgC7/jO4IqNN0TpCE9
CQGHck++liDmmfC6ZEudpD3DCEyPBbewZN1cRG2s29/CKBBGYEhzQFQv3Abolxn6cNGttPy7rAEs
3XdsTWN81jMy9tJel76uDWnbL/oBUA0EwevC/0GoVQk1kJPbqvXmZvM8sFRK17yiEnSuWpi47bFR
9Iw3pfRRaqeqE26Zq4XCZm2XH3UqxK1kQqb2ZoWJ455ZQhTUa3BQm8L/fq479TOWPhCSMxZ7kZZO
GATtpYRocdEXObL3mWeQjKq+tC2RUeokxjYeS1Xv37HZT3Ozx+xtVlXSTGCkBbXehvJmquVE1/db
pQltflRz4U4yEHCRC5aJndbse7TN9dh9+wRxcGRdCmbDaOUt77rhkr/fe26qbp4Iig0XR1x+rr8E
aZUooOEU14Lm3ccMXfuIwOR/sgiYw74kwH851BnWWAIi6p7of59YJcKLnXkzwSLdsIDZnrLKxsjb
qvA67TJw+fV3FugPuLoxkQxOuOvwup3pEYHe9xNaz6pMjiczJVbj9WXmX149XjqNub4xbDvSgra7
6wSjFMOcfxu907XDbc5kF2Eib4cev9sfS6XXQlo2vE35KFb1u3tD30meq4JJ9kj4DOns45gtk1gP
l296PYCK6VoGV2UU06eIOqZhUKCyc52lo0+7iuTkZPY8JcAIvGk4cAX8pPOMzJMjT+zq8HhXMpDb
01Q6mm14pQ9DVhbILLR+UA9UOGopl1ZvpQRU60D1Ai9ecMNqVMusjMUh1+nb14B/1QG7fdQEo7fj
/tqJDfqdPMNjQuSHOB4WZ/v0lINZwdreuISf5XwFYCLGrS8/OvSYeH93df7dwZEPuAqZ23364J2V
aXBXjYeVGckDiDShDZnQ/yKyIszaHknN5EFjcWILY+5uQBzZHq8YoU2UEpQRdYK7IepxXkKu+ksG
qIyQ4UVkP0rUixC1nSs/tn+Ta6uktEaz3RLnMUjBbG4z2oFgk3V6szazeV8nTDNHJduBV0KhxvHO
K2BnpibXFd5fGrrL63vy07UW579kEpU+AuYIZjMleSMm2U0BuDuSQfriCmFMC3b4x6ek2h8IJsSB
z9Z6+is3VlO8kz0E0Gmxgnp2y+AoSji6CpUEG7L+Hn0sg8kanFG3yor2U0ALSwn0U2XOxEkHJ5kz
NAdUTm1XpWpn0jFtNmrFtmHkt4pJTvaveJxrdjW6Q4yvofDS2VCfec7BTdjfZh75u5cu4ay3Zv1C
8OvvNNbD5stdgAwsEl5U8oxWO6ltx8VMQPxSWQ53l9szd3mNRt7natH1f+LYdowPsihCSZWAMKLg
bVhrsnjLrmUIroq/i6Qc1Okz+MNJ56rqf4/A7wK83pyYnvbxonHyjwQ7Ap76GZkqPzufCVD5dloo
zpS7SVX2hAqVD62Cf2olNVt1PgUpJ/G2uhphx5Ro8goQnKLYtGQOtmTm0gB1JgiSU4UoN//5BcTh
gkwVCu/bFdPeNVZcBV0e9nitlX31JZbPBEWA9r0Jlj7tMOGF/rLp86Qz6KZahs6QMWSay6ldrSqj
lqil1Jo5dQ2i7gc0pd9ZrSpmHjeFf8LuCfT3dPKZ7oMfY23HlJ/QGN/SMA9HiwXbPPXEbVjgOAkW
aoF/pr+dgvrui4GAhiPTAyLNtlfUIpOsPpMipEWAu7fuRvBKDpP13cdimgpOXk6sbB5pcEImE+Cu
sPpcW4bP3JUVMLbcNwCLu6DY/5LYykuMwr+l43TZeNCmRWLP+MPQQ7RFCVrrzlwTj3eVdQx2qiya
7mvbVJ+IkfQrBXePJBFrK7rLb9NRzEsDtrr/BAAN+oSqL7HwYE+40Ct0HmBbZKcQquzT/8oPOHPn
cJt1N1JtyHzzKE73fB43yS+aXuuqm6sM6QqEru64BvNq9xfwXI1DeLPImwx3v30RwYwtg6YPiYWF
oJvvAKYnNyn4Maj0pXMFDtI8/7fl8ZTR1TYb5+cDdgOeL6G7H5rX90SVkn2xNJyxWNTYwy9HNc/r
iyyNbiXiUP2uC+aj9iqEL5rtL7JLBmHC7UU5yKxzXRQKfZz+oq7xXjyp8rIpEJp0EbKidU8FI+VH
3ACEuStFACI7w94YkRY4lFEsLivOXnbf36pwVzkvst6zYsciQxBcQZPS3pAiNf2HrePKF+7bzWEC
Zbkf3/6COHGtFTdxlEH/XKTI2Fx6+jr6XyCQMRrcax7IOUwkcmzU1PNQ8S80s4G467FnHIz4Qu55
6p4A1f5M8EL44eLHXx5ASPvTmlo083YovKxvawBw9MRDh87juq0u+bLtg+DYiyPjPv1HcSOfH8Ia
9KprnU07aUngGLEJSt1I6xzlSHb8HDgzZnM4+YU6ALtpMmPA0emNipo+uJEsXnaxl372mmlYJa/c
FbnN4uQnh6m1BRGIIBD1U+/2eEpfJ1dmwLGeaw8vOqwyF4K0HWLzK3MRNvv7ri/q+x+JGtNHYLhn
foLU830GONbZgdOOutI4k4YeoU4XzWQhiHL5VWELX0rl6U5gQ9f94f0G9GOcP0DFpaiVb2ZTEmYU
cG6Re5vLfqnjuAOKmPnMoe8KW+cgJsTCPJKDInGCpHJ+2XEn4/F27qqdJZGx9cJSN7m846CrZnJ/
J63Qooic5FrytlvHUkKGlF6kt3+imaArSBxbePHCmg5jocHjBo10XumqSu62O6FZWotQd3ywHX8c
YC11eHTk9z6qnZN/aFWON0l4K44WHHFU/nx1p6Qq4R7iuyCsTQeAaIJ6yQH2aTgLsq/TE4WBB+1r
IeNxr2bf2kiIBUOuceB4ZLSlFbi3iYWY/aceoxhIPNIfNYvn1MUNCDJnppY+CxkvvHuRYsacfepN
rCmR5oXlCItM3hz3ApIjk+KMZdiJWqMF+pfzjvs5C1zmTqVFvKbfoCnPPLikpFojVS7CZOSRCcKT
sDanO94ScIRyWelmlbBRhwWuQClWGTkKaSpXVrteiiajCVstR8cLvNtkzGyTIw9bfj62G7YKoDUd
YYXG85GCOo0/y+t0JpKq/asxV9gzIu37SAYI5TwWYQa8VCxtp9J8MyfSdeCOpvqlG5PCKfqldtYS
Gh+J5RYiY6jJwbVinq9+MD2PfwOavdmO2SJdF4krBbrk3JJbiKoX5aJZmhF9JrotsxrcjSVVdt/L
xjLZ4pwvpm8BT0C3Fg93l9hTD2n4+2O5gOCs7ignM+ol8zzhmW8rEZo04wNbn143zkUaAOn3Lw3r
iTgyCKFGzZdhXZU3SD3l/gdZMcFFb2ss7ABlAhY8PUsewcY+FqttoNtOo4MzrF69fpdLQzZVlT91
d5n5cfpZeiv4LKPYgME5gdQEiPPYH7g2m0IjplqNEd/DHsuuvAGfdrk/7mc07xeJD25vGpmt5Cbn
X0FT1s8E86IgrFIidyCunHXRzLFer5P1s4TzcNfheAKWVKVU9vpTMJc2n9svApX72KDYk5WAYJ3t
3BdY6W9aaVrsiqkBU+Zy94ZQk7WLiK0aKfTja2rmZH/a0UyVEBVe7rH0PhRUA4NFroJTn/9PWs0p
8nhFUI6WYds7a/+dBawzTs4/2tVodRUMloXWhnI/khyd0RQBTQzt/rNkaPVtFKE+6gR3B6v7Xu5E
AOz5mHUYwS2l/vTaL51lIi5R0I2h69bEWtgxGlllJAG8GBS8XteuDHrLoW4LMQFrJusdNvOsqM+x
1zRFqXSoY243GVb8jeSVndPMOCDYJGTMpAaAMNhbSDpJRRQXFGJjFlrGn46z5eKfuaDwwa1yML2i
9+HgT59Nza2VYOgVGsAvyFRbCxD/+iGfkj9itgv8j41EwuFSxp+sdEOtsiX+52Fvi0EBr1Nu8EvC
jlgn/tP2KegRjKb9UkZgb0A4HMrbM02BX13qSCsofFOCpmcnaops0v01FcCnCSR5toblfsREkfhe
sEYYdhCp84fE+AEg0c/fQZd58ljRmjq0VwTVq9AxeJNXZoefQZvQHlGfeU8O/1x1V0MJ3nT9a6My
srqKp+gqnv5H9nJ31A1n8/1CFI6XNUPotH6SpIo1bKAB+nKoTPkAVCf8khRDYq93+rqo9+77mqKe
ozbi851w2Z+NOXRI4EIGGtUk/PbH1lDaUEBLI/d/XbTzZN+qZ6obLJAI3+8qsp1clbN4DFDCOPIj
XoooVQZpdMLymPv1sQF4JtIE+SJPP8aywVgBxAHqeNndh17EfdyQNF1j27PhghcftO1atm7gnGWX
OMkON1SInZ9i8+t/XRGEc0lkuUPrcEyTH+80WaaBHDJOPHNLeqj4c9oODLuzPUPteG8WYKqCxI6y
MXgzEwhtDN/WhCw9c7TZ1DKV9GsspXunDbfqE1iqMMAWca6QmVVdwmJlXuSKN8E7Mnqz86AJGKuN
/U/IQW+4tRbdaL4QIZCnT0jVKxrKUBMxfN/S1Vqmjpz1mrIn0DR3EXmsGUf9NN80ECgMtd+PzqPr
3D5Qb7I7IXGLFr/vN/5W4T80oXFJUiFesOS+CEpCPduhYJuL4uT+LqPhUZ+1qnusLXNhG8Eg7wI4
fHIoZAH15smdvUFfxKX74UNcmQ3Fg2jRQXVVk2KdyFWjrhN7/FoT6ZiKyWltH3y/QAUukyqGBA3b
H1utXTO+IsNxtKBMaqLOKSJblERVd7iCY8Ixg8eyHzcqZ7DbwMsnOj9kZs6eLsEcm1o/n1HUfafE
wMrc6eBPgNB0hlaYcLgpHNjUhzpexQBGfS04mdxHCUr1yYfJMuv+2X+r8chxI2/S0zc7HY7G/GOk
WAT6mZQieQhf2toVQpK89/ew9Yc0dVcI2su+NSx78ImRlJV+nMkjms6rdV9VcEsQj/aZcK72eBYr
jrsWQ9n+fTECsQ7YFKNDAaOVFZatBFkPFJWPg9FKkcDgtDevVfDFJ0S5kAEYynl0ACi9qvIZ9Ewh
YpB741Spp0hq9b0fUBEzN3HLFaNrNaTuOVelCs+AkTvvSMY2iwtToQqiZu04xclBDvcp+MpybFdb
frSa588j1NsGwJBI5LXEJ8Zreb3YGwB2wtiEwH/8OoBtIQwevkJUmhIMC1z4Y2vd/sBExdVozQEc
qCND3zMyh4Wu5vBhXw+c1B28QsRMNhXxs79vGsaRSEwEsXlUdFz1fU4u8XaIjNMJE1+O1edkxQhB
AVTQws7CFgnLLpsPWhBSpN2/ATYtHgzOiIJ+U2YhdzJJy7IhyWhR0KnVJbkvA9dlgTLAgyJgwtBP
vT1XnFPYKCdC56ksLV9kDO3UUZ7bTZs1kVW0XFm9PN3dDvFOvzMzSfa6pnVNxa9U61ZHYtczrwO6
GHKmTE/mm8/J+yU6i60RsbGwnRX6tbHythfT1/eQgMcGMwvAsOZ/53p9F3NBKiuiGhM7ksHmZzka
uCVjns3CZMOVjx2cZENG8IDX+7tdcSX5+5k20/7ecE1bbS66Y0kILfVLmS6EsKGrVtdpB/RTpx8Z
aDCA0P71xJ34huBP5lVHl0Ytj1h8fyVSCmE03dAXv+gmhxAFMcEg6x1kja249GWbKQTt0bVQ9KUh
zx4LDCINBb2tr0eYBH31Ac/Pvf17KgUSt42j0K0GCecp6d0oEWjljlut8HZ3xxQKRJl4qwmLxSVr
/RJlY/GJ8vNHKAbXKPQIX4us3wIWiB0nDvU5EGx7knxURU/OZiRpLBotf9TYMMODYAWA8n1gT7z4
+Iz6VOr66bwbaanlh6jddumwSFM01crbTbGBNKvyDLlOmBXtCrIp93tLMsowPKLxWsX8A551LHKZ
UQjc34E6QB2AOysCKvVOqONFatmLYZ93uDxk2y51+S2uSb3+A5cORj9OO9g4eCWWLlZFTceRLGHs
YuQSmKAzEinQ430EfBHa/AyGiHFX6lUZMlW0DWbEWYJOVcz3WvAFFy63AvfPVMUf9tuBuNFQRi1E
Ngzj+qj8+8eyYVb/0xR6ZZoOsbGUWgBskZE3ZJ2fb29zAZyIaF4jU48tqbAFPHYPJQaqz9Kchs9L
NPzNmBxP2tszk6zQ/BxnIJ6acrVPxmw+XF0H3G3WfTcgyvJaC90+tENQhPIck9Bal4Io/ZvW3i20
TLzTIz9hQKB70HiotnK4B6rSa7sPaBy9aHZ+/ZPEyPpTUYVOmC5v721KsoV6hUWDner9KrrJoCbM
xOL+e58MRKEtug2BqAOLRfQCq3R8wb3nzBmZC9FONMGmBQN3h7aXpX8CrFPP/sBft6c6LGV5zzTU
HlD3oCgs1oudonx9ez+hZHjBQMG1FGXnLB+hdkfftmzNMv/uKaUj/StH26b+syrAw3vLeusjD5jM
1Oqtqk9IqfX6s8p7K2114IQvHxhmeWsCxVC39uQPidcn1mPz0TQ/tMRRe7NMLrt+ie9F1Oh7wMFj
JWQjKrXjNtAmrTNGqTdm8HW/faWaDGUyjaFN+TMBDF3Mg93PrPF31dOhTn/49ZOCQ8OXo5dmXQbo
qKJzMiyLzCV1H5swmLgcgSvCXLKGcduJHjYl+CS5bZewUM+vygbBkiZsOtZFu/LosqgmK8hxrVAP
D7OeNsmAAfjkKMGBj9LhBQk6+YvjiPNVuj3owHQQkQwO/zR+9muLiGSIeoHk9qPHeMMxn6iS9K+n
RD4N0RW6WqBCSSZw8YmPhPbPOT5onPlPy8/pgbJ+vwahRxAlpPiI6kdGJAM6WbKsDLbDXKtMTRZg
bOyQD1iX6aDgGHkoB7ceZt9Y7P9GoQU0Uvr/nuijYAX8A+qnt/99Qqs+dvsszWWAYRukmu+hjl/p
tC/ZlAlr0H01VKhZJLbZlRRHBdozRNkT7qTwz8J1+TaoZtfm1R5zRfflbIKynBtRp7Fj0ho4R05E
UJWECBOy9yWXckv0OLTWxix23KKTqdOJkdjTF8O0Lutqfz/B7R4IlvTIEcioPkDx2/y7sMCW+FdE
4wlfL6mlYMlyY+xK5UAUkY4oZXTBw8j/Tv/fNfs3XlOV+G7Bc0yadAxWPFxdL+CFK871YDegFopu
9SmqgLFe6mG49tiKDEnWhbebqzx/HuYTlSxJ1+IBYGJj8QNHJg85XH6QFolNty9xDPoabUUZIwWh
nMa5/WwOTJOLRCzat0gfoYOHGqIL5UoZQ3lNIumM4zhl2crOqCnLsG2YuW1UwPespKEGTYSxRSmc
jsC0yc86pwozgRPA6uZ+198uVN9yOkASX5K4Upg5lxOOiVagVmQEbI1C55JsLhmHQMxmWnNybfz2
OgH9/3hIm3BsNLETWv0MfpAAS9PJWesK6BwchsZ4PDYdYn3SrE5ABY8om+8/YoI3GV3PCCYPnu0I
wmH0WgcdT6ZkitEcw+77keuV9o47d164TTANvAKVAZ+rtLtE+cKxcyTzX0xivJBb/Yc8weK6r8fI
9qVwlcqDKpiM+c7eozO12rSVVYAXOrxhOQ2oTMMWQRscbSNnJcAlaksTvTiMbOmX3RN2fMpjrC0j
Y8COD+qZkge1hPF3SkVnqKCnBEkMk1Gsfsm1HwY3nPvONHBQrJsdmEvzs0PxQt5++nmj/Twtp/yv
jfGYEwu/fO+93fDbAi6cGfz1e3PvVD8MC6JoIl3FdDcqY/CdZLMtU3rrE2aoloS9vB78KTG9WTYB
B0kYvJwBWNoqlTegsqApKzRAyqzlOCM8edo7YMYmruZR1VHXpKJchkl4fjAuv3Nz8NtYHjr8/5nm
PZfaHXCZxpMOJxbOvKaAhh/fptvlPCayOdhMCmRH5ul9ql6vY40u2GjJsG29YSvzMhsiLo8bUyZo
Pj+TyekgnFsK0ny+IGN+uCAAs/YDeRZFUB5F/6SQkut+dQKR9EsGoSEIKSTT9ZSuZTgEzaN+0FRG
Hx904f0JlomHf6eoFvIT5SZTulHKtdQ1768q1h7Dvs/vSV6m5rkj0GrMoRT/l5cad2aUcnL6rexn
wxN7XPXAXqnTXE9eS32V94hCKqgaxRULEZ0Lca5nWL8sKRd1t3nheuDRaILlzvDlyRj53K0Q4sV+
m5cTR6/1EYRoH7JakkYGQWZ7vCGv8KldSFhmGzAQtvbzs9W/aBpyF6g/l7iNmbFciNoX4oT3z/at
odsHZMnxX/+X3b1+b/TAleKCYe8N3wOLRk0lMs+UvrtxKMYWvgOWd7KJmaytBoh3SevVuPzDbuEr
qJn7PiV5UDRuoKvOx4z3aNXrGcFZIbRrgVLYOQZuXO9HiSH4MPzKlzpr/qZoH/wSipiGaO+KK6jt
2lEezxl+RRNB+wSOJJKmrQkhEUQx7aeUXaYfcc1uO9djZlVJdM9RTAvEuEfhRgWssHWZQ/rBaW7a
XanugRzQsH4g3+4vW/jctnIlxgrq7OGckyAVklophjBMchUSKnqss2dTsl+qMfwwKFxtK0wFDJWN
MWL/KvJ/Snpw/Ww0MWah02x53Md+Ab3dIZe7phoUzKfOpOY7p/mBilS3yBM0CZbTQPV5gmwBdmmL
MjsAU81rC5zMbed9wzNT/c/6VqazcssHbJi4dqmNqDTHqWmawVpNErWIU79vxuNcdbuf8vNMLaZz
FImpHH4XS4HL5ScxMYYiLLIACPmwBhWBvaZIsRqN1zb4I/ZnlU99dm3TPeVWHdSXyMvmOrxk8HrT
mKIc89g6htwUqMDkNRcFmOSNcrwcIrWrdBvAavui04Gr3HZMtHY5VjFP8aGYeO4uUfFmKSHrK53K
+skzcK6tFXzslON1yflpkAxbiGk/ZqTQhkSZL28MfvA6YBUD21vJ/L6Y6uG5sF3czF0bEiwZ1lMi
PtdBVGKprBA/u6ADF1lymR6pRWZ0XrSh6KowKrm5nM7kTCB4M/EeVnUF3u9uRFI7TvPD/5kvFhKZ
qOKx0mQFlfVMqlHc1Rrp8yz6ep0EaZnrQV7mPvFwjtRIlkXosDePedpKHvhItcHaqqA/qPosZPQb
4DZLUPgWI+2lYQVu2597P2pbK366xSI+RolPG621sGdsTHq7I8eCW/99mY24aLuHjJaK4BBWBzkE
WbcDYPLe6lEEmO4jc2SHdaDztbJf7kaPh/GnKwIB1gUANTdF8Tvj3dqWa1mxOMiYxmbB4odW+y5S
vGxpE8JVUF819dhNB5Q56I76ak3KBGuG0LfkN6D9qNfcOYdgHBDZt49ASv1ATkWKOlMQsdVb3Cbb
iyjRh9QLT5yFbqTthy+u8QVcOwaPiN3SC2giIw/ADcBT3TCmQx2yvhE051LdjDE5jp1aRIDuNAt8
QlZzChTP3nuOdIGqysLr6B1V/PvPZIafDjzh52E2/A5mSHdMiRyR9TB24QprmcYMsEB4CyIKP6r5
fRvuMVRXPEi94zLAAkVil8kBIJapsACTZ2ByopDfZMkyHGZqIky0dxT+CHfxs3jx+H2OTGpaUMXi
874mvugmmpA27rJ5ltLxHwC4IQQyhEDbdMk1QgrXEYyIYveLU0KPDgxpzXX8iVcXyMTuVi2ujun4
oEFUE/jKQEX3rKlaTIiQr8OiRepOUw7AAaVJ3W1ppOQ71ZyUJ0gYRjCORQCiXdcCcBPMogZQG8kA
vm1Cplr8dbMnlkrwabqPqEfHJRQ9a3JYdnrxhg+C9WD1zEqtTb8iFBVqmqmhpTavxqRFygIkpsoO
azHk/oCLpwtKU4lj88Lb0bKBYc/2sy0PZDjmDxRs+yO/s52QU4WtHpMW3+PHn09KrKpNxw5eqUI/
v34z02bH74uoZk5KhKmLMJMvUbic/VCeQ28qujRPVrz5ehI7ts2D6rrI34Orz3xnEAW2dZaw8/lM
CtqRLeIL406+EWXjTupCEKuHBiIapuHvtlOj7CJQNDilQ70cbe8yEItN4y1t1CSGrzwU5DDFwtpx
fINkjCRN4clHJdNNb/jmXtsP7NZdQCxKanWdu3X5j+7xei2QTzZWhvhV3I0olg6vOZD1gEumWtJt
W+dGRDl46J3bATJMlrtkxRvK45+ZoJbgX7Th5wl8EK9RIOksQeOf1SmvDjZqc3sUTMQohimr2zQM
F3WlBf//K0zrcjrt6XHqdTmMbj74xcdEhdq51333RRGsyFC65cONG+S0840OM/y8zeLguj24nuof
lN7FYi6QAJUY6IZtueGq0iIueNmLVUpUkzrShLHOW+G0qH35VtR6kOKwCYilWhCv8GrEIkKRp2dx
80uLstIh06XYfcVJ2FNRKz8smHOra3MjkySpYZ+fxLPbEI+Wlvhi5i2j7L55+m4Lr6c7CFGhRuWV
XiOykGUMYmYA3OwZEyNwaXNuQQ6C62kf8pJO8IWm+6YiEEapJ44S7AyLVeKtOTTybPzVYEDJaBXM
y8weT4zbPSusiicpztNmii5E/kH4W4U2mkR/QMapZde+CbpRsv/JBMnepRFF/6a8XpJG1fD0RlAf
kW5tblNg2dvRBOmDyUalpMU+Cz4T70f1lifqwY5XBLlvuQS7aRUmwCLhVp5mENeKoHn2TRKinBCf
KKozDytFMf1+RRSk7k0QKc49isSXEmZcE5tG0b7uvrCbSWUfZ0YJm3Nw1GN4NrQ073EL0tGpedkO
ONMNq9YIm4d/FOdUMe4vl1xmnGYgTW1px6EiT/MvaT4uCr7uo27db/tgqJK3+GHe649eMhVVJTnL
nf4lW+lVhBnV//msu4ecuVX+W9A2oV6XwymZZ4FS6VfvvL7tMaH9GOmJiOTBmi52Kr3zFPy6tAK0
C5SEMxgTRqNJGBoNI1fqoo64Vqi1v5bRvN+mjWwxi72pxBSoGG3+YTqPgjZbn7lNh0XdJZlhUpFD
3VjCb+WW12Q9Yz4rHEklVCT3853v9FpLjJBZ9JegDY1Qy7/AC1jVlqE/oV27fpBkmWDE6VycijIu
RLZAR8wQqiogp+ZBn++quNrs8HumulcH8CyV3ImUX+V9KQxxOfO3k5nQY3I8ArIFEpTaPNzYc9+a
ulgQ5nv4NQFpk+ks76Cr3TCI790riQOHC+t02zESYSPTfvptp9lTSyrZSecZT4LGAL0Kp1k1yXUV
U0J0icNcmog3ahN9jZkA1PR56BJRFUttOuChkzAL3tchJZ1IyfJz9p2t+95zDFKAERDThw0nmrSK
V02mzPKcZ+JrHdfrjIQ9v270Ic3iOpQF++uWQAqbWDdeyooMc5DnwhRlf4eoDkLYeKqI0HPjrsiJ
gTLMkvJLBjEKcn6vWXWfX+sVwL71vXjxs+b4aQ6r3k7iULvIDysYEDEcpPqNjhQjbtakqAuivQal
ROu5CGInqDv2oKo4G4xUzLHBN8wF9LyFrPhyHtDZy32g01e2fwfZ88ruUowS4Uoj6iwj2s5FoEm8
L2iJJcBP0rWXCAeiFsQXUNyQsCGtbH5YXBbqxWocn32zoT2IVeM1Zd/pFILfuFRN+MSPX1jyWc8H
3g6fb0H8sM9aSZQWAratFDMF/Z4kSPlIVJ8BnpDAwn96X51Bcv3iPztqEnT9LPSXvWGKYmQ83RE8
FKsYSqJZWNqbM7q1ojyLiEcyirb3IPViZZiZmSqJQ15qYVpFVXErFR93UhQJ8zKmQpdAGMVMi576
gLfdAMChwVWq5Y1ZiAKFdfC9ASlhazE5N+mdIWiNa8GCwCQDi75nwqZH2I8yb7mqzBum+x2PrfQc
a0Dw76ilCbgW/dz19msg6PryqUo3D223HJeu1GfBSv+KjUfZstpzbIt5HY3CSQRVCpKPAU0L2F1Q
KgSbAMS0L9RRovFqvOSGtk5fglq9UcJ4ef34HzgnVMNhQ0u0MDjMn8dpXJeBVxB+SjA5UuH7pUey
tuCQTOoTDF51qy+9ZGx0PizLkPK4T2MpxEcF/J2oHzPrjgvXqF8Bc2t7VPGyYAG9s72hlwcc446/
S9I8SGLJan4mIBeRt83OqqGc3fQz4LcyZY6MvQtrV94E6oGb6L/jN/N4wyqzQBF7uEA8e1PZIX7F
vYkF9vPLhpqgwtOgUgt7E1dOdX3hMpAmsvUFVoz/iwzDYTO0TSv+6ig61wgFdaQ8QQpaEmNaG6FK
5o7B3JPUM+BbGOqdpyfrToDtUoTPOMnMmDz2K029dveZHPC9WQCVUzjgvsr5qoLjRMUXLCTm8JFn
LVGVC2jxLtiruCbEyZCT5hcQhLZIA27IzaZC0nXLsr2n4hLPp/L3u0tjYtqYxD4Ul5CbqGqVNHcX
mfW4wAcSCIbJfig+C7b3jH7F9fQqo605HXqS99AjBvEpn2DLV8Bc+zFVVachpmwf8nzLSLM8Yyk4
cdMstVnohG4JpsUGYkWaSHNXOoXk9EuuURIEsWFtu/U2U8Y7zVQGcTiEzSBa6SrdHzJ78Kh65UJ6
IAliFRtEeZEKK4ycC7S5IBApTnGm/V6tJYazzfpCYjKC+cmGFdLZSyA4FkG4O8c141b4uA393cqs
sRryIuELj0XprLAUIlGv9W2zk88EjbAIECa7xpUtLUHW7RsNjVHDwSjelyl1n1ocsh+9OQyRHmfE
zgkFPUrIT18Nsv9DgyP9uqTIC4/FutnGq7R5+hAIdZVRD77+vNgRQ95obcBfkXvtQ5TOrLHR74hx
ZRqNdbSOIiXEyhakcfIzIIrIyQqK9itMkKiq6hU7ME84JfBgCsRRRcwG29BU5A0SgB4sgkpD1xvw
QFWHw9MX6q8mWZP5v+uDEHnAfBCxew96bUTeeHHYGLjYcJz4aoV2uPJFf2RfbBSWm86LQ78/02CP
DPGc4b8aGoVJHKJn4QtWAs8+GbFBTjdTlOKpRGK+7OHPJX5iKgXyV2+4vrmq6GkgF1iebYzKQ7Zr
D93COT5r3hEGvpMjoSlVq+BZNMMHBo7NKM+2hQ1ujjPUAYWSXYBsgOl4vh03jgvp/CYGixtuBau5
LLQuj7XPWqAYyyMkbXjowVXCW8vdbcWEywl1pR9MxvpD/5IzX2qCPfdBu+6/mVmAoXRGWYFUT4MK
RpA4q3Me6B/vRZOibUVpJoHKNPpnhntAH45iX1r0mTk9UajCOnC8051ob0INybmDCg6ckvgFZGhe
y90DL2ZaVhJspIpG4uK4vO7ftuPUH+Plqad1MgzlNuwgh9EzZAbYcukem08rQqseIKx0M9DJyT6c
xSGLx1Rgh2ShMwwmEIFf9cVQkecqFZf32cz2tkCOscyFyzs69rxUr8YV8Jp9yNT6Qq/Y43ndMxUz
6F9E+eevciUZvWcUXBZ1MiZjnvNeRzeZoHoh4gXYtf53niJEtJMCaTA4pp997TBB8q4Wl4FDqQWB
BtkeoRsL/mwGCuQLgNuohap3y3bLZUZX3BpwYWG8EPxfwjmqH2w0oUrxJdQb55r4TxiM69eUCPiz
hpax6tmmEpRNEtOe6gJI3Osi2A1b617WP9th7YDpvBuIjIApYk8MB+g7RWyKmemGlGGa+W6kgmTS
M4H+X+8YBLlzK6cV97YkLEOB9jN8qQdAhL9SScFugQjLyojDuWUywaal3QyeBzHhC+1TyqgKIYjf
9H6xYfEVlKs4EZCunsLpY6QI8G/i0JJay3LXJkN1Z5GPCVbtLFO57XLaKmAm5bKe26GHToHN5jjn
djF/wQxjk9piGOWyE7CsYxfwKwTGmck9EUh6c/fUWaJHf03VBmDo2Vgfcsv4c1sfjaF0P/f+qPZA
c3nL994sMxdl7po5mGaHF+mRZbj5td81NAC+cBiQHP7MtjYjx88jIwRIlpX8CGtVSXT9gea4PsaO
l3Sxz6eSjehUg6qz2YBBQsWsmKzOck+sMzBv4s5UqNLoVYD/o62ll6v7dD/MsAfKnv3SKg7VWFe3
A6HwFdajFIo4d/uSjmD3LvyVgChDFzhEiYzfQ3uFlFl6xrGxS99Ii+SvNegMqZzHU+HIaQCkPAge
wv1CcnaAC2c5xaAyIZjPP46XCpO3F3r3QyRfCWh//0xbPDQ944cO4IAehBVbVQCW/NsHHkkhlmHQ
h2iuq4dF0djrjoazr/IOaHdsbkn1gW7jmdys4M78Qg1jm+IUxbqjfB/of1vPq5t/B0OYaALBX7ME
O2TzZosDv3vd/1ZktJViSPKSuo/YBC69Pykbr3a6wfLU37xzUjzpvIwQMCKPS2J/Kw2xrZX9XM3c
89cf+65mGVkGiFblS1BDLf51E/VBKAA87govqjw+Fj35u3o+2aTenunv0pAbOmQEls3nLNyRFxLY
vXQkPul79RRs2xWTE2hXde2GhiyFgThfaabuuioTdONUk7GjiZlyuzV1GzcW2DqLAUtP0NNJcYPa
kpJJZWroIXKNLV+45Fwpfi8b3o3WxzfL4nI1LIFkwsbvPO3EVCOZ3NChgvL2onLLxo124Tcex2ba
mibz+1n8DQog6OCpCCJn6QdClkDruKZbw0J/ifQOj7vkBLLRvrykAznnFTKrClMdXVKu7q4ziv9+
wXWnrspvyh74ce+GvY6IY9Y6bUYEHJmGRdQxwF+tANJbtUX7EwGfRyjMD1vbkP3M/1t5nPA/+a53
26lTd/DkxQrphN220MU51K6DJfz33r5IJzBdmR5RqvJK5aTPNysbE73J/JhXH7i6QGi8LHJCyhC0
gpShG8IjY1HRoFMU8oC7MwoKqnvhJgDFVtg/dyxvTZxEK+Pb05xspBuXwZZ0m9iQsIDCPvNQ+HVF
JPy1OH+VLDd01zmrOJnvNpy/K8es4zKTrGVOYqFiSHOYEO/Any0i+2BtMZDSu++odwtIw/+kI5XG
mTwaECwJzhOM5MUuqGT0J58lie82pMTVVs8zSy4Q3bxtXbxQj4hzb20LiKjZ3up+KJDGF9/Vog9n
ubx2vEbSVB83LQWcy+cCCZfDwKO72yaFWYB9mVvLRfaJdtqO8/Vl1RNwjYsjjlWW+ELGcbgDf30S
jgf/SBJ8JniLf4gjrMajqW+juXRBKDp3DYhwEE5yvXUDh6KGFygKnjrYe8QKWPc5LXwCwJEmmE07
cjcKdCW+2KgdfxL0foj7b/0pN/eVcaTTdqlF6VFPPqm0Z7e8rttCz9qMxZF+8k8p/R4C7/xXYMcT
k/+f/9UASseYiVh7DsQG7dKcY5mqK1iaOM268QhvXWRWrFQP1qEjN9tZKBQZvstTZVPeZzHC+pBD
8p86v8ZFCd/RmWNG2QfmdMqva0q58BQNKawXlP1PpPPXopsJiPmyGu4+xnsU388LAnExincKox0T
cbs6ZMuXru02SDr7vpRMNRB2eOPePzTQejFmx654ea7n7xFZq62BVOm3ptwOBY/9yaB3V5FsAouq
9AM0g1fkb2kingby6qrq0vXzbqV78nu2JeR3stsUiA4Z0LVEzMcLgepY8nA3mstn3lrRs6xugGCg
SVQxidlOuUACkitw+rKhH4doN0SMnsfeNc+9u4QKwiBB/3v1peMe82k/89McBJGCOCoitAmMNnVt
dIsufhLT1BEkk+ywKohiLoAimr/FBTXkURU3RWHpYSwYWoNypYEyB+prdlggBdi0gaie9NEoFcdz
KeNUu25VuqbARuabTKMmjjwc4FcjZFuo4fTEJ8Mm5nGGUIDu5+JErwpnmH77h2FX0790B/PxV9pa
U5VtHUstM7c6gBuzADLq+xV/vlbDaHOflU0RcH23kqrb5l5uq96bLJUxdQ1JbF1yq7UeyJD2Omwr
lRwM4cHzFsmCMfWiU11w/EPSk7akzkxBiU/3VJzEjSMqG/QPKg949d2zfk0qLs+qxIfnAoPk9ceh
v+07q4sZ29NNWDLxL8M8/oF+2RS33lu6XeNaE+Gx1dP41s65i73wYRhcd4nDNCEv7SHwgCh57ehc
hMwc8yjAhE8/1DOFzMXM45pCFSgPcwOUuL+gDi/Ih4/IShD3I6E5/PK0SK7h/wKEpjT5fShOwrmZ
b6E9HaxdWWqA6296WW/PDHLGx2KZCq2RDzITkrlRrfXM+7jgFrYh/wi6IZGsHEQoiS9SpBkfqi7y
PSlxWyZWpuzHc1D0s/A0LoULWD/tt6eVGDh0xKse1iQWmGtooZqDy1BUPYGjp0vzCJDGcswAW1Ae
lF5MD/s798CRg47wwLHI6Gsq1tRfN+N8/x7CH/j11pQ1FiRH5W2kfdfrsa8Dm1BuEBbI/JJI8WmC
MRPsXsL+7ZmBWH5NWbLWl2UF6p4j7mep8mDHuTFWnoRRlbRzP9sEUV7KJ06ULwGSpPGXoH73ln0Y
duaZHr9r1EnqP+tFYQxd6xHhTI1rs318HuPOwb5BIOnlpMqihyajwmbh4/XoXcHa2fIWsDD96IuD
TCKcIzbJdSD9ZLiTLvqIYi2ZfpnZp5D9LLJp0qmOJ4doQzUoFJCZGu0MpX5NobQ7V0gzD0lr/2Bt
ZA6M5+Ii16/EALJeERTaOFr5Nlv7sx75wPjThCYd3OMV0rkOehQC+/mt29vmJjM6l13MqYPnW3Fz
CCOd/t+j4o95Eq3N0FW7ic8kW/N7yOpM7KjrZD6HYDaKPbEqb4K6eREtjmzUcnxawuHUNjndchTv
2LVy3TwH2gqCmq5HFbestOaj4duxUoAZB2Za+Je57sZcfKepYo/ymisZPOkNU6SPrqkR6wMJWQqe
dUBLJAHWxWug6hAUBYWhLu8rd/NqxZJT8rVRkqOFfXAtWzsT+BT54/SENjdhwlSpwR8PHA2DV6EW
z7En7xO/GexBpjeOYFEV7mD6CcXFcyfw5iMcyAIMxKTvNnV808I8UVyj1aANbyVhbMYc+UhfNw0l
uwVZdfITamTYTTLQd5fwpGs+LPVCGghWXAt/CDgF8iGSioWUV47qX99WtXj7vJ1EZ0fSZWeGmOgI
lYN1EspbQl22m55AdJ4xjMU1bIQ81wVeUUwy67QT1Fl7eglBIkeuRYB+pT+Exo5O+6vpdozR46K4
Fiq433vUYFgOsyInXTZBtS5pHKH4ikVltdguqe/YOZjxrXTU97l1zq1iYhAx/8R0ehFHZw7QQt5a
HLk32BggVM+CsasG8G3D3kCrwlzpPRyZ00BNPZbTgIaT3XKlHVj9ns8FSeUUiwMNj3q3daJ450/W
QYBs3mTDBRBbAQN7lPe3CQFU8B1eid0nPQeZP30748s/ZEsoyhkZlT6kLTLFLqn8VNQ9yvS/rzXi
TFYtPOp6NYVWm6af4dA/tTbpYRoHqDe2qGgbpF9WdHnX8/58PRhVDtvlSDEhS7zOX634N9lDeK1n
zwgNQ894/t+NSqh10/fiflKSxB2p/mLHfJtFmuSKKilkLD2H6QuW7wWi8aFGANmXm/ZKaqGd8Atu
HVyGv943i9W+5K0WPoM+KNJlXs8VlfNxkkgzouj/Z1jwbEyEqzCH/3jRZC3XCXvIDAbHa3t5p6G0
1AIOkxFX3HM/w+VFGERGWCtK0YLNYGyGZJq9ATkbEvkLVRLo/SkicJWGCHsqK1kthF4cbnEcECTv
GIQ70d1t3VhwOSFvZ/DoK4LeRUakZAa76lMTd6c/CU7QLlHroTNzuAa4wg9rdQoSLlBWwX/78S9K
BGDu0ZtUFdipHyL1RF+Wvf3iaQ2Q0Zrumik+HrzhiMek2IjG17Yl+Lan30dxADUh0mjyqSZ+4zX2
hDPO1JGv5hAY7RAg0Gi4kGod7JongTuDN0YFGqTHXoDUL+MczizdqrF8/MlfQkXKc0OToVs6Ouyp
9WKbSAREH4kwqcM3YIjnnob1BPmR0QAQk7nTLMfZZ1QOGXM5gnDUIjQSElUAhkUPBvdT8gpRybow
LCrfEztJaOuyhsL8ATjeCtbcqLtluHh6cgvCvlAtCabsEvC08RLxturT2s756MFgENb9/bubGm2q
a7ILgupC9Y9kcy4U5KzYGbAT5kbHjhagZuY1u/jcmzDzfgL7HJ5fwx+ykjtvH0z+66fyfskn/ci/
nNDXohEwuMx/JPyhHphUvMbNy5hj8qzkEMfeZOUgpdG19jQkPlYUCeTbWD83cBsoydsLJuK6Yidu
JAuxo5Ru7SadD72+bFylGBCycF2MOnX1cLBuiGQwPO02m1bXOFZgQg/kAYh1YJi1Gy/k8aYa5hlV
dDJ2i3IwWesAmOIpMn6TUzZVHfQ2YwCkOp4MZfuvMCpZ4WPEvqchgh0/Uqft6cvOFSXqfpy9KNWG
eWjmpLfXWth9p88vKeUtDrlYa1nBWD7LTU1iDLFbHH7HnVwrbWAYpWOAKfLVHGgf7jY3AOJUGr1H
Ig1mHXbCKs4PbMrNOuyBdNXCff8l70b8PI07zXfk4XcvxxYjDtNpG7r1NT1J1dNcr+DquP+eHEjO
405rlJXreZas+SrNTy8YpoYf98CBTmweLwJc/v5k0Jbw5BQrCC9KDcYiwckW9ncY/3WTBh+IGUsC
tra4IMfFLX1MFkx2THTW8mTLt9f8qQNComFWUTP1nXnGqIHRjvSQ/A8mVh9opETuvkA78TrPCa/a
SnZ4wNt1Ao3JmrnERvidU6HE+Hta2FmfZPhHk7M1vlqQbVrPhLKy7SpAg1pzPE8s8h1ERwMFj4/S
C/e5sYpvFPlBC9VqeGYYvdgM7ekKJxQMKGHxJKDcchJQcD9Ab6OVHu8p7VLfrLQ845KVsaFbVmOR
UGXxs4l62qdKie3WESz76EihNZ87TDekZWTljzs80qUVqQBJiniIDrk7hEMFef713qloaXyUz/r4
xyYXxYJfWgYYRg9DNye/iVcfzAa1DFnILgxnFUu58631JkmXJzg/lX//b5vmRzRaPVjkzCqkpLlb
kRpX/u8/oY8cPoevoJdDGB1MEZPBOJJ4yyB9gw1cyudNKE+qp1kgOyx6br0/huF+Sdifv2C7m0bB
nz1Mt5fvAIR5TgY/ryblFzK4lX2Kj6Ug5kaddV3Jj5A67sNPaM7dd4yaQcRn/86Vwa1QasGHUn8J
u43CX7f3Wv59Rr0rXE4MtTaJ1xk5jU6tje6esubQikZDOA1c9J+4KhqJOPS3Rdn90lkWMA7AQ3g/
Ob4fkgGzqKXgdvRH5qMOuLm2K0NKsPSViKmpJk99RjKklg9AVMiFw+7cDfwhFWaLO3WEAhdQAbMK
xMP60fOOkS2mroBUtCGFYqtYy+uQQp1iTGWOXJxLvGPOVjTJ20P74x6t36X9HVzk5vnrBEgmFKtF
wb/HlE1wA8ZpjFt30kd+Td9UWxAYXLdP+IM2c0WmJe1u7b457ngcujAHqUZfgggEqy40k6SE9IgK
rbtIwD2HrLZBnT9mpSEQYTfnLGrvatg3s96rUe1V/zNIsPg30/ae+IszBnkjMJEcGptTfxVfXIQW
/0+aqT3Z1UFGuVfU4Gcq5gjrSPfvmLp0ScHyzc9vQJv/KBq/57fkMBXFdHW7kmD0bJDcqrnTsH+V
c7X/4tdF1sCX8AvBQ7AhzcFtZB9lvPJbd32S3psShaBObFMy/cFvtlwLKEhCzvUOpI+nKpuyxfqK
SQ9ckmcBYw3BedK/LA8pMrfhNT3OrQhvkX57+xRMZY6N/nAJ8aiNmoL24HPrn+tim5jQ48F7NcNx
VidLbAa4PWUCrt9ayPvbhykzJvHWMSG8i8Hfr41IZi+x2L7RbOTmpFxmVzs/deJSJAbIpxV6/T9q
jEff5DBcV3HU1PY4VYIB1c6yVFb1yEQuQ+COGgHO5waOw+KiVAn3r82mJ/g7sexijgFM/sSzqfs9
/ywHwVDaTIBaRTux6ezMHtgVCbmDPaeGDtRWDrnFKPItbz7/Ye02jj1Jwwmbfnc73jgIbIfQn2Uw
fg1jtmIqXTFIHxqMyFv/IlSj0R+Cus4ITGo/wOi6HJmrz4tT50VYZ8tDYZ2aGp7lJFH3bw35TUvP
SNPHUb9jzD1L5cugkT214cRc6oN5Q98EkRD2mKCt4KW/ExbLDtuWaBep8R8hJzaOCYXF9M0Uwfbz
98nlSS7nbDtiuNR+A6dTNJTAT8FGpFDM7sjJBL2t2WRq2qzPdnqJdK8QEbntg6eAx0ptLuk74qI+
nQa6LSQyM7BbdxZS0ZP8pDaBvnDLODEAl1u8hKPx/bQ2K/yvxjJPZX+sBsbY37Y5F1nv8i1zLcQl
z521SWUEXqxp6vrXLvU3EEYbEgJkhJky4p+TLJLMcrcwKt2tkLI/6z9Hgsx0Yn3npMez/jY+1fjb
gYY1wbrxSGCfX+3SKkw+4Ct479PdrawYy3mxaaV7pVwSmUOmaQdsrngKrmW6UGV+xghlHMGEOzoN
JWPi+V/1To86Z6FMeXQcgyvCO4MfQ19vvADfmuCdMVfCTx9hT4Pv8ar4ClG35uP29u1vafYFqxpb
Mw8dexHvKUWNqHpzlV0DHPLy0qfCHJgtWJnXkP+LCD115/fXuyB84nQR/3Wfcny5oSHW+XYMad8C
9xdch7KgXvmWhN0k4AMKPwEcCNrYErdLQO9WyrDmUH8a7orXhiwMrop6Q3cCXeMIC55s10Bdimlk
dspq/oJFHWz11NLMTiSOVI3Kh/o9bblYzpevQrq3mN/8H5TwUevi/jnEjcQkZsas/grWSqpc4Jg1
R9j8F/8O7C1zhM6pD9T5Trx56QsKX6YCYr/9v1c/9M6evUGQaYB7tl2QifVIBq6yM4+JcLtwaiww
GzqvP1Gk3KdMchrexUjpTs6azjXK5fScbTn8+q4tzudXlNXLAR6lPvg1snikXRqFCr+INidfMqEE
sfTJ7IioQLGQoRrgpdgAWdsXkiWCMF6XCSfWe5ou+Qq9Q5JcE+eMybEtG6uszqSfwf7mm6bVUZnn
6VRx9LSnSVTAZsSTvS0vQBT8a2xw4d99FHUo8G4EIOEJf46E79XLDhCDnIqgsy5X2nsJXbFuVH0/
epTztbBFR/CEL0+d7FrLHfY8qjfKigDAdfH46pR4QsbYtT2Ms/YYUTEYA3kGgSUysy9+iQRZlfmk
B9P9Wt2DJBeXWwSo3AD6Y/AtIfJ5wipZMCnKLcFvkoDb5mWVfBA77cHidh+oEcTgleD7mErkJJ3S
qmqEet84gRglJZlelJ5SWBRKCW+aocAzmLKfBxZ/jPkNjeUxhmU2iOWsnFc8Kfd48dyvCA/i8Pwz
6DTsWYE8jRMmVDSyS2+9RyBhyQxdxRNZZYpHrjD5IuAWEaCvIozQbrbh+zPYDrEdEBjmW3gCmPNs
ALEx6a30yRhzb6jpo90Xw2ccelX6ht3zKxf0wln1jySvOYX6oyJhctmrt2MtG6KUu6Gi6uz9Ci5W
GX48lgymZk5zWNziM4/4UodC9orb9EPBDI10CLmuazEeONHjTL2T+FsnYo7KOzkrwPPXTNzSndmd
b/Le2Z/oOPm8fXEP5UKXuEz9Bao0uprTeffLnrvd5ExkKYrZhbR446UWtiYo6O3igHYr08zdPJ/I
BUmu5+9OjZv5lp8HbsQc8WmjSS3/fhJnq5Fdmx9sUxIauJ1TkdYEPn/PiHqbMKWHJx35qBWhvQ8e
SzzVFAYzpWq4sXitsu89MWt8fMsDQMMvWX+QLHof//w52/ZeRBhJHdKUbOj7lvnxAIpgmyo/XU8f
2WPjsE1vrxIV2PLff9/xPeVg2k0qjPHhWL3FyYBhH4Uj+KhA6GZbK8KZpiTFv28jX1GyFFM9QToF
Wy2+qiGTE8lY7yXJqPDm62AZGmndphjgyQOqpHOMUQlUjXP//kPakPejP9EOgAk5kMz9ML/74BiV
8GQ3JNzFMFi78qc2TNLTB8A9D3c/nCd3fR8D7cF+i/ZP1PMrmf7RIZ7x5Hguv0ZvFwq8/X15w+sb
56qAeDbe96/sqpv7TZFcZkw3FOA0nYSwEkRxM/s0hoerW3hy0gUpFMQg+37r1vggMImBEWmn7ebz
mh8HgkVi7qDWUMBTkg+/awKBklE9COhXwNgl+U7zYcq6UF8RhMzOIijewch4tdIIGptrJcAqBxyn
zJM2JooPYISmppC/qtB99Qhi27C5Qo150efkofoNiyTBOi8Vanky/V7n1C6TFUOJ8+F2UdPea5yC
0BcxFhV2TgMVDy6PXqyE/Mlr/RpvzTWswIm7hEA7UnCSJXendHT9upwcj3/sR2BYYsXODJAJYtkW
5Jg0LHZ/PJMTWfAmQGDluyeQQWzufO/ZdMwtBY/EPLoE4XyYS5VLMsWPpgEwsM7kJASKNWfEGpUK
IInWhuaYMil4XNIBLaTBFtrH1MSmIAe7Js4Vnv5N/muTTa7Yvoy7EKJzBkpItXHeGLqw4LYf2DAE
4buTgpn1K5GEhRYc6PsmSB40o1YNoIXDyhEEnC+lVZBNoVRCgbtXWCHPBlrgKT8L6FZxT/6RVAHk
WIIcsoyBRXtr0x+DLD3+bQIfqRKFEiXdvdYLE4Gzqn34pcUCdj38682ySZ0XtuLdx+dRLRHN1ShS
7uUX23gFV482H46CG5wMCqibHQvOexGk/x10iObNqsY8sDKJqWU+zuWoSbbrsDR8d8v8F8N26x96
gaXsE0rsfYr7+UV94p6UAgmLZLIcwtUFckpHkcG93B5qOOdpe0bzLnLllm8fOp5i/kkQDbt2s7UW
1gN8Q5PAoYNuHoNYOO0jXlT7cKfr1JKmhpChBXi8Rcm+EiAIvjI0A4HKhBgr9dICAeLaPSsakcS0
VTtwc//GgGE1aefw3kZFM8AcNPMAYzxcb5HhJmzCwEkgAowPq87iLHgvM5+1R+LBDJ9jO+c9FIwz
Q04orWjYl9eOIhYrQllJxMENf14/pPLibHQH5+USJUh9yJogNxNZXrdm39rPkZSI6R9ZOMPvQ+ng
O43BV+DRtzpPQVVVrb9k5hR1+7CezEVydbmhQa4jjN8kEgjxPD4mUnNTWueR9GtOCSwik6Y0iDi7
v+sE9VV/FgFaKjForoUmCTeCpmvkMhO/fBeNf3XC2a0CKaHyv6u1fhOchdTlB7vpCwXClQ1vpYcx
68YXFiSxpqOf8N727aL0tbBW4YAYmdBBPtHll1KOBOaupz6F9oBNrvZ9WShSkGaoXNjRhUiM/8O3
im7ObZvMq22J+IzRZXCtoeM+avJpsX/xl8ym0NZam1u9ZAHuwRVyv4tab0oT2uu+UBjpsqDlCVdG
f8GA0ENLRWwTAEkCwK7XADFREVbMY+zCIcDCBSqk4Aa9g1Zbfw8fkIwbKnn9AUxMMfCxWrCfUJfX
W8BYOrfgeLLfYQfcW2GjB7GlRqP4i/bANKa/780H3Uz0SEwHicfw1Edxd4To9fGLzvZooXGehWd4
6b0MWICnuQ4X0GZQo4Q4lSDaAPBrK6y8hPPfQqkD1mgNt6ffDcXJJYCkEA9GZNMGRiK4HQ5YSbn4
MprU7qtAhfHeh0EyItOG3+3FE24rTw8Q/YLoKfVBgSlKmYjJ4DDI1cEosQXFaOhCLUu1Ht/iArUW
ehXV5TTv7scDia7ZpXjtl8Ca/HXeclUsyCPMTX48ycNlZ/m3tLr3MqkQtVrNkYCo6EdN5B1HTs/Q
ICJCX/FKrgih7fLAT22dt+Q+PS2ub7EES5hk//mOWn3pHO1Id0yvOreeLuvG1ouvr2b7ct2g1mGz
9fIBJxN0A1rfNC2xIIdrGuyVDhjhlR9xK+MJHK2sDxr77/sTvKKk9uqymTRnQ5GfYpfNnbdO51+F
00jBYjCApt1Nla9WPt+I4LZK9HifMJ8f5GdiAN6vTAXyzEnh2Y8i6HAt/nHI6ME4/ZVROe2BmjQD
fRUz7sDqQQkeh5OH74tEDW3pD7l9FPtCyY58EhvXjOAWGerH5lFIMgCWg2QCsXYC/iBuMRd1pBRw
5TeVVk/KVrnmGnGQyoFR0fdscNrMILqzC9gad+DmPZXeSX0yamvRtaKdDOOE0XX5wn3WmGgboveC
MiWYvYf9s1OHe//OOGYcyvLXHuN7H3iJUuRAEcjzjC4uI2DqzUp5o80jgkWPodr5nj19FWq0/Sv+
43q10u1eTz0kUBMI3Myc46eGKehX6ZMMFwAphwYpu0Z0csJPtbzuMPutP91MpyBHMEGSRh1krbvv
ZWxuqe66tekeukOsIT8sZmcW5hIU/2H+bnkDL2GtkNPbpFSoG3fV1PTRm09OvVhZvjI+sY3HlA5C
SlZUIzHtT09rPtN10yc52qVL2puaRsIJp8rVLjS+7zPgQsVfYCRVXvkUKL5/rRJ6LegfBN9q+gLI
+JCPqzpHEppPC9vFBxeB/YakBjQhgSx/lg46AUwlbCprHMKeCMzG1HPbTXN5q9E78aStgPofFDcF
H83G1ljhDSwMCc/kLzjledsT9b4q+h8xYFDKiqTh3bdEfS/ppm10Sh0sCkbfwH8/UnzEwrD30Eap
Xv1wnOMc9izjvLPmtztN2CM1E2cu4dKjE3+Sg12TQsldrXhRko7CGlQLzgg1JGRBLfkPiLSSzb+s
IR0dow5qlzn3wYx6xWK19QvMdBHuO/YiCEN/BccbxTFYMU2gav9DeYB8OKCwDga7iThKjuwkxpG+
baoMwQ3io9joFC6aqpB16H0yUW5G16H5kBNHJaU0iyFkDdzZJ2LcD33BCc0wMysdy5wcNaNfEv7n
0XA0tbHGf/QBeE4tkyDF2e6kLHMXvgg2cqmFPHYLENlCPBWmvKKKyt0dJZzQmCRPLWWZ33LjyZbI
yPgeM3JfO7QnRtQ6eHubivosd30O37WtwCi4vh7oLS3jVzv8JkxO1uJjMkkIo75EWRAmN3a3uSeN
JVtpSZGlVwGAeKGBEVq4kduvufmU4dJ97MRIG3cIGxFQ6ie7akcaPyXGFH/SdMZfcpZslXGH5G6L
HhCB9Xu+81iVRDYJdZAn2pgoEQS5CoeV/fhvi2vcexlfOi4IPQ9ZWU8TPWsniMk3qd4kIgrSaENC
s4NFQ9FAZBtRjBFxpP2RI+AzYHQcIT5qUhihoa4P2sykrY4EwxUkyH8eKHE9s+vyy95TaIKNTLDo
A4AtvqkHYlv3LjYYjQmernr27stvnEHJlxjumqdMAe6Rqk6lsgog0XzQw8YrsL/mbZ1K2Kcj+Yvl
ZoHT6lRBtjHauztSBUlGULF/elsxI8OLbOXbz+ugxTQZpjvKU8JPQebRuxa7fFzlN0vbEbT0rQP2
Tz1Feb0zRylEdJIGT1GhFs5mq8t9CdaV1GyFV5Hqr0TmRGqUrh4Ki8H666xB8YqaiI2WIHhtFfrN
PvMBvtfgAuVCg9NOSVSafttGsVsn7/9A9DfehlwVBzt6nA4MLtmY/yi2whPCpPfoWrYZYZkFvTZO
jPTsMHlRDKQNsCTJzwNAMQOPADODFLAdSFp/ZaTYmrimMJexYSNgJ7VcBMIDw7WQ9/Ubd+E/z+he
gUGASEa+7IatsNsN3dM7aqHanL/WOlMt7ApdO0IoFH8KQJcHRBtms3zCsD+XkLzO+ePaWmjN0FAx
39PWslnd3KsDSyiauI07YDoV/wlslfVq2bVZvcKmJZ8z8kXplriJKiqtDdDtcQ3U9FLalRfBcZQO
+ccwBQ5bAPk37WBK8K9uP/PJpD23srZbw50g9dMgoPcpzudn5vlV9DkUpse20H1//IPDXoYQWwJH
Xhsb0QfPQX/TGhZIninic1SCUPCubqXD3dSnQrDnv98FzrUZcSgCfuxz2YVTqMSsfxxIQyzz07DW
D2cqG5d8pNnAeH8OVdfz7CPN4esxnaXe6lLRHyh57c4cNbpbR5YzJE0T5SThGzP4//1O67s1cMtE
IQTUmXgnpAqZKJWI791vgdZD+3tjgTwe+sRNoME5hO2l1+LYZHmizE14+AkoKn988eDd9W4OqQqO
bsdwPSwWcPa/xiZtUGTlV3kjH42i5jmud7zgEi5FU6wQZCtyZ42rMONlCug47brf/SOLiDQxcjNw
YR1MRpYGq9KYeBL/eunlSYOLl8FQ5vU64WsMrJ1Gy9fnAOXpNxSrHscDuZZS6cdnBaIFYdu7igNP
6f2gNj9RSh9kkBzH28f3Tac1zRkHRQO978DJwer+BO/J8r1uiAXfiNAU+s2Q0gBGS1EodSzNZHbt
Bv+v6XjWl+vAXbt3scYgwfxzB7P8De86pbcALAPyXQ/+0xajYQ2cw7WAghUGbkOLNwz9mD6BBrlm
Irhty5qCJ0YkeDa1n8n3iNXZcRpEhYJ2jVcwQ2w9gSrrndyGwCzHKMdi3Vr2H8guEOVESNz0bnp2
Xm2kUCZb3gmZltyYWDbNbdtq3WL9JeQ/DGFxZfTxSoHRHcpd6SQ63dERyZhV13AZUow0R1nh2cxD
yHX3xRPFeUtUoE+sHL4F5+9yQKz1BHWGRUeY9y0lXguJvYoSCp/MLlYHEC41Gk0nBMGFdN326Xuj
O320S8FPJAqJqpAzsInxwG2AXkss+/FtVys8qVgvzkMcPha7gbyEAZ7PNAykAGUXxpQc/YZPplGV
M/re8ZGqO/0Dcri3oXPEUKLjreSRkcYrQ9fa8rO5PhWRJxtN3+kyBGePtOJZ0/y7S2V/grFbP6Qs
oZNS0+Qv4nuoMnxNhH+tvX9neVOiyRISOBCvaxUN6jXfMFzqhd8bMNVM96q/8opKQSzW2NLuViuR
Oh/GGyYDFsuE2z3vkSsoRBDcgyeiNO5YPy29O9jVWFOFsBqzNy8g2/tlTaMnMJTuYbtOto/tPbgH
nNmYkSLEHrdYOhipf9gY1Uxq4etcTQd57wXVjWmqdJURZAapjyrzxkb10edWTa6TB1eTLS7ava51
b+C3R4dRpAm/XSkc5gbA7/fBAcuzD30JL+dCkTqm0pXtcn/KMXQyadpNyeTm3ZeNAkNtS7L/3dZz
4ORSwbXJd2DRVt4b3kqWoAzItJBm+ExezLum/AiBZ7iiSPVm8cCnNh3aRP2clnaXJ+I5AGass5aO
hZKejRBcB3HH8mnnPGBnB/m71z8eqCNY3nxePXYogy9HFECjbx82yOyf35FDaOA5PwmPswl0zotr
8CaDe2xF6/ngWAt2dO1YY2B6KB5oh5uLu+1jL6xjJ2h/5o30OrsH1fGVR+MfSoIZrjiMfYQqi+hZ
pcqmAkpKhfwYDZCxBgYr0+KvInnGkPQ2KZThWOagW+8vBcUuHp9QeFcA1K2ucP1yuRYekM/Oe2F3
WJb/IDGdXXJBqryq1mWiwQJWElfp1kaQetAmT2J0lc4SEiwLqH0h1216D4ePkKg2NJDW9CHOaYWt
FlwdME48yEMXJHSk+LOEZoBdKp75AzLMlZo8hl+pvfkWrj/Z655SLBUinxkeIFedCXm402nL9UXT
vJCOkYa1E2wLoT4SibwmBWFLSZqdAO4QsOvEFOJYYVJCRXmXGzxS9dimRnV0SCDYWlBpMWbh8Gqm
OBTUvg2cKfSFpEeLYf8vou3jcIvhf38ENZt1VQ/wOpOmT3/wIUmaQrkSpPd8+7waAEw1q6bk/5Mc
29SOgv2y1mE3ByBwaufrQAY7AUsQVPK8NkDbbLhoW4phnnbJ7LajLBEyJ5p0cITKRlK1ABvc4Gwq
RkzwQpLGJfs8EkN8k7UMFARTIPpclX4aYnplBj0Dv5rkDjd8skPV4+q1u+CMQiiOkLjetWpUje+L
MmFyAxvImEF2RY2arJ/uNFB0FYp/sWYqHWCLDgehQip4gZjI3cmAcdbv98zpVmlJM2An7dOMObx1
JeOtr6yoypXeDqLgK9AoJIFX4w0+0TMVAIvFGT0uWXsGXFz53lnkFb+CFpP/7LtSXo9T5YanEhis
LSDzTlt3O+Wuc6rcg9CXOaiFZncHVjXSX8PVsAyBq8ODHVAJpqvXSMUcxRbGGhQdnNlyFolrCTlb
Wqh3ICGSay9MTPSCiZTKYCAcdfrbXhvUBG96eJ97lkZ97ob72JbHiP1CFNI3lRPLHEwd45j8NGQH
1kVnTW7YeXEN4Nr4VlOkhI1LFlamp1Eb254W+FRLTFBmqroL7Q9yHN9GeXLrxkoVH6Gdbfw/X/5D
8CPSjQ1cs8KnpEazaZ9nYU9r0p6Pm7hSjSzJv9y6S5bcoKsrkaHJUgPC4HGBzFXEL1DrcoXxHw4d
bP+8akOfDP1NXbTw6+ZFK0nu5VQEm1HVxVfGXOACBpi/AnsksEUeCeCvRxboaXB84Cb0oK0H9UwI
2POwdhVwEJruE8Aj45gCTWl7/r6FPVEdRB0S7jr8hShUNj+6auT+VY+Bk1ZjIIue70H7NRihXQ5q
hVmFXfq8yHHLlMsK5VTDmUXsQ97tprySqRzrwnilhGYHg+zT1TGLA0Wgc5OYzU1Y1as7ni1NrqX7
gI2FOndgGY0h6xLVaJyrAvWuH1wHGyvvDNdO0GF8chGqswa3MXKyuPASQimt+HNkMFn517ecTZ46
JZeY9zSEaPazCJHm8gLwm6/ShjeUHQtJXjvKWkWMHcv/RYXF016IMqk83nKicsv6zjC5wSWFuFq1
fpfa7X5YwAve0HBeSdZmi4kHOWHKBWSAxUOO+uTulURwzpxmAsdHlHCjeeAveL9ow5IIHlJorgaF
A5U2aY8HT23UnN32+xG/lu0agQmF6mtpuIJzw6Qe0j40cbFGmCC86MmzHQ1acGifhH1+itXDGyVt
aqeUTwNlrh5Rbogko1ohsaYadVzC4tY5RBvmfBY5wgl7x2GGLmW3iAYRpxWPctbJM2QywRcihxL8
hUOUhB4XT9qnwfX7WTdvnKQeYVwH8lYA63JhZACiqtRMZmeAu2Sh9zzi+eyLbEYta/0CYhEC3xVd
JNmcc7cmQKai1k24Sw30i2Mb8ZFikrzQjd0REan0k+YSyHpVKGt/VhzCQDOL5EGb9IjG29BithRY
fn8qpjpiiBp4mi5mkf8dBlAV9Y+Kc5VwCikqPkB15fuvdx8Txx4sA2vbNPGYdxVhQun4BJQQqV7d
71bWy2ht4Dfbnl8exlzFYneu8G0iMHnzwAeeXgfKe3iCdMa5TMM69X3StkFEAr0MV6BO/3CpwJDZ
Y638nSIxNZ7Rvc9x3riXodkiGF90581F7xK1JYXu5o8ra63STX2mnnwGp6073U/NDPP+ReWA4KWR
FWdC/fQkmo5YKGKjOpjQqn9kb9QKnBS2BL8cGdyVMzA9+hgVu3Bj4zdDmpGX/MG0Pv7xDg4r8HdP
w5TJ2GBmEOABD6Q1SnFZxKnzwEMqHNXf6hoRxGTIaXH96vx7WI9weD0Al0dG2YoV0bkBQ+xDGdb8
eGYwCQEBws9dt+KCiOJyKPBiwb3R0myzvkZxoGYIOtniIpO7IB9VYo+V7Cc0EMqTZCN2nApf3d0S
kjJyk/24EpiU+uMRnda4F7j6UBRYvoiJyi8THY5b6nS9Ijp/1ZmRf3x0FWTI+7mgts0bpC+p8t6v
F6wOzDRsCAq7/nJNCg1xOZsf/3vHUVoFhe8uJoQqgkKvPIpnJe9URjsudaLLH3zARe1AkhzthzEc
gj3klXPXySpKdZcx+I3BiGzK3ehqhLeg6QZZjlcH6jrSBCNHZWo7OPi3MwVTZOvGdNX0RE7V0r8t
gpBWT7rzwIkL69F+/K7oDiyfOBDncIQlYUG7FoamSmejhYMzC/f9nR0v/xUc5kgBkg+vOLCPrY0+
LuTmrO+0kd5ENbOFwAlo5h8hKAwOaADcnFquZFBen/b86/uKyH9Qqt9vZwqmJJlL6FieIqgp1slS
/10q203wu43/dha/03y6yj4e8H1z4ymrNOQAuRkFTb6YxdirZG9e3Y8+p3JefA7CNQSJN+mexyVn
8w8MA2lsp3ImddyOLqxH//VwZxSw3e4BVCytEzlmJJgTKhucXIlIBW46kaeKl5sPPdMZd0odyXLH
+JRuMYoh7BsRrF3wYDbPfZGSm2lmnToKU6jP4zF/T7gHfKxj9OevlUkM4j9vUJxeK9+yVVNH+sQS
QNi6AjIG42/TbUGGv24B3ZlbjJC/HVGmsxlYUXuZ0azFZXiz02qJE/noAE7JIGM8JJw7FFThP/yl
ul+vfiKt1sFKCsQClWTFgsjqCxhtewIXiE/lp9o6/agN03Vk+Evq1YUKbEAwlnQ4XVTXuiN5Np7Q
9CPV4WKHQX+0GZ2Kp39hWNv3EkhcFHoet3TslZK3iBF5Hy74rszm4A6Xem3CK/nycM82zqvVYQF+
WHKeXKGykVeNSWMOPmAwTL4BSD+Eby6DJ69KmHtE1HOg0zDFdz60IapBmylU8snv/QEv/6DztmSx
uctdy9yLnQR7boWLjMbd7jQLTd6EpNOTQzi7X5IcNX6JR4EYSqg6n7aqFWMD3kaLc3/39TdE24nH
ZjI/UrPnOCrGHLwbhcDvldN+G6upwpCcHwAkjuT3c+4UglKHsBGPHvZwum1GYo+4nkFHoDnQxRM0
+vnOMDVhVevPaN8AQb0SFSnsjA9CG/h5qTxlYXOqLmQmx5/eQtGTB9Ex0LiXYvdV1cVZqqCOQcVo
xKGmr3PViBcf3ELLDV/7tjuD6l/PU4xXNLg64mmZZ9p3Hl0yK+6aqRXh8S0eTOlf7P743Fm9Lg01
ZKCLRTfP8IEU4IsUVof08TA+Ve54TKhipWPUHbAf7aRJZ937CnTjTR51o5yhHSRX0J+3V3dqkle0
QNF7Ca2ZdlXEBmGi3Ob2Tz0hPkvEqU6KnuDfCUqMpMbeSbx7/2yIBwngxFdzOZtu+GIL6VZ9XZPX
gTf8Lz6g1x8ZiEAGesuktnZGw9pWTU835YdYHdB7DQtw1lMx1r7Vt5Jmxc5oUB59gCIiJo49BXzy
+nqtHTG4RGa7ovVikhIcK+zaB+brLKZcBTzTQNdMgrf4LFgrz9XUWGOEXsh9af/1oek+EYeD3Tma
FcV7eNFj1q5SzA7V3Uv11MDB80NdS69G3V7J321r4G+IiCYZi8/1ZAqC31sdRCmKSUdgZlRErUtS
PL8SOtarpu0VMakQxHL3SfSJkTBiMB5aoLl7bMIDNEkIM9pHdlsuiw+HmXLDad1rjqmR2bQ3BdMS
s9AsZqV5pmOMmT5/1fxlUXZPpVlJWf6na8vdrDPFdQhQXAfOUNGJadCxfuE8zCZeKf6iEklts5fH
Gj79pGGFQSmYVpdoK7HNWot5Njif4638yqaZMih8i1TFLCVTVXoC1jNkJFWaJH269zJjROZUkUlR
omNqDwMc9Gku5STIQ1p3Wv+Qc7R6ef5zCOmaKVX8nnumoYFQEpfbkdaHHCiRVvPYlAlmFocxPg2X
LSKoXfgsT2CiAsfpLRKZML/K4/ipiPtTm7uGmif9d7pP6181+EVJ8A59O40h9Qqp26AZXHmLS6q+
eXtRn+WqgEaH+AdU/5Ik+KSCrZkXs4uWnQ+5N736aN2cK8McIrcrvUq8TG25BnB1nSmM6/bto98g
+S3AyTQP9Eo+AUsGpzU5FeKCFpYKJS9ua4Qq+k27m4Qd9KF1Y2QizeELDIQkx2l8uK5I7nyM/w00
GoMhTNpuDYDfvN4zOKRpPPYmBgLME0yCZKLaZSmGUx0vTudIBsCSxZ10He/Vv5slbFj5pjp6uBRp
9Soh2tFOXgiDvfEGXvsJ+sqHHBIugXSnp6MQPACsotJOjYi3jQu4rHni+/+gjYaP2+1FQd14XQj4
LdXBuHxk62Bvc78PZQ0nbhqndcUxp7mFHffaAMwHxhF1eIUKJcK0EyezxviTurKfB9wXbKFZ+QwR
R/2tyWsLGd7vvCD/Dyz3q+bHyN/TYbK0kwdq1CcjVwDktNxM1CH0HrJlzPq9B029ATFrGMJB5sdE
kUAf4NSduEYe6dRGp49syjF9J9YiWsyAv3p69Cfd2gDSd6GCD6T2YHWT6u1aPL5Ua4nV9UfkLrK+
45o3NJqZP7F7pCOLqeBay5MfpJzvmQRRrYuycEaqEL37AmtIdFgpfluR2sTKi+a2MTclu2Yy+KAq
F0XmBauOf04ABYVtzmdN3WgrMEvtt3tu2HqaEikNvIdTsexGivWdgUFi0ysH8p08aKGHk8cgC1nh
S/Qm7GlXV6TyN+f+6782IqrO2BOdKRwXgOpOwecrrk1SxLn+AhgnOhUuk+zV0k8oTRrEGr02V+c5
oF4wxRicm99b7qyLj/FGVAaK62QVMUJtwpzLi0tt2om3HsP40tsenufdC+xe5uDs+j4y+2v1W+5P
mnYkvv6xtlsi9BZ4saNKNw0mw1iuG5063TSCJdudZOPVRDvapGA1X6tXEHA0SdomUYOoUD8o2d54
m6k8bryPdaZECl25tepqKAAme3SNm0t84qu4OHF+Li0ry9U5fAHwI/73++y0egYlAvnjLDdhh+RD
Or2PrdSQp87jo+tOJPvdXlSrvJNyKl5yk4Y0wVQ+71lwa2s62wW3RrzSrrjtfJFFyGBaeCBxENDT
mQT0dpfIqoI76wqlDhN+uRgXjTFl+q8Z0Sz48rJn2jIIP37Y53/j7qamOEFbpyjPz9f374tEVAEd
0R1mISB1SAwxfGLyQI8ZWTES12ZTCTWz/odpqNho7AkowdoKzGbiHVcZgm4x9dAXBt8dIbRkOpEh
TXYO1S8gTjdtPdaWuFTKJpWV8sbzI22A8Q61Dl437Aha8qMmC9nfWYqLKwDPBwUJKI0JHm/eIPHk
55qHRB5pbSe16dQq1CNDl2AlYvbjQcZFw/GiRtRNfVIlwQB4S+cwYKKI4+/U/1Ks6utzsizmWVMc
K3O7x2/CszwC3kXsmLVswCFnk9DzVlpg9PcbydfQ39rjb7pUGTNmc8kuDW3egG9UfI97qBPzYlW0
i9VTy5/dRbTQwM6p2uCdStBoH00GFWrHD6T38mkMgeFmV2UFQXFKNjAWEhI0f5qVN0cvEwMGq8Qu
jIq5arlPVDUSPSf3NsnkMIy6ph9lPB8TsoKx1x+YXF9Ax3jmrjKuKxvted9D8NMgF/B7WhZgq4wo
C6PN6CJsnJ4B6KP65QICXI68bdDbh6kawiHThE3ENbJNI2T7f2tqQAQoJ8cJ4tPTh/9RUPz8q+mS
rb9NPzoYDWDColY8B/oP5sCRf/o45ACdg/RSzDnp071TECV/0Cx4K/IlbG6T6v5XITrn/L4ibKy5
Rtg7lb3cILaZeMmuN3eLHVgxisYop07JsH5bK//Z6bZ3LXAm4Q54m+pxcPN8C84CYqQ8CSf4FGNc
WOarRlXXFRAQglMM4LJqVree+/81+tLKVSfFoqi2VjplzLmmu32soJFuCKXI7/Wyp+ektk9Zc4Dp
2hJ/5uWkIbQ1+pKFlGJb8kxeu8zezWfW+hto9AsAGqwHI2cEfkVpsk15TZNhy+rOGsUkkR0cy+Q/
ZEIbyHHP3BZVKlJmf31F9G5lnhPhaaptDfLILuT0/kg5kQ3ChuNLOQne7BUD5/8cCQjNz83jRyQI
3neBhjvDKRCAWmxTIj6DBseG5QgpVnxcmKTYt+pnpSnOUzpkoVQdNA8V9lhIifxikTERbj8YcJ3u
vIHOZj2rCIIQn1SHhMEGzB1qkV0dCZf4tRk7F6DJHeasW6Xnhbfvmzb0QdQWJjZqkWt3un6X5BCQ
OFvI4fYCe3Ekbk0xK02kXqugvJbF4ote80iB8c0P161hMxfxzP+FyFeKcFtMibDLEA2CsxJNbdYT
g0Tc58biRCnEP93S585G4HA4IMbhl/OyFIzaSs3K8mtOiiKBo5KLjqBDgGwT5LfbwNWclGLaU0MV
9luQaKsMGQpWlQhzUAsHL2Tba2mif0ny1zslUvh8AtcW0+rtGOqgYKWLbJdKKGfRpC5PXrZnVu3w
TgpWGAwFP3+haLkAGlrTIeJCDmNEQMHR9hEwMrT7gBK1uuWgzhWhq1FmBOEwSiNSQfvkd1ttF2SR
8M33H5PMn4arla1agMuNrusjOE/ljOTAVGfGJ/BprTAyhsQyO3Z0tq1ZO+jP+VwPadKU5R8Mt8Gz
Ff9B2oq4xOHDfCmScd8MSDzASJKuyie1lkJdi+D84G9p6jp4lKa0hT5+AGic/E8MnZ/jCt2yM+oO
pBLI5bCyg47bNWIprhnWvLZN+0w9V1y3FxPAt1Tb6nOz709U+nFr7u4eSqaxhE+asLFP1rv6Xvv0
1/AfkRiPfzuynd7QO5WwQuaZZrboT29vuZk/9ZrxgWgxzhdDEwDuLhJ7roCCUJ9+/CKCunTwGzGI
J3x7f7lzViLENaGVCCAeO4G9dOiDWlijEUEla7dtDfSQaAPdyMtC4qycQMdIc5/AzGJbqV+/wAFv
mWqE6Ms/AydmnHfkHYT+Bsaf7cYX/XyA8oSOK5ufLkbwr5aV1DJTI5IefSiVOnsiBlRsWcaXd6Ef
aqUWq6Z02MS3JI5c8+i+sSZaiIaZE6kDMfSTtsOfg/kLi44N3XBYglr7lNDt6Bl+DE5ZZPv7/SyJ
O+RqRN4na1ZucS3BRxW+QLztfo4F9DVSfYZnQR7JGfLWm1a+chQLfIW1dR9ovW84FJtAO9eaFbJv
/QGJWLTV9lWT0xQvQ4dIgFB2XqDet/piJ904eXn+dDoUDtIIBXzA82tyZVK5vgEHmlizfpDq8ld9
RgTqdBTVOaizSj+cv51RA/JohNFxaGYyKkM5uUtYZUaIgIw1FAFTL732HwNY0kYEqNdYCxbM5dBz
C63HoE617TCc6k126FYjKJwIKjCn7ML79d8ifGJdWWWyfAKWS51P3KxXC+RmRiuMOljOSu5Yu4Il
oRvx38/r7Vy0ebjcG6zi14iMoXFeic3//spR2GJAikJ8u1AJPBRt0A+uUlQ1FSu/u/RNs/EZcGPM
ZIH6teEvI9TIxMK70EGUQ3EmDkK8M3Jw9tTJdWICPdD1zpX1B3lBAbrsNmSWbfmY5NRttiAtB42P
zgr7bgWPwKMcYvnQNadjnajPN/KZzQ9aeu0Tk/QRTDvU7/NcYQJ9FwJhjYZ3p0Z6DkMj1PIW8Hj7
biiAS7+IG3FMCfOrRRdrOkjvF4Y1j18WUhmxFtXHIVdYoUF1IdGRCBM9Jfj8r6CLPLxO4OMBr68O
7cl6fYcoujLN41abRGAv2tpnulrL1CFqADELpNGmzPHeHQv/aoYwsUCKQISuiEx+o0shEQ5OZTZO
A9fVHdIJWu0izYBe0pVnCeefu9m060W1yaG/IkOri0Gi26ZSxNBatuYxEsJ/dljFrnO4ovmEEE1/
xJqtJxedTUTdxOcqur6yvuYs551dFfaIbkb0cw73Ap2PpkOt2kglmQqrqlb44zA439u5DZi6hSY/
iLatK3R5gu3WGocGdRfxYTIIcOkNKAz47L29gvE6wuQIuwdCb6pYMuOX14b/67+lj+HAqcEtc5qv
+V+SMizNX5BY7hkqOKCM4Hperc+iegQqxh5jiCCmxO2zc+H4Wwg6xt+erXDyCsWgusIFgxLvh4O/
Qf75IR7D3RqIDhp3DK2aP7fevgFmXNVeJdf4XqhDBbfa3+M5mU5TZkqI61K4QXTuCmS0Y+YJP3j3
i0UBsvmrCyoScjrMrEADbNhduBWut4Fgou5Er8rBlV/vD7BXFCWLcBLK1XNc2s1o7z3TfT26paaO
gpnwktUMXDaOnsV+41JpPJa2u9xKf7w0v9fFq0cVfzxO9LZ2thzP1zdC9wucqQV/Kx4You1Ui0YD
KbOvs94XzoCXE+ErkFUaylacsWItoPS7n5QFNmS4zT7cJRrkukOLzsH1ZwP4oWiu2vZKuAOOccGw
QdqC9hoNeata/FvyqXrTr3TTWZ9hcfakp83hQjiwV38NzCzIK2YMkPmF7uINqpftCGXM7IXf1UaU
6SzEzBDDkLK3T3vZr+osuzGQ/WKs9PPuW6Yw01awzxhYywGBrB4CnRUi9RdH92zxWfEw+ydnQyWr
M2F4C58quxfpogMrmyOFRZZOWL0/wwel7+g0xSbn7nvhPPaQkxSTMLXqtuGWDMoiblsnNGMgsv+u
SsSs/J8MwTB201d3N84TePEcdjBDmEPM+m9XI4GEfZapY4FcvNScUeqXdZQfYpjJMfitqiohWAZu
0HYeRfXdKOzqnobQPvtd3ZgkSW3arOuXYzaEjHwVJ11NqJE6YeX2+Jyq4t8ZDwssrYdRNtoiSubw
NWpf4J9SPO+x1VPqmKA9SfqYrtbh51UFj87VA7z873Xwwz1+TKzFasG0QsiMp8EqQsjjAH2ujAuw
DtE2CFV2hqVGHyAdNJjVojzmZOzSzxsKcxftA6UDQMj+10vSd+9fMUgfHD7jDop91sBKX9dRA00b
kBvAv2GeckZTlZKf4N9KsMBuwHSWYNKM4N1DfadHdYQ2V7OiStTb1uuLFg2ICSMe1iYG+1WyxPQ1
HVbVFta79OrOqyZuo26n+Jx9zmzdLlszabht411JzIIvIBLSUxtRmU5PtiYIOK1ED3gDU5KNq+Tu
pWF5N2TfU+kjHt+EJlGKvHF3n65jSRtXuuzlN8GKrU596dxrPX7DedBOcTz5tjsRxhqZh9jGEmst
tQ0BLowaAifmPCf0806847p+YCSbhTWlB/zu1yavBK5/QB0d6cMgDE8+7ckIFQA08hdQmZRtwzzP
WbFLRthHh+QDEK5ngWkHaLcC7z/stgJpxBaP+Vxa/kMomJJorxkg4qu//0LdMP9yk8fCwTeqNZOI
u+b3nXx2g+FRfqSDwGr+DT2ij4tijZK0/JQzczQ8u7IAMHTQtb8rgHfiz3FNhXeCY8HNgdmb8vrF
MDNwpQWlW/w7e+WCcQP9VMDPoRUc6falUMQxK06m2/WFu/NvXsi+zDKV+6pezOgKZBoAt6zFPEOk
RyHmeSC+QznnG9lnr+0JsYwqVCBwaQ7FokFG/YdJ+fJm0Pyo1wM5e+6pirM4CE+HwHREG8+jMsZx
XacHaWLS9TNC7fjj5Q7xZgN/NoFCZ0BTWkSCMhE2oy6D7kLjjaRXHmZVZB/5pKj/VtWXIwaVzRs8
8KjfYNA6tVc+Uh4BDOTlQklyGx4SMeRT3FwZFQu70r6hykF7O1RKY0OZIADDEGpNG4uJMRDle+ov
1JpluWDdblHOmJqpfffW8SBIALMYd49I7RpkLed4CRYNpW1vOJxQgKGo3yiMs5wC1011UbyK1fPs
n5noQynqv0yelixeBpqkRJIVlmuMt1DKh+rOowRDln22SlqGlzpHXHqQjQ/WMo+jrHSFib+XBInl
MCUbFIJABfT2spUF1mT81FANVV1wDuNSLnwgiImpFeB/0GZhhgjrmBi+AwXzqlEu29VeNoh+Rvek
gOcCDB7thEYBKnxq3YaBGDsUxYbg/pcmdcgLgGtSz99QlH5L9inunHM/1Y91m0TYukyGdF54Wv6M
oDUMRC2Re8ow/VAPnhukOzY6bV741rH0O93ZCICkUMf2Yl7/2nqyIVP87BlH1q6Bm/MN2tU6pQwj
Anu7/KMu+Az6+5emfeIzOVJHQqPaW0JYVZc9pnIouoOeC/MzE2GCegxdYdmDWhPvifr92Mv/1fHz
T5++o5mA0E8+9IsfVqfD3lEt0ufS6kj6HeUcao3mpMlkWFMDyKYm3YSa0H9qta/yhxg73YnJy6+6
MQUwuxrVDH/kmWPQkIUGrA+LOmdF/VXz1lD3tjuV3HoolS6TSKKQtlsS53qdn6ah1oV6QXdoD6Pa
CBqBxb39V83nGtnOXIK0SKSuHWbqex0r0B2exhLDC4snjoWuy8HrArKvMqRXrg8UlC/2Q0a4au+I
xcpfNdH+tZgnZuLH5tPciu6Z5ksVQqCUiYiqB8hQfP+K8V/PJdhSD1SiYmae4SXXR+3D8q4mTQVs
gzZIOGFFKNa5EVKjEcXrgbqbrvUYPjylnFKDxVmhez/ApTm1SvqRQY9Dc/seo7NNcB9k6zxgJH7l
COF2r8/XAi6liznZo0jtcZoCZoDK0xpKcgcw0qhypJn7j4UVlH/MTbtS5Q9V+LNERGyiy+m9KhA7
Bx9vdH+dM5Mw39Vwj1fyK2/1tLM9zjReJKa3g4UvBmsOwII8bPtvIqxV+7o3T5m/OA8eB5vjHF+b
BlMpkdAVtDKJoz3wJ8Us+4XXch5Ve4OWy3PsC0ciQ6ypWOV+stn7XeuX+OMiHdHaM8mwlZY1lo8f
raqY+pEMQnautpgTRFAlLMUDQ9qJNq2pDMSZvduZcoPOLqVyFQPGF+9YSG3Q0V2+sBsIQrm7NKwO
YHzJtYjAEo+FR/kbgKlZIZiVaiFiOJlpvWmw62wQsw30mDkh/dLvCYfcO5clC0EOkKRb9cPRMRfa
XUgIC1AlDIYgIs6QVyOtGtoymUjeQbxN7VKZVWitW77S0MCxsf7vfeU68mBDFtrNpQMRGMFSo7wN
6f6k/hz7gZ0WmpM0E+ibLFCCbhX40X4lHqeRe6s/cQI0op39WRFMmCkemFXVgmePgVlWi5tVaEFz
uWFczHuPuHjqYaQeCkJLGH7UWPlMZHNazw9+KyYPaMhUYXDWZJiXVGxy2DVTJMo1Xok/LR0Ktsu9
16l9xgWMiQpIqY74zYSHSbHYR+8k5TMxC1t4wtenmupYDZnDdq1jFnYyE5R0ZJJ9SK61fOdgslu2
zAYT4OgoYy2nBASjFex6qrkpTYWawPng+GjJpWo36DpWj6LT1j2p9VsMqFEZu9Ibmr4OjHDMZ0/q
mQwxiaP3+RmvWRXvMkIFXfMqsR1g4u32AfqFE1whP2yirxT6Ewr/l2LcExTnarIcd1IWt8C7Z/UI
lA1s86+bTB/hsTItneo9LNhizjxjvjDwP3cEJQb+KfZbfXRkTkhYyUZk/2yZogeZum77y+xKZrJU
Z0Gzyf/pfAPzWlfHro//hwc+XcLZoxToq+m68be/nrE4MNQ87Dur0EdLoSeOUhPU04nDo5J7H+lZ
Yjs1MZNxL08yPBgJ7eqyz/Sis/VfDvG42TTAuuvn19qxpuEF6RIJUDeHXY1vi6RCCDahaQIeBmyz
YzixJrYBJJJGOiDiDJ2comJCEoyXup3jRHYptZSRq/XgLjsdl6utApODHAXOUvNQJ5GGpKGoLlQg
MKRibWzo8D4PvUs3ENEWSQ7hznvFJgKfc239xk00R+UNREDA9XSGfwFmz4WpC7eCafdj+18fAhOc
bhnK4e2z9At5tCGkFjmRrgfD+LKFvRNUOpekn8tTTDcRJjyPrIpd/sYTtiggYabV89QcMCC906fC
A8ZDSeLNkcZ0wl/R4O5qSJ/L22QqkcLMAuEzKcLA7Tip8jN5o0nNlQ+M8sUyiy6OWaR5LRsEhvBf
pnHtSdohYEQXhZwPNLiszfQQUo9eFqlG1O6Ho8HfAE+p89xop4ttaIy3w+ni3miUsMfMo+N6dHGE
7UUoNYZ1BV/Qv7D7so+kHlzO2NDPxr1QcA/Ai3cZ/qi0LD+qdHEKEsOmJZ5W1EZvk5Invlflhslw
hYDNkQxH28VbQGONOf1F14zy8jw5nn0hQLUjzBJ3CwYf7LKZEDfuAFxykntUJDs2/b8B47Pd4Uzu
cZvNTD68DzgmSerhZBsjDIG9z+ElIyaPe9hOOlh/Ts2qBCOpK5L6LKzJlUQN5a9eLMy57OzJBMcK
/DT1Hk3PQOkmZj8EXDjS4SFJWgpWygihjU9lFcStLW5csCKKdfjTQQ6dl9He54pSA7o/6sAJkGvs
VSSnOunA88D4yULPwgcXKZCymR+WS+E8PYTXlvpbHA0O39Cj4RwAld1n4KnVytfEr9vf9GIW+ylr
vHsjPQEDLIQch9e/YIAbcglXL4K0soc2LbuL8qOvqBc/NQrOHAQdLOVJfNo8agz4vMQzZy/Q2mBn
oBA9g0nQSb5n4k72UCMxemoTk5Giq7PyswlKT2DNJtEBO3osRMO3r0dZOjdq1aFs2ytm0HH0LAI9
Nw3GGVdZSo05vsFAL61CWL3f779UkUVW0mow4Y0M3YnRvXy5SbJeyKa7jzTrqxfe85r832ohiArB
OB53ZLgUp6W49bHSqwzNkvCVCY0FAl8ryyp/BDtUkfd3ZNBzjyYFICplZwSwHodhiGz0r2oROigO
HMEcA4eaKJSxOVt6Vsbu9vXFp5LYkbpzlxUFQf1/Rfx06sFywLfehpWKI1pztMDvmnWS53pA7/B4
rELtoXLl3wK6m1YJ99fPa2faMFyCRtYH5vvl2FhIzXf8C/S+3Kh6lgJMsOtnw8TXjCgHXLJrBSKj
t3M3qKkpEEslPSq8XqBFZNexmPuMxVyLAMBDHbATTYezQLjJrlDqDQfvOzbeGoQFN6GtMybvCZ7S
tdQ88tnc2K8znJSjB9irnnv7nRCxrF6GxkA4M78DpoNB01EVkKZVGjlYVec5WTTEpnCbTu0plmhD
KjHAc9Z3++xvbPyf0ezJFOOSh/pLGgcw+bvfiFMzBedHyU9YqGmm3xgpRozub2SxwV4qtmXqjIff
5gSxCGFB9mhmnhC3vL/xpoSdz5W1Wqb0mOOJQiWBqaH+gwxvau4BELYYdPD/go1Eyrk9KTtpT2EP
IiaXPltM5x+wv3ZqVxUHeIIisS68tBEVuPVY489UaZXTyuCsYOEMXWDENhAPDNjede3IKUC0Yhzj
Ee0mOCnL9l0lzG1u88CxZP0z47N4j8ffoo9tsQ3NAYE2H7/xJRpvUaeOffm9T56gXgVHNParNKUj
5RDM1gWn/2SZampTnxm3tKVYvaESGD9RxhjhOxl53zXR+8nX4g9G2TqjoowQQ+YshSDBlzCwHUE+
71aHhB9NHGgmCh6gL6lVOE2Zpv+fyJ/ukm4PzB3kgLWejbLtxsCjDpZ9B2kb6KzHspHACj2sGt9z
rQn1esGPIEnhOfl9ZMn3HnOfRXLRNKcmLEn/1+sXMYD8mpGFDXv16JZKxSJ8aGOLlwoe6ZI7yMLo
19mYIDvzRC9qPblI3tnSUmYxff4uUnEb008sBZpYC5Dx3jd3JQe1vBG8Nl6ALBk+uwsprbK3Uiix
/6Yz6k9m+0qazZg4rla2F9A/VMaLpVaRwOhYFKQZV9DPh83p5E/uMu73ufrpsgIp51UPnBK0GDr+
khhfb2vPI7xRDYrAsQuyv9ijl0XTf9bLiY/vrQlut5lqKT741UJZ4WcfKY6wAH6Ddaw7l64EujKm
7uj+5ZRoJUcVFKdpdXnG3eOKfvsxPARilO/PJrSNPAUDC82ZPzvwVZG/Dc3vGNn5zdUQAcK3vz9L
PX3LjP/rVTRLLY3UvkGuPvWjbiOxOpB/1+ZxqogCcKImAB/dWXZen/jMRW82ZGFRcZSXSouWeh0q
awhhnKrzwdbHut471pM4GI45RWeGe6oO7XhgTUH6/gtRa3QuT+IKRMqpVAx+hStVgzlPa9i9QY7V
sbmrL7V6+kTl+elaanm8A3LWiQnhhW5HRSkfW5BSxbwzN3seuS2fpD86eNrkFISvTKCmvMslZR6v
XsHbrIhaFrxOrvGoPCkWqmEBWSxEhQkz5YCjMMyyqaNKLNVtHa69Zs2ET5+AM7XjrsGV5iYVnH3N
6ZFwScuxqx2hofb25jknpsZdLAZONRQTO8m3F7ao4PPnipNZmI4l2ndXsma0x8eLa8OstJzzWnTN
dQIQhwATiWQh/iiMm9xKXhzG42/cRZGXcV9jYyBK4QhNqykrYBg+3nMDD5mb/oHuuPuRVNepUogZ
3qo3diBQM6Lo62p2Q72RQvmUOqPjZY8o6l/bfNgdG5ANm1Y8jUk5ZfCR1OOWl3a2Zf6lIjF4/mnm
mKwXIjPrwhcpAGfcTUJAEHbfMTE1+kqFD4alCoxJDwZ2PIEaHvMe4TsCtj8wHkv0MtumdvWzuJxX
wH/RSoRCyVQHt9c6nbTGU/3KIs55/bVUf/YzCBxv37TLFtqqDct5W403+PzdoeLL+Ho8nVW+pbDM
sDQCeg2VWntAzTZzJRvRecUfc0X2HcLfyOhzibptkYjWhJY87vU2dv/oY+Zt1ny9o8rL5jWsrgNl
caVRNdybuCm/3lUY/3f77T4hVk8sBF4GRUz+08G3id9GK4P4grJ2kxNCmpD8pX8E5aYFZelR0CQN
fZzXFppwgM0gm8nBNStI907KnU47iW7sWqp0cgsxrg+xBzZebA9+Q3c4aH5U4giJepNYC/DoV8Ga
sCtSVpQnYbAjiWCkcaWKl0VhD/5FFzxdryp9Nv9XSBWxkre+33fKJdwS+7UmSkWIIOzxFq5d/j3z
lejfiPoODsKdb0n4jIJPr+trrupBXEEiRjUyPPharPlbiCG4Ee9ikF8hN4LRc+2UkUKPLzrH0rcW
KRG2l+UHefAz5dBhUb3SQN4t2qfGhJd1p9ejJMnqONpmAbcB5GWxveK+oxXJy9JQBdcg/OTu9mj5
ULM2WyG2ACTxE/5Lzib1ZAsW44ar0TzcBkh193N97bKkzViP3RP1b7+fxUsr2xPV5YM83E7B0Xrd
hT5D/z17iJpchUCiVFUEpTL5X2YPF9zxj9hZ47bb/InetiBhxVyYhoadtEYLeEBErYzTw1t1ecGQ
INNmhHe2MflnOb2WcGdFhK7J6QQOL7FW+tQjzs7eBJAIu2CyoH/ck0Y92aIluNBiAsrjh18ecjee
YWfOwUD6hudaSbzSWQf/vsKRtRkGVOOv/eeCR6+DDJDwPtA5PcCRlZa2jJhiF9HFI9g+b0S6ri6f
F8xnTDsm7oAHDNrg3wtNv9Jyslm+ZhDvXmI0DmgTTUK+vFIvqkor7NIKlMPW8nkG2pU4tPUK/fDp
kTNtOLGzkSmL5r+KTIsJ1xuweSm6h+xMcNLlcXFaZPqG
`pragma protect end_protected
