// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Yn3tTP5d9kTRPQHzzuRVQTw/Qlo0LyBIOpxWwYJqPcC7ex/RlMP3VRonCNTwcbvJYdx7R+Hmsl9b
XRY4TcPTHjtHNFRwiJciyPL02RVES847MuNikORZ+epfXPP/x5x9/29ZR/4Pe48xd1zYieeMjiaI
T32xKfzhs/URQ8QLvMIPegtjEin3fz2/c8eaSAQ4Q0uWLT7G1bMO96f4FAS4cR2EV9kxa0ZtBeTx
L3xFE+WzVOTRAMgIh75z0Psh5sGEbzXLlb2ukWhLTETh9oz5jLbFnMA1bApE2OORQuPr9D56q08z
W8la6fDKRQ1GIJEXR171N/P75rdvCcYQdprMsA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
m4kW/gUX4d4KxdEMw9kkeeLRjsLqkAlx4i8jHwDXVn0J5LW31Hu6UpQ8T8SKI+16f4jY/8Eo9uBY
8bk1vHBNoAFHxU9cN8264uMxkIXGLi6WNhygGqznoKQLa7rC4JOf98sbSQsRCdFx5/zNNAz6Vyqz
EIcbHpL1PSJrbmxe+vCv16SUlpVY65wKq3omqn3YNikoQtGIdqqj05kWvzHQmC8xn3rtQxp7WXuV
CX/Y5ejgqy8wUutjQIfLfKtfqpzCMVYNzYqySCDnu0zd87/I+xQXgCm5VVyuci+i3I6vAPuMJKch
l5pCRLkOdO7zZhJaaGWaJEerzXYhvKGLgg4bwX4a45wzvUWRlyZXnvMY4Zl+Ui9IQpxsJLoCDJj4
tI0y/Y6FUV5/AvobKcZAzGrfKqs8eeZ5cYdynRrYydo8GhgJKewcKRzUC1cJJ7b2xGTLl9P+kUPm
oehMRPk/CRmHY6rZR1WJ3RVPPwd6J7+Udr9+4vhqTUrPFWd3JZijU4ddfyWxK9S1/sY7rfv/1cng
1tU+nd9UdWmzZr6Pf+NN45DDX2xlERF54ZNvi0VOoO4sVw93P83aLzTUYHZ9lT/ZUVFmA0ji5XeC
ddOjAZXLr8ASR8M9Qt470uegqwphb9IkztCu3SK/+gSmJLLkpz+e4vegq/LSFaDYhFzojLn3cjYK
/1FuJiyGbTDSA+nPgNIhiqjeoBjhAaeZp6FigMVFRk5406J3zoFVRHKT8kbw4Xd3Y1l2Zb3AGcBl
8d0cAMGIS0FSoOJv5obUinPekF6RBkbKc00ydrC6TsVsfNrGNoDpWm/hFvGZlwaaJKIng984j1hw
XdX8/SdJU7fUtrX2J8eEjPiGt64D4sE4JKhBgrFHZbfc5EkQB9QqEhnkUqz4YUiqWaYdOqZrO0nk
T1Fryu9K7C29MmX6QzqyPRXEqoknKdQsT5bLJlgyvHb3f+V6rC7l6cCFzjoNA3VXexFFx+hCWYCH
7L6HCUQo0Mrsfoksl5ojV0RwOoEnDJAOf8fdUNNuUgWePp9nmdhs0HFG+dhtEO8TmT85ibH/eKyz
a0HSkhEIrzgxeTRaFPJol5qwkGWFVH6XRL4nxX5YoeUNtYeExeL2A/6llIBhvCIbPJ4QAyw6kmA2
GpQuTYB7gYdDzBc0vQAzk7m9K/sQ3aRxKGzxtjf8FCMGopCMjHUEc2srixpLG2Xvrre0RvwXk774
ge0vrWkR/gDU8P2n5TVvCUqNqHnfB7jtbzbBDjtc2yygV4mV0k/3T6yrK2weLIOJAOG9dQYETSIX
Ho+osP/ja/8W5XUSnzf4JR4fdq6CAUMX50kvXiWD2d4pXPQYqZAQQH2Q9l6WuOCO2Ulgn2zxBQWg
klkWTxfUUdWpIyhBXNA4lV5fW9cVpEDQmYdJIwgnA4qXbPu9LK0ZxEmOI0SEItHhON/Op9jmYZiH
eAyiVVvM2R2uzWu8xTEYD41WZHyajCko700aQi26/u2jWzWsTQBKYcuPezJOHp65BiwxikWTJJuA
Sb47z06m2eN+XL6hJ5FQgVroSaiikitT8ojhozIjG4K/+giWPsFGbADkwDIefIzeP8eIJ8yrsORw
WeuLQEgqYw119nFoIDUwxOhnd1HVWn5o30dDyABAS79ygODsmONIoORnm4NaDYFy2MMnJ8d3wdOH
dn7Wq9zESXKm5N9qE7w0zFhDYRenV054EgDSdPH1lsLeC4utYu4mA0Nq6BWZ4S7b9aanI+EJ4nhx
0qLiOX/auUdmH92Bz5OJJqNzcztkBh3z4TyAc2THzrOpreBRLQCYo/Ax0j+W5CMzHm0fg5KD56PF
LSIxHQ7hxzXSoQC1OrXfVwsUK6b2vxp3GtXhjM6ARLebhSXYqKm72vvq19yKxqHtCXGvZ4FFbMxV
ntDAWU1ZZUoCEziEvswa88ADUKH1BHkVjhB5j0eOACl4yO7BSe1R3XjCDe2evfXpyvzr92NuouE8
HOOZpe9C+L0z949hMGKlRw9x0DRspoafx62b59zkrXBnTMlyp8xL2JmwQ626pz15+bdTi4j83NiI
Noq7u8XlG9shy3gE6osh+xoEnpmIfbnroAVCFclg5cOYJLRUxEYLZ2xgtdEWQM8eATavYj5SLG3+
RMnrGYb2gEg0Iif53VS4v31WqLWWuRR+oJIwQYs4ITimHFm4EIO/XEd/BxiT+/XbbwOKWlwi/uQ/
vYYRpNFvDQaAmR7mDyUGHMOvt1ZwXFhoCxSDo3Hd+fCYXXnFYvjd2QxpA2o4aULdaVY3NFTB3aJT
FRXI9iC5hwzipLXXt3roXvRdy0rm7MGU0ShLyfBarq145fIb4ZT+iaOIwD+r8X/H9B6zW6f3sLaf
4xeVGw11ho17JnbakHz64duiF5wiyEBZG6R6U9qc7B36uI82D0Ppv8LUcuL/LwtFQiYtgqmd/5DQ
DHErWlA+QJQYynl4bbSjL5QuX6qblf2UtRTe91wVllLIWX6oXkbF7tO5f3ryIKDkyfLgqmepGENo
9Uau2m13UOZs4bypFA39v4bwD5RFp4P2U06UDcf/Mc6BRQkossS3ndhz5W9V/eBc1iLES1GpnhlF
I3ZI+0e30Inw5ry9kjIQA8jMKzfu1c9I+JAkuEB1y9mtd5IDzkqiW9LhCJvCrX1AQGHMr33Dq2Ni
30S19pJbYFNLzlasCmmSfembZfBn7FVrnbBqcQdohVRINEP8+8EN20qvt8nCm36rKMxAc6YJ5PCQ
44wK3Zqq23QsbbkQvQZvr/sdAnATJjgumSTQD0gTYS8iJufQb8ZNWvwsv80Y5ObDVtf6CK3hOrW7
i2gvjMiSrn9VPvtazZIYJonYKSEThw0eVezQ6sNYNFkW7GEgkt5MdJy/dFe8868WWmQV7VYaC6ms
WsPnTj1a5Keujz0SmfGFwgCx0IrQusMgxj+tGpQhUGXa2U/U3STXZbCwAaVIKcELsgplMbGERJMn
FMBZqaS7MlAlVIBjC3E9pTIy/q5Q4blqrfj9fnKuzTEy4GnO3m1/LS88/witqjuUgqg1jx4mW2Cc
gF3hHtE1EasyRnRsPBrAhJE2LkcG5kZiGiRpxd4AMaMjlI9kW6VZgaEbnBSIrcJgedJpA1+tu7y2
5AjHN0gYgGtZ1+GVO0W47/HqCD5fslN/Bv3si9mWbFga12CNf1lfGuBtBSTmWvObI8iDBdYSZZif
l/0ppiPSJbVul1dCBbxyTYeICtN5jAlBu/ycontEbtZgRVDmTOPQA+FZzY2cLcyq/bQ4YkDf82hU
6LkeF/WUX2MahXQJWEznYYJac2IiJfu27Q+PEgYPEzjndjuokklWo4AVvF9Y4a7grM9xkotM5SOu
XLyd8i1D3CH/zkYBAwWQFzJDT2zMomQhxgN7P91QrOUa/ygkRcrWReVIWVHcHYcTeIImv45OIe99
Stc5zJaeS5CudyXkFbwzsDViyZoUUoKA9aqtLTD89hlHjnnC442Hje8Si5GiRqJ6D5vRBF9gD5cD
yVAZx/bZw5wdL6LvgfxQgJR5D+VpFKdXEJmmMgww+FQPLoxokqn/QHla7Tpp0L8qvb6aVqyWcSmo
xo/G/dOWi1h7r6DoYR9IFnPimx3BFuullKzTDlhIfe5L2cFlm/y1WnGvn8bxLOjp4lXZa7moE/fa
o1kQvH/uPT2oeC/VUQca1MjNKAGVFHiARfGXVe86qYTRGC+obDcFBTGHRb1o8PUzL4/v0UmVifkT
Qg3xtbY2QCzs0BveBCa5Eh7dIJhaQWQyOyZ4PRvlEUpNuKl3dpH5m3nTMYg4MXdxOP4ZPdLTugAa
zj/7ad3KgMOW9SngiOMW0jfbCpYD87+RsUEHXvkm9jD6JIAwjX3FN918spQYRTUHLImqkMYSC0Mj
Up9mtG2SkUt0WhcAqgA+Zmvg21Dg2GNRbLF4ovBTZHfjip5uOP2ZlI/OOAVFY3Jm9VDMKmlHFhBi
S5enmo4oIjU3NWrdmDQryPYRA5xZ6kgor1qFJLF/MoCcfTikAKFtWYLzGb6oh18bni744KZuwn5v
VMs39Cha31dU0LmcTacGjdTLAY3JGNZO4gYCRoz4Lgu7d/jQ+NecMOvMyElAEfDzxUsSa8wf9NEe
fFl1IjZtt9o5L6eS7ix1d1RDqHTX4hvyf+v48RCPafxnpIoCAf+bcb/EnUm75W4wvqJjvkXhdg7t
zaQIzmT+6uAm28L1j0O5mwyogtoAzVagwnji04G8KsBa8JGpOgbKRadwS0VfKYnhSz2dEGd5N5Yy
rai2wHZFvWsEQSMllcUnoFPIojsLZOec57lMKTsd1UG90qAOrT1ZnN+bq3H/EUZ1bB6QUt0Cax8j
CSy8ZFreg7uPC+9BQAXhMnbJEWhVFmqRUONMXM1hFOe4nlkfq95yTnonnk7EA53x7wbDNYQCKB/4
BBtOfnauMSBewijzMe962S8dJu0CDHck6vnD6UUADurJBIjSs6QQHzivYdiJaIhp6bsCSHQcQOSM
k1/p6i4caaIDb7T1Pl9nqzWfaZLHYIXHTjV/SzSGC7F31AQtJ4YYer+fcNOGZZ5H9fItC6YOR4wS
tysczLlhaV0NcY1fQWUyLvzN22GR71Nm0BsQffTXPZvv8OlNR4AKjx+aZ+GCz6J973wjGzeHA6Tc
90EeHDl2UwaP43CBoskrzNavxeGAOeCII+FwEcuji4zMw8UiOCDQ04/erpzGD6rGssZqnDhXiId1
79ZbFEQo79FH4VW/mMJkK8ZgxMH4IyqbXXHweTyQm+Ej9xzTURkoWAykjVGdTKOF5b02BuKJ4Wkm
VEkRYmV43iYtEXA++E3KyhkPgFScxm3lIqEXpTwlPYwGvL0yjb2tk3aQoybgJhRZoT47FJ6iFW20
xP0tuKeSB9TtE+JxTraX+MFtCg7zR660GPGRZ26l7VJ/6fF8UfMvUt7bWcLc//eU9S71QgYzT3tq
87gN0f+PVMTEbQI0jOWkSZJcCrLXAQL5EV56/ZhTeBBOTqWJ5lozAed7X+0URs3pmlAf1C27DT+8
yUxIrLe2yRu0GrTl8z/p9JcOkGKRG0VWaroFUS9Tn0zM1LrGRQrxZS/7TVq/yZupEgV6HldgGtMC
snFdgBpV1SwUsp3QVf8vemTLN7oA51VK5ovbpJZAFv3sKhz/bPKi7BCr9F3jwPFytQ2010qBNDfl
VRe+ydoMCfyqUvK7MC/Bf3uvNisI72iFh4OWeQe2KV2KeB0XX4qBwQODDRFgoyZXO7atpbNZ0u8L
WD/F71ZdmJYl/a+6cjy7vZVZC3LqW5m1jowv8ySGFwOeGI0fauAP4bWv6bhKXOtvcDgk55VvzSKt
4ujdDv3nyNjCWA5dUQ0bMVb3QowjAVW96tWHDsWYb+GVUTzcNbm3hJtUy5j+K2xDaGQFMENTw6mN
8jN26l+9W4EE0Xpb0EDZ5xZDutPwD2KmNLjHs5TwpgZ71V/h8I1TvGwbWCOq9uxJB1utWM3aE57o
kzmk1uIOEqY6Is7+f5pnEn4An03r6HhNSwk0BrGQd7YJoMkzS/9JsuJxmcYLfNkOFzkobVgVuU5q
MI9sH5gtvCYMdi5X0UhtGE+lMsuvJ/TEHOIpL080MeJqiXmzp0iFiwlFTckwlm85lJhIUkufresp
7sqb0vgqE27p3gJHRs8GrXHHZfeVkipkKTIPQRpDyzDLd+3GNYm1q2OfC/dVlpWyJ9cKFtUKbYAK
0fR3C2xw5Md5p/sP1RFdZJj1FWNS8+70JoBnh7jf1IiBPyaoWgyLDDuNbUT6sO1yaOQJ1+HZ0GFV
QuY54HrFywxdxgibD1oYTyyhiIM2K2dC+ipYKRSN1Og///crPzSeTjl8JpVe+BeBCMmWGsvbSvaL
+QC2IvudZ7ZGppiPi7VA19zb0gzKPapEKhuhkyTf+ZE+uzmeLGUnuwM0tnuoD+0L9x5idSHm1bel
BqsLE3fV9B4P0hqm/wgflbzRPly4Vbfk740mH70kChHHNS3uu2CFRpkZD1H9GSIshIJwCOJcpYIS
qdzLzEJeuaJ0Lm6sEtke6ETfJ1Ko0sSBsbGiNx/tjmqVtdrW7V2ezn4zBSgW/hBFujssL8A7zZw4
QA3Yo7ieYDZlJf+Vj4LZCZYzw1JXEe1ms+wWVMnoejWqoInjqcMQUh+SGgoTXrM8wR5rb/QOoWDk
5tQVCfRkXeIQb3dMFVGuKN6096H3TRV5Q6nG0owMN8YP6lfwObzigOYUkfFbu6dPaJM9lRRV+CL4
WgYAwx/5Y9oYrRBrcvhl1T0jJswjyjfwbpAApmEBIi3+mcgidx6LZDu3Zqat3N0iqF9VB+27KZWL
R/qDnDSrpR0PMNm0XnFEMaRak7eUTCAeu5ognJ8YsqnWpOoW5eiv7U6G6Jksao9XYdoNwc+i9Bwf
WJ2832QsUkQaAWyn90JIJicMXucKfc8DAo7/yNYqJFD5LxGjugLptm9tiukGTNNaPbqv+N47H2pC
beXyJvY6I+qxrTiOPDwwVfd8miOF95UHbNe4NNVAQ8v91bstxrJgTD812HBP1V1htzcHB/q3e34V
VlauoW93TpaN7gYfkzC/zjn0Qt1oHV4eTJCD71pNGuAc9OtL7/pwLJqJuPklQXfUzuw67d5bHHxR
ibhD8r/3dlDabJW5L+CQz6AAF71cu7cFWLUrlkG5WNFp/TlsPqQCwc/a5rggpNtOtyubJhkV3D9y
TWCnmUDOR/DL8wtjJirVAvyfZwWvOPZ292QPs7aDKmk0fQc87imQbx9rkt4reWRq4kai41snvLc+
7ApN2thPP6wuwEzrEhaNyrbFvEoyg55MJjaru51F2s8H/Jcm5/4NMuw8487cgA5Emv7gpcI/Ja/w
l/eirxihLXaT93FG8dDtYti97fCTGpdOL2g1hx8c6zQUwys/G+eLCfP/cr26sMM5xFDJtD0ygIni
B8SaqpOSOjLZkpRPog97OGEIT/xkQ+kWpqqBog4MGG+ZC/6UnPt4QnmWrz2yg4ksnZ+wSlFnT21p
UVhwRmEwQJiW/2TGMWsbi+3i/Si6LbLFF035qPUPE1Zass4kp9nEQrSLRwWZUhBnbox/lvup2j8E
ciJO/NdWfQL6BJMv/VSC3y4JL0RbUtt2ConqYf3UQIpW/jbw7rnW+AqAf8CrLJ0lRuy7tZY36z/a
PByERITrv9+wTxZNOEDjJItdO8PPIy/75lSNxProfzTyJaV9tKiCk7AkKmTNYjNRdeGunuIYVz+H
2kY/FNFSrCr/5lTDDytaBsQi3yVLDaznBYFpgPPxtaE4ALNt34b1DQQRivsLa8w6UnQy1jtpLyQ7
ZpNaDz8gg5a3SnhDkfnRG5FYCnjZwzrlH9DlxteN9LQFQiYkB4OMeHiTl5kwqqozmPXw8SF0/sj1
Hrr0jM+LllN/6ACvrkJ3bUzhbFcKi7SVt51SMtQFJJUxTajZNVhLiqCQCb1cyK9abykzXfEWtzwy
eJL93EVXMrE7pJPGBJZyWLGsCClo6YNXk4aZLfcF9ntoYVx2wmKVl1aajyt//iICeLRi0mkC9dMM
7szgNADQ73UBd1lhixbZewP/1bOFZjueBO07N0f/7+mpGi1j3QzOmSkijWAzZic3663RAHNU73ed
eZSSFuoVsxDhMwSrc4WxsKPmrekB4EdCH26ogEmIeJ89qadCDAmovvcneWGval1+KZHmsPr0UAFm
Nis1t6efofvB+qlRBqFqKnWaPXykJlGwSA+z9ztcNiIhyRYT/VZIcK4bN9UYbQWiLuHi2xmdtOvR
P9bhbIGpSGPKNGoPOe7RmQEOMdGb9zQCspWmu2gcwnaIcyl35WVI4G1NIIV38yWhTtIM52jIQ7xh
M1E76FZVQ8KLPmok+2nCon9TlqScvA9o4ZSw8MJrfwXPtBaXzYxg7BMntwSOn4SCoFvnCv7XhO5C
QIgBgOr3IWvRCPoFNkCw8GRXFnfvWOLk16Fe3B/OmAk8NeOCPwvI3PxYjadqJsMhQQRgCCpJ4oo8
vabXE5MXlqku6xmvz8A1kkDv9bm6KojZP1mf8m4uchqBlr563/nAj6Zw5fGuuJCUdLrqQFXltr4L
nhxJyieQsAAz3w479TnZot0eKqEyj0L3B07tcZ/KomSKlyhRLWPBwk6FJEeFnFjMiZLDFTCXCDYJ
bCjntPuphn0JOVMoL+hGDLg/hQdvsNzJaW5PC06469B8QKm+Rq4hhuPpkHcw7AGcd3ESz8smKGiT
88S0/g/hllJ3zGNC4Up4H6zU6nhvXU5wS/t5H8mCfp392FCwiIRmtKwqNVER6fnzk2vTDlfp+7Gr
du1mNNz6VhRX6T7J9rTo3IfSG6LZalui7sNuJNgDU6LhZ8zQ6maGGeIkR/LWcOy3SJrEWs5OremI
UfDlOk2ealVon5q0gUkAeePE5QwlJYAFM+yEwwxsCEmekANc2CnkUzrLEUD0ZjLmXWuKDDe7vQC5
vGLEbIKlH/A+cqZwQxloFpYSjLYOnmTuxlQTjCe3HxtPULWpv9i98tOmBjsL0an8Oxs3xeSSpZHa
7KeT5n1QZzMsPk7v9K5arejH2hcD4nDjINtiaDRqM/6jyJ8gRAGRUxBnIoa+269VYLsdy+VG7DTl
drtRYJ4cAW0g4qceeqDbBT8yj5pdwGcPfqJiYoGCaUcTcKLWksRo/sFPrgbTnA5b0mILbLcqtvfV
15cCybfepaHLWKKtEHkXZwzYPdXQk7e+NqNYBZgXILfNttA1cXnG7k++mEwLVnUnNQOy9dBG52uw
6YmKMUg7YsqQcLtF1l3Gu3pSHynfKdBgWgNP8HWwvd4Nb9U1IcPNdXy9+CbEi4rptwHwEeHqB+Pt
JVdw0TICTo7A7HbyS2UmP93mx4F5ofb0Gk8e0ht52pTNBfnhMWkN7Lxiss5rBTrSpNIvBOlPFfRQ
TYZ6q/mf6EUbokyNHPCqTDwwRh2DIdNmxj9CB/vY1DjaWYWl0dhJUWkkYjzDaXFWJqEte2YTlHKI
IWPiM/bCZ3aOkkNMlqjwmGVwqUcTOSxocF9xphsCjxP0CXiZBioSe54HIhxfFw0x3HvuTssIwtnm
QIl4ZdAKoi6JqFCTglEHbpW7BDdZMfheNiuqG+kKyZ7myb8HKQ4piGtJ5CBe3Br50RfgP4qjkUbd
nDtK+obOTSruAgt7GfgzzAlXCnWMveoYsOmXx8o9dBbQ1e6y0qICzmhy53bEhfA56qdy+gyY11eq
7C4+D6Djy9IO48caS2sw9z1ECbEIBPHORnQgLj4KytI20kORV9BiBqVXTBi5QLYzlpozCR7SoUqd
T/8WdnSn2O5iYHC/KzrsM/TynY9YwePt1G0bWpSnI+JA5PHS3zEKsvZylS9tvHPs018ivNvPCNeb
w7yLm3KxXK2OdyL4I359auXSyniYgI2VvOYr7iigWLAQF8C8z0JpDtrYOiseX6z+7KeASd8QmT+/
LklqKFJ9eFmFZiIoxB0fYT6xLg1WR2AH8X1/+NpuQeFylbG+6fRPufXnVL6I2TbHR4iRu9E0b3pq
wEDyFkPVcSB3dFs1VFEvPHOzF6uFOdM+7BoXOnttEkcIUb/cE7oNgZrfRr/0pHdN11/oPnh/Ir+1
2Ud+owoeG7Ydqig50s40wSttq2/29HEC0yZXkBCg6wlBjPIwTgeFJJqQxiVjz1CciFZqadEVhQtc
WAD9fv7mLNFRJ1e36ipNhAk6Zlf2QI7c8SPaFl4xOBbhoaxbaUPaZKvIev16WKxiov9m0hFGvqyA
xjWTxM8Y3eSZPnWX4OLQDGxmd0Cf7kOoDdrHGCgEZUwxbN8WB2AAaIYa7Y/DhvEXMv0tR9r3/su7
3lJj4SKlGo9NrGVJmY9JNaY49aDLQmcyFmpLo7EU2pm6j2X++zFDprOKsO8OhWK0dSKYwlno61Zz
bzkWRUgYp+ijNgHD8Ivz9SFzxgUpiGk+gjrrsm91ws9t19Vchj4k37e41WBmmubGvtb5DbT1gmxn
yqbpTlqWvIhcb580ZsD3IgtpYFcJBrhmtm9dmKHK115iuPwbqRRZ49qY7O8EV++DGhIwvPLzZIhs
bSXmh7CDGJFI+G3qALtwGgNWhLwkJkN4/0a1i+QzsuAf8QtGhi+zM5eAtAMFWK0TNuY2Wy+d4VAL
JpuRRgFjgQxBj1Hm84Pk2LaAAJPQJJfzspFAC/qx60xIpkd2vvxXb5A+D0icfJIONAUK8Vl+x1Ut
jK1kzg2ChDo9UYLfbHPmrITwkO74m7nVh1yluDWGZeRkvAaAjNa1e+qhxmfr+CeVdd1IsIPapAlu
2oP0QkY/3EUkfvMmjUGpMybD2sPZ0g62K4VzEgA/0jnOI5So5+Gc4dgywvDqOJIpPsH++tdlzFue
j1LKZvHhYi/AbBTqx6cVB4l0WfQV5s7Ejwsv8Nsac0X5WIdESl7Q/C5ULJk3qKV1hArZXt05Py1m
XeS3L9ynpTTYAKyur/QwJKs2sTaS4gVYuUGrJ2Qtcz7qG5rWeGVlJvn0yrZDohzTQsSx7av7ijLC
+UwDWD5GL/soDdWOnoMsWEGEmtgxTFE9TQJmKBwZQtOXkUfWhavNP4L9o5wFGTrNldIWjSqT7cSq
BN6sqdF6PAYKC+YsYmkObUXwYmZx3T72SL4LCyhCFMmYZWy3+PC1/HyZoKNnzvaKBzvvTkVR+lha
aWCLwsajLGy9qkYqVjaxwFSEUGhN0+2/ZIYqPM5DJfNxxM+B
`pragma protect end_protected
