// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
rjzttB+gANiczavKfYOSsNEjwOL9QOqPYAJkaPmqeECBn9aiR+asq8Xq0mqDsproiaGKaOi3yWvh
mAAG8irTaCgHK1jFT14swS+3d2UMqsqCWmCAbWGgqZ4bQ7ekzXkGyRacV6d+BtZg8NwRyO1GXL+v
5W8rNe5u1JrGvi0K5GwXZB7E+72IYTmTxofFa7JSfxbLQd7enh36+Nw0Nc7Nz4bUFGu1mI0xRy2n
xsd3zVOiAS/7krPfsLN6GFfL+xvaOTBcyLf3LjSHkJulmamlJk5dvQtcuQS5VhshTPn4/k8h/HYe
kD28zrry99ULEc7hskdpxOIIuEH1TYc94ivF9A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/R0KgmjGClBs7uetOmk/1XI+JBFn681UMH40NMEzCo69J+rOAXFu2lhqP1NAk6avCAYKrCTiP1yd
zDg+xVzsjV5/u6mwtNmrhss4SjPwmY5pKHzQ7dvLDIyB7TUOsAyniak/l4QrrQ5D/H0NMpMDd8SZ
ng7Nzvs1LceDh0zXQnJPHxmM7CsoUhVhkda0GXkNhW/jbBo2lLOJxpmedZ9yDJprxDqDV1CI/nab
nq6H7eSXlrQxCOtpMD2H+WrXMoFQJbtBlrWbWR44p1CoEnIct2sM6fg9jV/uXyjTSwQbxQ4y8mYj
AjVPSTcKH+kVGPlhR3zWOSo7g7Dgvc8a4puw+nrXt2hiN3/sB3SxdmVKj5k+PJNw8zQHaY7Y/+oV
5TQG8Hd7VSLkUb1CKpx6JHkqWbSqug866i+bBonlabvS5eoxmeBTWplYrf16kjwDwspG6SN0URGY
+twnttWJ7TquJN6fp0KbobFUx2FmbFyvi1b48BXcst2j01bAS7uhAJofTRW7rqm1NrqvM9QsgTx/
EXj5m03m66F1PmBr5Pn2sExhNQ1uF99eznDSyq7SUtoa0slxLKvh/x7t9Fx8cfEAi56NfasExp0u
SNJtnarbjVlI46l/8WQGLMnzN1P5ctwdJcgVi0BG0xcUd6k59o9XYy4pTqLjKDcg7qMwiqauTNI7
SVpjfInA/0+4Zy/mje/nSd2Ye9B2FRwYXrFA+L//U2w6JJcxNIXsE72UhB2Sf1i4j+PIRaKdU7AE
CV673h2dewv+VsPIJmOz8iyeYITBT2SAVZCrBUu3I79oQcj19OuwZjMv4apZauwlhI2ngO3M8hZ3
WtvVr4DJx5TF5tAySyqxFirBjfgrQUMbuTbG2/tEcpOTcq161zHvdKeoXMwDXzmtGJH8ZIPvWYWW
1fpB7KLdPyjKw8ukXpVZW52g2rJzePCLpPkbHlNkHwIojiDef6r+C2Itpgx7XamQkn735LLFSsaZ
SMZt4wMryj0FbXB6V06Wc+rq58OhWrsd1yxPd4fNmErYJn2QaxziuHnkL/X1zRrAWye6rVxV2bXj
9IgQ70jaA6O7EUlPlg8W+f9+IJg5icx366PiTbdsmxDsaeY1ZIHI1cDpNu+oJlK2h/fKWTh/+jdv
JVGwx5nQh8s5l0xV/aZh36dQFlKtMZEZFJN16jPpU3Va2oXtyYdyk2sMruEvo/KXRbBT5NDRCF5O
MfkUnM8Joz8Msn20E4HwJXakyMmuFbSdYT7ZaYRz4RSgkEkuunUweKsVDtQVCZydMfcd1xS6D4J8
QTNBcUm0HEwClItJgqjMLFLHiDvy39NAYjB8NcODRSuuAEBlUpLj/E/VuKMnRIZNCIzaCi8CCeog
12S9xn9dgi4mASoJ4Q9m4g4KU2eL5672Fmr64BzNAL+ZYGkBkeQABlVhph7ixCJ4U5rTUCK/jp6V
gG3HPm9uWNWhruZBQImOiNpUPyW1aWg4QTEtypMS3J3EqrLsjCj2AW1lV8ZDRDb7GEkQ1j1FKKLS
wbwLOpwckEmIsHQRoaTzz5Myt8BZlMO49m9yf8PRqMup0hppcOruXZccoXbrGKDpYcdGr/hDukvZ
pIJp7RAABYZj8z7iuP4gEozGG7nvLbJLniYUtrPz0mXlyuHpLgu7Y5fN7YKt7SRJPSImqyxZeXK2
2LbWDLfX73QRhbYtmuilr7Blr564RNX4jORoBd49F4SJvNKZWlUVH08RowpCtJf/3iIZescfDjdO
9SXSZFpceAH7zprt6DExUzPjgl/QitkjNZ0D+uUltjNldUkbac0Tbg2sDi2IwtFVIKp1CcoFjsPD
U0D3rI0KoSSPQcV+tbNiiwFU36Ey6WVbwKBE2lABD3U7pjf6f4AzYft1/uGoI8emws8n4zDGMzsp
ismeHvoTsMW8OHYIcTRNO/HxeJ73t1TkHUziauEvpbF9K2hdUohqrA14uCRcLbg1I8Tcd2ExRVVp
9snjW1cATkzSUwxMiHJ+xUHQEfTEvymXmdNNMgk2fCEdfd8Yj+HYzmlo5zYJ8C+OIP4bLOaMYkj8
IgpW6X3TpCO64OLDl5k7nOWsX1bv6bVLng1mXq2EtVvdZu/WMUzZk5jsyxAtRbBn3AYPPAxX9PHf
N+w4F8Jquk0iyp8Q4Izwzj8fpmJ0qxp9ljkHUVK5p76o9ifqeyj8fkeJ+UjrvyBpQYIJ3d2671bQ
8Eg3z1W/UWFuejl3S1RCKkbQqawZd2z14YZb7ry98dZRWLvv89u5voon4cL29L2R0gxRkpfWmAAv
AeK30ITsnDKTtTZStc7O7PUGhF3/YATRQNudZ8mi09Ufolm9Y72MxcxJyb/ZytbY+xK12GsGUO89
M0H96rUhWMaGTA25qGXFxkH9VSnnbaeaZ+MVoly50auYLXNu6q8Jlpi1UBoHIzSOHw0Zf5dHwwIv
R4D2UJj/nDE/73ZyIXl9dB2cuhPZzMMUXdr4ZKGdOgbVgdcGf06R8iN2iyXDKmsO96p+8uFMfiO5
DRryME+yE/KwX0H6H+snOLHkK63coPVXw9d3U96nbBte/dHZQ5eySIFFy5yZEqpWbww7HVi9rMZG
/ybslYzbJxVgCP9rtdQsJdHZZKWRARVkJAYMjCyq8pS2VXtkpMnHOj8EPXldznt03lwSaEpLvSd1
1QtIulLt9y8wbb4cXTHdfisWKfp8u6ehGhH0ZM4lq0eGWlYozVFV/p1Hi73ZhIpsP1dlcv0xSfP9
Xh7eQ8u+7gO7M9cAp25JeIy1IiOizKlxePfGssDCfGLrZogoetdrKQlDXa30L3x9P0fYLaVozPqH
tE4ABzF3kYSx8ewQGEO6CDuU6i0KAtUAJr8LkEO7Hg87EnhqYIuwbCphhPdl5ShjrdSLK8hfEea7
GX3Ab168ZMwggk5GkkD0SNchkBkRoOW/l/JhkUfxWCMJAyzf3vMGeaa4wgJtQbtgS1yJqF8KCJPM
qHX8cUn/qalLnjaI+//wMEgur5cWRO13Pn+td5xI1RDzWo/IlcHE4Kogaezn5frvZ+6MSLhzH+QM
293dy4Q8HVExmwAbqr4CK48NREOENf0k5K9QhnW3ful5hwlrCSLAiTlUXVrjQv58PYf5W5IOMwfR
82bHt307554FrW2NKhe6mz57nhtTuthDI6oe/Lt0P4yhOH+mbVvsOOKDfa3tu/m1lIEDyT8wGGEu
k4O08tIriyJupXbQFR40XrwabJCXsvh3jV2Gz5Rf3TUL5cDNHms2rz3jIfuu4AhqhZIUSjBXV6aR
0X4gpE2RwSAQ2NG9B1u5ZtGqE2lC28kTBYlNMBYEjYrytfo3TGVUuA1xG9sRb3ufiCRsD9OcM3Er
+V/pYStynj4bnzFDwzXL4e8mZuymyR0RY8bqzzAk+vAtqqvZt6ibDrMqhpYaz3IB88rXyDSqBZ4n
1WoR4Po3fcEe6GgwFzfGm2h0SB1uHzVl9iIYn3jVmzkJiUjQ/VFNx2wHMnyT40MK6gl45x5/kWgA
E+BkIpJDjm7xIehzA09nWZhqvr9Q1B3f6zP5e+jKFEy/TZ1ptoPpIuZ+s+eQR6rUPW5OpirrbiVM
qsoZZcKtJ3DASTOxP6n2xOQRs8YeObXHptiWxra1pJ50wvMM2vP6YyG+ot5fbWNinsvo6RLMRMAp
1MP94fmAyXfGUdMnqP2o/WqnprQdW09G2mnE/kmSX3p8lBDr3Wv0YWA6ml1Gmlhw/L+AjDeXRoVv
Q2O8hwan7fKYnfuuvTUWzM0XWtpTy95S0tmRAI8lVQBFa2PSNOZ97wnoXRu54La2szbroR7+b/5O
0zsnRFNAKKnVvluCkMxkssPHBOcZ7Gue3+Y+PCmq1MlSv8ivmuBciPu1gMfMthHtRevhQYwshiQw
vJFh9U7+C9ytxOD7wogAyKpIaaZ/UPeSyRT3ArQ3Q7iXKbEokZbutmgB4Vdl5/zh+dzj/AEW7j7T
DqgotQTOWczIlorxrqsX1MoHikhCWqJXI3zUodiE2zuX569YwFK9A6H6AgXoTfXM0H4Gm560hJTJ
Wz+H9OHcPtpxJV3iNSgYYrmbYRFS1e1dxG/D2Vu7C9EMIseLTrgcnwNtIJG4Ut8hQG94+2dauWxO
S+2uskT5P3gxpJDD/8KrBVyGdpLsobm3fJ0fjIuwMDpruYBjx/kZJ48L7ON4bAOuY6Tve1T0XnUE
4CPflaGoYOAwlj72u6VwF6qE6O8YgzZY7PmOEV3BxYdD8tkCSy5BBllK/5Efcp2FUWt7X5bRQkpO
ojzZCW/pNxEesvyg30uA3zYesDVhrTDHZ7ZbfLoBsUDyVlYn2InWDDX7er0Wf4b7dQ6dmMc97BWX
+BPO9i8/9G8MVIou6OYZXRpVv6TlvGXUkKJ6dz8OJRrWCatf9ltZ5X3DmIn05bXnbusuxzwFvCao
StHJreDneeYPGXRXvXPtP6DK/qio7zk0hAQt4W2PliHN+mq1/+LraEMV9MqWlAT+a9rBdKYRNJU9
QpvvmbhocaG4E6fUZ3WXBQ1r8fbDi8x13PC0z8aRdHY00xqdoYjIsDyd0Gn12p4VpdA8rDv5AolZ
ulfJfTD/oT1sNyIRaB3uMpGNddjBkp4p7QGajwK0LexDe7UEJEYBwr4iNimkplurzfqlWRctxtdF
5r/EEHdUOcz7ntTOUArlJlclKo1+dTqcwAYMM8HHJLvyw+cn50D1/stzUELIV9+3eYW5U5/Td4um
u1CLuhhInRiLws4iS7mFS9C3kOWu8fT3lqnbAYK9yJL33H9QDG0hiV7TT23jRaRfrSgqH9yf4y3J
KaR0BpluTfj+nC/M9eZE1caQFx35SZXC5Gr3sdfjWW7BKyEA5KsNdlZDVwY7MhnocscSGOZWv2J5
CbRRDuFhBSQmNEhuODhwggBqFnmUq2A5zzvgN/FQ14xGdj03+RcPqjGHeoHoIF52UxgyLflpqJQB
+rc4fqYXFBlA8CE9oLko1oMj8xPevTtKV+b72kUPVo+iT4SrFBr6vPMRV5k9hBxnKascG815iXT/
pJNKDf9soNcnM9ui+wtqjoUFvh2dEUXerEtkWAjRZygpMV4E5jDUzZpCT5jAQl+/ulqqiFNXAl0w
weX95XkF5cGQo4M49bgRpINbUHYQhCb4UaLv7e1Gmw6YJoQwYHPhC1Kk0xbsa9F/3rpcS6YpbRVK
XWZHPGCbY+xiaK6iD/o7tr5MWV008gnvCv9ojCPwHJ3MbU1zi1mR0MGqcHCdUIE/Uq9PchQaM+h9
foH8JgKsks8WYrpzrL8DMZIJPvy51NTqipUcPJlbqD30l6m3aUTFKgIRp4FRMbbL1LbGEmrBFQwH
coD1D6qso5p5GyTE4c2ifir1L07THduHehZmhwvBXZGIJMyekd5YBQUf9aIUFhbA6KAPQhPiroUr
rXuFQIRc7JKtLeGWFi8JqXzuHYavOyDRI3H/HH4pyYh3EyOnqFHkVO+DFWa/5Kq6fnZvwEeL8z+/
YEMXeOwj1NTO9Nf3RZK1AmIx5NeGg2642d7NrwKAJLbXJnWyy5sTSvad+IWJ7pY2DRN242D1cTM0
/R6MEJ8eFYB5dfKeCNmSuCtPckCbnvDFmLwSsC0Ehi5TTp/XgAdGwaJJxhYPQeTi+5lAFnx7jtIM
4u6WHM6JwN52o/tcF21Bm+YfeTSrFfPZG3sEFP0ckBGuI0Cnju1nu9ZnH6lgHT8KbGI/MuiFtYB8
RxQ8TLrPAsxsJovbwW5nnby7yto9QA7XFjttAXBnIUFL/BvU/ybWIqeb2UZ6t0ztUxIyveZdJ45t
EvZHtkWI7aAaRAUC0xy+1OfsVcEueIVzbtyACgDI8n5vs7ytwUq6XdhmgDt4EgQx9VDpwIrd3+oI
Dus8DHaMbCC6chpdk9vIp6KI9SKV1RCHWeGvvUE/RHuzet1VN9oVLbHg89MyRvYPCbPb7O5sUBuk
qR+0be28ZADhIxcAyXmdqGzi9HSeYR1mJ3IrBJmwt9rfx56WcMLGmL16EsVxXdGyMojb5l8meS9a
WqqRxZC2qFx56F/Ml58yC4BZVO5cAnBHOKMO6pi600iDeC4tzuRZY9W9DYkYV7eGycmTo/R0NEPV
nPvsRSNgN9Wf/2c+hlqV5E453o+98KmMzMkvcHPJ+GKYcgX1LyDMudj/DVPLD0xzm/rEBTxOkPmV
oOdm8otGI1oJRDEP4WB3ER2yHOlwoizsLgMAw3svylcZIqN2RfFk7osNkEBLc/fBSFt+RcWeTUi1
qFvOUY0ixEN7+tLeyQ/sxmhwcP1+HX8t7f9zC3IA0vVnOlInMzd77e2GH+CRZToEf6zDJq25ydde
PAVrO23wkW45ixHnw5ObbQitMKkIHzKBb4IHtDpsbQ3jdOAbYFu2DlvzjbuYmQ8YUiHGmM8oLMse
w/5Y/I8IlqXJc1cYa0aNXypv5JrLIPqj4MThWtssDE074vqzWRQVdy2xjc+4OfYZZl6u1jOxQMJK
USNgwEvXYTb9WdFTmZ1mECM1N11hNlpR32cuCSlFfrtqMHQwLBH0ygpBYNhGIS94UVNRDAtypbwn
IInJlLwFTxwYVC/sFCOaFy4Rjr4m1kDXwXdij4JAI9dwuHrSjWLG6Z8Q+3n3o8dDl2MIaNsSOqCh
jhHPRrfbC+BZ6DXD/tasQk/87X1i6U0VrxhveIln5an/4BbZSMoHHGyzXJql/dywnemC2886MWKi
MdWzeYfjQmH0aGfv2Ngz0D+QRB/4GByKkYRk3rYUCOdWgrsLSfxbpj3uF6aJY4V28qSGJ1/zDTnt
h0ErHem4UCU6j7LS4uffQaDAviBEvlHbNjVbzPbxSOkhyCU1iFpXdHuSpLCzo7enpHL/tSiCX9Yr
/wf4wyHpKONto2WCZC8CAJyq+3MJIHLWw8DfhIWvEhpKXbAxjUgpZh/fs2ga7iAAVN4jjqzq2UbR
UZ+PDsHyMItjebcC4n24X/NSdV+AQ5BhKuzjjRX8RzPXf/l3fsTR7C7z5NbrMFGT6cm2lH/9MTqc
36wSao2XvZkL4PW0RL5DqkSGDExCsdqp08ER8idWhBqV096oZlATr22o5njLHSoutOkv7wEZZvIg
Wqu/CP16wOm+pxq6YIv/tJQIUachLgbw0DEd5aMVO+mgn+tjcUjf2gn0BivjBGZ6k3dEFOnd9TvG
1Mrf3dPCKr+PFnlKnhANlnvAkGbSpHj+hBSUWrVlfari+9qYmvVkSMLcE/R2XfzU43Xs1z3xYf1y
n9kW778xtbCVg7HcDhoN5HDwdscN/tO0HJPFUWQgk/TXFRsT9vBly8EGZFD+y4wX5pRAp4cKZV79
Lai73b/O25cDor5S46kLD2zBFk88twgfDiQ0gMz3svA9tRw0gurMLobAk111ix3tz1MSeTfJRrG/
qu+BQN6nbSwmqh5X3fEzeYNknZEs9tWMgCaOXXHHWpyfOLlYw/A6WvpVDaBgzw1JjbqFKY5HL2VI
iOFlyN1xpFmlKS2unopudOC6gaR/xVXuM1XaH4OSJ+Rcgs5hz3LYWfSC9nZ4MDlpgTQs6ENcl5Gg
qCHjV4EsB3XIISO4a4Z+B+j1S7TLalRsH/6XwOML46UEQZw40SfXTTdUsElucG5CEv2L3MAB/+yC
e1vTnoDJ5r02pyadClsQAayItyaWlIyUV7PRgZrjDn0qfS8t7h5OnIC9iVf17ALK26H57FthQOAb
LuZHhjHT9WiTu1vBHEqdZsJ+jFtn0p7v8hwD9niGRs+D5HfHFbjX6usurdVyDXEJoCLDwKBmIgXR
oWQSnS6lUsFnEFPUpcgLz7ebaI7Xah56+H3dyOHRrTSTQ2fQXs00PZra4iJbJavLP8m0ftWmNWtR
lF4SAMGvRf2z6FxofiFbSiqvgXugq54b6zvQPixoZuHVpijUl0fmI64iooToxPtiil7OKFzYGGZD
J64z0zmAG2t5ejx6O7flohdWzwVoEO1lMJbsVrAMZUz/3L2uLi7G298D9oo7UoYqpy4gSeLn5axg
MRahkt40iR9b244Ys1Sm1iXEbv9grNPAmPyqZCWr29oM9VZMGQqnSaoS9A5NG4P4jC/kPoVDfk9d
Uz+Ow5zz6oSB8Chfps2GgQgE0VYnnnh+XYzuGyWN9qbIbruoFbwUMv4U1j35gRo+NPkej57bFeTH
OEnzWSDYqzw47IewzDxvGjHP4HKNtbmuMElsbRwUoehfHIAlC2jvkHk/asdnB7KhLE7D2cx3O4PC
BgM+EHtVCZ8xaaoVJFclYZMsmDiDhK89oSM8HtGib2Fn1tOBCKflrjzcO0PPzl3CWbrFVEhrufby
yQ4ASjBdmdjaSYXmd9ogKy+mlkbnDRfwzfiOGD9wXrYNO3TwjzhBtUkj/hTSXEvnIg99AgQhrZqc
8BriRcFGnffGJHaWKAF9tD9LpbbieGyGDCJyCmy9J9EtoE1jB++qiHSIfamzKdUBBHEOsbcCd7UP
ArL88aUmFRdxmaq/FZwSfvolLeJNth3Rx+oaurwss2UPl5aWi/u2R6johSi9ZLNVnSyspTV15xFV
bAdtNaRLtQW70B1V4FKWGwJwFu9yJlKBESsuKu/DSWVigJQkH+psZ88VBdjYHZovG3Ov8lanluuW
v/Q6tSV/FGMFEjhJ/5Tx49N3rBO2eBbW1aVZUlk1rpFd6s2qofsbSLm9iGJqmRLetP+mSlgW9MpF
nUZW21zGbyXC/yPUQ/OinAkRsFrvuqeZEXSNKk/JB4MwMvoU8epFFvDtvNFC+pjvMyXohvivY3WC
WH0f/reYANwUaayoJln/akMAysASIB7BTEE7SCmOFLetMjNHKq0nHTqEtDsHum6x4hyIkUOYgGo+
3FMcVdZO2UjoQ3CNZM4cg2qcecit1T61cIjrAMgc+nPe8vQlBKh/CsigKkcKJAoWe4lRsP8F0xns
hLE1suXyZfQNBvTuCq9SoGbq4RTA+Eo+WTaD0C0VuvDWKqkxktuB2KLYhsqz1+JxF/1DeuTFcvqG
fwyfHZ6zAtYynQiy1E7btAdHIvt5QYVHXYOuu0xQ9mNlEZQ4i38CIMHS0p0ySWjEzWxVDOnh4TDe
JCo8bSNE+MI7veqk6ixYv4ixorBj+x+B8nsJB6RPNAH82Kr9oqm9WUOOoxyC7xN8Ub+f/YKQOSzI
+lA8fA5tAMel5yyrgFiVP7BlfA5uLX0Okh3cinkLGGrYbunz/EQyVxj1JKc2oTlEgpL/KNLERggs
vm6PzoWkLBQ0CmPIeqUTHwbEopRlCcJk3btGhYclemLQ4FXuFAfjWCENNYRKaHMLVDtzDmZjtKfY
7COSsSUrlT5xtC70sPpAHKD1VhvmT4C0hesre41MTknKW/nNeh5yV31EPM3IezcOeRJkcHQWuOwh
ICFkAVxV3iunGiRcOHow/EKdtN+7lQNLAW4fUuhTdq1mq7RvXH/vpiaRWnj252+/m44hrTUrlvuT
9Ax2A2fJEPEd95LZCuFs7crfOk5mORl9rXwIsWn36Sb2GTl6uQAc64h36GTAT/d3lDKkkQHsWvq8
WxewIRDWQYBlYAcy0Y3Q+tAolpdQ2JpJ6JfDXFZkp00qEWKsXazUzbTa+0GLDfYEIoBC8Rf5DpBR
aIRQ2IHvb15jRnVQ4N1vL1mGO2oVLtFbnCIYjDaN8BqIORlKCCy2AzbVSD1O5sVDsaw8XkQ7JOZg
/XrhzZQ1vdMK36bkQcV6aWDYC3y04LqdpCUCvJ/sbZvdIpLeQvzy/ykDw2PHwT4Cg/87Zpetkrdl
6hZenohKhUyhbIPN+ub3sQPHczi7btYG6yXhhUQXSUIlJZvNUxxkZEiROZ6lJ/wYxmtrs4MZ28Mx
jxSwSgnX8LcC+JWRuHjLZ9RftZn3+m8yzJ8aik8Snnm74+uOpRNcnNHynY/+OoowNpcj1uSsg98i
CYEKS2e5OGdM/6JZf1ocQnh7eR34A2rDdzzZwobZnBdkWSk6e4S7lzazO6DqCFab17s6OgAfHLCT
rRpLcHXK0fRhTo4VFP5zc3cUlb//q5SvIfya3njM1XfevT7SK40PzXoTvNSzvljpn1ef47nENEoJ
yVRPlH0VZm4jKjHYygIbN+7H/zk3Aetdf9MhCcvUknF8FGfJ4Sab6U+/r6OKyxLMhLpREYBhiQzM
3UwHy53vfS3j79tGY68/ZLQ50FOuhldiRPbBHwN2mUTJPArSkaw+lhCH+hn5zksGUEZ/xDDNHpQD
OraaeRj5caJDP85o6s6Q1f+T6Sh+FbrS5fYExDZpiyyeXiur6MrGSDUCJTvkrIjljX+Kvi20voKt
PuaWcNT4wflws8AIjc+/x4tPozKb1rKVWx/hBcAAjtiOmUF/iC65xncdtHNkl2kvDCtczXC/SZGE
c4gNYebjxWkraSljy1mSFa0HFhPupuVa3RCqOrbBvy780zXV7kT6CLxag9JqvYpJilOU5nIz2sR8
T/OWPosNPgxSxpXbW8HxJ0AbTINswBZxiIQt1fZGIM1e5BqVlSN9o3N0H+H1rhlE9ECBEI+55Lzy
NgEs/pcgxs3eCjkhgkC684l2SVcWzbqRFtkAYDOr2+wZBFETRdMSoEQ6LuT41XiFoejGmVAnh6qx
WA7NnJtZLXf7677mwpdb6hYkmRULp4xS/INlniXrel+k/WZJTpI+4QDJe0cb7SWdq+slhI3eZkCq
DfnaOKUONxMUXxI6FRjOecrAJ/esegVUTBkO670GN8E/31KSrk+dztNQ0FVbXLSkUpoUFyNCmngR
yKsrLNVQkxiMr2e/Q/ZoLk3L7dnAt+WFwZ47mLBC5Yuy0R/ilcPw1EOylLmfW33Hj/zUuAHrbJk7
eiqonGsJsHBgN+TYCsXiK1f5fPHMJwCQ7aZrwehAHDQe+ZQd5d+K4S8VD5IhAVfouVVYTLAl2cOC
IQDo+LweZMgH9+HCnKG4IdUNbFtScEPxprqLzptmfhErhLtD42ajTD01EcnwsCmZnC5INyHOihMv
JZVgktpRZylWdnJYY8U1Yapi4MDk9Yq61LWhOlmzbJ1u6pXmdNL6qZp0XtsGVxUaTBRdCnET6YAL
sxjzmGEFr1NgJl8S/eP43uKtymPDgwLZmxKkxRGKq8lD8En4sT0rVu0uVjcpRvDi02zGUa5GIt4b
Nw+WWU0jXQItHWRR2RB29Dw12RzoYsInYLsfG+8RAld6qcGLp7Ey5j0T2stVppDCiu35/m3bsGIj
rL1jkiUQMAe4Yp42O/bhEoWTmeqjUfU2WlI7n6yqMuZY9wSUGZKdC3JMDX0niT9eKhLrD8CfpHJn
3+eMFwEu9uq3K7qEezUuUp8b/kGbJE31fUpHxczaebVJyMxDYOAvjYDG88oyHshQ5r/91ba2HV+r
qUdE0kzbup9GSuJad+xDvdK1ma7Ea12egtt6Ash7S69qJETFdouNif+JhBsTgBNK+Pq4giJ8fQF2
vV9YSTwsuQdYbbR6fNXYMiGSOT4Cul6F7tp5ljC1pHUgqUZ3WGcNcQqjuOG1rPsmdD2tkm5t7MFQ
PCwxdm1XCN6AN9/JxlIgj9CARRIGTqIT0QhLCnz9GLUXTSTYW0ANirxv1qnrgWFc48oaoFTEp1gg
V+YH5Bl3vcj1D36kYQPrBDWfsQFNFPPPyTSepjEmE2uL4hOMfY4pqEaiR6jWz+dVWu0A1gDNckl5
R2fo6yUxzeBZJ3LwBWUSlh9Mxlxm61a4qBskKkE276tiyrqfQOaovHyrdJVODP053ojRxNKAFkf5
KjCPziT8MtnTTiqPceQ+q9Wtmx2VvvBtSBAxB5yluSB8QptALxldfI4L8OQGs7Y9Dkq5I4zhVHo4
Iw6DGkT7pb8SF1ilNK1XpzemBYfzGqcvax72aXPlS0b6i2Q2drGZcL0dJ+7fMu99P4Ahvjk1zCPe
8CCnVtYELO8hRB0NoZmDGYnfLxnyR/gzVSXw3LsNQ7X/jReXn0FRJhXa0zp8AmLOpqKDO4iNWInN
7u/c1YKwjFbvOFfHT2alPnYBNlMkXHfXxs3iaPqVQLBbVJDKkA6ujPfy85NttKPGBkKBiM8Qxmy1
0l0igNr62ov97PQ9Lj2zkWJALimyU0BnMJ3etizc3l5FYoBVXvjSt+fY+sOumCtbJFi4jicgAcKJ
FPHzXzWXvrsmg/IV3wM44esskUgYD5DgZPb90CvIUm09olm2UMG7SxBvEe7fbhKqXxI5wT30ODIh
ELH9r6BX4krn5Av6Mne0ax0OVjPxxLE718HV0oSW3O/z04ThzH3NOoc4kKSYKyGZ2lA/UhxpSgOq
mYQGoKVLVhV9udItb4qRhyfWfaVZYM8+JVD+r1JxgqVtrCgsx/BjeQ6Ooj75IMKvPe2cPWK9Xn2c
P24nnMip7fExanzosI1kdcCUtrTuTsTrRGZ01QZ219QdM7xblNvusaKEInXSMfjryPhOyfGZEgle
omLSchemu/Iu9xk6AuXe+Arz31YIDGEVaet1PJEV+9kijCiU0N6UVIc77x+QybuDzHpHJlHTg8RX
tXRUo6hF9vvfej6BIhd2vvpj58PC+8gxrLbO73QJOfURHj+/nrboL5bWo4AXN6azTaLKQ+ZMScuF
l2iApc68Bhww1kh89x4m5mfPOYxe0evK0f0wDXE+ElFO9d4EWfOARGj/2eIWrHJciJl7L25ijrUJ
S9ZdNz07o/8bQko7lKAOlHvH8lvDyvryzqIGfQ5Q34QubrvxMQDBrpzIqDL5jh5y3GfhFVN54hlJ
GTmlbiWePDM3tAK9wmxZPd2DaiMcJFb4Nv5Sz6TZQvA9vDgMM0AQIXDfjJYT+PjUxFE+cyp6Iv8W
8LwHOkJu8ZrUYFI7CUM47YPWzScKfz6lgvO1h/69zQ/ehiE0BLxBzMCRi0Z5mMB4AXVdNqksXkQ8
u+Vyuglp4shS9cLTtqcP+sjIRMno3I3+x09BFOqC0SZcn6CQF0B7lBbhSLLrk1LfcMVM9TbJagmD
ZvcspBMNiw101/THdsH32UjmHV7wBWcdcJbKm2r5CItRlRQHdTlUl7GtqLb5+wPKTxKF5TujriXq
fvtEls4juJX4eImlhek/KAclx459RkSY9Rw0D+zNg1x804yEB/Awj5P5IwGBcAKhWomIaDB3vEqc
heLZLTeZ7wWbHMUhFqIbZDMPnfz4LA5SqJejoFjX8iAnm3cCXqlAbH+CJ2CU+4XhGcqrzDECXwqG
udNaxSkteG7utLVZ+qHnl0mXEfshVBn0992q2KrV+vtvjOGEeMlQ5dXHiYbRwXHEfuudZ3FlkeJS
c35tGMGnnXyPpOptvZcrzxdV4ezngk7PzqHVB1XRnfMbyVESXwGWTlDcc/cwIplFtxUmKlyvaDI4
MEPb5mfAmaV14k8j4tl4JAl3yKjAf6JTgRAv7Rtl3HbxWYldMhk5/PnR6Shag4/+8aH3MGk4ld8H
q9vQC2GJ6u6yVBEKTkuGfa4qODYOHiB3fXp6iyLfqGZv8r9leVziWH5VSzwGMc1hXugTVReDhLXa
kS0POGPNiXd6eAUuVlsod/s0OJI1yndQ+ezdH2tEvrgNO5aC7A+aY95nVzzLOkMuvyvvWiAj/c/f
cYtngmK/QRHyuhlQnQxbaopUB7w66v63JU6KgiybsnSh/FKNX+onfujv08Ab9Eih0OVLvQkbWJzC
dFQp+6csC1ifLnug/dh9jC+UEqU2IBq9XIvz6kYrJJB/6CBWct65asrbtclX25lxhQrHaqS9AMyW
kzSodBDkWvOUarZVWkzfakHC9WcaeSx/vCXe8oQmLzTHOTVL9spkwUEI8ZbBdN2E2cESMZ5ujIe6
Ds1K4mAGZ0SBZUEweIucAO60owoMnrU9+D+g51YpAmoKvI1+5B9U0CP0oWOtxFnhEf8PpDMPXOhD
1ChrFloXg9e0+Egqtn7tSGpSll94k6ILgRq9kmfee0bM0FBAj4QfImJmV4khF92NYWPS39zqnnZD
+6a4sG7SrFy4sXSbQnEOPb71cBYyXyWJVaFwRfPwww+t+vubYZOI6U5ZingM40PeWUvZYUYmu7lP
JgeCMW9htL/rQghdpaAIAu20zMoJlppyLxjCulKZ5TYzTd58rgqI5vttzESTze8ZqWiTvBSQZC8h
FQ4M8PFG83qYxGdz0DDtiqfNJtif7zxEMdg28M9JVNoX0Bfr5dy9mY28D9z00AkxnbyUQFHehi8V
+eGwz+oyJ58oPv/2Sd0MnRKfvtWvS4tqIogsUz/yRPgKLOv1gwlAc4m5mpB28iNhCjcfS79EUZmz
sfs2RQXuaZ6VB8XnlNz/VCbLhunFLdPvP27PwR13dNWAurAkUm1cImEJl0uUHZh+9AIYuxEoiy9i
ne60zJZNdDSyMr0Q+tLhQVEHCzOVndz2VRwP8R9GENkbMHRvrPNend1PqjcNhHv8Qnnsu9SH64I5
AWEoXYFVaP7x+bz7k0RnDYJw+d2BVJBgIlocCEUYj3KUDJdc+P99YbWRhbeheG1UMHogXLwb3S1y
jllPeUCYpGGi2Ywvv2pLpWS2wKpyYoX1qGCOzpSsVudADh1DG7DCEHKXtL+eY+PfHvLlBd9SPH+v
obPCz4clRD11j9fRYptBSogWk4c9StGoPf3XiHWHQ+wFjN1Gpty2aiuODFqw4SsspToiq2hRwCEi
EWlzB+2ejpcpv+/9BEwDc4TGiAcvhoWshh4QMF1SIk5ouiUzX9zx68bwxYcsR58LwEFHUHaE/Obr
3+5k563Z0qI/EBZS8aTuj0if37CTUyfaSBKSLshir0JRU/y838eDVX0wesPcRkSZKDKdRRlZ72uk
FfLGfAWDFfn1igZuhG9j9TNUK/iLSnqhbimImjAVfprQmqMgpGGzo+GVcuN1VdZ4BjqxQVx3VEMd
WhjIlmW1J0oZ8bOouXEADCAyx9wgB/O6f3HH6Suw5EQbLOzCr303CN4GmsKMvUbUtK4hsZJI5l9B
WbmBdvhY1rUeq5nwdDkaqZ8socZTHVpKYvcHEKlB/JNsxj5aYSgpHbd91h03stGW5fUkMjSHZsKf
T7988XvSTi5JidPm+D0zb187JZAsUWbmoHRtOnnp9aN0HbKnBMLCfWllSYuL7Mo3GVr+OHgWVrb7
BmZfz2wbz2u9PgO7IqlmO3gFM0pP4RVGEkwqQVltfJBV9QH0pLfeMUluCwvikFP85a/Q5sqR4NHj
TUqUXxRqTv0EVviu7CE91OLWCqbqH7ovA4xHkHRS/GXO0z++a/Bh72E/VN+4rg6cDU/Xfe1hRgL1
BJCnDy71oI3ak+jWt5Ig70uQZlCal8gsBlA2Bp1mT3hjXBtmTAm0/LwSkdpsGswFCbdMxlEnE504
uj9KkQotgUM5oAE+P39Bl/8bDeasuO2HutzFWRDgn08VLwBAQ8kYXxw/NMicz8cY1II4To6c6vTe
A6qkJzonEx7B0/REWEBHpoBJyQgEeEH3LBofX8u2Rx2LjTqZ7G6cJSB4uoUYYSas5Tfro+Yl2MTM
1t3eh8zWZexcy3JHJWIdrbM1SNdZsgNSDljNCr7S8bCtF6Jy3b5tXRHWx4WxC83/R5hxaBKRqlY8
sVch6qm+Gvi3nbuLvIlQ3VUmWItVbMNaOqoU97VOZGj+g5hsn6KGdVGzKztbqhEVrGOJRumQTZeF
TbhtxrOP+f4xwfaXEypBDxdqydyNGrk9qxrdCOK32eXIcQEc5+EV+f/QWo3az+LuGKa3IzBkUNV5
2dT122o5EUFCuTKdc2mM08U+XgOiovYfXRawNkGquBRtTZk42HLXl/xMEJ3+D+QFhG5zM5WN9oQk
x7NUzolAYNsAwK1c0DBrfG4dCh8AoCbO95X1t45o0ziyXUXiMmjhwmg01rb6773wzasmOm5Z5nH/
jqaBhebQM2nGmQVHGIyloXmVHPkIOoz/0VxYMWdcV7MGnwL24C+iQIhZMHzb751V+PSIyiYjqvD5
3yjx3je4at/ol8NVxG4PGSYiKsub1/ty/Fr1BasOfyl31bSByG4Md6lanR7MFyTuZpNk4aiLG28k
kmlYhFOHkJD9oCRqrPSn0FLBynhh6XYI5/MRW3Cya/t+aRRj6ADNassqvc8lIKDNJlCWDEgCs5id
10FtwjnaLPQEwE4L5cFHb2MGPweU+7s6p1q78KhxiLzEP35VfqKnYx3BvQn9G1s63br5IF38ogBi
UI0d+L0kISJX43sXu1q82fOwZQHj72ZpueaU0KjsPaxW2uv7dR+ocJZMIgS8oLc9P8k1yO3Z5600
4Sr322o1e1PgFlUOom7zkeZ33uNNHWTMW2Q9+ol3AmJC+0PnfiWUH4marctBrJokC/JGao4CYThR
2a8OikxEcjkavCr/ehT85dCwcRfydDVbnxjEfhOEQLVaxgfOYWS7PRpIh4dAXxhzm2ZZu1lG+7yf
VqdJZJqn+XZERWvmxUygPRhwb4NrfljZV4VF287HHWsQ0JXB4oOxDyMFVxzDZt/wihHY4+yXyLkO
MJBQitS1CpxUWbKTCDTlOjBAwBaAiqbJaB21HySKFvJkMiZnV52L/XqbV447OeWylo9eFL/OfjfN
i+5JMjkGN9eQZtEV0dlo6UOtH1aHOw021eetU1VH4ALX9e/lOKe3s5lyGWtQZXM2z7xj/DTz8YGE
r3WSoiqXFPzClFX0mODjJ+23NLHkGcse+CaYlNqJqZfABY6FAb9Nl7momKuN1vmGNre5eY7fNTjE
rKwdb4SvAKJWXV5G7zMtnT0FEv1QChkzu+icUZVckgkaAcvAcLDQH8iA5ZeSOGvCfz/BNN9OBfpg
y0OuAh++W3rxfRuXGTPYTmPwPCsmiasX/fSwMRlOnvgcunEXh2xHytx11gg9lPlvqOOUmidlLEDp
A3te02bg5eJ3VKYR+SVUPttKEoyjU+a8V5sIJUviiq2W9EaRKvNhmb3wZT7I1sxVE9bQZIkvs9yL
hSAHMbbezptkGynf8irGXx1PdpzeaDac3ljTjGxmzAjRQS0d+6CUv95NqVNjVJkh2N7HYj6+zfwZ
kgIJMO1PUAN5J/KbQ7J2ALi99/32Ki2AJA0rQ4AzzeIWryUXte9EkCoUDy+SsZbBRN6XokCcaOfB
j8moPGb3Ejcseaike9OaHXf56q6/wAnIC3hdDSpSCLDz+7dC6aGjReenNGwJsgt7U2cB6W7SqmMn
Oo0IdGCnktvIByDyDz9a/8giDrDn7LXZ7DM9qRnq4HWxuW0UGhUfcjF1GhaDfnfXpauLuAFAlO9b
tlibR/13S0yyMKE9G0EGxk3wCs3PseLRIyT+/FLv+U/ii829r3z4169Gde+6VPRT9p62qBr2VT5d
geudWgmEwZM+ZCKSw40M9lD4IPFfMmlwSekJzmWLp2swJq0Azj+wrNE3AcPUuvmpSdZlIQtQHy+z
Ytiz/WBxwoC5YSVOeGYNvp3K+znB8+ccgMrjp5kJvQVExW6O6LWaoiakuaMC+Rvrzc3HGBiNiS3S
QWKN2U+MI2rGh9gEVrkBGc7SXU/6hjgILpvqTamTFn81Pbe6QuC2imDGCasxdwR40dIcpgQwyXmB
8kBdc8Pvmk+xkamfcU2f1wsamadNLyqk1wYCj43vj03Tq2h7BcKfBF8dwqgdUcKPjTSzDkUlwvme
EAl8DRrg22MIUvyDCqkmuiWWIy8ng/eYB7KHiZcO8hTolfBGqBA2bR/Cg0QeJYYsuhlyuSHcT+wc
c8bS+igbGG2B5tqon1W12pP1ZDHXhnGa1PZOkbf/L3lWpkWRp/uB9VeesDy0zXFowrTKfJHnUBdw
30W3b7ANIvqN6Rw7+khPQlNIpKENyJT0J25Zgwiwvs0jBza92rSzaMj0/6eaHTGFLvGg+is/iLXh
xthbBtQyCmaIpzZZu+D0cZn+6o24F19ceGtLi3QfD0/S28g6eNNJjHVAJKmD0MwFNoabacdqxkI6
eTvIqxnF12+nefzhivLKXrGLI4da8wOr/LgrmnhgR66NL3F2vSLQz2vg9dxD8dv+VBtIAAADQSRi
FZt+e+FfojJRrAHauSlnt6Elkutt4ZoVbUmoCqay8amQCa0yhNPu6POkOqG8VECSwKiCsSVXO8rd
l3pc5P+vk47XTWay1hXd9QFmTUK1iFyYfVEVMs+iogHHx58px8LP2Qcrwv01qeo3q8Wpc4WhKmAT
YcuMnehh+0/W6Q7/bhfICGsAbmSaJWUqFm966qIHBXIkbYFB/bhOEXGzfP3pKYA3iNwQeoCd6ijT
mZq/nU9Oi2AqPOuB2vAqZ8zHKG76bYxm1IC2rmX4eWl6s31jqrCt51PL6lRPVpTuMen0h2zi8xvm
s2TuWsBKh9vX7RLeMF6F6vHRv8FoPXUmt2iiv+fogUJaejovoE2v/dyJ7vvE7OSj6qMpwllVzJaU
Pmdbbi2u/L/ISRtzNoUG/7MmxMGuQ5SfIXAlPb/isSEhNFfGv1qRWuQG7V5XJU85CQVoWOC/QuR5
GmnEIYl1S2SrCKk3dqygI3zF2j4l9F9FO3/92NFF+thT5VmAY7Zd14bMG4uJi65SINXL0pP3fZ+O
L/aA2c0XrzWAK51s6lYIT8lGdGuAO3peU3BpwfUpE3yDVjTg2oQzB/Asj/TeSR5UEahDUXsUzmSh
3pRXbHUirpVw4XnfWKxwyxcCBOxyFkNO9HKNg7Bp4slL632dYmkU78vlcKTLtBuNVYTBZd6q83z1
/7Mlr8tdXNr43W4AnyNQAMZu+ONGehqGK1QRLPYW4CSKO3iApWYGHixKuFqkyFk9T95Kou+VZU3q
uYxAkC3s3kyD2DDlbDmr1QDeZSxf0pqmszlWYSw9j3FjGEOvhbkqPbmUQCCbNymjJbLiiHRipeut
S3IOVngDL5sILpPOJ49kJKXgIgjOim4zdHKWoXVTa/E/oad/e5rEpBepkKyvMNJCyz3z+FYNG5Oe
ZurIFlPemL/hOIS/1VMB9yMj8b8hy8BGrjHzk4pKjqkJTUFdCx+Ou89T+UvR0sze/Ysh+acd1Jal
tYkqF9r0SdJUiIhrIVquyG9/7gc05VAnf896WXiH7QZxSe7kW46BOjts0rj5mg5D1o24dG4uPyLg
AQiGpuUrkfMpJOsgzwlwJ1fBT5bQkz0U08EYe7Z4uLms5BzabvQ+ZD7rUZ4mLxtRW5wOC3hD7RD7
YhtMxyNvtooeWi1DXyf5OVYyqtbsR1AXeXIq/PicxeJ1Ls2keqG4sU702+CQbjJz4bcgCN612y27
2d7tnpTzlJI7oeojNQAES7krstk+csJITZIw1Xo8BzlMPYW01dQ5BfG6cGeoJXYClmIYeA8jPlAZ
5QE2D/PWTOkDEx8lW6J4mYgQgGFbyPmzjsYBbKydV53YLsbuB89ZL8uxPNO87L8J/UnghvT9YmVI
/HYff0cc0ASBTybbT2mLnxFAOfuAS9bsSw7oYnJaEWrZ6i+zXYLJsau+Tf3pWVJQF+HqRiFwdpwy
jjR0UYZ0aefgi+HeTm3/AE6Trqg4EFnkt/P9bCU+VOx8fIp8N4y4IevqwPm1RNYO1Mzc8MckCY0A
aiGkoeKNVTDwTB2njpDb1h3N799vSDluEBrZlaieTX+zumQ59JgWvy+hQX7XKgdE+a6fRDC7C1KR
OY8QtlIqBvBETqqhI5oWXjR8UzN1N/vnaR3B8EQmVsGiIymIzOgMtPxef818X3lgBIv8n4qppwIt
bmclttkH6oSE8ECd8XKjk5BcN6g36zzVHY3QmNq4Mm6/P/En3C7dZIcFc2xA9m901923ANj10Zgo
51CJ9pWneh5caCo0gdLeVZZ/a1oGEnxYpABda6S98Innh3xfEfOuEPtAi3y9Bm+DjPQ6grJYILCT
mC/76WsJpM1iXNNhO/gmv3jgdIwefQI5rUFWrgyw4/QWREQfFkQ70x9ClH8icTADOxTbi+9rt3Od
dKDbQjqOYJ0F0VDyEi4sHsmfNK4hNakDn8UCWdAWOlWVzL69mFt1xYvk2O6bhn5gLR3tx1iJ5MnO
Iu9v5pOLKFL/XNoUVYUIyEFIfSGaEDBW3JKuorJWUZ3lQ/Jta6bbmYY8wse0/IQIzQ8d2wsX1jRA
SMwHSpU6w8X1iv6ksLn6Sn/MmgoSOeean7mUb7m5rnGIa/njWYU1y0CKvmSkMYwps2ad4OCnxIZx
aY2nLqPYGW1vzNFDFG0BlLjY9wuHTyMd6gH7MY5guEoaoSHQ37mj64P2P9XyHsgjvHSG9+MnpHtu
d4g8bwEPilX3wssee9U0z5S/cJVpkB+HBRQvQRN0cwKcB94SJhKp0twAGpXrAmzjM5xmYjmQCw0S
3XLyjgB9AIpV12sBqZjm1PlXbZQ4XKioOPheQejrap1lneQ6uA5Ds3bWjL4dhJfFMWYd/wsXWPWd
eb5OPYFbyuEGU577EKEMsiYqWmSZklF20Lq0L39ThSp/Kld/hl0IALjqP50z9pN6YSrJkRmhW0cV
7qt3m3JgIOxON9t7mCukrUHJyOIzDKGDy6PaPyP59HKTSZkMpkAQyQQjZoPNqq432QAid6M6C+Fx
bjgMfDMzRiU2JawnLIGRlY8dCXO7lixCYqgVzOz8jY66/GC80hJ/SY0EdGLKAZgF8SSwzBdvgaoI
Y7xupuBGXVucuTVYy03G3WshbvDrNf3hOs+AMdaqPz/vwmosCbuLdFvJNh65dYAH0/V07GRoM1CY
9AV6xSgORRENbtMSZI21Z/PRZRY9LZnNn0AoQPxV4lnmeIPjN7sRMjU4PzxEM6sHvQVHtgvtU021
i3bGOKtqq2YDvEnnrTAOvKOfhV5VSsICmcyV9FUJnDAI1YbMtIQIvq3Fw4Moy7msjg/se+U5vgIb
AX8FPYYEYJkk+6DtDBifJpUTxdNhWDVA6i0XYO/Y4KeAfHXaOQtR8oFMHBzz6w+kiRXQadwMRP8E
VsUMQY+Txv7mTTS/mjvW7i27tKX23ZHf72X2hR9hcMTQmToZkR1DYRZrnpVnY/YO0ehatKPlXmOD
VV4gIEOUqZSuMRlCGXj9XgKt/TyBcHEuXYDqjKGzvm+HyGwqHLDH8+FYsrSrnGuVzGbpcytj/0Mj
/ZrqQY0oKJxd/++n0vHAIb/+kxxfeZw9KcQfjBWRnVmmZX+Mt2DTNl6vP2HC8/wBW2agRB9FtjBx
/kt7jle+u4UjjKNx/tpHMsYCch9jpeYW7pjAs+DMKmUnsS2Y6TST9mlxjuszHbfsfAgzj2gSmW/L
R8Pas44uUSF8gaq8XvtnzOIiJLC4pjmn7iGewPaFhuwIkXeOZTH8rnNtTKun9ZDZSKmZEzz1B0k6
Q1RYqpD3hp+wdlfEJ3uBLNr1j4rh60qDozinWbEDNMZ5oC26HZkX7wzGR4aHUKnGEK70duOh4C5e
kM7Tq7vbQUOI6Ljhq0twqcidMAfybZtEs3GerIaFSUZDGvaU2CckfzkTssRfXqe5kZezO2iDLoah
7x6iK7Zr7EwCyrKtMWXU1+mmDdfAojpx+R1A8xzeL72Eufvk4yWF9FKTiQKpKDQcWPGcvq19EpUg
vfT0J4/X0vMhtQpdtRR0sB2/Ct4a5nMFdfLy0Wyv83SK8OwTu6WjjRfbC61anwAdeKEHBU6G8Qnz
Vbp/tg29zbldXSKUfZQ1quCEuhTT77Bad/x6NVVNLazDkbvRMjBrwFmq6Ex7IutXAXyIdUVSJRNN
qbvYROVhd6D2oWTi56OzXuNSS66oBlkE2wWy3x9/H4Nbexkqu/h4kHqnufa65+oaxKqJkaJFlil1
Du/bER7kMHOk7wtZHc97UXpA8SDquFj+BvtgVBfWkSottX9WnxhaxaRKJmYBGplvEGGf4lGGoVmC
oLZOqmxq4BMcj4NtQzYgWNBeQYrsgGq0ZMA5fVGwUVe5Qic8/7uJ4q9aBdq3FYVhsnXJi0B7vnAw
gYDYPnTnfLbKq5z81WT8tYXVTWUG7a9Qx3z3S9+1aj8zQjn6HXOwHo2x5qkgPkYCXBOal+sh9Ll1
sF5FnkWoFwbnzIVSxonN1hNSQn33PjO6Bz1KZDkIEkUKrrtMfBUBowZgPQGFzvNgghIefIoUAlvY
SPR5vI699y5zvZk9vNPbfzGBYHxKClHtpccVQSFTfWuu8MPAhSluFkKWJpU3KtwvShld/fHHDCXr
NR4x9qgw5AUyV+4xZQEtXeO0jsCLL8QIoGYGO3GPgaQ3bLaznecewkRgQ0oDjjAHh23oR7aJcl9o
ACA/i9LiDIZDqMcgSNoBj+y1rsWzQMM4QikETCUjHfUBN9lvvUL0TxL4Ur3e4HYwvcO5/KaIrpsg
67mgqwhWdp/iYo0SnN+5ARIACmXgkOMQi+GX3/LHr0k/qWZFo/rFPavhNum8zmx48Z3p6y2sZ/l0
hXzYyY7/B3zeoG1p9NRIGDc5KSBDMDFgyOHDY3LnpZAp53sKvi08K1jI+Cbk4I9sUi2qxiWBBssH
GKDLzL/NWB06LYWvN5korZRz7QqRssBYlTgVpTYe1Oksa50peHqVPpDwB1gtTmjejv+f7VDjSCFP
xccPMuY2spugh0qaZFUJkXhuMih+FXz/l3d/WLZ6qwIHpQAvojn0If+rY2cBEJsYyihjH5iV24LG
DriXLLN/nb1wpB08sq4FhiJ6Dz5YcQUjlxkps13Cx1+Z8vHrGieWX9ha/GFsMQop9bOLXY63XG3A
1R0p0RpMbmmLmvw+J076kJB94rb1bZXvhH9ttppX0n308JJQBouCwRumRkycOPNbFzCrLlO/hckT
nqU9XD0AyyPSy7h//qM2CBodoRvDV5Wq6zHTb7A9/Kp2QVblUmIlHJzalFfzw6ZC79YwIBXe80lb
KmFHNkRKAAjJ4xc7jcuKkBEzY/s2E5ekNFp19df0wAIqK1dfi+IiKsmIr3oXKafHvUe4o7TvANYW
ekQ1iYsNB8C3BpsMxFlr1Y97HFEP29h/kppDoeItivZsThZ4+bL4tf0z9h1Vu6MxIDc3Kvw+D+f9
fgplKpPvAeckPA3CQDKAQLgsmJyNJRsu5s9SxiTQ/nb7hZ3BKjZpce4s7jMLOburolO8JF24YfFg
XtCZN2wYiUHNXuVVsTUjiady8BP59sr8iIlWa3d+ZQg7tgFZVns0W6+4ECgOV0r0HcuSA1rwRWqI
Y8zq80f80rwBTjgZCP64hYnJyeVEyZ4FwFrQUZ+k9Ss6yAPKSRu2t5ts8q/L0W2U9CM0QGXRR1GR
zW7xGrSFJW3hTlxJYeZGOdnYaXVrxglucnjsBEOeKYDsYAUrMs6q80GX7eVbHPqRJUciyazkyN7C
vXArWbTmcy0QXBym8vJYiLtdQmtCtJy8P6/QUJ/BWqnE3Nx2oYaQp0eZQQfQjxqEGjrfP9MtnSdH
jdH6jT9EYt6pX54YDmu1AE//6BdIAaLy2NmMejQNA/H6cQh0hDRYKMSxRS5CtD0CPv9IuBHRjMVb
3sRngV89KM1fOkoH4CnfCBy2h6767XLJFo0lypPCsmpc/8DZ/YUten0lm6RaOJ5ouZ5LArh22Q96
+WXd1jg8rOfc0Zb3wUjG2x0DjbOZOfUKa9SaLOFChR5TD3sbA6flDZP1/lzsTKS183YjC8z3oSSO
5Y09aiIhfXng+zQt6bD1zvUSerUTvysRPva91RomXe+poYhTHwFrXDrhXtC24Pmt7Xh17Ir8kVNU
2xe6GywX2lQ6SWCZRrTmffQckgVjYXAOctqC8Rxg+xXYFmT4C1lvryKUpGjXPoWTPp7UOmTg0xlR
2k8qYZ1YYowParGYJxNNogwKL6cvM7hsnvqqOpkpRkD1M7rQ47ZyjcfcVmWm4RiEug3cUyrYOYLQ
O3CzHDyElQw78FidKkjl/XZiSkQ0R9xo5qTgpQu44VIglyeNPESiUBL/DWdXDlPt2L9QBJQYap0i
FJ8cEWJD9/i6sNvxaK0fMiP0wHc+JKtlqEGXgm3SNaKEhZJdVyqTqQvGftQhTkAGyVBkXfRX4wmZ
JPJdrAOxP4TazyWFt8+DUZFnAvFz/UQ4gGWBC+LcEmQ+I2bLBXYwouGE2l/XtthhITgg0hh27+jv
Uc0EJ53VUVgteyzMOwwe1nNevObP82DUFCTmGAyMjdb+3eya84JRFd38V/rRZ31OhiJvAD8M7tKB
jCJ8zF85UBmQULT4xTOrSQ9++/zTH3Kn3wCOf5ZcLpQrZJA5iRMFmWekSGxbu4YIalfQIFnRUd+T
XFw8hbKouJ7qappGe5hPby2qnGQpVQ48Id3FE77TsDbEi/ZjPj1e5Qgm/3Bx6+qyq6tmif/LdMVo
ZefNCErumvuEpGY74OrFOBCHFyfhSxWTw1xa9tErVuZe8G6u1hhqrN6hT+xyRFEF9f9SEqcroGIl
aBEA2LuQNtEHKvB5wdGbSmimBSd08X0ErA23F8wTRkC96UIWbAIjmys8vamGoRiNENwk34Vn5tyf
PNfGxqH+iSpujDFrR/6CONXQiD+0aDsCwXjl5LAMJ8gG46hVm2QkOoNHKXEKVhTsNSqO+xf5wBdX
XOU6PKLIZ+1JL70qBSBu6lC4TPGghl1W28Dzjr7PxEKJB9H0W/T3PcjBptFqDMuq9nvLfjd3jaOe
RDWuy1iThWuMtsg7t8rOuo8deR1Ch3dEbCZ7KWh5IA68rTE0YiBvc21BdQiNTq5xe2crF5XeDU4C
lQmMWLYqum0y2FJEH8/BEpk0ElNFNI6HW4E2wzRD/UHxEWyGkYksdLZjnvEVx2MwlkQwiw+aaTK9
qw7LD9haQJaTMMKWwbG4g6WWTGO0zSOQqu4leauJrR/fclP/K853+EuiZD3XgZHV31aeHr/8ciR4
aCV6GvxrPDCHVTUalGOd+a5e8590rR2qe/ypl7Xo9xFFgVQwZUDjR2hAo/MKTBW5wxBoGx2UweRr
3+Dbh9C0DJbXw6s9GObp1mJzluUjK4mfs+LAXTuQVK/jOWmePlwkkHJeELoJFdNZlREBSWAveF+U
FHrOFLMkjNbkkzesUHLzLgb5WNMOOyefG6QjCTfU9HlKVlVLAXKwM2hYiNrFe0AkepJAEpJfdfEl
nMyfdX+x2P3MNjrWUwOy4K2HzY38YPMKIhLINFXgHjPkuj/sg5T4waZR48+RHXqHapn/Yhy38U7q
G46Tt5A9Nsc26+B6VH/ZRriMtvPnPaV213L88fyvgq+5J/+0U1L1/jFlcwyb9Fpbc9zP9QWM1bKT
i7mdCdyZE8HAlsP4NdVblI68xIBHyGKuIg/iRL06pE4W87671GP7v+NLZLPvJVXFNxqapXqA9J5t
KSNnGtAUL7pce20m9PU8yNO98c0+tq3ZjxS4r7LMhb2ny3bxi90mf7spMR3UfLUAHfkAIJJzr724
sFX3rjeb+U8yXvPXdfS4u4sJ+TjImfTs7Nxoa0e0F2dRj94ZDTRkSrNDb/htODP8JhkI/acXfkW/
SXnosnUzWQKV2Gue3Q+WVn8NkLDWPr2Mlj6IOs1F7++s0XW58N5Y7PxYRmE2avA7F1nnHI7LcvhB
atRdrlcEIKXqcpb9HRV9AkLJEp1t8m8MjbVvLzkCcE0uIZe2BUCZMp0GKyGtZoKC/5+fGfmQBKV6
ZxyVOvsHjOXk/0RDRpfwS0OFYnyLLrO/m/yd47aq/Zjzlcvhqk7aQrSzfwd9Gx3YilfbstpMPIHL
o68xiqanh1T5ASJR+h1YaJoUhbduarwSU50WTOb+BmNOjkF4yZE4fCCkvgRcuO/VjE952LcirKoP
+Up8QWE5QgS4Yd/L/8QEIGZNYcQ/mpvpIwj+KkO5VUm2Iv/5bszkCbfdP3iKaKXjAB0ShIDTvDqz
SjYnMrAI0DoNWsyb71/zxlbvS247KUjBxRcYmuxw9I5nyO/L3d1epPYAi0YAlU+0xk1pdf2ujjnx
eq1Usat7Vo5dmifVjC0gWrNo5ijB2yoYlr068TAwpdiFrzSfDM2NAaupvmqnMQ7en0dpWqkEwj6h
ieXjRRzoogGGTxMCeDTbqVACWldv3LDAxOXEf650fLYEOOCrIiVthGgTIJpWztlshHzx3nhR5z/5
vc+s7709JwHRypuom5MtBBshrJ6L1RdQsVfJfTBTYkVoyruYV5UlyOdNqNJ/JrseAKve+YBalAR5
A1UDsHvulo4+5iG3ZuUv/LDkuzHqyYoFl28DB4iCcHeKjx6dLY12sM7l5pxjBFPNYG9KT7dMUAnY
FaQk/L7XhIuQCIrbdatk8eR4BxkGS6oa8x6RdT3BEq64o0A2bj58e93A03Npx6wsk9ex7sxUTRG6
4KnQe6lJjV5wX9itFBGNrgSf5DGNLgrGw2C/WtH+y3Lz37PMwX7s9BLh40miaRp9lpEeIeuBRY0u
fc/uyzCbNnKJ5/V/bmbIgN2P6Dop6tYeGdtaRIC/OF0/yccl0Jp4qHKQGR0R7LOMHHh/l8yeAeVd
znlhECnCWMNN9x/yE4IUf9o55zVzSCTH32I3fAod/6DviNVGuqa6C/RLgWK9pXyEZcSGlv2R9Zof
GfWDzNlOrrYviRiYMJhFY8cFTHPwhJI5pryfvOaAj8zQyHHsXlqJU3Fi/i6l5L0zSP8pdjomu69V
Jc4AL5v82Cw/XB+IRoUuWhXoLDy+oF4ENhXF1WLrs49P8Ywjal9sHNwvZjf9Utmtx45UxNlqvt0k
DtaY/QMdLTHgVX7FKU2xTHHA/wJ9iyWrzOgdAxT/dHldLA2K82RedOM3jCiTyhUtAOEC2j+ddycw
uwwXearcIvDSmrq1Ep7eIVfaigiuLKvG/VRbPQbQYEGUI6Ef8+00aUuVbuyVZgTpz6tEDoQKdrjV
MDMALrdFiQBoAnZ+9tVH8SMJ35rtTNWzNq1wMcj4u7gkYKjI0ShaVf5uAdObbHulbBngw/0x0LTx
8Ps7RHI4c5PSpoX51b0xHOgUN1T21kgQ/L5MF6LoF0YC8Pfdhat+SHINhWD9MmQ3tkkIzZC9Qb06
SEUziQgLf1v2GGhc5BlszaY9fIub8S6maS+CPx00w4QqKACMnTp7b+3yKXcrUE1fVscvA3eFO0VP
lYi19wTovxv+6SGWhNkat2WbI/Zlh2DZ2oG5byv30EMNzYTE3JEv4rFfMKXDWzJm1xhCcI+SU2ZI
nTRD+lQCQr6k0XPjc88O10N1D0eVKC3T5Wu6GqfsXl++1NHLxFBjd92esRODjAsMXBe+UKIAv3Cu
km9KrC+nisfnT16CJCZJWOHtItlH8HaApQEIYUNIWzHuAs/pJMr107HZcPYZHifqz+nThGgNe1w1
jwIwcwz5kGKgIt10fXPBYiX5kVozli/021bzgqzfl1bHV62BJQZB5WA00Ppgk4zfYnZZomzCGvMN
BGc/x6lZ/qDeKuLSZ+ik3V32WoqDU3id8RcyLqQqQFdRlHxyN86HiWFSoWCweQGTxtEteKku9g4F
6lBTg5uxpwAr7eSDlFhmGy54DLJpmsHkm20/JKj5ogBY0rW8kHThgiRP75F1PHox62E4rgPDsQDh
wcPUVmLC06L5SPtPNjV03TBvHoyF7HGu6OXjYVtKFZnMvgU8a4fL2fgph/IO+ysTH5P7bRgWwnmY
ahRjA1TLppXrj25jd2EoIiz3Depm9lOoCIPTf13WsR4tK+Yaej6wIZWMQo6ErzX4EeJ2xPxI9d5a
bu1YCCQKVfhl+Fl0n8SJ9XpSbR3dKn2bUml0bV8u+j2ga0gOCLd3gH4v04ggDQ7nB05iH2u/PywS
st2Y1sZutqER7bp5AZKtzqEQrc2whi5aBrfaG9QtXDvNNs95U3fo+WiIFUJDXyBFeU8MibMYEZ4t
WI5jwcQcYPNOb32IWD+0YCfHQoKMgBz8TMUXlRq1URtZOagEkNvXQO9RLQM7Qaot/lshtjLsgmUd
ZcQFyHFjo1q/K1BDtI6bIFYtdZUPujiv9tuCz9QXEBaUW957ch2ApIrrAEd8T0b9h6VIGjW/9FEy
IZc96nveUbZrFtoh7GJo/yxcncMUZzxNi0nGBK18hn5SiRNFyMxPLuqyLqj8KFe5TKuBK/bgwDoU
N9x/Bti3luU7soIIEMsbZ7hax7wBou0RLoWCmsJ3fRmqTjDkxrQEirTAmn0WZlff63Wh+7rBOM6a
2rXCRG3N79zOLwodzNcWcUI1+h7z0F83vqXbO20W2qlnIazBqKuQBrd+bh6HYfg9fE5oHSZaWw3N
DkKEqnGsTquCi1qvHohbupyoNu/FEGxEqeESw7JGRYQDaOg+5kunQ/+aJ48uodO23UJMSsNXkH6Z
j4ZeL8iXCe6l9Xr1KTNFIgEjG6kPxGeY+6H/KkWi4I0UyojVALgZvwPg3Jdg7XjOe8LTBbgAV24W
zCN1m5bX0dYmJwNah8GE2fWxBavkmAOrCyOSWoMY82oZTq0Z/p7v946cK1CbWpXoB3Wm1aHsqOzD
ZF7IJ6W89jD69h2h7xzWCseMwpAu0cbdjdlWa+0x+NQrrdJEVEr79KMjNZ349VQKMKdNhZajSvFI
Wps44vLOCBEbLnFQKR/T+Hp4usmpHQe0rY7S5yzr7f95D0CsABjnUtHpKMixRBG0pHQKGqOLSSnk
XcDra32uE4FN3TpHIYfpaNplgOxGVwH+HKUczNH9UdWsaRdd7Iiotr7NKVAWGl9Dv7pt4YGXfPut
yF4r0wpFEFkDO4QHJlpYCeZhz/Y6qh1M0g6k3/GG71AmvQkUCg1f8z9eobWAEZkb7QpYvfLrGyk+
4MHPfWOnhGcysTtZYRPvSJiUPZSP+sQo78/ErMzOX/mg+XBLNfZaQkXO0/Fo9Qcd1qy9nTwVBcx/
ykpr7aVVKWloU8ISkhP5kmPp+P2o03kplviV/X78NW3TL4UlEuZn2aa/V56KVBI7+7uJ4ogLOIbJ
W+DybL7i4uEct3K+dRYAHthRGgULcB3+JmDUwv+EoXUqqN1WPo2gu55O76/jaJmY1IaPvd/1xTaP
WViu2fkUiAoQnLrQ3AfTUvrQlheCVKYA5asUgXoZKN0T396rE58L9cinU3RfuycC4iju/kegL7cB
kfFWBAOBaVU6rZ2HvsZIXqn9+WiKqcNq2eGvSk2sHlobwnANqW/rRQ5T3NBZTBJ/drnMh7Cne26H
WMfHhGGN6UX64SlPeDst34FvAy0r7Z5LiyTiUPs1hGkZYoMGfxF0C/HLhwj1mdnD5L/o0t8d2K3j
Yc4gTc2hlDR++uSr5X65Dyzi8nbLcclwdHg5rGDbBUp4roLFFL8mrIPqXi8M2L7WCALz1Rd2hS9B
34H6NeO6scsRjgUR3CKSa6DZm3dhV/wkWi++joxv3NtfEcllN1qAAhhmRoh8ry2ImQCXbSnMMHYC
hlAOGoK0kaFQphEg1EGO2av/pv0qdYdVrY0OAIJ6yTF57cTZOUk26LH4Nm5rgefnLH3gAN9cGA7Q
xCKlGjwKWYCh8UbmUXPXM9ro89eTsfmR48/ePtcJwuXiNexskJp2SdA164uwCBfFWm0PIGBvuoR1
VXHHfjZu/gxga4unqlDIAeUwy22E800x4a088x/wRrtbHZ9rYyk9TeqPPlglx3Yj1GN0hxFbU/rJ
ehIj23nlTiPdrOhroul2dF9eaQYsbL0TRHFvkcB8qHERxfW4ItZTEpnty9TzvhgzkJwgbrGUJ7TY
8riSaIEd758Qgl7Ao++OCND9RobgyWFMLQ0HJ/A96sOmDFswcE5qryNzWeJRf7TVd2Ldk4CjrIBh
O/K9dan28K58DbizsMt9cQGyT/Y7q+3NR1GK5q5gQK+imkZ+2z2FLcoWNu0PxcAZJsjFvEsgsMdw
w13GNoNdbUAYGuyEjxyBx7ZYeBq7o64/Vbois1TxNoIlyByDphI0lRhdXuYrbZduZaYDgOrw5chL
kAITqrN5+dzJ8rXl5coMVVZWg+lQ2MKUJbleB5DwfuGffSKbZQfmvHDuUIe+rCrDG8QDnMEH6pph
5C1gargX6iWkHYrrSS7onfU4nsXuR66ZW6GZ6uVqqTyo2XKG9+8ZOVBFOKNKjWTg7aQwvZMtfgO6
XyY+rsTq/edGj95tgT3ZVQ3RmoUSqhhRJF55f3/Fyg+aL01VLcQAvGFcWUb5qmhBkIjtnB/MEiz2
DlyM1M8jChDQvUqc5466xrxcuKTVksZXIv6fbNHv3BA8VCur52mrIiNzbQbL1IbPDbat+EU3D5EI
OcpwMuL9ffJjGYYHilfsCcoe68AFkw3Ar18CEkEToCyWqkokon+fUTV//wsfOUXqrEWAf1TDi9wV
RJ1Un3r7XfohzudO4xiv7AVt5toIBMNSYW7auzP15yfmwIfvCIPMghXbZZHUt9I2ZpyL8CkByRMT
0XWWIwPpql01PAzkGKog9rQNbrWfpBWTXCzcEpQ9sM0DSc81MyQP/5gem8w7uDb6GV/+2nJRmd1/
/jw4A0pKev/7NfYhIvJQBysrXUh74pXReqqcDqdUGFV+8ea3PCFcoczNBPtmnBW6AUrKL5TXTdlb
9P/NEri4umDwwMxT8fXpLhXbqUM642SU8IdoiTUVDl/STR5nkNkqD6IrWSr/gk/bMMW64t/2QAfY
XPSwb1HhdeklFHuYeJwb8SUNKQLkT/3KuEFkTCeZq/aIDRsybC7bPIYZqzOMAoKSasAVnraPiyUD
zzx9pe/iFnWRwhUJmqy4sFRDykxWUTQ69deU8QHaT+I5n05mtFwEPSLEYH/MtasGybQvycfDdqYK
qzlzvWMW1kvFXAw1S8sp034XobdRpV9PlC7AWiwtY6JjIeTTqbEdE4odEH/i/XSEA9M/2EJglHhI
XMf5nzL+sY6Hjq7qfDtYu3FR0Xc8CF+54w4CVPlSmZGjn+1ht1iX67gnmxzxrI+Hr4EtitNz038s
GBg92idIS+SrFfKcMlU62DCNywWPHcjVkSu9fEiVkoHKT9jiguHFOTMu4YOSWSGQwS5S/8Pr8GIm
USEucINMVa0DQ4fFJ9n150mpoej68vxKh2qyhOjbzFW15+mxmZ6KoE/m7lmX+LtZox8HUI899hyf
wSrgdxfOXK7YkeA3rOskDjImp8ryrKVTxhXA6Nkadvr4458xQBVpdRkDXWsnTh7MbOsMttqHezu1
LVnix9JKMYa9+h7QB8ZONmuMRw1Yo2ln1oAOC6tipJ1wNag8AzML9Tp/jZmqzKXx9bygRwS8P0HX
flVlX1FjsVzU8ZTAs8yX3V+gBk9zlEtD7xkEqLL5vjsyE82TxIvlVigepo7BaDWHyLt9yIH5oVad
dxP+h1wZVdwhdV5+3VBy7vQKLe4t2tcN91PnslHpx+fH+ackrMW4EzhK5QpbkLp0jkg3CW6RyFWp
9Dl9eQz7rbvN9AKyi4iqWcHEMnK1VAJvNJ8/qX+5MFM6OI4Al+cCa/1G6QzIzAB3kg+jrKrUZq1x
W0N52L7y+YVu4Uxr2xaeQuxJ68FPmJlls4K/9fMY3LBa2aUOhOH/7kKqqG4NNAkU4FqyrzNlEOVR
3D2HYmFvElCZbwwAExB4nnvME1USfcQYtBE69z/84TWgRar+lpUqUsZQXGE30OWeRpHywXFBZMvZ
3oYsu4M0vApD6YbLDYoERN7tF5qhxlpNkWsNsh3hEQZ8CQ5PNbbfR5HIMnT7w6DD7qa/9EkPU94m
l4CKYHWGTihV97UVz9CAQOIdqT7es+lJRxgYDsFMziljB8SySlkSatEnfWJbpThjoOqfXfLFELqp
KUUDJGQBC1XZ8lhoglk+D+RUnTErLC4p1XtSltYczDDkvUNAhHyrqO4sGTWXubmewBg6MvJvQOsO
AJgXZGtHATwkfJ+GIDb/IZRkYAmqYjybi42i9MC4alBSVeP6gtSvWrlusncO3kSl48yyMo1nxhGX
fUwFrQa1Q8mH/TOzb6OjViRiCvShYKtGFTkjXa+GmOVUvsoRzuO6zRPm4Dv5n62Oy97tTYDniG/2
v3HROb9vtlGWgucA1ily7++ImQuYh9tDRXYi88E9xIHVm9Kl8b/QcxeYBw1D1154YY0YcTjNVKWf
jttiMMA3cbO8WAgo+vXEvdEJ3pidR/hLfL0KU/kitXZVlwMkAxNjZfKpgU4fHHufl4rQIqCOpGfl
NG088Gh/fY0l0SMUWyde9jrauIkth4tnUMKRPdRxnFVg7OVh3MM7P3dCmQfXO+I6wNIdfGKCh9oO
E5+1u3ESQgVyc8DJXAxr61N4M+qO14qrhWwXnff+5ZQdYjHoiuh/fk/X0/q8C6hsu1nDtnaTLkoX
fi1nEfkGEGspNTLrXnZvV6kKBgabQOVhAaIGCoif3liu9eEqMcSrpelskm/jRCfZErQh7XjXgYEp
qC3BRSrTTPBElz5Z1iVfYYt/Mi1IkTBiSJ7qu7TXUDMk9XDj7OR5zcl7q5mnB0LNc0zXtSo7hrnp
k97AobxodR1RazyJrNiBT8IJPHM3inXE38DS/xh/RFtH9lX2LohwgvX3F7i+riCRMnyp2tR/zP26
sd/CTOuQd3iXwCijcBHh8tiTRxXjdrMOWNwvLMinjhdkXoJjdhi6z9hfPhfED3MwHNh3BCs6SM+n
OaYZWxx3T0sh5l8nHWmeg4XdobuIIVdcIdkzgi2q+mDqvcu2pSJj6l49r0VkU2EAmy0XPp5SfyWB
ThrYQ5cVvpcqC1nmQ4lkZpK1vTFAjwaLFUXYhd5P0CRc3wcZCjAqC8HlZC851DdRKorRt+/9Z3Re
P81EdeU16aGdkmMN+RqcLc0RXHdxEvqz9GpKMVcHj53Sbq3o4kJ7gziFrLuDKDBiLpHSar+K/Lm+
aCDBww6qY3m17mXJet3aKhIc+v+JtYG59sKJystDfVDX53KjeXXzDHhxTv3hD8fcexlhNLBsHXm3
aw55L6P2fQPhU6nH9QnHylOPOz0FU+KWYp18FbLRmQxBcFM66uGhaBdFjztZpGDU9mBRxJaHKZZU
FE6frDDv6Cr8pgtf34rvf6nziAa93MxNsqHBomaNNCNSWJHesC11/ObTs1U9yh61N+afC4wFyj36
YKaJH6FpFayegibz+YMvv+ruJCnBHiDcAs3zfNjF2ohvlksloBPlhHdNe8tgT28Fr1Xw+uQ2KHGS
94BzRc2xbUxV44EiMQHDRFommrrIMgx4TiM1YyWD55jUjyas282Lw89LWY2cK2cIYL8zlhGxn54B
DT9I19Hz5CEUur/nmP9budHybo4tOw3GiFM3gcTX0yx5SppZMi6zSVNr574dhB9R1z7Ka4JT1v8j
BozSG5HIXF8WXqrKT7UB7582+7F7sf5tqD1dQ8boocBOkMYhm7FVg3UuVxRHbDVmFu2NAd7dRvpZ
L/OogBO3W5tfQlOTcJ0pgz7CGmq1x8/9XQecu41eku6eBQTkdjeODV6zRWg5B5dq8lk1AaJNL4rc
rhuTzD8WYvtsWualaBtM6imnRuAKALABWo2VSIV9QbfKXjnES9FgGepPW5LHm+9Egqp1MUwjkH4w
Ws2desQlnQfLbXMoDOP/mqR7xSXtvi+VllyCwIBQSPRUP+koacXqzuvCivvzg6IneNTPyBPqFCRg
tu9xpBJ10YCuPZye7YGLiyvEbHAgI0T3DChb9Ry85kyzYTmqbTtkpHKlpAr3jPzpdXLg5Pe9bZxc
0RW0CnAhSn8uM9+B2QrDAjyz3CIDyC2S6QtGOHTVFpPRxLFRzLaSs1fBQOHMQi12DfJr7SwxX+Tz
ivwl4SvUI0jaDhUuozJqVeI21OeFFJvzpJgfUxkWjPuZm0U78SlYxWwotRPJgA9VcMXuC71Ra6Zt
4BbCVhBqB9TvTgZlz69EGPGNTcQf8pI8bo/8gFt2PrG9HbOYIdap4bRamn2yvDTo1CMGZ8bFF3zK
SdWtQlmICMUcjsMp+FNldiS+K/nCEyndiE+KQE7UDMch0RT7EYhH5CEilxL2qGMR0Jjurt2pAA1I
eKPCM3FE45OpJ/Rjmnw1s2jVYYk3KIHu5lU2UQRYSYYs9ANHzpnuhfMFkUHWFZcRcVbo7iqxvzoy
sqCbEwsH5OpEJZH+lWT3dxKxjNqpJbpVKAN2tZMhhCsAX4Im0laEh6CCm871zCn7lOe68GJioDsg
64TDMkGBglqjd9mAIJ3gldn48rOfHWvMavxHYrQOx1jhZTBZMHbLFmKvwH5mL7f4Cluir/iFVgcK
iZ0hfZs0WonjvkTmY0cFiyN9IW8W/94iMRopXIYI6sWLfrVAssRnRMldGg+mS4ywQRivGXmmvUQ8
T0SmBEKFzlirkD8dqFIV9deryP2WI4Iig6h+80d2qiwJbFLThfJSNlwEB23HdaMjWhwWxgbpsfvz
+If9MrE1PSrALzEWZDR/A8cMhqL0AjpYkh1Gkbsm1FiwE0/MKSbcbGQAa9sOLaH4ubH1evIQEB0H
Ntwbpxps+h74rHJyD8VCDbgp0KkXb0b9iF4doR1F3O1wNc8E/TSnRDfoszrMXJ9nDyiPhQmZzUNV
BUeSzJY2D1W0S4Act+vDow3weOj5onyA7n1wbEkR3YzkuseUYMdbSwyW9S8V5QTvmWBFwOOgkwwA
WRvbvovzl790gLJQDyg0CXvalFaRAbZ3udqQA8vsI0H8aRD3gzAhnUfJuR3r+LPkl9IBS8CZNYzI
hwCp+GKFv2C1lSj5Hk9BRUjLvqwAxJl/fMN1vep9WCSNwBU0Xr7cQ4oU9nklBvadmfwN8nyvfVYQ
z3cpszKA69kCt2S+52Y7wsmhBnDWDh3+Es/BF5Z2IZs6PYllWBlc8X+CR103cMDFKKFhHuU91YBH
SnroQ8gAWao1hMjKAvR2EKUOHmOtCxFrGRSfm/STq9jYx5tmuimU3ger8BdeQNHiDsKKyNmONfUN
RNb24XdjTW/6Q0Z2z0ADgHIMjU9txqJm/2Ygbaesi5VNaXNE8YV/2HmjIjGV3XXqU4SFdGDHfzL+
0diHv2BehbUL5zXQr1ps0kDekSwqLV2OymlbtW4F485inTgtprf/HyDQPOF8x0Dv55Cj6Or2WDLi
XRWS/0a+PxMCTPZKY4pPmrF+LS7t9rdBHlmHja3D0YRK4zflkw12yB2T3WgzaDxFpah0XHB+FF9d
hEE4G7G0WJz3KZtyCxS2bEOj8hYFKOK2bwc2aq+TJmHN1UHXgRhH7M3MGCOc0qawtb6V/qnvY2xK
QZ7TXL5kI9pPvRCwpXfxIpC6VAL/yJapZz5eVqyaklAu8pY9P2BSr9FwqQyICqzMl0I0Y20TAeTr
MdeKz4xNGuC56G8vOMB+HYyoeQIyK8+dwOrt2MEEODoKpURT0mzKt1C61mSwxKng1poaKl95eAxT
jjz+9Phz4mt8AaJ0GW89H2JEy0UjMBjwoLs5QHpNK5oUtZPS3EEfZIq6Xk1dJv4y0ITUlDueS2xn
2790NLGmlOugRH16DSHz+YOTtx6U7T0hBWtGf9snbo9jqPCWT0O0g21HmZ8Ii5uO8K3BR7IDdqm5
os+78WEgWOZfaG8q52KZoclvIn43ldAIpTcgsPqVvlwkWJnPWF5py3PuXnz0Ep3qzjp/hceCt848
ow51Ou+UdBIA03iPdJSvhQjrUtVdfG1CKJgWyttswoHrLrDBiY5RmLyRSZ94gmO9EomZy+trL5+z
ZMuOnvezHtKRogxFx2x6H8kAkqRBqp7WASMDOhoVRq/HmbMx2iBeskkCv0Uf0tAKkNv+yluZ3v2m
pVLGA/3e52XCghp9TmoShmLsHWerNzPO+4HIz+fEDyM0Cu36STFawdEWWcyxWF5l6QtBuWxMp+V1
Z4VWnPRmtJe3XxC09QGS93UR68gFYhwhGoLFksYVpelJa4pxpaTdKeQzk3dwATiiLjvfCo36ng5W
Qqt3OLH6ax1tii7hmbyKKXDGqNdFpI6xtOyl7W7cVkQa9XKIvIYbm9hFthkve+afJ0bVKqVLPNl4
oYisbw/Wj0et5RT74RMDZ2LrgjXNEXFCXR5pJXV9tzUoxCZIKMEEfwHT7PH+SZjtlY4D5WtsO0pf
VuMbGqUaE1CrUqScl1t/Hoerg4s+0BdQNV+NOGJMImAFchhO3Shy9ph/BpEwG5vP6xrp9CAPHBvS
zIZI59z43EIvHXlM75cyidadSpRknWEtRD3/YjWMDs7qUP2QAPTpwovQF7yVsCGZaIyCMxV9qsDJ
1TF/L4ICIRGVZY2VTeoIM3bl6+o/Rvft/XKTQoJQYTVzHO+tmKJFBqHY64fP3w8VdcTcnghrpPTF
un+RuBITPQWlarZnvuBDDeD6kE8DZuv0woKV8YDMKQl78bHiU/o8jSWA5GVI8cRATXtvIh0Uzhv5
APTGvxX17Wg3ej9c9POLMSAGNV1msnJzNiKzkZt9DRGQv8egTpeN/NOmOnXVpjO09Tb3HmZisi53
WP5c8etneq7j8kyB4DR3aFVyg7/wGhFjguVlhsYUS7O7dFuA8X45LxVShvbOIjuiqFuv3sCEnGuu
tgpIflldwQV5cZUfjUYQIM4ajT/4HhSFu6zWXcPKUgL0PKhLd2+n3FBw9kQsfQp0wDbpO8awz5lT
saKav47W725zdlV68/FeFVFvMmi1Nr+hh9ScwkDVsoYt6YnrTMhCx5P2NmxrVzcri6/KrIKl5s7R
p/QGWTOpLwP3VLw9H6mWhjj8o2/RYBbEfxL67Tqqs254feGOXYZN+PO3QrQ4bzBo+RejgFq0qTk3
FgySro0Jio+dATGaP5eIvL9cVBv8ihK2PPlDvJxhsKpiD+rbzH/1w2JlvYdqWKyBfNdWZvMkeOqD
HInwHYHUYLj/DHAeScNNya+XzQldBUsGo0mrIlzWISrvEgoHU5ZAOizSlTFFY7+oUZt6sbxj/RNT
U/DL4FUGaJMsDzAflwuX+nlZsvE8DDoZkznsb4v8iohCH+4xuYioxno3FTWUMMTpjefeDFbruupl
J4+GaoG4xls7W0dFvgnQo7Q6IhphiLpq86NSCphY1JHiovSl9Zx/C+lyYCRNOyvFdUlJ5oBtpwWv
zULpbaIaEeg7Oveps/olBfUZrVGMgYnRrkf2szdxX6886GwGUSImv85UhmuceG8MTVAnQPex22zA
qXzLBF0S4r9GekX97foRR7oKjNjUbCKlIOlnqhNjg7ZxvVt/8DUH9srasWQR8i5xltZv7tgDTYTE
03PZ0QjFN3HczGkPbl7OaAaUxvIYnpdL1gvFwmVnh/R1uxL/aGHn0aOuuWzdrA9Cw6WuuUNT09oy
dMpaKJlHkCAjttPro7m0PW5CbNGFaTN0cFA3Qvs+pvIn4aeAQZdQF+B7VqXc5HT/kahYpQsRUaua
gjI3JaS9eVE7oQFjtkWx3lrzRshoAL0Z67/+u2H2xYtQLqR1R1PD/f2LUAFGp7JS250lDHH8G70Z
nL1IHDxf6PviNhlDFZ4D+jt12RdQy1fLvdpCtNePpTFxFgyCWHF2s40m/aaHARCyQZIBC2Z5qvuM
bKEQD5Kl4sGvwRur+WiNUuSJVtg3IUNblHWO7EP4vZN+hhBjUS6mrPWS+cBQRfJ3+FIoF6I3SK0k
jTO78hyMq9TrRU8HdFHwxRI5zT/VLXF31Hz1UDVM8wGnINNjuB8hh3VQRTX0wiRAqgVvxWRvqr6a
wjCvhh3VyhibsJkcuCWDQk9izF0Ki1Zkm0cnbfJa5qBXsi9NVmuy10h53PcGCBuWSC/Qcgmn6ElN
8kYyzeC1h6kL6Ax+oyF4qBueGuSllJ0WkyGxLL9sam64PA9uE63hTb6/eZcYkgVkB6nz1MiVc7qn
4mVfmasvFoAR6hjVHi8T4c8oRJqvUqsicyRnbY8u2Sy9BCYL5/xtCXS53D9f5zRKfb3d+0hWEPVW
TBRntJe3pDFrQXODMztxtaj7nAm90pU4q21UC5AgQdR07Miu4g2kaVGnIUA+vyRF6IH38XwaN3YI
jhb4ggE2UoBXjTy0A9V8987cdvUHWSh7IekPV2KLX4a5ivcKbE1Nq8LTMq7DSAbuJqsYAU8lvLmv
ITcUDTQw8ZzeitoLbQbTwEcb5ZB3yU4EUeSikU0wKMF1SqflffmtImzbZNjXSyOnmODlCbpM+x8M
JAqpEYS5NIQOVGRysFhEmfbHuvLnRD2dceEXJ6fXk+7rIP/cE1SpMU1oQDQHVTHx1R83xjQGCmB+
oitkKHPOUq1OG5lufIBrEVMp8fIHKXcqRSvOlPfQlEET4d8vEGVoWzJbLOMz3bCmZH0j+IzLEUY2
2Ftst2baRW1invpNHfaNJNOx4YLFHmkaeCT8UW7rtSKEw2LK20ezO2vwAtX6J7Pe4xQ83Wqrn7uc
RA0zzrV7Jl94/gmGyqjJs8qBDK674+HInoqkSV0rwAdvB4YXbEu3nCpO9UlEMetazIJBZsDoo89R
XjVrYKJ0CMYTIacr6gb2YcO/0eU+E5IKfoZX46/+SsW4eTWeGapvdMVRlwAiK3eyRQgxj3Xq/pTe
ShHvBv0bjO+QJ6S4UBkd6EF/vgPe3tEA386c3ixled8+kskdcC50K7kuF3qQK5vWZZzepzD+yOEi
CzeyzjedzJeMR/LNT+Gl7u9kl6EO/MIPie03vAYvqF1d3ue3f0uxhJ6J3LaI7YNLkivqkVg/CT3N
nCywZdFjXuaMcK4kSZeKysSR2MU+8fX5BroH5S7gsOrgH638qwhPl2zn9iPn4plKN8MJ9UkgHYBX
oZ0nRrS+4yxPpC8OJ+s70k3OWOUGz8acPV78vm21m+KSqexfAwOIyxxDnjW0M1rxw3Kl+KHjwYN/
FS3OV/a+RklKpV7QAnOVgugH1rSNaqOeQHn2HoYPuEQWpHVJrJe+gkwA9y8VlKSwa8K3OdBWoi3I
hi9ZJXGhvSZeKBOOo/r1YD7X4ZE4bl61AAgs/AIVPzZcuBl9IxBYbRIOql7nQbflgHCdLmq85ghg
BlNvPD+f4Vb29B5Z4sqLbtJ2nZmBz7JA4LrmbWfA0d4EfBBnLWHNF+xLdXjnj+74LpRnQoZIgwj+
0T9b23KKWpW9OJ8IvKKC+1kNRPPFqMwc1OpsodREBWkKXgWAX9rP9XMjiqiO5lXtlH1k3BpByTis
ykDH3R0JUIflS+/Ehb9G0YN4iQHfZz4gHYvEjyoSk+5PUSbEgSbh02R06yXnNtkjJQmpUSMAuX4e
+kMXyKsfAYpReFDwM9fXQBEOEztcshWlarC3rcibwqeB9ZPTc/iXbmzjpFGNF9ispAkLp6tCS5WB
Q6BS80XmH5CU+vqMzvFP/2rR3YwxktbZ9wy9Q9Y6gH5e+qsD/0H5gZWKvtz2ueZs9/ua+KArfvwK
Ln7hsYm1WMT3cciBoOhviNfJWMtSGfLQIbYeGJv2+DJwju9Ptt5ShffoyRyq/Ud6qskS+gKYHTp5
LOU7xg7sAt1Mu0xS4tcK8mWnnMOy25bf2vhSykmUjS9ca7Mec59FrC5Nd8AHi6UNkBQ/JdhwHWkk
kYHF6N0DS+oQ+cso82LKD4ad5ErWGsC8Qqql4iDvma0v45qvjrfMZDk9KMB4pvtAJ4D8lX59ocXV
TKElxvpnxjdd9JzJ4V6TIgvtYkz/2uOUJhiV6HWDPnw+05h21XcGyYMd55Bb1EsOPaW0XAXEdWbx
UiLj0NvZzLH9wIknnCvkAXyUXUmuMaOzpRjhFl7+e3cyzXsLsxbAhHKRIdt+Uf5NWhZYKFGPdnEe
HdAqikHhYgiYGJ3k3Gyu64a0QZBYhpnZTu07eltXsA5zNJ6iWZLJJdB2dYqBkefgYkSbkDk+8Q57
z6lhXD2n3lSXUJoFX9MByL7Nhfss0RzdE+2mxw9cUYtaCMIOdp13ugFrg2ukS/NxCWYsmVLUAru6
c0zljDg3aPK2qmbFe0+s7yhwsB0Gls/oalPIbJO6xfXM7fq9bVaFJdFObQuRo+Jc7+9/9Bq0NCRP
eKKYG2VM9emNHg7CL6GaVDcwZvZGCtqTgt+7LA9hOTgZD36gHY+UXCF2GSYV1aidzmhJr5VNFTvy
OK7KcdhPdnq/UsX5f6xDmVYGoX8hO5DUl6/5uKJihRZTUcJtooyhmNNdOGa2e//eOWgm1hifkK6G
vLYhq+9BZ6RiBuEgFoSSDRW6v9Q69a5c2aISWkIoEOPiPy2uE7lONW+yklt1BDkh/l969EGV8msi
uZy6oNI17uCodeZWpHC5SjPyf5ty6AE6Q4j1DZjzZ2F6ljdBe6Ou7VbgPXRcTNumw4FGi9H8RUVR
wswEUKNlbrd7zVmjHcDCWLB60xb/xZ8ELL7yi6jNcS6avdrCci9blDCYbKXxhSwiXn1XqRwhr6uE
P2Cteed5ktiJHOv+zt1pD+n+UT1S8ArKD/eHN+2pdYf40nhzm07GSezwyTYJSbSKTHd9YjZqieFQ
Rgw+KjZ0OUrAgZ46s0fCXrpL6GVfMJgV52m7z6fbr8pyffITnlK0nXBwPikwIjFoCGoSxZ+KJRXV
De7jnEfWroeiD4mp86j/qIxJS/p3gCBZ0xh5EwVt7pRNPin9j8octypY6/0Bry3DMuiucIjrH9bD
e3zJ7mXvl6817PdnsmwpgCJ9XNlwS9cM5xHRaanTO6MdG0WHDeNFTJ1sXYVeyBYxTugWHY7dL/C2
NcdEjQ8dOwWe/dhuyhITbermGr1JowqzJMshG1E9ii0Fti5aVYG04n/qTyC01k1anyGRDtvVxyjK
BMB6nLgxKI75LJDrWV3DB+0OCKZLBqBEdghvlxHtG2jtStohh3NlWLpMz0ktJW7yyGb4D7M8VLk5
/8gPN6FZn004965CERgzg8ldVbcEauJ9OO/S6i7vpsOogbexBQFKciaPHcLHQHG6n5XizLes9x5u
S5cQ5Qy1yJN/GBsT0hymtQVEWgFAacnhDZJuQ7D5LymnixMV8nYi9WweaISesN9ByNpubgMUJK2g
Ew9u1ticfzIuesJNzhWupjr212Bjt6uMa4Oo/ge9FfXOjgj6+3+G9gHapQoI+8u14xarIfNcLbuC
X6qC4YhT1BOdWKhl504iMoJg7RI2daVy8JeYKXamsrBsfVuQeNgtseE/QKW9fHjDd7/u+PChDyPo
Ex/xKsjLdbw/YBgMZqNCxClS+lzexx0CEhS3PfBaXvwCMkeY3rEQ8lCFnwYbHI52a5xqFeAOy1ri
DnnOhBc/nneh4Y94ExTFLB20P4mlVo7ld9LG0MBKC2XEHzZx+uJ3oGPFfgSZB+IutkZN3Cpncmv+
ge/8GRCJo8h4R83m02szKGM8nJk3M7lQ8upfq7/gLeQ9406zYvxcXR3lJPBGWc0fO73psZoxJbPB
8Dq8TkE0ZPSsWFz4Aoei2gyTXVgIFoyuL/ZnRJ6DeIeFAKvZ4j56cq40Igcsx+4QyeyGJKyHGenn
i9Gal6yXc8JuW8Va2l2Sk+t1hIEDJxuWZx/GQTIU/dZ7xC+zg4fyLcItIUFx/six0pYZIU//t5fQ
kja4lHo9q6c1se2tZ0qq5kOasI0JNPr015kf+K3wCy0nUL1W+grsrhLqJVBHA9Z7eNEvpa/3Cdo/
tO/Dn8qjQ/qwzmUsyCfsselTcEJP9uQ5G+Sx94zQbn1j0fWDXV+2P2YuYhPH59hYdl+ncPVnGlNP
7+Hj5cbVcMLZrHnEAg6fkY6e3d2BJBFB/JixY+ysyQXN0C/Wv0JjGdkqtmKJmJcrHpGLTKrIW9eQ
pwI0R5oVml1yPz+A17j5uSKPgG8ebBWkm2wocOtRRaYfXn0dyVqymo/EGwpAbN9qvcpHOBZEnWrZ
xbcu79gmAXdHfTI9oMFm2nTY1cuOP8O3ssz+4g95Gnq+EXQcSuQIGFB7mdR2foKQ54lAsuCEW9o3
H+Q3De/67rvdTHRAio3IXBLSexCG99rspywPRPgHnPg1OaWF1kPsnnNhPwxCuX6bnyelVUKLdUOZ
KnCG1nW9BeOMxp5YVO0k/hA3AFvTuvdbOWO7cZPnkZVR9WSr8x4OcVez8JNllJ+Y1UqI08Wpmz83
L4pzCt4ZGl4EFuCFxv6UqxlqI8pEzvI8YKsJ1r+mhWAuCQsLUhU0ddzsju8+BC52YpZ7nv98Aub8
1z3Rxl0eY6wKRov0VbEmmBkD68txZGJWFLY9vpqrz5CiXNdt5oTxm8SJ32wEAoYO9NB9EV/Fi5IU
ItS+/7DNiK6Vesio3qiy+ZmoqZSDhBAQtAL/T/dycZPV0NMIvnN+Uin0Zi8CLKUPIVffzG9oquxO
ze2Hf1y4RuJZvl2LpPelM+SpURI9OZ7mYz3RUEGH/Zsc0mM+JMJYhvIhQgqjirYXq9r5WdJq9A9M
PygUtjrifrM5VSBAr87sy9ojQ7pP1Mi6DRsbKpUyGNxav/WMsNjHmq9jA8PYaGiT0RTU7PUmWrLg
GKhUiXnNvp8DSCPZTKyo2S/R8k+rweSa7/Qi8QuBNiOPTGKTXJlDJMB96yLORfJ31WUT2pE+qZAr
EtH8Bfm9s8Yd7DjdmTuIs8O4rH0NYMGOzYplG68fWmi6fP0ylgrpNjQU0oxqMxomGfIgTZjH4b1m
b8PrpZwqmiwM6u8n4i/BgnmZfwSY6cgyaZnAd8TfVg8k+oZ6mikNq3IrcSvlNgqTGgVTD/LatanN
BpUlSAldE7rRgQ65oxC7bwrfmCzWUcMcM+9wNT60iAMfKnRCBEEjvIE98zwWBpqQLCo4FIi1C4Yd
xMJBhFfor0aCZVu0qpbMGrb0ueXpSEZEdzMNlkNzCZ7mlfJ5FIrg+HQfTQqDYvfIUR+poQ7bDZ5T
DRuYeAmkP1HZTfoMcZJI8uaZEAkJA2uypVC7ikjLUm0ntTEGEtyrOLbretHWO5rdG/mhLr/j9LZx
vc77gqCG9SQpj4hDl0yGGqTyA86CQjDE4PZR0fFigS7xXL4VIvpqJAX66ll8PGvVYVD/4ibIhdk2
Ix6P7jfa2t/To6cRLK1TaG0nPy04ImyVuFeDQr2FcFfSId1w3X+FavigJ5Q7+it1fGeAk3PcgjNU
wEpgzzY+OV7RoFlctu1bWraVO3DvLK811uSYpQ7w/0Bvcu4i7dwHy7vNsFRM31H6S7FUwE8ixfNe
KOlzhVKroD8sjgXg/xkj2RuPEOuUXytAsn28s62mZjrcIHDLlYbT7tUnZof1yYY33kJGkB79DQV8
nx0GXrRaII8cALhlf1ovajkXQk0dqCGJ40R5msy1KEkbytyXijxIo6DG5GYbCDWnApgOiSdnNjMM
2zcTPw6h//5f2wdqbt48KxIjoMY39UQOHIQgCgb+1WWrAHJNc+5UXicNNL/jtEJeziPEy4Q2S1gS
PR8OvmToGuApIYcr9B1NXp1rAwcJPHhORMLQctjADOkKBokqCcGoqGuiXRAUHGML9btLg/IP/h3F
XIzqOn1q6Zh4asSTs2VOW9gbUvnN7l11REPCF8GCLgdLYGUxidjqc3jO6lKDszQDh109DrPtzkbs
fkZ10NJ1ZImtcOqg9tg+LfB3ve1tnabb1QMklJUYc3ahvvIEUNGC4pGIguBDa6RGjOETsTahH+12
7PM17HEQbKE301HXHIExueiLxM6SxRnmvXAit/2OxoE8XDzrWuzcOf3tpbT+btGod7U31p+yQYlv
5Torsa7e21D51GOMe3GIEI/XiLE3yjb7KOps3CFbE3GBvSqiPI8O0jZCB9/JMd53npyu2Zow1lxB
kUCoIsOiisLQyfY57XSmeC20DbZbQDXJJUMDwPwaaKUFn6LYA+9lCQ9ji/v1926lMSrOYPTMkLjt
iFtU8UtlB7Mt0kIChi+/c33x8tHxyqwqsZguit/vVZyj8HlxzimW8l2RLbDqE9zfMokbPzcizbkP
RNvz0gjBUnec9PPrEZOr/15Mqe6lyfYJ9QtN+qb5fn129Klyk0kSH+vcVZ87ih/5qFdC1Xl40qR0
UJu9AS3nXEZmTRnd128z7BG2mvoiHIXjPoB/lrhyGL6/G/HctuFpNoWJEQ/Sfp+9yBPfCszerbII
k0lqPBTocdjoJSY85T5o77b/ESv2UcYumoCgN8L7yVQrIEET459p7T9mlTH3vWRem+nHreHB04le
kW+69I/QeWLCLnlUqPR1wcZ2kEq21D8gxZ+iQQNJtsD4kpeF8DNW3CrChd+x5xpg15TzAtjvFaGL
mpqVPYFw+5UviQeGiXeibFyE1M+NCeryubWgOI0eL24qIhYsfgcwSwk+xpOzt9uCyQGjDvZni5RT
Iy+nVUoyvMC4WWnwyWncG1eDjxsDbcBqmONkIUPRzyyAHigATWYvEEO8qkzjeAoQGLS8c4LA/TyR
CucaoUnBKvzwJeX2IzhAJuWhptdd+rUIrM6fW3pnC6ArvHC8dsAClhqSsjtrAqnA/66CwKl2vIxQ
GtzrhXxCuh7KyOjNxSJnsvTCJoeSbx55dH/RiGCAGZgfX5foD4BZDAcTKiPpuOPV2it0W/yZCOwv
mRJjdT2KcRMqoBkmCjETuE4YXSCyRuzqz5vzwyWSVaXPdALm4VHmc6kglzfbVord9XDXUdigbO5g
um6QA/jGrL+EIyhR9lLc8I8d9hfQdD218caYXKvcWPljJK1LMpnhRr9bmSvw8ynzvJabwQncD6mN
55bMd7MnoUt7P3EK0H8AOy005j0YoD6lNYFS2KB2pZviksRGoK6A4FnC9EgoYlir0RWjxEptl06/
rfYvPaOHd5rb3r2kht63fp1i87k9mPIWhjGHDlRsRkJA/H5MgUEcwVh5e7hDtshky9vVXIenPi3O
615FbGsXtHyOb8L7ats0p86rNC11ZuMP/ToRouLSuetSezwsR3y4eXTVPQzGHK6KMnZ1bgs8NOYc
0iVtmuKXlW5ClCd4ZB7nd7dvgz1waz/3Av8/a3w6CQImuSZ/9uzPUTCLl2fhRaTiPwRXx8cbZmug
dc3ZK6UdIlgTChByRTUZwUaRhM4EbCa2ONEt289E4L0h11MinsxJi5xkP1LjbViQfTP4hbQjOXRi
we78RJCZOveLX+nLq3Rzl54A4QL2Dyh3WNlnSpapSOQUoHUhDdqhUb/9nhgxnLN+G32srUeTUccK
FZZeiJ30nFf0uJq6ONfisMRjA2o2wshgVxYVKp+c7agT7GNrmJzkRodMIphVX9rdLIxrdw8XndnF
ArdsROyqeqU2yX0qi0uFGBqKwpN1eQz4zAcX11bY/tDFgT/I0awyyNS3ajtfc1y0oenl/Ra3BCW2
r53xYjl7Fe78cJglPrvNvsDJOITl8P1pOlMp2Q4YNgf3N4tM88YU5PB/Qd2eO2Hi//28BBW2Z7PC
7amiIxw33DLWgYZ/cyBnekaJbd9tQDyPXFi1/Z/KG9PZJBXNn0XXwa6f3YAoJx7+n4GYpn3mKX6H
vLR6aaYoaWPD196EGuohwDNKKaCv317uFZgXpdC+tUnF93s1zf1wh3dOInmtOphODqba5BVZdjb4
hKoiYw26TLx0oF85ulifHaJKGEnCMlqd+e9yPU8ZNn5S0YLAC+vn5j1r5CPVEcGaXUsOvlE1XGWH
NE4tq5dsIs9+ymI3SpcmvaagsrgeiggAjzju3oLEjcQ/WaO8A6L8lWKBOnFeK6VV76AZ5wCDsvWS
TG5nnWK/UqIKkI9T7jEMka/kqeUtZ0o+MFw7oCMHKlnJfr8vbk9esAcPdDArr2V1OkvCS8tWBJgU
T8lSgaD9WajvfxXBCSb+dV9TxCwoIVhZdGquvVG6eHSoW2ybVhiootF4v6Dw0JixhF5BTcIMsoYi
zbgcKjXGsgPxLwGLKCvA8fomdc/nshjiqkyw34VuH/C/xpFhloEcCsN0ywxTWTUW4WEAju3ywEfa
IFX8s6DVi6k4b5AImXh0kpW96frTDS9qZckF1TDJ9ZudrlnuEKuDUnO9ItXFiYjEqhsDU6p3Atan
qMsX4q3m2YTMn/YaVFnrEum3sIwYOnnJ9ahbaL8W5gwas3QPUUK0JRk6SfFoKpvKqOXXxOykTH0k
LjE4oW+1XVX/nNCWBLA/QHzISvSWpTTJ7WsqwEVgSW5rYDRQjSxm1i/arZAqldXm62ZfcQrjfHsZ
bhv5e6LRBlImM68/tuvAaWjeSfg5sAXgEzeyJUmN9q+3goCmvF+cQfb28hKkUBY1x4UDkG0Oph1l
U1fdQZSp3GbRG+mVU4SnUF2XhCVCYDcCV4UAHsndj4nunQH0zg2CHFTYsi1hP6Lx7LFUuxnCunyE
FkQl8YaXPY8AuZXhHljxOtnDgCDwxQUmyoU5bfHzQexnMFbBNPUzUO7XVyWO+nqZoSev3RBwcw6Q
+/jvanlDakArEP3XtI2MjXoHf68uWQRjh5jDR/8DefpGd60qN2c4BDXJ8vAvVB+BjvjLd7u7s4Mc
A+FSBgpmf0KrXLFDQaEF/CWwm0F1SFx+GCS21C0zgIxX11SpYPoF8klz8Kx3hhyGRPfyNUz7oPpn
izMclllhmzEnt4HDtmMnJXiIR4TmI6QfSmaZgKH684wsrFezZPDNWV9v7KVeCP5UfcoQbgUf9+LL
dBRb7WH2KuosDmb/qGD2VdFbpDUiov2cjHibf5VXHSWC5WmL/WLt8JPYrt6RfJqEBSsbyV1LxeEN
UR+k8yy7l4RBMK9sMyqaC66GhQOunrHzeeOsibKPeSJGKXx738Uu8ZDZVqW0MGGT325qV1C0Wx6X
ofjMU/4HBEp3O7C3Zou2yI7ShCqi15a+/hjWL4YC+IEfdunKYeUXRwSjH4exsnuisNyQf6CB++Fe
FWTuSfpTjsZkp8HlL9uDt3PcdICxLBD8BEa6w5jqVrueP1+QK9Lo7yPZ1IdX0layjDXf2M00Rj3T
xNaYAFjrVRgkzf5IUma4CKasic2sTDyo0c/OTOXAnBgZpCpzYGwtWlrEluAbd6RqCvoXd7Qh4fsP
mTBeuEc/fElIZSFmFwc5eJs0YiYtaZDoAZD+3tNuBCSxGlvOgXIkzRYuagZhStcylQ0KI1kL3Dpu
Wqaf8y8RgyERoXxO296mxZ2CmXbqIrIb525gUYKYVQ/9FR8PKg0IS2P8gbYI/LmhIeXq/1COkONc
O4P87ly54FwgAwZZ7bmMy4Cm33U/KhboDRjON5DDuYd4x2CcMOjOPC0QuTXKeG1c6G4nCpGJo4a9
m6i+h9B/WBrwOT7PkUpsB9mQaL2wwEhOCa0tNYlGXbEere1xiW2taFbfgWCRuQ1vTDrwOl98E52E
e6Hw+kH+WcSxXQF5i8ZiSLG6hpfDPoZTlWQ4gwtKIwHKYAu/mnrOgEzFYbgNev2EL9hOpp0ew7Y9
uLZgribRiZeS1nuL5YsRMc8H5tv4yjHxsa+K5GAmK6DGIEjQontn/9i/i4crOQiw1WSHxkKzl99w
I2UbKVbG5Gw5q84B+6dMh7lql/BwWuI5ehIgRDTIq2niP8QMjEjdcAKHMlVBh8IH43KlDt5nReUt
3u1+QQbfsuAGHoS0+1APRxXs1BdDbK5wuSUJmwuzqzbuQ47okMLT72w+ROs2AsuelJ1VDmlott89
DTlSnXaOA1uWFY3FbntjGTDWDtqghgMdkiCSOTfFVJtWf4dX/nffjnBmvLJamjX1KqwjXic3pYhn
VkiqBiDLj9suB0shBpK15HAbM8Mj3q97BdNNHVMI1+LhUzqB5Iy2xqgfZbEOWNcK4sORHQpC8kdS
u1mvI9HIFQgGeMUELdu8JKXg5D95RL0Zo+YRn0AQMFoLZR48pDfMhK6msV1m3XjAHGWu8jyTTaON
krkdY+HZ0rzEmJMg2F9C2bXp4FhutvUupFFweUfHlSxyFvlWV1paO7gpvuKXO72NBOIM2XK6NAfw
upKR/35yIRWJYnWyegIEfbc3nPvpbshr1UJg1q2Yinjn2SmpUUPhqzSxUQb4n6ZoRo35Wx0r27Gu
uCmoJC3BlUika+jIvDzdQQB9WrttmONwAvL68Xi8syEFeUIuiwAW876cJakBhcdTN/KvpcjEoS2C
giAx1+wu6onZ17sUgnjrZy2QeZNOuq85wG+yLvxRY1Bn4VwEuLh1KvST0oTWaJOYAL15qfCybotK
awROL/1tUIWDXQ+jdkF2boOvAJEiYxaFJgI8nHDPUQuyzLJITX/PklCJp58W2ktAN5G93JqfKZR+
NPfwmwWUb6iLf+8EzZObhVIFkUJaEAs0HJqHFUHGSXISGlZxjwp8gpw13Dff2AI5CJqNisezfj91
wOq/gOoOwsqqvmWvDK+frzx5ttN34gtuZsFVJo6L1ABHqf0r0bKeEYqZ4p44/HlF6wuVh12NjNvx
LsVIybF6zcfHKEk++0H9IUMBcMJSup+uzW5WoJT4wrZLDznBSA+2h+WGReG31e8HL/iXlbWvM1b3
Ml71ED/ZAHf//fUE8bU1cNDFFdGUZH8m+hTduLfGGJJKEYl285iNcoev8czBkLFNHljxJwmErzUf
1P1jbkZ1AJFuoMN4ELtVINFvx9oYPiA7GlRKbGDXsoaw0QtRGhQMXHr54NkEBOBL1C4DTC3ogGlc
Fhdd4/XJjFSCSB56ScQq0sIqPTiZdFJFHQJ1q3THuQ9RGBcney4zIw4Fp2YJpNUR6D5O+IgArzt3
VB6yKp+xd1XTiuC1ylYCaSQjj/BbwXBGkPrS7shlCL5iKl+N3aqnQIV5EkmYYrCGCEuL7WszQecN
61fhwjO+XE4SPFZZlL4AcVyEvXiu/oHMxoMgAm5dvkB42IVpTUnhcAQxAdT7osFJAH7SdodgAOD6
vuH4LziBJQFbgI2LHwH452eL2OXydl6wMqQ9AJI4NO/BAoQjH2sXxBgfoDC9GXMJGYDxJrIxcBuu
dH2OV0CYq3dP+B7Maig0qNoaqRQLOP6UCoB9378n0fKpD4XM2Xc4kD0CFv3Wp/KpDbTX5dOKCe0I
pBbO/WcfHqtpGCFEwvwAW9p8VVhklS0VA+6Pf+M/nF2UmyUwfgZrF6nd1aggpozE79iisiJwzDmw
C/zY1/y7j+m7URYiI5KvVC9yIX8AlaSzkW+97VQRO+SUiLwwnCN9E+al2Wc5FFpVaHxtAauMJjNf
M633sNExlA8bioyyTGQxYPOVoi0dH6XJ+sagQgrdE+s5pBvzJ3u/ozmbJPiH1Q7vurOrdnGdxT2o
XkTz+l3IuZpc1SNOUZQF9GJcVAqONNnq0g2WY0NYSRDOEPS8Yp1X1PhcP7UrXqFSE2C5lTdHFYeg
EmDrR78DzslOGVaUCLNOtTi4T+9VSDsp3eTWxSWS1XFYo2E9cVi0MomXxAdLGuMnqg5o3Igh32og
OOoATKASwDZus3mcCeUGBv9sxNv7DSsZLqf87HmGzKeKQifaXF32sku5K5UdMtz8W00sHz3VEchA
qTZ3YFLkAvsVI7kyHKdjLwD9zTrvmkoS66QO+xlg+D00+G4otaL6WwZPEu/+wrAhs8tLZ89WyaT0
fdfgwQfviWrjKxQ+aXIuvckjBYK9rWaXLvpYBi/l1BJa5sESOSBtjvyM1Xqvci6JoaN5KLtrywZd
BLO3BpMMReLNxyCk6jUIcY8sKjdIn5ohFivpSMvt9Y8FkvBX4L4mgtAlu6O9aDOmfZIBQVB1+mTF
1lKD+3ivIYvRbQHtjJUjWclAjdUoCNRcPGCOEhllJ6CslQE9gFFrL5RfPFwM+S/4q+6gX6ieKe4m
I9r4SxEuQNTcVdnxgR0CR5oO4giVRQfDWV5VxQBfXbWh2VJZyoDrDxFr6z3dgzK6hZzGil2UnYEZ
T206TnCjI3QTdbnj3W10O1Y44GdvVMMQULstXyrYfZApzz/8GlmkyD6Yp2t5Be9sPY0o/L66k9Jl
18vxsdNz3sQiCZ1PuzdpVWA3ohEWGKoNvHIdL8DuwWFsO25VVi8CljSLIz8ybhSPpd70osk7Lj79
kUJ8wARwcaxDLI1+dVZZpXktmcq7CsHATXTy29A3vTBSgrhpXAhTNlFlGOkHaXBvHyiZAY7jqMKD
xUL7ecmonCBehfDHpz0FVif1KjEFI7JhTH6+auOdRn9fzwUnMpCSRtAQ+oDbVT/eu5UUxZFSvzFT
TnZxBpy/oT7B+sjmGBZssAM0Poy4sJVLoAK3U90U9/lhAk0cMDKtuDUpjEOxweLEs3lIMM3Klfs/
HD50A4fY9fHG2Y7KET9Zl73JX1gWQ9Ml9FNgaO8RQ5Ytw7R/WuORtfM4rmzeyBXq0omgOIJJ9O/o
0XVdEYJIEH0B5/zpzSMXqEicaN4yDDaFx231Uvgyh798Xm9A6dIf6LV5io0CX53+8n9id9eYhnO3
ormjtAomMRKhFbOpdHBRf/3uv3Z04B5EJla1PYD+fWYgFmImSOgvcAGSIEtJPmy2Y0Zxwwe8nG0O
3/lHFUpIMXLf6DKghnEIlRe4dHbSvDc2EVkAZZjHCfGyu5bwvcZQ6JjKgOvZuNqj0Es63AhkADqI
N3EcLqJsQHZoV3oAhsF2IdY7KPHrDFSxfVUNcRJPDA+mRccswr9YDpwi2lprHQ/MrgDnVEReoqZD
5h0R/nuY+bjtOUYGCnbUmGrW9rEYUzGZyZlD5mwcFl4J0bW6MWfTX24Kq1U8jwFzgZU5L1SfVdhe
pwjikZhJf4hTmqnF2nid1yk2pY5rLVtbLRjp6+pP4Q6QVaVcHLFxPVqE5O9FWJQPC1HwZXd3prn0
QgWbanjxeWIMJGQyJVD+y0r5SviEGM31kkpzRRye9uP/swT3My6o3UfPgbEtFt1af3xyff9CNvWy
lyhRRxYuCQrMtcT0wrMIHJckjnXioaGH9VyDCBv8NeBpgTfZDwmUOMlQKnN6NcTMoUo/sKm/uxA0
71BoAvy6P54DRWp5k3Tb6mORov3WcoZYl77E5R7Hk49nFXwsmhAzNrCXlb2tG/jZBGhOOEszHtyN
0o7Zjmo9zy3KkASeMGQXAl3uoVU5Z3SuqQ163zzycT++zlEaTyQ0frartn7MPjJ7oENqS/rM3lJR
LflfJyV6CKhifgnv0YSDAe4+4EJCWhb9y1J1J321Qo1eM2R4bE2i9Csxhxm6uk13fIwk1S2prskr
1kaH1K9H4r0hq/P2KtZhITK1ZacQJFFHyxTfzuuMvfG1KqmJjDD1Bezyms+tDhC8xVXSgZAk+Qur
za9cdGnV50QlWG3GbfkfI4L2t2t3ribHOzaOiqrMv3CGlFohObEZFHY2wrIReyKVAqM0OHTy1Y5T
w0/f5sqK7Z0fVKniZIr0PGsolKcOcCqdsaX3nkavLXbmIRUvslQbQ51sdn35Qi5FM0wnQsNfA+1d
0/CaJOyBswdEDrIg8z2OitozrjdPWp9gTUGq6afyvPfLGpLwZe6GFidEqYDXum+u8nI0DAqxnJyE
IKw4Sg3qyFZskLhiZzuuOXOJvSw6rzWUGwZFZqaqNBR4UMHMkAg5C+KcTnEk7k11E/V13CShpizy
1vCsLci6xQS1L0wr8AK7K5lRQHtqO2BmY2SP+H18BxibeEvEIzXL9sp894k3FaYjkcTMrPVCU2Yt
JpmEx3WLASqoXoTk5eLkJst5wjQEOBiVskO5k4iYZTcgaFEybGE8sjdbm4C+fLgUJ48UWgtBJYAU
pX0ZQA/Ciqx/9V92VnF16f4tkJqzO+sMp6I5dgXvGBynVscKXZXA8MY+pzuohTazo/k+IU2JKH1V
N56PG2SO/ol+wwO5dktjxlIuR60TdSJjKn4qE0eA2BHjek5RXfxd/R9pwLDzgMQYxs77BSfZxWXT
/wjplQgB4iZMQCBgntxGyHcc7CSJ1lvasBeghmjaX1z8UaztzCTiixvwn1eWwYIJEyPLKjJLAF04
Qj1DP9vr5CChxzEH/Z6A9aMD5zGB3DIMQX3uhSz8f5zek9rx3/yta4+zRvOs1bg/oqCiFtyCkcck
83GGkCMm7hnWezgxJrn0cq+bUuHaIvHxQZC8eXVePxrPGGwNpApwhDomTbLbnsms+JZoc0znjICf
iDSWU4MuMVng3Wd/RM7o9S2HDsQDVZxRJBcu9Wsm8zYpZ1iCpqrm28cnIvn0Hxykb8WiGYL8oK08
8FApcDsIhYgliq+Bxqe8PPRJ4QHUiLkq5+LcL3iwjyamjsUychCer1xJCt92hV1nqIPs9YalRIbx
wYk2SyUcwUrJHAvQIKtJRY/cLJGUZUIhUfqhUsj2xSDjK7Qf2FLik3B5pzDr3tTDuB198jOwjh3H
3bcmPyGcYC5FtNEqy05xH4vNNDQrXkbJps41rEG6oRx9hxqet6RbZRA5XXrEk8JDEixwOAIpr5WU
M7cpv5GVmZWUV1elrhtaCxTrkKkZQR87Ib32yZ2whaHKFwAe3QordVo02VLsB+9lrCdF1NXz46gw
5kcMnRos1NrKWp0Asxc5tcVP/wlas7caBW/0Ll7mYrA7b5pxIKaRUtd+NoBNpNlSQk9HM8BU19I3
cK0tmbl7rTZF180FCVg8iJjkWLU/c/3uWZtTK/sUb6eA0zZtE9/YtfDj6nJoExrnQzhEj/NgxFWh
2tJH4OQhdXLhjBMcKw+LkcGhx1E9EWTP8yDmHBRs4fKbbQoavIRpoPq2B0UXCQ4Rn3hctwaEtWoC
cxrbpGUPqxIqmJMXVfnWn3WhY239LymxXWfx0Xofx7PY1nJ/eB8GMIdmEtOHISjEZ/zSkj7i8qw1
LMltKP9+wmvIzOFjpwBgjuISjUsbGLcoIfmQClVSFq1iUAYZuAnUopxlRm7uhVlhtfv2176qGf3x
TZTrLy+i/3Oag6iroirSOpY/y6uemPVX+7lTB+am3SaH4Y0bnqQH8iTlGBP3hMkKI8g6lttcigbO
xmtLsXYy0IUGcXSLu1YAVh74U28Ee5ngFcXJvHYtaBRPwXuWqFuo65kDZwCqtDWTJ0vcq9EJC6Ff
rea8AhwZd81L4DEWzOak2rHdOPa94LCP0+6/EBIghBE3UnTm3HPwWgRAbRpsRKGy/PVp7CcMOSu+
zWhAHQ2fXNFhpw70WJo8YxgOf0yyd7MuFNtW68BxWqjQlvWdJ9AtU9RCIssMtLqJl8K+N07DQ5Lz
HoN7zsvOns0OG8kZ6ilX0W8p0RQT38b4JmTBnd4qPKpe5D2gfXYXW0NC+FWUOLFhsLzR6eeSaCe0
m06RdkeDeHY+qBuNHhrBxC1RdVSw1Y8k08/1P28rWZaKSC181nFFGs4jRB5rU4i//6wu159k03VA
7inx0hdLP75IdZINVA/eonEw5l2uGFAFuJmzVw3hqrm0SQr9nRR0+dPTdOzjTeeRZ0OxlyVyjHeJ
w0Y2AllxWQkpMudBdwVDTksr0+2QezWKW7OA5a5ha0uon6OcCPulZaSI5jypfURttnRMWImqp6Mt
1gPvXvjtTEMncVrM5gWBwexql7SpvlBBZx5BPAnTO8Uz0WGH1St6DD+neTZtYEJgmphpW2A1Na3c
eW+II6MKWSoln9j7C5igDnkJNONf2zTHzIz43T31sjBib6z2iKfnhb2qLxV8owSvC/QmZ3oKMzAu
cd1bwBh6fCcoFHue2PpqSnasYB2neJs56JsghZlCoRV9GVqR3vUdjTVkJ8Bp60EbwQNX8nEfY/6N
y0YkmVTJgWf6BET8o6PhuJ7LuLgTtzxHOoxlXrmdsuR/sO6mEVZpbAUv2EgP7eq1Uij1+G05MjD/
OUphbBpU0nihMPe6E1y8QOxFRk5zkt7SfBjnGWooiZtD/vI3VO7fN8gLa2kaaeomPFEvzn7A5XUE
iJ7Z/9NngxarZ3B9bnLuKdqmQsuPufS9JWSGmDC+UpDXFcmZro6pxUcTGrR34MJufotRvJloXybz
UDDchYtzTnZIyrVeMC94LjQWsYnvrgJg5BCig54WupJGD7Sc4OJ4XHZJJ5PpnadcGaltR96JiT/c
cKLV6LNhDm9K1whXqkBkc4NmeSYun3C0evCxsIiSdNs8ZdvqRBNFsHy2yFfLO1tDbtZJeuQa86/u
+V8tvgsYwbK8ae2W3rmnKgDtqBJ+LgnZewgnZE9eFNIpHGSoktQIQ3E5n+cjIzWaZcAdSlnNS91M
RQD2Pz0sc4SbZG3c3FbHsURL2J3vp6Zl8igtyt5+w6hQoVQkr4wKWp24re6qBaMDA92RCppzth3N
4G3tEtpsQFsYI2XpspGJTBovg4T2uOvPRVE3zDP5Gote6SP7z8NJi5FOQPUOhB6lZ2DFF4TCHSfS
s89DLEAGfVUsrY8mV0cd0xZbG4lP73WCLVtMNNau8BJODqt2JZ9bTPV8C2qHt8uBvwpJ6A98HWOO
HW+nCHPaGu01HniyVbaYT/VzIMQTM+7nre7SBwQOYjBRwSWdaCv8MSDpXpUzmSdsPhQ+vA3Gn4Zw
9wSfrEDF9RW7YHxVRht6TKZIm7RdCH4KlPKtB/fZ4SbNl745J9eXja+DmAwpYyDMtf3eWUvqgRD+
o43GZ2t4oZLUJIAv5uvjCPN6bzb1SI3+BdLG+FT1iMhwumfT5fd9vWlhJQKYdNAf1mN1EAelR3JO
OozSitVW7eF4o8aqF5dCItZkHlDUuJ0OIiBaYr0nSr4NVmKOJl8tvFCF+lSA6M57cp7o6JAPKLN6
IKBrL1y7inom6i2otoevbT5vF+4vmIxcy0wFEFf/otPEFvW5Ug1EqEJfKYbx2WzbAs9+lEeeL/eZ
vdYuNjIDNYUdX0RGnTcHwf8O1hTK0M6qzNWao20NqcVybCYIfacEDM3qUbm/wGjdV+qdnI/VTBYk
4j/p/RfAzEXG8JtMlRsa3hK+sNx/q8gpdfPnHeVoGyKgEi3gAtwfp+PX3SWg40/1ao4XRMH8wBP6
BZteTfg7VSzwXCyuc79hXbaks+qMbBmokm20COvVrHx6qYZFKEekKws88UJ/fq/6v+2IG0Nc1rvu
PfudtGPJ2dLLjidCJQqMgYsJIANUQ5m9j2D+p/DLS2GCi0Vuo1THzTHagu+yT3RqTyQI145QdMhS
BV5WjAuPK3LGbtOkFgy7WpsgA3RCcYGKzZKFQV6mCPlssRgh8LE18H8vZRJ8SDte0jkykstKxjjy
a/75SEwPiRcDwfMVO8/nW+yonQlQRj5V2SaLddpyjI9Zo1GqBDEh0L/0/96aLyiFmhblNiIODqlR
OE/U0kdrUqlzINBLJlm5cX/sI+rjLAOT2LoGHErBCcr5yzs3+VPzkdPZ50t/DPsB1BFgy95oj4+l
MzG5Se+Z2TE6LI0T9BwbA5xXRVzK4HGkqQmD3ofgsBERstCI0hFhvooew9C5DfmS7OyKDGq7DST3
K5qIC3d84QQS4RQ6gpit6JZnLl0LzGHq+3uXPKFwLKBIbBgNNaWJ5EMLMMjNgW+DWqd+1mCmU9LL
2d8ut/G3wnMhEe4mRb2d+6VyZU9PGeWrAKgMdUXyNmgSNgqXy/ncMuUQTdb6NbpXu2naHg77dOd3
PoD6I71x9R5KRvRAEXXQYwQ9EeE3VNW3UkGy9aHKb6eSNEXigd2W9K2Y44RVu6oVdQLftyXuzVcX
uH1RU2opVqBRqQGCnzK0ZiHobj+/5ZESlClAg55pKO9CWkRSVq/U62/2obDgm7+gTs8HJWobIg8C
ABqjQNKc4+os93yFylIQMrf3spu+dguoafE0Kde0yEkX2w1STXclt35DZzDBVCtlxuh7bisIAtSi
ijahHWehiNnfKnpv0puTtqrhA8kThZyPYAu2G0ttJLfB2uwyqzDCClCKSW+Fe9U5WGVot8XZAT54
kRnUwteLtvVzN+dqtVOWyJB0UWIuChHCjUz5M3dOklO6bvnxVklDTPQJhZMLJX5L469DCrZhoOCL
oMoZgFiVMRcgXGZffPihkzz7Te7fepIkPW/q3bRTGiC5yV0Cr6mQLN72eY71Krc6r5P4CDLuVyEK
x3nvwgoSFLmaB2nwFfUAwU3iuGHecXbFJFBE162hEKIMUvjNBo/6W1bKi1eJ354BUzCsiVS6G8V6
FUNGP2Q81fuokpIrsM1KTBOi0T/rwcD9Gm5N7SjJqSH0r1OkjAlvGj7A6h8NLh5t7Snvr+AixO7c
cIPXqBbO6W3Dr+KXAktQwTT3YAydRfqu2iSv3rk7SXDyH430owLfTDmfh99JhdN8YtghgGBUt1Qk
/ktAHZsGFjrbra7fpqEBZZ6nxNdO3E6jsVnc6OD87jIheHHOJ+4FMZBzxxPoo8AwC0rpmEhef6i7
cfvq05KSjKhsmxpBAP7GtAnVgJEzhfHUTAFXpoR5Omin8Kq0pZG/IVZmlba7LJ3Qc9E7tEoLGw04
wGhRqyZzys4W59arRDAIGb2yOHm95kGNvBtYQ0ogV6zXj9XwscUra7mwv/PK5j0h4xyDdF2zd4BL
QLF+fiMMmWKthIoaESayzrziDpCmcqqbgimYLYXwA1hFBVBH59QPQ6yJMVG4ROsusEjxcBB1BcvU
I7O5sdA43Djdm9q7E7CA/fgvNXQXa+2urjrihXVVq04waxuNDVXduYdBhT3DmVYGD7WSN5t4arvK
M+I83DilzOsfjKDzG5X3z+AiDJjlpYIUpaHl3ViIIo0F2pGKbW1TL6V9/hXu8afFe+9OWh5l5d7d
m7P0YH06hUP9tTz+RpTlGsdHYE5UuP3uXct6FMqvv8WuUyA8UPBcr24x6j8VqOe3rcCDqWEMHljA
wt6/XRl4Yn3rE+khLfUG8rXcuNdqMtBQUGYHFYEP6edrjXv6+Iu2rVKgMiPhogBCwYL5v++zpLsl
77EESSEmYJFYjKFvBtiHccMW4/CMM6Ua5nT29DeV9liTGrJ3nRP7D6K97OHw+9vlhKLwEuK3wnxs
pBlhN74QEPWqN9hAQuKkWVTqrWj/s8GP9SewT9ZxoJcAC1Kq7KcQIZRkIXVvpWEFWW4EvchEefFn
PN7jMT7VoJSHYLft+Ik5NQR9qMRqPEMmvUje8jzFlMF9mYXXMKgYWtjWueA51p7XLQPEFWLf7D2L
yVp7PbyBcptIsW9QEWbjR4aVJNGgQv/ie3pkadIDi+H4MUqBo25GGDVDHb9csvfwfmFq4cCN8gP+
UFcIXPFFp5uKm+eQzS/v8voJoh7drZxQahIWcKnr3cMub2d0rCfhyaPw4+XGKuCJ3jBtNP2xFQ9J
Avh9zamYYZS7PdpZrBqSJHZSH8xJvqsVQ0dwFex2BZmz1yLcJQ1QS2KdvD8Ww+Jm+sqCyjIYS7Hp
K0E2JsfiC6+JaI28aOX3HfErF92Fq9dxYdrBScIRPbD9JLuM/BfayNjuiE5crSMw/CKduecP/qvn
Ip6ujPucuFO+KAq7sebW9i0jUfMLPkhFXFtnUEavLLEEHmowXqYzfkZYDo/73EJcQxrohTBMcvk0
1IBmEpc9AtroxjELfdWjmqmr+BLboIwSKNOKGcReEWhVxjZjnjth2g0ufd5GIxPzTfpVAIHR81om
TOu9+E96ldDeWqri3IAKI4fYJFi72pRO16tvBo36vRAQIy+iVwz7klcQiqDWtEpYEZDT0aV8gx7e
aOeZcPsSNls9Ihkqr8FHbOhAAU+9z00Ao6ewK2HQU3z9ZoDQQnqAju/A6VkAbcHW/CnGebg9YfhY
eLxh7X09YxzBi8kcyOkNcHkbe0VfjJgNQVweqO+vkLOrOFTrHFrN5a34Tg4HKns3cuikykQxXjRd
MTVows+Jb5nTFart+qinrqoIJ0xVmj/EnuynmD6D9WDeKGFD8ASShwvTiKUGcNySzkURdvJb2uvP
f6zZB4xlV2nDUBmjmnhJY34lWjXDp7boDU0i63BQ4MrwV5MWluHUIyaSYc25fwJadF2byARnqhlp
3mH8yOXoQ6rg4Mc1cdlFgNoC4+/ltlHLQ8ayZeA4m7lz5AfDcq/CjQZmtHC3pMd/B4CkVbPQ4+BE
plh9iw4gWvjaVfb7TqOjeYPZmvU6S9BQ0Gj3Jsq35JIJ1lMOXfOliZmTOUdhwqpn6lup9Ea+pNmI
eU5dvONUDmvujUPNFVZRflBEMe25zZq40Dms4qNMObuYqd1DgwaFhnSh2YiL0/x8OwhTYF0Pdb+W
FBdkn/iYbnVGJNHVgzCVgIBowvqrJXLVEwm7vDs9n63kwLpvNqt1VRuEk2ZGGsbGVumL99hk+mf+
iO0APXJu0UaB2LZWpu1Ymusg2gyCItUz+TfRPAtsg20BII6suKJOySgcCM+cowoB+74/g9yy0HUJ
EAXnfHaSre8e2ke3TsfCevvxLbrnaEk+l7UArBl49lnE8dwDd5KEMXUAy4JLt76xx0H58bFNurQf
MGrpMlOKJ1khkikUvxSbUaJIGud/KrTY/cTNEvhL+crJb1FxVXlWcqfN8FfTKy8O495eVod5M3sq
GRn+V3/p5AYllsiBQ5paRu9q0s1h+QwIbl+Eaa89vnL9xn0BCtnNYvyqRQFgMGfxGE0RhZvF1mIZ
azhDQVwyQ1WavB7Up6I/K+YelNE5q3mmyTX/TS6IKbAY//OCiUIyRvqXoy/pWB1N77MGqtVJErH1
vSvJ3Xhd8tbfuCbH0LcjQ5f1DvCBlYUToFqDTUooWL0yTFreCY8IIBveYIYZdYmtqeAMWu0Z5Gd9
P3iwe5cNOCM2XGtvV/6wW7dl5rwNY3re78CIe+UGHKgYrjx2wxTRezLY3wBd1VXjZBIAVdL6eEZx
Cw6ezuYJRPw4gn12WTKxnwzJA7TW/kMiYOisg4+T6pklJr8qVkCgQIeME1/0RZ38hgHHqY5TKOUr
UPwNtZv2PMZb0c44YWMf2B0GWdYhjVvvMhiu7s+jWf5uKtB7yo6kLlG3z3OY33CyEgcTaa6yQlsy
s2AOHIBWTpzcCOcXdq/lwTaQVCyOP7Xjbpqh/Z9TmQBj9sT0cH2XI2+1miD42PTkiq9w5UzAp41d
LbcI9cBvuPTce+Ur+QU0ZKuKV4QnkpO4zimOQ+6JwHJ7ezI49C0kziTWhXOz9fcoMNzeE31Vzva6
rin/Oln3zcpS4O4h1NWRi/Wkutc9LtRsC/yxjHVYC9FKXNUFjRQl5+erLzPcOBHBj5PjmajzBNd8
Q4HtvufoST0XpIfNZ4H/acABtMMpWh4nLq1cLR8yrr3uqtuChHZSEnqnOamwzG4GmHTTm9AEbidK
Oyyfo/a7MdukfktzJUpOMo2maTQDCAtKhrvWHQr2nOyQ4zjnhf57Y5QYWWt0fH2dTGdhU82g1D5/
3GmtWeWL0p3oq/xOjNsGVdVkpkcBMyQd9PqcrE9CE+ur4G835UrPGSTPhPJAVE9TI5EyGvoXTwuq
6HKqz2u9HUoR0nd3aIi2ow0VSWNFQLalZkTKOOWeu39w9hFXvhFNSuStlc17WkVbAdwLitdx0hMt
R1T0DFcNGy1r7Rkt2Vp11aps/8DRDH3JFxmbnRtPf+tiAkl9fs+v7Ocnnn7+uxCHKVA1GFxSiGsr
caoABVyF45h7paoWBMfayP4lDUj/5+Ql5Y99CwfnKMWW1l+2DvprIz5/T6+DweDjB5l6k+ljzNUM
ZZvg+7MZHNq+JjnszNTFaOkS1MYMwuxzQ2kZR++UlCRghAQjRosIaPhQm3CmCaE+aTh9UV5CaMJ6
DecUqTfx7VlH5zeDnVUWeQ3Q8adrpWoEu46XzRr8QKNN87odEWFB6RJjS1uEi6mYDk3U9Vyb16Bj
l6rM28zo5P+hfFxq1w5x4v87xlqnWmbPeR139nOu0T05nAPo3+IWbxAHjI5yD8yhMRXXyaly8qZf
3mfmFlLTDGrXrS6iqYXy5bHpaIhw6LLGbzY544939Ck3lVxQUFX/FK2+9zwpgAVfyjvay6n5bL24
Oz4tJPHPXOflmP1XulC3xW3eEkRH8fA+C3hEY8CHEEwIMYq9amzq1Bhm9+t3mPDrVUuWX0+kZj+J
KWMET5hHEI7JpuU087PgEYr+F2Nu/tiLdl7t+B5rJi/GptO7rsk23RCXSHUK/7KufWIbot5DRMC7
VEeG8m6gUsIzYiiDcP9ZB695Q6IPRjPCGTtdlk8PTbSfLVrY1L9k+rJqf0KvvQpBBbdMtDz8QG7S
CVIzWiXatTJCGf1dGjQ4EOlxc96dih06dDR2rDcZQFtXW1qOCmMh4bR5QTxMFijuFvSIPPDlJ4Mp
gYdsl3RtnTIau02hD++++gAZG3SrtBui7mctauX11um0agzpkOuQ8yVtZrn/g68clPFqrbTjmT/J
OPPcbVU/r3AJLlW5bQZ/6D9RLnd514Xj7KwLLVA6Ta7Y+Y0hlBJO/n558wmYyErKzkeo/Z79S8DI
AY4IXv4mu+pNkdPWr+hnCvVNJppxRaO4Z+Jc8/ErCLhJ4KI06HHg4lckP2g/BOQRQLqPcqzx6rCb
+y/7cqvD20gpA/4E5aRv52YxkVXZ8rdiTiZj/XyIo/BGQRuC1Wz37yf0LYgpaO1VlsQpKOUqKwze
YmjhY0gR2HZSa4EYVgYs//feNJYzyKdPUkdJdcsQ61XIpVke4E00IUOPKDgHvktTFIFhpkv1bSgw
l/bLr1gpMMiM0Q5cp8he8xYy3WIQzoVnlu05YXMbjxteZBrvd0I8fhxPOM03k/ZFuc5tDIpi2n2a
vnuDfXreP17dYHoy8FPTHwx6d8qm0bnh8K7cic7VgH4T04p8HnSrWTEFB5PNfTM6mZkk4fpiP9YB
KNx1r7biZSl7sHQDVHB+xvjGtszBw5Vevsp1bkvwgUs/mG5mY+dzNDeg3tA5zdYimwcsgCfcP+sl
nvhj81we1xJas42EndD8ZulZbJysxU8cZ9WfWDxxjzXtMU8tapzmYx+KxUvuOns6fLDMM5NaVoFZ
UtywBVeAcLaQFveC3hqfdLeJuUmCeS+Js3IsiiSDcNT7FEKRpfNzq73G36nkhmy7WopSxQAttKYE
Npne69+0PfFiD4btL9hEkWc02fXFc0g5Gto7hxHwhbBV8CTPfhi+RtActNGc4nCjbiKWhPXJ6dQG
79Kd4Adh/8sJxs6wXdO69ujNaMu5k7O+Grik+a2crlleg9poD9kIJOeSLkGUzk+Q+7uh7mGXPOUF
ho8Y42KudkgSIDQf1zUkZwE9Jb9JsjWmRjqSADV6Wb2u5dXoo0tsd7KAOtBhfriA4X0GTkgSMuJE
q3VE3CPIBg7v35LW7QfYKg91lVG1+f/2obqGyPq3hg87G/xTl4ZNAEqj7pSRk1Q5nE5G5pp4OnLD
0VHkW73Lfe6AXtcR+THM9AyK3uHzmdLcqwYUkA6CepN52KY1shqCW9clwv3GJhqWvN13UG7+/pnY
3gvyi894U5P7sT9jriEBpveHEV/lzGaOHfkMWumeaQVOUhJ49GlKw+nXVm4KSshEXoSBsn6plyY9
vMc40YGUwJvD2n7xXsHM6pf6D63lM6jyW3fGbysqFa+JqskLWhHwtFHhoshi1rUthTW+rmg5PGPo
7azZeimhsmvA2P42SBjDNCtgmm7JFvE61OzuPvLA3bRs/3Kd6uGhzTO8ZbvVNCDdeZMff4JjtVFl
l6q24Ss5qkmfqJqsKQ3RRwmEcNRSJwJIw2+EKaeZDCZYzYEnmtxOsJVgfji/b4Ey0keH01UtkjtE
N4ReGjdm4mB2t9gf0OjYftV93/fI6hSK9GuWTkeyeize1nuy/NHvI7JKmm9fF+CKP15RjrijRnb8
hnEwu8H8ONdWoqPwKpDZv+mgxcuwyq221u+aXjCeazxVRIM54IV+xycaWnogTU8cm+u/gFobOPPq
2gX1B6ava1xE4ap77+V+mzcCW0iZNOK/sBafncmtlg1UH2Ml54czlaR72xJaCP9Z153AsRLymt9m
c63o9NXXzc/SvxWVEHD0A/nkbyUZYAYz4uJA9ItSqp6b6k92f5O+ktOBR18fcNMER1ubsHV9LErq
mFJKa3bsx+I2XY1jCkJf1PvmtLUHsr/hoPKGGn56NttiONEqNF4DA7kn06ZzT4622tXpjRxsUQ0Z
7t3O/xkpK4+vDSkepyN95SmRzTUll3Te/vr4wJhrpR7n381WutvAgQrSjQ6G4HtCoA+U8SFUAJtN
tIVMVmEXmObVkViOBwrc4fVipOrqMS4blEIaTaeHVgnK9VGY6r+qtq2YwHdj4M/JQxCP1dlNCOKc
MSeAeJMQJ6ZP09i0AWv4pqYeUfqLNZ9sL6wah6aKSk1ImaDpP0JnK/+bDR0s9lK5DeSOnAaYKTF5
8uKShC4a7MLxwbQ1iTrh/TXGpzDAp/j1YYEs82X0e7xB26MYtxBNeP0TK9aVADcbk3BDWZ4uz24W
N59rg7x3ij2t19rZUrN4YwNg3pufbg8PC0Kl58fosIItyqCmehhfAozS6daX6dERrP/8v+1VQWlZ
wkAaZVf0voIqTRNsY+lor1OhRNNbh25fQAEXA7aj8q6KTS52wI6tXKijPpk8Uae60uqXyvXiwl9W
B3d4MHpn6ppK9tKuKw5ieHWMstujZi9CjIu1KQlgj+HRkegiTZAy0DUab/2YBn4paPJhVCLPSIo3
nT8IiqXx9711MTTI4Rci+XhwLly8BPWByu8jzSP3scWLOfkQtEb3ZyydiIooVZ/iIY/4NXn/87PG
LJ9hGnE9lhS4pxFu3XrMgzPPXlbGPvRRi0KKtNVeNoCHZ03klFIcfjUaNF+1UVYtm9VXj0nSGWFS
m/xLfypupHYPtw0gEiaT45zaNv9sm4YpxF3gPIVtAwp80Q9GWU8yblQXlMSjQgHGsvDFlmlig4or
LiOgRGKpS9dB6KWCDmzDbWC2JokwU6vmVfdu0HNLx+mGbGolMfL5h8xW/+qU0heRE1uch53G8yPI
xrqdtS+i83BS151fC+i88NqJ+xJUROAlx0bdzXvF1m0zQVPsU6/xZ1h2ISwI6ibDsWmY2Y03JVne
832ZCtnCned+f1RzzI3dBChTF6vDWNThHPSctBuanlENb7xdng6GJZRjo7Tq9Wfojn/F6c5Recgw
G2CYB37XRWhY6YxkPCLEzsNs8AtGDIyjk6r4Vb0/u0FLeA2aYEykQ9Wf6f3vzlwCtYaqLxeVqFF8
uLfx0c4L6tL638pDWdjEHwpYx0HAuxAPPucC3LXHUNvjQdgf+iubNWSjSxM6ii67MQwPSNY+troa
W9Lwu6J/AaQoyR5sFxcGH/3L7DwpJqKn8DAR5/47p4E2fJRXxzTvKHec5kUQmJLCFRkp65LVsrRw
rRoye2m2/NATJrOP9KorLbKfp94bggyDbOjYy2Tx3Ehkw3dvCP9CIqfaTK+n5UigUAuJqu8YONpq
dmQ64HvntLfv4LLz5kIeoMho2RZCpayquihpK2hY6dlL4etPstw84c8qeq4mhHO7vqvElH9E07EF
36B7Gu/CAfSBK11pqNBGaFEaM8yDmJFymu8SRQ4506YCMGvkH/CDNV4Um062HmKLYicMdr1OM34x
oCPCn6wQFCF3WQUzQjbgsyNL6ITu4791VHCKDm/N7PXmXa9khd4kjBWsoH5rB+LELG4KJCIL1ccH
4LVxGmkOJzxOgoUFRuXs0jbDtrLvBmso6adsqb2Sj9pCfkY+wwY81kQGNyWnPzE3yKHb9BUlBGYY
ggQHE9Op30YDzK+HcQVvCTYwia2zj9F6piFprLBk502ttZ8fQzhwmCSxRS2AHXVD4ffTuPJodywz
U8joOxZ5lfRZI4b0j67tK8eQtbjEcDum/ADtstcAp6hziqDTKcCXXC0oi8t0be01LgLM4T6ONGay
1xOxeR9Mobpp0RcAwFP5/QQIXFHKIrt38WGCSBuQl3/5V3puYzwJvZS/fT7MUfRBXHwhIRqVPTsR
RBtsdXt3DZe6kC4oBvcaqArf8/1cklhtMb+mwp+3KrVkQDTsRdu8phsbnrlOb18PlhSVhlNalKA1
BiyIJifcaI+yXRQDQGgajizQGalJ1rOV6scPVuSgAtWPJjhuX5YkxVSBY9zJUG1fBhGWsJc92I2h
M7bomEhWvc1QjBSZ+lljE3TmaSOVE8phXH0UxyUsD39v4Bauc4nE0DQz+AXnGNdX3KJNlEc4R0Rc
/6ZPBnbDoOJ77CosCNd5paZ0m/+GbMTtC9xbOthon3195W8pd9FyJ8lAU4OyvRm3eLPJbpX24+hH
ffHUdTyVuujILRASiLWADzxkkAdO9SU4BqE74Si1rwD7XqgzFBgY2M+GRBth+INE+VszGthFC5og
BrwyLNAINwWyhDIM4c5q/h9ZCDONGH6Bc5lr7Ju+rBP4MmjqmwF8ShkPokWm6cYTB72sNWZNxXxy
H49gbMlpwVjFpD0AGhFG2HY+52Cr+e+G6r9IoloAiYlreAihDymMYlAzTs+IiD0Bktab9FI9nYWN
KEDkyjdaifWzbXTrNH2hVP7RYnCzLFVp1LvN8dU//xD8RU8/Gw4WE/pJfsgibEZcEk2LABFJDtcE
ndXHepk5ZlBlHBV+04XrmuyXNAZL1MysGcLryUT02bYQtEjEf7YgakbsnXlVFfzPMF34SvaTJkcC
Fqp4rdR2AD+rhOYqE82sbkqx7fxH3ieKt/dpabO6OlyZV594nx0mBw33ApT/Fhu9n6bPyU43F7R6
p3uVZc7mUZyPvOjVpHAq1OhkJAV6AsAejTRcnGK+KXi5N4VIFOWiH/2EPoMLIrR/RasAANN6WwqW
yiRu+cicOccBi05VvO2uKevmLytmN0381ZL92d03mA2YDD+oZQIv1OsHYO679cCkJVEAzLl3GFlu
jxYWuWv5fru8EUNsM38Sf1raClt5tzI/jUzv2w539pITplGSCq5RfEQ8cX4+UdjSST1LOcBNSFka
MuDJBHoxOi5nZIMDNOdIHlzivYm8aE9gz6051UmByPO3pIBl4yvi79hPnHECMtCmUx0xlnLSVnYL
ORU8fNxlPZPBJCErYaafXCjCbkrMs1kNAaHfEZJ8RLfIPXxo1dSkEUwtD3AlakjExvz+J5imrJIH
pn4sl1UvoUG8mMUKm6FwMAbM6nkSvutVWmCVnVo632G/KB7FXyan+SXiSs9V349Enf8fTxgvf4ZQ
fP/hCJSwqs6Db8X9ZK17uau45thzDXxaprhHWN3VoKKRBS+OmGK7fQ7x7LLYeugFxv9d0dzdzp3p
gGtpeFlOIPRR2cn1B0+4M+vjlQhbOWGWOyHfSRHaEiTo/6A9XTUlqPrXKjmoU2aPFNdWhwbAQ+vu
hkDxPIBrCRoWGTI40WcrUV7KCjI4BDDUpW7MKTB1dSHeSDnNE8fQV1QVUltqN/pzS+yNuQWu0R+V
BLXQsbiJUnGoSS9uhoyjz0dqCkzQt7bPXl9jQMpU/UhdgXfaPZNpROJaT/G4OeelJNJAIfJLw7mX
ZI0tg0K5h8EkkHRphAk7CIeVVvk0QQCTDuFJvx5O28HNLvjmE0R8E8Rq3INa0RYU7waKK4bCJGgu
/4dajwoxDF8AuzykEMGFBbbuPpJmRfMi7FU33kM4tIRXUlucn7fvKVc2GWC6AJTEJ/j3PEmscWkv
n+BWsTmIDEORjmkE4/BFiw0UP55d8SUPe5qpnzdVz3QnkS9Fuc5Cd32YnAHw6DaS+WmtDtPkdOTQ
Jb9phim1632E8AwYA3Pm14c1NUTt2x67yr6gDS5BBH16p1cQeB6USX2UlIPi3yBEQT6vWtfDccYI
Mt+N/wOPSBMY7drohjKBkrnrQqNPsx1O4Vl6rSV3/pYK+cu6V1KGEz0jqirPK7WzVJlk3RpAIX7/
PZHb53FcEqLvp2qLz93RKCKuUTC4ucXod8kv+ArWxn9oRZyfrpKprVo85sxTFe0sK3WCNho2YMWU
2L86CSInP0VW0CnZ+bXwBSz1ueHdTwZTq3Q1HFdciKhbkei+Hg0IaZcAZ4KHyAgn/BIVltjBvaBJ
awGpCpbLTBbrMMbPXIactuf89DOvHynKP7mx2Snadvz5DrLmOh5SVBMGApSiRbKfFsOYBrkTytf/
Ym+EiMukl+4g3ULuLTm1gSJgqIw+LwJBfvRtID/NPLe522wpS7RjqHICL8NQOQHgz528yZ/QbIjr
VPakmPXcTQPeXbis+BRLAemu/N55WoEUqAxkASfgx0YB5DAOkeT4HB5chSr91FUR0tYp0buxSJ1w
kUnOpD8FhbZNLw51xFI58jp5P8ZJw1TnP61xD1vWjJ0WG0sRpOo5pG6/1EHpuJ+BImO6XxoSomwL
rL5xUvE+BHta8O+BoCynvIWEQQDyHuzTrTzIFI9FO7tZTpSMvs1qb4I8T+F+Bx/lnwodh/ccUbEW
2dJmaCswqI7NBxJrRpX/jCY8S4pqt0Z7wLf+yN/c6kk3iw2I7mdMyju6dGaSmLc17V5xrGAQl6yd
axtX+Yh+Hm9qEG1NWA7SReF++44aCpnJRhv2Y/beOWO+8bvwLAXYRXVN24gZ+F67I6GSEO1K8NxR
IVwO3KrHHvR/But+4nygA450Wrsi5zTst+902Yip7wk61HgVDDIZ1LGeWDelmV/wlNbkHSKTmKGs
zT+zAmFzdscXje3Bg2eqSR5bZfSTD2ZBs7ZA8/XcMZCH4hB/jDvvawB/ip2/BHkXcPC+6FdjP2Cs
rj8SCh4HoyvGtgocr7WaWP2Y6yct2azh9hyDtU9DpdtLGWBjjEyralnlI2gisbWQx+hKhkJlmHVr
qP+m0KyfSvYoQrIjqjleuIr1hXFYbpYH14CdfqcZZ8oVA8zr39nO6hQ4QDhUCGwSt7DNRp1A2Y+5
Z4gWYFDaCunyiecBOlmMI1Ysd1YIzxEJgpGiaYa5oUwYYpRByKWRloCd6p98bRVrbJXMtSiB6UGW
l+rkbGULxy0spkspDRrLrVlfE1MqLarpQCWWbi4T83Wg/sd5RXFgNfcos0RWoVDec1UruhhUyxAz
HC42WfHBXehj0AmJwoASP/XjamC1lMqqUlfJ6oOFkdXDUjGW3HvEgiaLQz213nkAHO7ZdY1rP2gU
e7V+I16esnUVINMpPIEyxGFURbamRfHl8fHcVF/u874ET+Oww3Q5TAkIqubGymvkiJuXdwBId8mc
2TBu52/cwBoKkV13q+GF8s3ZiThiGLlE2hSRhKDnIlBPLeZ8Q44A+hQTfVUzjkVc7JgflMAg0Qr7
MptP6J0QYORC71D8M/VmeQEQJ2/YZL7bX84UGagVKeLC9CjjQFScX2TkmoGLPCj5ijbDdruVgbOq
yQHykxIsV2nrzT0Os07jZbyPsN8txRm0w3eY/CVMm0B9lzpAi8rdqUWSP5vx5hnt0PfYGCaQ5SRN
y2/sdIXaSI2OXMw+wVw9ikPAWxj5gfy94FWJc4W+QnH++/iquBhZ/+l5A7BVJVU2iacmkX6IjTc4
e8aqx4HXCXQLm/0ro9yBA4sIxkRdFwYjxh/LrgmwFF9n2n9jkQEoHUjqJUsFFcxzeWdo0VVolFi0
B9hiD7S1xy6F5OF9E29hgSTWdV8nV6ROMfaVPVRB6CCZp5XdXND9DhYZPqTQaGxIqfWXc/FDYjgd
IBLNyQ/UBypHTCNppU0jSM5EIY6ccqsQd0qtWWG9QW1EkLA8l/n2xXR5h+VyCNYjjCNIOisXfULb
8oZLPgmq3/pHZftvuH1bb6+8rAQufZHkjNMNDMYB07zgkFs8gFQP7wz0JR5lf8gehA3xeMIK5HZv
rkTg43mF8CA1/1jotwRAUmzTWf5Mhv/n+EVsuswsTwSSVh1jW6sv9Pu//poPL70RuwrOwsr0HHpD
dlYPvEfJsqXzobqSw1pfjFs+xuweFNpRnUjfGwrYibCgj6zVEZpHoSu6DPjZc/VWzHolE2ImcrDg
QrGB9cFAPKRDWsZVzfYE74S8MuI/zL2dNCKNWUP2pIYnUrPWfE/RvKx9OQJbFqKDbbiRab7ArNcF
zHXjRU4MOm9wG7Ijdpf7IgM+CYKPPgqbJrOOHaI0HdyGrv4q7Rws9ywqHGCcP0X4+2DT41Ubm0pz
NwtScNcaBZj8RdtuRVcIL865afvNhRCNuhtze3myE9jJDF0rH45T8Mcg8ywb+rm1jEVYoIki/Py4
YZhEAFv7GymhOJEKX6swDblhBA89RYrA/6FE0fVY/hRApYtQngDv/QnKz6hoHs0VTi9PflHLl9R4
XFeHLAs4Af3BXTHIak1CADqhQnBilWwj1SsIkCLiKRVELtxXlScqOCwnYkGaqgSEs+AubgUS/9sF
IYe3uD3gcBl48btYopgMbFRiqE7FA3GXV6Gsu7FLV3xrXxxk/8+gExBZc9XhpGNrbs17jZ4m/zoh
yaxrqf77xrXPRLSDUSvA1BNHkSW61PG5M5VZXKETRSO4aEf3USF6ZPWb3gkAxsMVUmYnDjTRM4ne
X+YP4IaCubZkgH+oUBF6pvaL0onPAJl91bip0rpSvbqNO8pVgPMPHIK7V8uyzPr7Y1Q1cM3CMGVc
OJMXfHSSEzlfJoIhGNn2OGAhcvzFM461PUbVUlj4ZisicV5xPmbtOlK5qOxofpp+dP22mpwge9cV
jHbdb5tzT7PWuBEQ33Ts5bH08XjkSK3giOtpqMV897qAUjH0djP4V2lLt5gSAPP3toAWUzt85rG0
Ap8yi547jPiSoxgDd6XciNAMSCOfarh6Hmo8R+hfKUlyfz9Ly8zhdrjCBU3sdV+ohAeqnCs3ihz1
GQ5u7YNlYY43flZavkPVir1iakHKWyFMllRGKMt4VuJTyHcA1Cc90twp8VzUh5GkXLNTaVV+O4kF
20vsej4qrgeUcFpkZRvisphMvXJDQ0VtGKG4YFMU7MhhHNuhLyfMgjmWONlA1X0T4FukTGxMVlIC
LocOw1xf0YKm6D1WpS7JVfMQNFC5reZDt17pU3l/ZNYUFTdjBKrhi7XdPOE5mZrIyblaAiRvvZBq
+pKyPsbfJarrV5Mhx+eoTpsLsyc9ZOPBmlxnXauSAA9/zFmZc6wwVBnJdhgjprtFYs+ZkGUt5WRg
b8nrMdLwayi5UE21v6HokFRI2boF1RY1LdS1jk7BxXbEj95LM6EFiZ4SgNoaLqSRD8nfINFUIi2m
cEyGtfNKCeenimSwfvNgA3FU5UBQS/hm44vsqx/oF++TzfVmZxJuD1YS4o9MSxwb+gTCt5Oi5kjd
1dZDQT6qdlJjZuMoTBs4jBAtnevjLVg8oKbajUNqcQt8QTVArSdC6nf589QJJlxqjJteTSAyBNnK
BA1gDoLC1nMIbQl8qGoz/R2LYX8wy4Ac9mOrbE/nwwfzR8FqvW5NITdssy2JX0yvQvpUcoUjLngE
kimNz4Q4mo7bf+NWjHUPMC6pimhQy5lmfFbV+fxKMFwS6p/E9Wih0i/4cRbHwV9BogEOLNwhdrf4
xJC5HriNqopmencBu4EwyqsdgBhahJ6BRXsjCEfMi3/DCGzaQC+fIoW2Z1I+6WHVIRw98Gmi7cN/
HLdiN0u04cjROOpeimLrI4q/Cf0IssQoa9btCG3aZ7+rHDX3AaVmL4DUR75Yjj1TgOO+S4z/9y3e
yyMiTz2VW+Hb+BwpEGnjHg2NUUdrBhzJR7JgI6yAafMe81JSr6hJ6/cmD+TkaCHWze+h1x7xS7Dv
Wk2ofLch40urwfTyp5LQk0YwXZlNoy4uxWRb0275neWvFq4vCHYIMA11vF/z/OMZlHb3s2ek5foc
VFxWJjdQil1uH7fJbYgevl7opZHrwpIgBkoqZPKytl5vBprOwevBs7rSAqFxOlL6yEgvtRYMPJ97
kxeHv7uNWsAB6fhPGGuvb64pky/9KzU8loUoxkb0hXaepSx9gmMg5uNBrEtfk3sZbQb2MOmLwB19
uFn7BWo58s+ROvtOrJO1P0lxHYvDMWGZtVTtKINyLjFHsdkgHmLogp36SMZG31F/ZguY0uL/+uU1
d8zPkxTTtYMPlPL2HuPDC1cAbgso2dbpz/aJJonSAlXKBZ/m2KCOncCbFPYrqEAvi4Qq7h8hNV30
ASjMrTafw3OiR1sKYnro0FB2Yzig4ga7D9Ke5qIY0rMPeJD32A1WAn6i6FAfJqYet4hcIdIxkrdA
HaJech4qDAki4S/YmQVO6UgF8xkcOrNyesGjh9dmxRAFu0XmWzk+ySU2ESq02p6MZn7AHFcUhQMu
Vn2V4GAzXkaPwrCsBlTTVC0M3EnBgVdGQA44Gt2ZmKA8T69p53TtgA2b/9I5fdl30eMu/YibIM9s
xVOkCTauW1hq9+CNodAfLeGt0TZbFL7dF0sYfcKDrKpBFd2UzsrEGcqXK1HeWO1LjGKKkbGFDVVy
rOES12wSBocpbGmmjqZ2MbPUn5gYIak4EvNc4wjk7cPpMjMokznE369XZPruxC9ysXSohuVBlDY+
ZsCf9d9u/nsIRpA7lQO0MVRAykdZk9+gwjQAAsC5yOaJeaY0vTHsIcr6K8Xf19mjaYSCVP8s/+9h
9SOyVMqQXQ8HgtCHrpLxroIhe/AinMlGUeuQYXsT6n4AyKoZmNdtFRv5Z5cH4rjYihudHx+mzm8d
VvZq4BuevAz/O3k1QrJniyhTCttQA8TR67lmh6bI/wkDkzVWHgGHOE4iVEd7wVAHpMrmkUp0ABtp
nrWIFdt5Iq1D9qSm/BL23X0WXIdFmONqdPZVuwugOkjoAizkH+JdzQJTB3XgmK9byb7ztILqXggV
o0bD/orui7MumzX3zxayKmz0jJdz+zLKGE0u73z+Sf80ICYOcNp8jLpgq0kOH3m6xPAjOzPqZdhr
EAUg6plug8HUoVRVo652EFEFUTSR+jEMGMDplUhOrMPvJxLhcC8zL+JKReGgpjcTtIimTryq7sry
4LTpGBZ/WQoCMFaAQGHMVgZUn1ldHG54KbDQXpvbwrDiS6uKcTqGOOufyKACtQH7liPxgYAikchq
/CuyzKjznMXLkzQMsbzw8VGVmqkMdIkxEJwabeIGppH7bNDOTZ0vv67yNzAqeWpHzTA54iYYuosA
GgCDiXAgY0FW+l/K4YR017Lj6yfnbbAB9zrkPON3x3ADrqlFK2EzeS1WEjk2FUS2TRPqjqvxGrmo
c6/z5OFzlQNI7xjP5Ejy7srMj3L/xaWMYxDIjTWlGkYwG+RSHNPZQ/OrE43N/chVdR62m+PWJeaW
BMJVn9WZAmsF9BUw3zu7+JVlIFP4xh6xiaMFCBPGZL7MieQjcnBD2uOvNktV2v5k74c77njYm99C
Xy8KNNFgBGmn5iaphHQn+AEEUI/papBjAudd2fd80wcPtZUaEg0/KASO18Q4SfqsdWATTSP6OhR+
VOOvMCX2LEDywaiC4S2WmyIxZ2b4oBtvRdQ456dTURmK7NOoSEj3W6HlLrWq3T/MTMO5hxCkGfSE
8QYAdn7EQjxXF/SadYV4LpPyDZwam1v9DgmBhZdnAwsNkcJH/I5XCQ8Y0ztPHmYKZJ3CNFM3382Z
81KzHNEUsWwPre2zIjwT/xwChk4NbgWbfMasgqgBA6tizoTUgeVpDp9tw9PjEvJQhYVJuX2bnR2l
5JWoR/ez/wnckaNY5EQZeXqxx7yDunZfiUtsP4oADBCMomkJ+NVDPp0wH1ew7kPd0SPFpVwrs2dd
JMX8mNWd3/1uO/OxY86fH1ox57kJYSGygjFLH/ugpn7KCRjp/O+8mjERSZDcAJmmq4jEv9EOBSE7
fsCB2sNuMxSleLN6yCYbmZNMADGv5PxcS9o0eaUgUA6KrvX19VZTY36cIrfz6jyakWoSXJHijyMw
/6aq4Srh/ybmgYfUIqz2k324HDDcde0Ao2KTWzSlxaG2ISn5osebjcgMgYThq9/WEvRSHn5jqsHK
JnqhF6swyatyPh84irhZEe7xYVuZSvRaCwZTy1JuFyJEe7J7MnhzqlEYVuHoqdZ64mReAPxQtNIX
RnLqvR1pKu9m4kKRpjtbTqQzZafOvxq79XYl0oA2f7UJPD+/vwSgYfrqiedGWF00pCkSP1004Ifs
ZVBFeuB3Pdvc1uGLGVovEPPHxIU84bvMpchUsNEpO2xxVavyEkTsVKSF97O8SVw6H7qpoMLkHuKm
gD4uKau5SSdm/GjihcZSA6nS7HJBmyA6SzelHx1bS1rcL5+fbQHRAjLmoec/braXUSbllT2twwuW
cCJlaYwVsFJFAi/ysyuAAc9+6oDWDObfjYVKIx1xmpg3c5t5cw2xxZFcoqWMYdFmGHaAHTi7jGU3
SVRFZuKuR2++PEmEFFNSa9fe1vsLJVjn97a42s5XrqqVALAyh53b+kMiCPbA/pu0RGNCllup5+tP
XTsCall7EPHercmUx9K68dywBRlwydzdP/cJbfsb20z3UunKVVuNPXI/p7zZPtB2MuvTCDZb326k
QjXySW+Kmdd21ZEXMDuGSx6D3MSfy3xsz+O5htfT2qdgjK3Uqm/1g1W8VP1d9YrmOLH1WXW6CAtZ
pafX3tSyJ7kEMfn2nssZXHBSfQO9ZfsDdmGmroFZPOQsiZSURga2iFZDId3F7/9caV6cmFE4+vjD
MPEACkA5cHSWJHUTBjJHdeyEnfEluS4PbJ5zVN1Zu80kY/24xVj56MyduRlnyAXXXjJXKJ/oGGHi
G17aIPxxPe1fiij6FhGdnJxvyXOtIy3B8s3i0gnocLQ2D3gyd6cp7cUVo4Elv2MwzDrp1MqKRMxR
DaRRD8Wahkcat0u+2ZD6blN6TE0+5Om3RhpEEKIksADwKykDCB56vZhbSE/Wln1AdWsO/EBzXaww
IbVlMZsY5yOiIJyfo+qbETaP5019denYzY0F56eh7uZMeCJ6JEnJ5F3b4DHBiGaNzQm0HszkovFR
BqfE5vBC4DSOe3oHxqMeVgj+OTtoiOsOPv5W33d8BT9I8QRZZooDe7ALTjXTq7XQrTJa0IpJNnhv
AY/8Ml2ZtqgwYS1Dja+AYh9KGHkhtUyaljYqH5QJrS6EqFLy/MOALX7M3kr/wRT8a4CPUb8GTANi
HTUX8CHsE1fcAh74r1BuHDzkf9FZLMC3WLd9ZSzDsosLGuvaZCD7fSYn4/hBK5INiNJZ7Jw0i8aM
HrmHlCKzM9ejhV0WCfVDXmgLJcSrLZePDvMhNPP86L/hdkomsPh9dYJCjKuJZVeQoDJT+UvgLH7u
vDraU50FdIevkX4C+Tx/YmRmbUdxs1xhMM2JJBjdTzQY1ZH8O/YYKve9JsJQxRLWiqJKvtHtN7tY
mx0wCw+LjvfPWat5vw0tChTcPZKfQEmU+EKb3RVOrGkh/v0AoD5HiC23F5rJKPpWIQTP1lQGRCdN
Tj8IWdRoqViHvDwZckz4OeJ/Gibtdu7LBljsF63yzHwZEApAnqEvoZwbu+MZh+9Z/42lEaDvzEgQ
NwYEzvn72Vzw6FzPya+xMa6NuhAiQrfLiikiOkxwBb1mAKoQcXv4fBl/tIeH+sMdTwLwc11OYsxa
64un9QV6KAVZ6Elji3xdTGLOMlkmNxPDeBQylWqpNib89K0vEb8M7Z3Rgc1Auc+y+5ma+ycL1+DD
NC+hubOWGeJdZgKM3j9utcl1h5u1PSiY+LLGE3WUlP337Ar0gv/7eebjhJ+OFQJTMKwlsCl4xVNP
gE0RLLDAVfuGdZjtUTgMqgnaC+B7oa/rgdMQI751tcOPuoh2AafcMjvm8GkyTq+7oQoiGPlZXrs1
DFRUIbCNV1NNluSffs0fGDq+Z4Q3Mlrzpek+jrfzuuItfqAjWE+ewSqTL6G2Gh5iD6TvSSUs/u37
5oJ9Bpxk8a7gF82u4YZV6NBNjLzHmMYYUPQWRBeC79o83UaGTp0y52kRXjE/bBNv1MSEk0To9Xpr
5flaApe9SoQmN75ArclJJblhtHpwMFDuJHtBc6pflZ7R22HOYnDRZ77z/9Pnf8IOsZvjiyx3qL7n
EP9Tfh7+yXvtP87KOvNQPQd/YLMPEydSMl5uYCfDoVavvY74EkTany0aiNTmgn2a+tGaHn53Bzmp
aa/P1FaEfMGagD0wrd9cW5IelTxoMLFQBdqbxPFHd0tP4zQwvrnIpR0fcXIzdb/use+1pd4+Mjyr
1i8nH0oTwnV5WiUnd9AuD5SoXja2CsjPYUpyvYR4nNekdCXK/ippcqyfmEQDC3KJ9MLlVzeqXvma
adO0CPMbVGDVQBbdjxLsUqIxHNVmaeRekZviL4zYzvb7U7cyfS8s4boQvhtbIpY9derGmeFur+0j
Y9KqG6dQximh7D1DjkQUyUK5VkpokE3tBwIBqmVvfb4NxnUH6nd1r+/woI5JhEHqSyYoGGdyDEzw
aXLrk4EotJCi37LFGbDDC6QRamWGNZ4gXPhITXslN7z3ETJZnxacsQ78hFxl2ckekxHSMQxF3dD3
tG1Wjur3xgPMeUSpVuc3av/2kMBdRYlKpBs2xKvCr+v2UJVq3z3VNEGd2SWrj9kj4xMcou/SsgHP
4TlN3nBYanM4iXGbE3RVQY+FKqaig7FFNoQ1dl9f41ixzoHfdqKioDHaaf6Vw2OAVRTYkMjkdv6t
4j2xk/wBwHFtYzkeKpPmv2LbBaJqZoloNrRRb/P/b7ZMEINcsqJafyFQkQLRaICv6RJ8ps6pIp8e
Gap4jMuCvojeQF1WT87KWfwpigB5sKgPLPPihB4dtG4iYef6isXwaeNgteAIrcc3/LNBfRNDQN1N
K7GtLtKBWAse9MNAMJqyF+OCNPcpzinz2GUWaSLJFiyHg/aeLiWpf0g6eK9CHG5Xe62aCsF0j2+h
Ug975f2+75sRDTBlaVUGmYKz+U0rQ8iZSIBwJP6g9yWie+wZax3GROYAaL2q4aG6dVraceP3s1dc
aCiGbZKA4TTwZ8tzVmo55tI2C1ztdukV7Al6MCF0cQ9ATEhsZgNpAPmBYaZEGrA+PXnFywL0ZFsi
8JYXNYdkYC0V/j+YUHwYuo2eIjBQz0W9mCTwJGoYdODglT9VfpusqGPztrZ9JThdchEWxBybinf+
wMQFWWG0ylzLfUD/cD27aXNKEfuL1VMKlp1lCATCyn3e0u0uGPaIc/2/2DmZ7e9jO8Gr5jDOvW+m
Il4k6dNgsj6tdw/KC/egM8Turh7oOKZmSS6KqrtW6cjvQzx+FjtuYpU/aOTA98R5jp022m8RO+ht
dy1CWOblt8E3Fs+xHoW0C2TRS+8nd0xCK3J3inNAD+gYuy2vLkkwyLVYI5t2aN+q4bU9bP/d1OAU
FzvPUAU55o45kW+hdSHVuTacM/HV0pulWhkgtMuJWygCzD9hVbr5Pg2Dwg1TAmQ44kMwKthHC+gP
rUifpqSmUa8/9uX1FZU+bng3OCfoZ3i0xqN5W2s5gHxWS5a92J+hqOorbU6bZ7omtaKzH+VZlKps
osaHKy+wzZrjryExqpoarBVcCZIa5vCc5stg7Aq2fEZOxrUhCB6xSX0PfBKgzZLgBSVfais4xtnp
9xFJPJxdgoUphBN/R/dAxMTm+IFgkTSI4W5SbcJA4YeZQswwfh6iAGGBD64+GJLvE9PHjs64I654
gxrHzR9JDnX7FKaV5HDReW4V4smdxTb0Op+oqLmQrPrArFxKppuJu5q/YIAJR2oW8sAQCFPtWNSD
ZGra0OpyiqHEDe5f5ZDLi/qR5HyStKj/AIp20a1T/62YiVcGXtyISsIFi4BbCfIg2+f9mdlqE983
Q1o7hygj2j3ZqU+v0o5alZk0xk+NnsbF+dQjU3iTXSsFg9ePW5u7XI6DIdx7FDqv5dc38qHIV4L7
nRqGqi7Ecfg7tJqPVfUsuEZWd6j3GZExMohKaxANvzTUH5EF0nb8YWj8eTtOvUgqb3FxBlrdNkQ5
fY/K3XWNtv0R5LCzUumPw1Zs/qVX4ytOJLG8pDOHCo6nksm21LcZF1Nc1gZBxKihuOP3wTk1XuQi
jV6wnjxjqporxvezutTBHSgp7k+gdwWbqUuLOeH8t131cxuLzcE81sbcyjEsRF36Rs6urgBlCJFB
pdaqOWm/RHo7uQLx8lt4d3bVGdCKb3noWeFQavdeHCP9In1OIJUqu6dUU2MRo9HyUdMMBh9k1GdC
4hb0SLgMck7SUs7bZVIT+0Ke7Pw0Ot1SkhvZ9YLP2qVc+rYfbYHQ7m8p0FHcgi8zi34g+XJrL8pi
gzOftjpLIfSZkitE3WvYT+V3Vv6ofY+zeunow3lK/tebA9AUaUmnAsDGJpNk5R+knqHDR2AyTDqZ
34Cb0DWCbJ89rCbAXr0ohZZdm1VgLbyp5wEvI6QFl1nDpbpSsN+9e41ZmOAXDUJAIkmTsUIylRc5
uCRLCQf3HxVCwiQ1rfaBltjWA0ACWz4KqS4TZiYKeToXFaR49WMhbSftRcwLh+hRBX/toF2WxC9t
S2k3TxnGUm/GWZEBSvnbglSvuzYK6lAY760OBHlGSl7gdcCF5u7PniXYUS+0Ir8YkzXv+CDv15K7
Dsg/gMxRmFpBs1xZPmnw1PkwLpaPe1NwPoVDp5pM2dzXTSFAOEyF7WkwIpiwk07dUW4/UKiq7FfF
RcFB3C0YJHrKTcSpyd8nOHQYu0Di+okwFLlY5hN1xifuo3K4/J9cY7a/YukhPcm2PCVU5dyfsNgl
lnmX/Cb2UXS3DqmeWbBtCGfg6hB+i9Z/3/bKlEA/COPqZ9NnGe2Ce+xfdKTIrBM2gZLzgMRu+ZoF
4lRF5ULE5ySk0VJDEbISDJTwxqRYHVUpjZYZrhQu6lJfPc3DAqBTeESZIF8cSnPuspStxGWXOCJf
prC4IPxQ5kVoM5kmjbclBMM4n62DswcCAfThZ7Y+L088q9tiEK6QzSMoyx1ai+Q=
`pragma protect end_protected
