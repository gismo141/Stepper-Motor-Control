// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:51 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
aWcsShX9cuHFbaRWHHppge3KxuAC5S0YDzC/1GwAWrk/4r6sXSZFC8OgVnbNTkYf
V88TA/CDKhwW7e1a9YETM471vqowwPLFZy3Zo1DvJIqHwoWUlRGHY19/GvP24z3k
jn26XXHz1tCf8rubo1bFAn2I8YQjTu69QZ4+NGK9gyk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57696)
bgYlqSE8Na5AWwWb4LLHtE8f0aPtXTqWzTIufoK+EXj6eXbmFevSFiv3o0LqEJnQ
+vTHdc6/YqkacmrpgBt7Nq9hxDmm7KAiPbKwj2h8jMzReM0NxTq1WVlDAAq4czYN
tu9xIhxJo7MsKLWJiC+M3d2JTrFr/kEUyeLkx9w5PY/W4z+vYOrPTmG4WKN7x3wd
GQoqObzbjK+czK4ZwM0ZBen0FdkspggXg45GHvixfVGzj2tq8mQr+oZ2hLjEvmSm
6QH3MBsel3e2BVYWvsAjZQT+CW/ZduphNxtsIe5krJfXPlK8F6jCCd0CjFScWHK+
NW824B7gg2uT86c0/YvvKKiwtiin+8l85hOUwYoKIEMVuCzDunK2TFZvEEkO+Wvt
DKNGx0gtYUXQgJmCsFx4P/knpUXT1PZic+HjqClj7QNH3Rl9i4v2M623/h4wSyM2
/ah9y1FoTpfmQACAzF/pWAIFi7T1rHB8BpXPFSWbIXIoyEUWFXC9MUuNo5oLYsAY
9eBbA6Fs2lXfx9l4ndpRsCumbhvOAaSGwX1QK/Oip+Rems1C96d8n7ZLkcjoD05m
MepcNLUPQU9qjtNfYHX+uhW/GVtyyJ/k9R4naVueNspa6l9M86l4FIOBS5NzdAl/
f7MatRN0HDJCRoif1YoxzKHVxT3fCsPtffLkUHwl565L2Jou7K5V1JJOZLg8UjjD
LnhROzjyTzPanztEfpLH2YFalfe5KSqZEdL2vKCjH61ywc8LnYmB9/IeuyqLAIhA
43bTyOfqeAfBw+QZk+6JQWw//muqruCOs2IwC1jZQp6cRcJFTR6d+tDuvgSY46Pp
FruxJ1Y/8o4wFXTt7ezBhqU3DdPLGgqTV4w1xy63LY7Zpnv4fzrpPS3wD1NExurJ
AkHBIAnK9PugSlNEZgaU5Mykqbk56WxIBMMz5aisCitlpsjc3a55E4wqfaP1sWii
RgCv0kDO1WcEnKZPN2y81BEFNHdhWNBNz/1HGGflqBd7Oz/n1CdIU5FwY48Cythr
K7Nbtyj0FnOn873ynJLzGKtOxBvVVxn9lVhSd4x/zmwTZ21FlVD/SReRl5QUk4YW
8Lc8dTip1vKqtN8Nq8xHbjBROXsng89HwNBsRRs+6jGnysH9Vwg7aloyIGbLZHFu
L10dATSXm4+g/wsuG4Ah6bj7v5fnSqN/tGss2MT9VAcWjq/3QXAHE9DMrqeitAhn
cQZOdzvBoWl607J2apWFe5F7JtWMNzvBl6daRJ19MgwkR/MQdcy0T1vaUYqQXH4X
8EdrEyEOUN+aERo6WDWDbh9Pjlzx0BwwwPNKYacXSpglgaAtWlClWa47l26iGGlm
fDs/NNgH1tCulBuzCl6EOz/XLOI6MoPyqKPAKegrgvVDpYJFZl6vfyPjxg+42BB/
fN8ElNDMo6iRDxRuyvUutdr/Lz52mzOYjw/iv4s9vCoUe+BQLkUUOfB2yOQrn4hv
GZxCkgotrvB+wLGIh/oXBOy10lsOTDHVYwuxC4cLuS6tX0C8Zs/qEnePYA3gyusY
P3eX6f47pxA/bJ94rE1WBWDMTx5SbBzZlV87RwHKkYST4cQnhp+6w8c43QPC0VQm
zS4wyFO4bKbbwrZpix4QEe4DiZHQsvkrPuWdiJks7LQHCSh7BpplUpmKVRulWQ4O
fYe+7jtU3xYI7pvPhnd/s7Z85aEFWVP0/mopqlhbpqRgUXh7PkzjgOWQnkxDjYjf
GxI3sVqk58CUK4t1BEP230HMRLEwifW5xFmE533SUE0+WW6KeQwGlc7dN9wB2S7n
XpoKgdXGMLJ2FDagZ/2TA5u751WM/2v7A/gIWsknDVywLvLlix0EG85/R94AU2xu
EpHguKIke0qVu8LuuJTClHfgKmwA0Y8bGrLqRI4qHNS272JP/YIGUguXDZQdaVjU
5fNLpOSQ/VZvCmwyJ5c3HlPhLFfYB2N3/kbXgo3+Es6htwBNED04q8KC9dBxaSrL
HbGTjJimBPjQPeQBwNfg5snWJHt3JZsqoMkYIzKQp34tUQdPTPZ+Kl05rVIuDKbB
SMljLyjw61hp3mnQxHmFhCKS5aJpfwAxSC5hJarjcYvAU8uQeonbXbAikc2z4RK+
JUK6oIJ7F1RIJhN5JeYXxN4bPq+sfh9VMxTuPYAw5vuRMTs0wpUP3OQ13Tg1R2Zi
MFIJ1GyMCY4R+tLrv/9QwgY3I2Elr06t+0FcDlQRPXF8if/duV6mh7M+IShzy1ZR
M5w8GivoMALQu7uatVl3tFRVlsddoSwb76lRS/SnL4jT5dZNZLcOZGoaxmHNB8fm
a7RwnanaeqDgj4o6LdlG7ZtCH2ttosmgAQVcSS/th2LfxJHbVMHrtywEQb2BU6UQ
vj2Dvj+bezi6HtCPZU/BSM80pKy8dO1G8dXKRPoYGNBx+Gbov16gdbERKAcDB6SZ
3bDIMz7+Y38YRMmCh1IX5txfhSLa5qNCRX1M9+eYo1iBNK+eL8Fxr8Y3CL/OPlh+
Xv6fV22G0C1EI5na92mHXYm6C/teaMYoTUofb+BDNouWu8TF7SiyC6bvzbRsMKc2
KtrSHY8aLYI+iRENJcmj/Ovq/ODBDSrqzYDYPOKfafoNRNq/JS0mxHsLAyooFa71
dl8PMJLPTT3fJ4aoNKO6cICdAkSR/x2vnbfDMRn3I61pzkohBrC1INhSfxcSHiJf
3ac6RB7a/sNpcuJqo4bGVZoBKqyboaqr+T4Tvf49rFb5SqvbLR8/gjMCi2osusMT
KZLdpBpd90AMGy3ONfbdnsEmbWnunql0+otQT8s4VYHCbVovM8c32dJyYk01r9Za
3nUWO0ajxASCBevUZvkh3+G46uo3/p2aqJpT2f3VxvukbINBZKEGeRyeX5HlWDXB
Up/tgkvXZjkRtfzMygZWp9W9ynzjVEVEcoJ7w3REMToD135S3IrDsxkFkbkLkHwA
tDzGXH/xgjNIDju1rF0Y5CfwaEY4tdcK1Yi1RPiDIp5+AZ47fsxCg18EOC173h1W
u1GUhpUt9m4gbLQBZLdriVlcVzG5kVUFtiVXlvhE8ftmnXrJlVzhX8XUcqyq3Ihh
exA1MJMj7okTQAv2CDd+zh/CzcPAtCH0RrdHCkTQolDO3wDjC003ymhRfSCB6h5e
TTZlEZu6DbiVYEuc+J8nPWQJGpMrJcYEXHM77hu9qG+5g7d5bwMj4eHTQeQlazPL
LEVaDK/7vTde/4Gn8HBGsrr9IQTp5Ln+NlQe3TfoLDG7vz1dczWqM3e9My06gq6C
GbXkwRSmt1za+AZi/MMDSgl5uUu3ljwoifjS4P5CuX+yoV8ekh5S1way4h4Q4lOZ
3QOJXb/OxcmzcAy8BbxMC/s+lB/yj6giRpOowPzkRLh1HPFb63Uo8mN7i+XlaO6g
kcQQLqwZa05ROyIkaDUQ2yHtVlp0m5iJt4Qt2t1ot50aAmofJgXjRiOPlJ5feXAB
YBXLFhw1saHeMMwfUUCheQSOdK3E9lWgP0hc3Ij7rMmhRI6v99YzS7Gkib+0hab7
AYRn1ZE3NBSM6B2bqeaEqSYQ386vNkCoh8bvvdKNjVdBB4aVSastsp+4+Qpkbw4G
Qr+YL3vqz+v3QLfqBOWiVXn8PXh990UePm92yiwVMm09eNmR8zdcN2tfq0xBfaMa
1lGJ6raWFjTQC5arMNqpb/umPKWVgxhELGqond3JYn2ZncoSy12gYfTtMYjvkOYP
Is0V7hPC0nZv5TQZvckGSOn/Klwb8V96dIAoOmSs6tUIGDt/A0ErEvaL5ru2s4le
9lA8KEZmAaytRGdW9/62tEqtYEVlcFqSw+L5OX36QWBqIFBaC3e6d/Vn4PKGOH78
6+/mRvO63il/0iCo7j1ZYYy28nBlhpz5R11KSGcreX+/94tRh8jMrNlfdIMoU/M2
3XGmOtC+j98w/nNEz/3qdRCx6ng3uh/bY98YLTLhJZ+xY6dSvAxZdI5dVLjGunDx
imEyntFqlJZ9gUfencDxPNOmNYENF3o2bCwTPM5ljSLcDd6jcP+Go89UniqyJ/cu
5TzTld7GYVv/56wp9e1DBXQKfwt/fF/kBo8yLsbxqkkt3gZk3qwlaHE3ji5mhaiz
hOHBiVteNQxUX2P1TYO0o2kr80Ob4vKhD/vAYVzN0jNrSabdZ/DVP3o7DEL1CPfS
TbAxzgt6Ss60kH49m/X3wka0JR8uCuLN4ZmyHIK16mDlvD+bFQn/H7cD+mWt4DJJ
FOy3fIq1mMLMTq7EvHUFVZypKbyDrWCeUwqkW6YN6G7lYY5AIDoCqam6ctZEAkVg
MLSxSKW0HzDVZUYRRhq23yTkSTi9JG/wPU+OlCHWl0nu+AvviDh2AFPDI9eUmftk
COsqM7Z4nIFQA8HiWHriq8U8VK2nzJf46wus9Q/KODmFYGnUpZ8XuFEZr0K0O1j/
DS5z+qNMkvVTH42UzbfR4vd84AW/oEEYDrdkq/6CEdBdXFnaGC8hL1E/KjiIFRxt
V12wYY3s3MZFOhAxbrCri6+ReD6vtRTb3u1TNR3ZUv02TQiLn0kmQIQ+DXqyuPGv
2VcvvuDY6MDsaQZYVSkVC7rLtQI41hjlIUzi9Lxyv0mRuQ0jSQh4Buga1pxmvwL0
AQc51+aA06BZH5/23CPhVhik+YzE0IeTIuXM4j3+J7QKkdjt0/0S1VjWQu5uCPTZ
mFZI+9BB7gKJGbxkZQEhoT/yg3yPCunNT243UuvER+90nNMy4M4HKPdqMTdld6bf
+zV/zkrCOOesQJQozfLfBaEeAsbXzmMY42p8cAIBbok1mYbEzmN95x97R/GJweWM
7jeaw8IoOu37tXLkFtt+AGd8sQXqapvW6o8vKY+PcoElGnMgYFpinOM9KM0dpAc1
OYPmMOD6JLTHNFsH9ZkXHXa62K76SuLAFvG/T+TDyt0DNpJYD7NIAJDEjoQZTjV5
NiFnv5LtRNwDuSbf3dYf7JVmNghtAnLT6WBmyUuwKi97J1oGTovEr0V5QDaNIT8C
LAnweHNnChVOEX5yk3twdrhv/HbWDUoDuZ7QXg3DNxyb4uV/3TY3rhm1jK0iZWe0
Q8F+zcU/9+WqdG61omxFvUHnxuh8ZK5be//s+emG3XKN18jHwmzLv4muxOhNVy62
iDXndOZNvU7dmERlNFfLDV/npfQ0Nk6bLWLuozjzzP52vRvVF31e4ILJbBQKgWsm
5YAAoYf8Hp4685ESP8+kkNgBCtffVG3t7AiUOduxhbxBauDRpDraQ4/vEVSi2Kcw
U0gbA7g9VJS6fmMhvYULWOhGd7D6jDyhFlkXlrtgSat1b3VnNZFH6gOQgzjnaD+4
SXdm1UiITWAohUNAi7h2dZhI8X147g/8RfauIgJmQS4fliYHXcUwg4uNQepbuRHw
K+ptjaKgzLJgJ5OsCesGPPuqlCZBuAWm9c80godcH/6RXMtLXCuBUZ7O669YSqBQ
AdmD5jeJxqB63hhyQgIiGUbEqhoE1/gdnbzaIGv+PGa0j8kWW5WAf1Oz54bCwpA0
1DBrnKL34iA8ETpd5czTzhbXzzYbxLngniDRmYi7f9mLFO3rli6kV2V0Yq68uBDm
v7TChlhPbwgA7Tu+p1Pbv2rAmvmeYlUkU6KaSe7kQu1cWIP73nuVBMXg2CioEcJY
4ecOjY+Hkp3Zuo1uggoChlcangFjKds4NmkWcwn65evG7M1sXG78tFIL49MW84Rr
Xyq6Nzb53wUIhbykhQ513L5s3ZgGM4RHYU+jVAG3yiYZ2K7HsvsTqER4JowdP2DZ
q/8ENosed+YloHHeWdpo1Wpw0UwecS3DTBI37/3H7h6jGQNNZvgdLcaw64BTX8nw
5uC7nqFr7r3pU18MWzgIRTbsnQgTbnZD0ZtCfWOOr59v0jW4cod8FsW4I7eNxYXd
frIJDA98YBltaxS6fbvtBsQPhEBmqp6P7l3yjp2dW0XhTPxA0wkgRqzM3w8ZWqKa
cnx1CtFDkw5e4sJmWHdzIdi08jmkuYe9OfuQ9Z+PFFLhF9sQplaheQwJIaO3TH3/
1C2v/ySItaZxJBzSlJnD157bIBxjNzOgK+eVPz0E+47mUezXg4/pDtS0+O9wITaB
LOzZ5et21y0a6Uu1xCU1eEIg40jG4M9ozCZZoLSCBHA/HHMPOVsUPrTF3ek3aZ8Y
QQmZfu72fzdjA69unSuawRAfY0Po9VqlWqsLuEvFBVKGrGfqMSvupMfY/881H9gS
tIJnZiBTsgJ7zW0R5t7LmpEq+bRPMNZE9jR+6674FISAUEXXLB7tNsxK7HisiNgR
J0+egdBAouK6EmYsgMVoh0+k78FBPxoeuCJDS6cWgliybgeE6OqmHt9OGOSHAX7r
J97Iqwb8E+pfH3VZpv2r2rdU7HgYdDQueqOUkI9q2MbRoyuEEMnFfHf68BZB7tyT
D9SH1OzOGPZkzR11foyMcVsSAmxuZi3WFkaRsD3f3HbrGC6UlpbKk5Fj43X4NA09
6YDjtu3/PLoMviwJVg9J1R4ewGCkOuSEG27ieZWBW6uYh706tTQdBA6DO3xehRg5
cJQ+vdjg8WKWEH7S2xBwIAF7h+mLhe9huKxHCkNDA2UitLBZLkpcQWRagQIpa3fg
SlFRtHMCBtrgRTq5JaVyq96dkyL8V44KIIxSM17PuVX1Aa2bQnOJlvyD/iz0QyS6
IFEz5oSGJDgqGR85lysaAf/VuZ7uqbbFoHtT7M+eIWnTPUyNS+Hecmh3zK75Ad+h
u+mTN0/RB9WZqBkJPh9/OikRWO58RCwr3MpMAfHCBG5VX/2QokSn0ej7CvyuwZ/9
xykqu98DexIlRlalSjHjv/UECmuVu61NSsoOnl942OHeRB40o7YZakVS0crMWDlN
HQAVelzzfihGy7uCf03mJQ46s7GEr0cpayfpVyzzal05gNhra2Z2QwSl6ge0VB9r
ebQ2pDJs6ZeuKLsmy+2UGjlmZ1OoiyiQX8xfHvK6e8AuzsmMPeosWSEyN2blWpiy
XTARUm3C8vCDjWNHF1TSl4W6bHqn8snBc3xroUvykhjWyHkhekOsMdE5l98sa+3a
h8WtSoqRVGOONzlI7jc6QY9Kc9vOGvrT2gKt9M+cUb8qw07fIYum4671Jan3a+0W
UAVrHBnhr4agZ5CkwTa4Sy5ybvoG8uhmL3FDTKnI+vpJK2gJwVgrb7zYoYAjxAnP
D4j1igiEdKrjYYYJ1dX3Ofg+Z0yf3F3JV+/GJK3auZIJM4k3OqnPkS3sqzNt4kEt
w/9TLI9Y/nlkrtlV0deKzD993FiWVphAsnONNrx/YkajZavHIn4PW5Ye8vPy1/2i
mB1f9dfZa9lEbwGKtTT+T+5HhWT/CxG/lBc5ZC9C456SSWn0tTbrDVRJI4HDtjy7
ogheN0BepiRUPgUqBXeNfsqaSE4+SiVV7UXBSqlroQW04Sxu4ZZAAy3YMxq+CM8U
WNatOb4ZNu+zHJz8Ne3MtQsAK0/gcaXIo3Wr0220+EAOiWmof4Jkdgi6u2hbmffK
J3+UAFuLpdv5i22Rv831wDEDwqVs3L9z0nvTbcDWDXaFpsf/7OZH4LGBEH13uYiu
ffGfBzbT3PPwv1f3/4AcW2SmriH9/EN3SORnFz3k219c4uJcHlCNUyDcE9Wen2ou
ezGkx7qE+l43H8LcEwKM5h7FdYuRkAUS7GGdrN8tDpp2jJAfrh53U2wggIFUlgww
X8SVKhJL3qUAWheLPz0KNZ/a/i5v5IKfHXEL/SzjG3Rh4eMfK0GrP2SOU5zKB5ic
zFJSUl7vm8NOKUdsouy/aYpXutCZw+djBFs/5i0FJ2Mn2A8dausS/050BWW/2KZO
lO6obQEu0jmHJXX/rw8ZtnffImQVl5CDUy6LaBV1o+G3gXSYf5n/8jg3/a8Zl1O0
uSe9Xvhf5i40NFOw6UzuwNOtKGXVfkoa3oVPmsi3JAhXvgPZsp2+6gqVvpDM5kTJ
JM5Q1EYw8epZfyyWp0WzHuDD44WWrlr76Z7N5xpULTJJH9kPbeDk9r+vpFnyLF7q
z1i3CVCt2TkOsHLJlwc1gKRVYU/lLaCeoOCsZpkgAAkVpQwp8FYYdiVgfU8eQPP1
ztGNhjLC3CjlIxFPyYJ8eugk5/UiSy4C+gFWagXEdQO/RCsyGumNYTnTt/Sug1gl
A0pwuR0Ld84P4Zj/uRJEpmb84ad6TKwufxIWenCvJ1dY8x3bLTwTvVhhq7wgDbkA
D0uoyrElN544M9Noq72yt2LRQYYGQNsAo4XNV1WQBL6XGBW8vwsmp2Az2/cu1Sqi
JBct/jiB5fykyv39dNWg/WNGy6RcoxNKBg/WQHzGECKxvc1Bk6g+Dhe8AAlEqRZM
1tn5Gp7pZS3i+tOrNvJK4xLpiX6IRiOaCrivfrsfbfD8TB/DZw4UXLm2MRfLOYUr
kHcQY5L6p0xkU0/wb+CLXbqrrtcZUnzf5Ps6zpe3EtekigMQ1D26H+2dCpJsgjUt
lcMyW6HdnntdglaR1WBHtL1u84531ycqHggpXaeRGZ8hNprbhLqAfbcykOiYCAfj
d7Tner6yfCv0gyrrZfHo6CnTezLRW7qPgrbsZ/ru9nyxmAVoMjoffzzNMtrpcNa4
WvQTuVfVTJGyKi2xsw7cECVXGl0vYkDIpbTr7QPcaQvZHGdbiBjRPWiVPagcB5Um
FBe4TBoc1ZI36IeHkuyC/AHbX4678ZLnvMJBEEvEAB0u3VOtXNAEBPrZjTPVFZTH
IPKeEpovKLMad6wiHGi6nKF2vUVwoqO44A48Srd1JoUirSRQoIUiZDVBw8NCEiue
SjhR83u/xNvLGMo5O3G5YeVK8cKHBK0k3lEVjVoVww3nikn3FoMiG+7kJBJVEDfk
gscDI2Ds6K8s8FGoapUGGJOR4Kj7nmYzIPO6tvwaCL50wz66Xa4RrFCEDk1Yg/py
F4gfZc6brUna3bx46N6KD32+N6Y01e0vtgvxmuvLi+QNVsULqniyQuVtiOezR8+o
WhQFEpn4KUmNuXbfxOEQkJcsndql3hXeipbultVRJV669SmPeTe3KoRkQIiavN5h
EEVHd0x82J5dmhO7azTZOTrCKfE4eqA6agDMhwQGfx4JQkS8qphCnVKGbeVY9/Dh
cXK1KlWuhvx3sAWx2KiNSoFzEHMZOK+YY8exw1W0gEp84XEjdxSENmRKGfYzbpB3
CQpaUJucFf9d6mTwZxFrrzzBnydqDpPAmr7O/tQIMCJqIxoBTlWPhjgCi2fMRfZE
ySZnE0gvewIV/G772XMF0QrA/J+TCc5xAU5FrUzF7woZaUi14BhkjnEVawqnRUSJ
wuya6/mcb+7TRpEwj+7yM0MzWY/dxQqsKlEQjClqwwFNVb8Ni580JCnOGemCugV3
Jv6od/yTn5gz4TW3G8nNkQmFD/SCXKcfPM+QaFp9BTAUQO3kkNaAKqST59VfTFsa
IoSjPlSZa085GtLRnE3DTKE5isX2yAXmSvEOvJ4zTAXabhK3bWPXCxCLR8qJBlzP
pD96WgQu/bbK6Xq3TLRuy0+blArntEC12LmwZR/PcEdDULEIWlCwHbq/jvKK7ASS
xYd1S1yF/uFWYgn3qNhUgHuLWT90BLwvnIX3LarmSAeX5n/qYDsp7KRwjQc9BxZH
W/iFloDXGAtqra0+gHmzAuww+INKqj6skedOfjNVTvQXPAonY2deRnyZeqYxu8PI
zWmytEOwwwMDEQTUc3u4ngdVQe8gC0SRUJ84iKf3Kx+DdhWm+vGuyrei5PNI5rHj
9dE+dk4DggCVH7vvOV2RzYNwY8J0H+43PshqB3KfX+FyxI99O8LyVCQz/eFDhE+s
A13COzXeVJdEBoKk8mOMmnPm/qLQk4TZ3WTEYr/lGlSyQZJEpuo2mDNffiRGli+e
nOH6mHhT+yH52Biuhuf6BwCB+WuL7rx99UqdTfoEMQAxl4okZqYuODj3L51tNYWe
zhDlHY+8lRqmYQow+CT1pFli1YZFXl9cHB8PkZRxYS+1QpvznkZIuQ4BAo0jFtIV
u61Ssft2bes+z1JAQc82yinDqf6li0NyFNJmhErskfgtWjpQpiZHXFCRqwdP7zod
rCd4iy8BraYPA/YPh+vI4tQ0hcfjIXzTsGMsgfJjdXtKds44P+xxysGv2tNT3RPd
b1S6DnywIKEiAwIhnnbqtsm9DnsM4k3Vec9POZ9JZjr4yKyziUZT0R332H73Twzk
haOLiGUBXFfh47/KSazoLrtC4DQ1LwK7I8zVehDwBAnrCkl8rl9QsJOQHgJs/DiB
4BvEPWNY/0l1r1drXVBVgveu4qDNVD1y03FhpyTrxxlX0NvJ/xfVrNfz/w7EFXvu
udGlHXdMO3mdNONVpZtlHCkBerGWUP3Jw2osq+XdPCevTn7yjnQ4JEda0cmN0XSn
wk5Q9mriHzr+k3Z29n8fRPAIsOJQ3RalKwOloQp2vhTOvBnCmB3mdFqzzb2qAB/p
b30B8gxbQi9RgE+itJSuUS30gGfJWOMRXslXPIML+1hif6YzNcegb8NuQFB35TN/
umVIVs4lBh2u67oOv4dfXCS6BQ00y0qB+1ZKAKZC0ONLKyAtEYuR0q+NNjq/Sd5W
r0g7iEEEw8G33cAOj7MGuKUlul7skVsxSONo8PjDtTbeVVEdqTi3Fvxb4kENYmG2
YTG7E8Dy/fKvOfwiDvoENyhiZV1RLpsBJQ4SBNGG3B0e3VCMilPxsje+oILbOFWF
Mc1snq+yX1pFPNiyZkOWsvT/z+kaFMSH0WIxlRAgH3O+sIFE/V7Mri+KRuvoxJvK
og/dmquyRwpMfhoxSHkB1Tr646o+hsPl2SV3cvuRPHKT1Olx6gpkR8+YEYKfDcwW
iyBkuV/2AxWZ7e45Ojphuwzs32KDlKnwgjJhBIY6T3wvgTRXYjn73WJFzB+7Am93
nxkXIBPc0b8FfbWDZ7TSz0KISXxNylqkXAOcOoXh3crTQF3TFBU83d+tMThkchu7
OT/a3FXAa3EQxf01RuxUvvrH05lpwvktCsvtcE7Y+YuxQm00Ugl4UPriGhFnB24t
myO0OSGp5zdHqBQYL6L45tyHqKXBTgGw6iirNbn4tDlWFS9P9iQWApRFsHIsguOA
sDgWWnTK5b59HhPtprq5F+2XyABzEkoTKylWeM1Kt9ouJsvVqwbJz9UYiGOlFocl
EgzvHEJNPkuuJsfnFpZ9y0M/5mv+yw5b8kQ1N6Rof7d2xQWfCnmlxz+TOttCvENF
ii7zUTHRpso2QrZdNRpGr12BQVrjtuRJfk+kpWpBm6KH2M/YJkklpYUrqeuL21ke
ZaYdeli8IT0leVQC13wyae+WmsxVJB/EoxeV3Q3ZMF4jrLwp6A/Ay52rfdBb2Ia+
dam/ayLkaXFw6caDmkeIdKdT8gpNDfI7LAoUK2SW9jcU0zQ+II26AyU2dKx65pvO
OWb6PIKWA1x/W3rJYBot5XZpsR7xHMP5OSleByvgJ3Xob72sMk80WM95ziUhzVGa
H63E4OrPXjHLV6GMTFDLwbLgdq1Ra1G4RIuPymAWYzTekVGab/m54omthlbJPUTR
FwgAd+moYis8IoWuIdPqLax/rgTdeAZzlyMqEU9Dkk3D72ghZqI8D5fV8M0jiEXO
0Chq0FcW71J5+YFaWtuEviAnl7gbEb87wQOKvoheScpXXNwVxmF2u4mRKfcahJnH
dLw/gJQCBnhXjBFtqfwyhYIlnwmGMoMiNrrWJh2CyBa33oZ4X1RPSqkeifHhAyUd
vKvjiIzyeiE3ASRjRGjWEwKuFIYPueCeuZyrXpG115xRRm/xoFtWiVchPBZIx3or
vPtAJi/1+esXPdcyMdF9PyqU2tvmKkZQvXHphjIvxO0N6qBaoAouJTVYn00JaZDZ
B0dzv1ra9aJDxOQNDEvJMfWCvqyTtiGC2eUgt32S9Xj7iNxuSdd9lx7KvmevTOLe
wI+4P6S31js4FiJhvmrTNXuWLhAjB4rbNSdnYd2h+iWpIJ483yFUNdQGSmHdub6y
Et2+cLXbizKnVE1lDCWtlVOQb82EDpYwrKZVcL2gRdpvlTVfD4JXfSUE1LHlSigl
PDwWQGyF5oHrM1R/NE5yTr5eqsfm0bM6FE50Ijk9S3wctq2st5E/0LdSup/VYmis
a1fkNyT6dJrfoiHy+bjpc5PntH3dGPY71V08YB6aiZLvWmgY9qI6jwcnwuGEjXGV
gMAicoHW8dyF45HiG6gna7qw7mCbNvm4Rzn0EbBMOLUeCWgVBQ9axbMWYQeS4Bn3
R/FvgOK9LSqF763nR3X4fz46runbcRTmRuURH9/FrhGurK5c2rfO2Y9gr/aPiTpt
dZdzzbfFzexcRPyNoMlXRw6Sanz8yHVHX4K9bgSy0ozUrEtMwotjGnenTjJGhX18
ikJCe3KwSZtPQCrsTrLsow2MyZfNpFvOtsWB+kGOlfy0aV+tKcCruDtrFdu4J++J
Trbu/AZng023xqC1S+Y7koAP2iOqOQnMOOexijT1CRsAnM1PwW3FyOXOo2cFleRm
miwmuUHLOkgvJxpM7D+ymg4+pvRNpAGrnpcwySbrt4gBsrFjEQ/U0MJHlS4NFTR9
GnnGiGO9tyotrlJkGlpk13I87vyxg5/9M9tzT8mMnNcVzxOAOXWBmAzwi+lqglOw
FgDT2gfz4k2fi0cjOqEyLX6DMyA72dgPM5Gu4bL58vCad9vI3vOvqpcN26K1J3Yo
ErFe1FhjYw7O2rqw6ar81XKWxuZBhpKCi/EZxOdszif3sSlnb8w+/+qwHM6rCKsr
rEvjacM+8YB9+LGZgTSGx0L8K82H82WITeTF8efpt+y9xap0Ewb0KspTOej1fbs+
c3/famVQ66PRxDuhjtOmx8ws3AwRdOfIqpVxKuDTLzdj+TpHgWceDr8QzOtEcLgf
OywCC1brpy00v/C55ymfMW0ttzxWpT0Js1r917WkpUjCSyFEgPxY9TdxvIF+4iID
0xLYBhCVYcF2YXCP1sUKp567fNuxDQXDCudYTlB79O7YXtcCHheFmkfxAoVGTN5k
hSZ/IV3Ut6gc6id1BIQZCHsmi7NI8QhDjI/CowK+iE9HLSywBGdvc6U3loRdqG09
WSfb5APsR3YiiiQTRTShgpTOIUFTyktMQYR5pbp4pYz7228aujReFWySBXtP6mRg
gdQqSd+jp/ppOACP8bvZpOss30MQH6HH2sKJSvQxZuN7wjKI0yDdWGQ2HxZ1YM30
3Qm9iqDG1LKyrtnRu/Fprap6hCGctoxef3fQ7SrnjffI2mUhhpc2uPAivqUvdcd4
Es8sqWzXFnG3db1BhHXsTKbco2xAK/G1/G1YGCqmKi9mFRRMYE4AvFNYjOlzN3i2
NpPAmC8R7F4CXHMptzbiYPoL71m8IX5LTtS0eg9+5BKmFM6DoAV1kQuCvlKhvQZA
D7yKbRWXbNc0ck4ealk0c4SCNuwMa6aBVhmVfBdjSw3MmvRYa55I+AcFVMwFLPeO
NzQCdfiiw2bBKP/5KGXx60TjywGc4lcvkkwhmhlrpcEgS22DnCeuyO7i73DMEctJ
0sUXEC6EU2w6kt2j1xE1L6ydUcTEtbgoAW4wuMGnrGlD69Y1adYoZVMpaP7g45FF
Cr+ukTWzKPzDv0VXe81h2HmDSsVxfxFmVuARZzehX47+CiHKUXXUjOKiY8Phsw/X
InAqLVbGJqMSxJgsgTEnfacXoPYFxYrVsGq7N/eLIFfpEOHqS7C4Dblt/FNmCH4Y
+30inT442wJmjGhQXANklnsAXhJ8KEAenQzEAKocPtOP2ML+vZlg8+PKNiMEtkZ9
lKpVhTSgDQaMcjvjgnvP3o9qKyq7+4xmD2gG9tIxd/SJIDd4VtsqTbqdonapyF0D
SMB+V+1eHB+rvwjPg8JfvzYf+53tlbqJKcuR8A/fK9eM+p8GLPxI8bkB2kdRGzCX
1iqDVPzDWtLaJwjFwCUmFgiLi68HghTEXWqtqlYuqm+g+174D0u539N3tmlWgvXb
Vo+kpMJXs7ujBt/rnTWlC8GhLjSbO/7U78wdq/tZNLHlHIn20a9rmvmwoZZRaomn
wWc9LmuLUxO8DiXgyRQA0MFUcXLN6K1155qd4X4nBqCOaEPLtOYMLoH5rLXeGDyC
mpuXWlh31VxZztkA+PrfDfcvA0FezslZyUOZzajObnPs2SAqG/U5GCdlKVdgJ3GU
lEgAl3NX0UKQufLAIKCn6otfxtxe0sZomixJh8IrbKGZNmyqld0UuLExjbViZrn5
Y4fbTAVwCBwDdkLG8M2N+7QdmO6KmXKR+spfEbCDIzwYvKGIBjcvxQ6urj7au5kY
Wjt8s/pA16fQ2D3WgwYrKdrrGWA9tYGkXFjPvSpyBUYeK7vWFUmSXfIXcBisPfmk
bz0bzLOU+xtaVOWJ/kRhNZvtvcT29bJBx1JGp09OT+XRIaq43DlRGfUC0adZ+YXL
+kmfI6lcYdT5S/HDiI2d94pl0LqUdPyGOA9Z6+KVnK23NbQX1FYr1zn1YjR/el8j
yVCmnapwK8VQWpZvqoU26PAmh1R0KsN57sB4VPN8ydo9oB0+ypTpR+1xUUx78wwk
TboWaltlUtzgPGxORZQjeK09KeRcLAOT4DnaBDhIZlzXpuAYEZf6PEuJ5Cc+Zi5J
KJE/Y9MJ+sOxbFAn+GV71PkSHJz5dilcD0wRSkBdT0XXsFrmNpxFh31cu7ixABYK
lefLznnIxX61rovi05u2DjwCKfe0JwRKfk/yPYQNNFhtPvzeZN6gqB/giF+rM3UT
nnTbJpSaJNtcoEunDa6OCNXFpeuMxR3vbEQoJxzRCu4x34MI0KomcK0cd/hFxUrB
VwmGR2rrTdTvYi3mIL6GBWtedyPYgfhm6Ua5xjtRQ+A517Sy2dcz67NdnThDL4YV
+vLF5iakGe+FDINyx9S/Ot4f6J/1KJoGtvLl5ApWolCs9zeWyjgC/o1HX7cGgMzs
TstYyzN8Rk2XgoEJVJzPKLyZsLzuUZU+yyVw8IINKlEI0fGJZ1RefOPN6t9bGbd1
XPwueK9j7VtKMRqnwhuAxlilOh4Vjy8v4ZdNNER49dfUZA6I1lXXE2XM0UOCDsfQ
IGAnF3n6+VRVdCNkC6qLDKHA8QWPgFQvbeX97zRuWblvIrX1e+MyYswPpwbhXMHk
M9aWQMsSOJ6we+18E5L3Thrxlx/AKfBvFatDr7Tro5RmJPdbDwA5bY7rWVNoSe/A
nG0umBhlJNrOw4pFjAv1cX9cHT0Y0meKEx3kE7DOpaypNmnorFZGpJU8IlCzJxF2
gi/rsptQiUUllFGZFMzvwnHR0qKu4KQvo5o6aFLugbj8l3YX+IdO2CFgHe38OMVf
l9CLwb55mS37mWM/QldfZGjAR7uT8MyhQ1OqMyDL2T9ll3a0THv0uBGNZawI3Zr5
pohmNJlJv5SibRgoXCbDxkfG1Ojj4zCEQtIxPnFRvOdEUaezNHhNeO+Mfs7dX1zo
ccuLHIoK1MvXBhF1KbWqZ23JoDpfLTwM9yWlGrOb5A6B+6OqfVAMgvBbGxoYF/9d
td0+4YtR4G2TLifywSlCFJwFIZ6cseXRdQjMlX9Vru8p0gT+ONGiPOKlxip/oDSj
Pp2/qkeLQfGzi8zy+jJNHK6/P9DEw2TyuAPm813ZFyOpRlwuGedQsRTvfPZ8zZ61
zmBBnoECw7tTQm2VpEUbNfHBL3GkqvAPKHtD+XAJy18jJnUAXEuQsgLiO6nTC/oE
+c7aEY4SY8hmJRnQfmlcxJjzaRLFaYsnQMimTJs9byZBOpdmTy7hquSWM2AhLqcg
mngMJF86PoixlDNHnGCEC5laiET7ZuqOx9BbhgTAN8KyuF3NnYxT9IMsltkScYsE
ukvIvtmeGJkRDVjpALAhFeJPyqba24ynWuMjwkZ5CpOIRneV6g92sWAhE022w6dJ
I0DK6lFsAzvBMz4Qc3b62SybmGTOOCxMVmy03vme7URTtVB2syaFxFmENquyrXKK
7g7l7OKhTtup91lMBdquenz5QW10S27JwNLBlqTGysWmD97eKFw8u4kZxwJEofiI
mYiPmrjoKEVzIUdqPNDQrNvcqBLCBy+pTbKplu+7gaPOY1aQYMpeNrb2nRKLUu/n
S7SIA8llHlRzKP6vdYPthDBzMHz5apuXA3RPSOjLfKK6/FOdZ39TLB+KawkweEs1
Ia1aaBAvLhdt2wEJIFS6bq5tTUb/IhtEUTdLTSDKqycc88Hxx9uWlY3OhtYLGBhd
VR4yyAfXs/HT2cL5OjMxqHsejEJXhOfdKGHKgKci+p8bekGUUpYwdYVhVfs7MCn2
Ej6GGjPOyC76LPahK5OpEUXtP2CGtVXaRLNiM9y2hYf1LfYZPwSkBRDTHM9wyzng
Cn+0fzBC7+Ob43j9JdIpbb7YHZoeKh9+rpkb8huzZ7e8XcFdC1h1SZZs2BfuQFJu
sdTfHjo45Ot6zS9M9fC6+1de+zczlCNCC6fiHzivB02VKH0rqiA4zpyxoflFh9BN
2apMTak8jJ6FEi7EFwBH89p0ZPy/u/+Gjc5NDQrHgcFhxiwOSqTNS6Sxy2XcsLv2
vHLRUjdLyNd+9TLiqBEzevLuKF346b62MzpW6OtwXB8GHLyDJ3jzW1hJHVqulTHu
Ocw65HL1DlgNFjivmpMIXBHi6vUwVFhla1aaDdVoBEuMSKyXqxvr8Zht2b/8aqnA
zUhONQDiWhj3lZ0MvvdVhdq1ddu2MMJofE9LZZiGmESah97rIgkI/gFY8wDM6XBv
X3lhfsq4ptXPgx8ka0Me/XEWTGNHyn5byiHRq6jAZkXeJO6pHDEEhBLsJc63wZPQ
Nju6UuGBETBgqAPrcOeffydHbs0O7eCmp0PTaeG+QMT1uwowV3mKT+0T0+WrphY1
QQufWkk5qEy97ufjYUGeiuFEU/qvYU14Z9jr96Mnm2CdPZ8Hwzh7489CaL/AbDdg
UxsTa7XvkrqlHPksLCpyH9edHnUQPriNsGFXXvuFPugmy2mWTyR/pBMV+LTSSbww
xungHpnoaqYKzqDJwAAvGaMR8TpTPA/NEWAryGDIMB+H62uyJlzzPsLM0Zhrc3sF
qYOlEjRNudypD/q7QrUupOmbseGrK4NZwZlP5Xktj49XDct+y94H7FbkJEehbNcU
QfQgkMb6l/SFMI9SR6kMmzoiXG3QcrLIn9BiSj9XXWfTMqGJKAU3Oky50mutjIo3
Z1r5t+cu8owBZPKRGhDyG19OHT4FQ5NJIGXHiEMj5H9TFO0ZHeZ22pqrgjJU4Z5u
R3nO6cDRiHOioY664jDP0tBulWRKYo4SmBN81i8TxnPMtyuLF9VbuOcigds6Ubve
uPnd182vW2At70HXWFN1LZsE72gRMI5LDljajyz5rxsmYY0udzaxouAphqwjzbjo
DhxXajQ5fx8A8ZpYYWfNIkwmr1MJMdIr+dXxEFKMftXvYhML2w3q1e2vBOSYRxpD
N2ZFUlBxXgYcV/sWj9Qd1CgJdp4M2ulavO4zBFbPoVRrTK3ZfaPi7/cOrUqmIQ+7
5hpogItSBbbJ1Ne0weXuNtoBU3gq08Q+/5WDhrEE7nRfRZQxa43nLyBnEF6Vknyq
s8oPOddu8ITZJ5toQw8MSMc2l+/TrE0FC2KbifTVz/vV3w4I2j3yLrxMPolxE1nn
HNZBxeaDVOfqc864nrDToK/0xfAUct70Qy3bzYDr90Eh7Hqk/VkBapBiQU+qhvJW
vBGxxXM6pxBbnVNU3D6H5YQ0kIdsmWoj7YuEijpy5Mm0q5I32M/n70FezPK766Vw
6MQCSJcB7zOIGGSjAk4OKXjuNfpZxKF1W5wj/YkFVOLkLc/+VILHZFd36N7k+NGr
L5Fpc3Dn7RBblrilDlJ+cqk7xMXMBugvD7/bcprkEsSm3dd43DOMDFekL/o6eFs2
UQAhkgdH/wkAka4ISlgr8PYGmjwcjHK6kAnCSTAoG2ebxz7hLpO6K0YxygcPCAUn
QNvSYjKPJDJEmgk4YHVoQEAMUJTxxkNzZ047+wWWHiHJD47/uLaeFQKkqA0VncuU
gYDzfJVrVAfYIXKiC/DUBPw7IFfXmYOT3bOfHgXkEwpY7v0CzqCk1N7fDDZAbzcG
lynamj4flR83TGX6GqacHknmXA+tBEtIH5itxUDeYtfDEYKRZXZIJj8qHCqQf0EN
Mwn6f32Z3FZTKPzwzoMw+1BYFQ5P+hIx/1szgog6dHRyH7HXkDfMPKVHuuALBIGM
BdMxvA0BGG8UQGFTcLyMGDhfiHlruHQbLKfJZRv9Tu25RsPQJXMJpu4zEd+8dEx3
p/xrvKsksgy30sCbkecUeGSO0HxrmG94Fts9axoqdrqITfO0E+rwH75eaCMC13hO
gvmfcX8GqMBgnS53dBKP15kBQf2B08mw+qat335wdg3jgNuZ4m3bGPwtLz4oNZVS
kvftv4p9TFKZb79gn7/rBc05tcXqYjlQtPtvLvYVMuq6ANyZLbyg28uoX1tZnksA
CpWfdjJo3WoeWQemX5fjchrg2RLM4VHjzet2xWo3Cqr2Yl6JEiXegY/9RcQq2TUm
++/NXA5b5vhtywwOOYnC/R4koOCqzG59n77aWMmg0naRwvIRY+JsuMPjhrHB/V1R
PZsEFxlTQYyz93vWSpCxIhyEybyeX/FdEJrexaiJtTUMZ7OHySr5RWoswhUTK+4f
EDGZ3S+574QoALqQWDJT0IQj60Y4IIbvSKIwhz8W5+yNCsOENlS9TSgO7nnOnNdf
8i+sOnraYrWhwSbTM7jg+mZy8EXOXBcqv8p57rVNknCnvGq0Vdv5w0jgkRTpejPV
W7Yo2xEcjY2y4c5NskcD6UVp9ov0+veN3AtGHF7caItgDFDgs3vbmiiAMj4oeU7q
vpnQmeMMyrDQkZmNeogF5TFuitUUOAX0xikgyIIvqZfDDImIkqt8sbqfGazsycqb
e2N8kEeJhzSaZjQUCxMn8bt7aKHhLl1owhBOPwB5jza0/8vFtQ+bhnTCglgHrP2O
t1BS+IYu5rVTorzuB77Dk54SZIAOrwhjUoFj6WWw00XU/5GOMWOSUf+aI9hdn8CE
P4yZ+1a6nZ/fQO9jc+VbDqAKbEL0eKlY7f/pEOdFwDNZnKC6VD+XD0jdxRa3gDaC
1Zl9DkyXk95gDqFU1E+frr9Cmica+dhI2TYpMiKyHSDdWiPIrCus0K7/u7/NTQ6E
5xIqkqXiEcHILD69pxFpPj8/BM2H2zKg0XRbf61oCXtGwTGObsYUh23+rUPZNI7c
hLM4sf3U85Cb188l6xJv0IRxGADUwMQQkfAQf43xj+BZlSX6DbkHYFEbhRWjBmkG
3LyClU2v9Up/124zbGTa8mhNlLjVTJbzA/3TkJEI0KuKXuHvgLYrPCDJqbNxLf0c
9VEmLquJQFCUYb/YP8jfFiVlXv1VGT8CE86ZcesGzjhu/Z9mtafk6iuixqAeAvBR
SmuBvGui74g3Ey1O+cyTWyNmuqPgS4DadPhMKyy9m4+L+9iKWEUtsOYMVOxVj3UB
Jyi/BaqW/BrIgrP+W0xbLtWcQ/kxHfKd3M9CxmnbbGAJbeje9LNVrH8uZJ4k6Awq
ojm6Ql7XpWlejvOeWCGnCcTCn3EclMXLbRWHWcLJsIfe1CmAvjVjUt/N6bSR6Y30
/5KlE0OZZevk25p+G4Pjh/9GW6/0bss4z/tw5X5v0JqRu0fhpwFfKm0xHxjEjThd
ahXAWR0KvQbPEsNFzgaJqGKy/hm6V7Pv50t+dfhfzSZhb4NGWXMOdUgFFJIk+a6Z
8XbIq1UMf/kXeiEuD2irPuoq0t7SC6QqecR5ATkGAgSRxt/SipnNdj5jIKL1mWUW
M0nsJN2Ci1TgWEFbb8Pn4acJxWQUOQPRaQYksRr9gN08oX2LO75L6qONoHZxfY+W
muASZycyVBOoMLASj8r+yCeN/3H8Ow75xhwsGz37BCkxO6icGHsYn5kQOPLo4dq2
DB32HGTM1qOcPPhMLZpDaNGB1BN/IA9z+UTmqmaFUfcJh/Wh76ayzSBNjWXdBusJ
yBm9WDpYvC29mn6pzuXSEMRyWUWpY1LNJdus/hpWD1eHpbPJVKPSGcc+9UlcIZop
kCShlHCj2S2bklZCmUIHo+e80vfd1tskFPGg8WLfvvdxuE16lzRXbVlnYQu+fuG2
dGPRf6Xr1M7W2JYUTgsVXD4b1aMzM9TRl9hTewwJv1cPboNUzGyW2muMjwHadMXm
CT4IQSgDWIoIEXik9lL9QoqrLlwB9v6I/FiPU7NPKtYXHVFlsb+vWlYbTylRWz41
8RnxauY7oj8ohP+Je972867hEJ21mXHHasCvOHHluj6lzZA20csN1Z+ZkuuNvJVE
o/bQcKgSxC12JISg+AsMoyNjV6Fc7LMauSZZ+VuMOfSvbXh2ayUFdZfQFZ4PYExh
cY9hDa43RmWvJfqpJAycQ1IRKJqzMtPoH1AdMGzwynboc8b9A5qjdBohyChH5IHC
wmvBYOruTHusyhk1OuGWZur66QBl8zTLRbQ8cXv8fRKN8NFY7+j10o/EI2j0CkTf
4+o1Vt8YYGvYqKiquFB+G+pqGza1dYpkv0C8ur7oAWVUFxOf5ForR/f3eYuIKdg8
d92AZzqS9WnMmmT67wA3XXgdx5nFHusIjNOKED2UNja/OhN2OVPNIbiBaAbpqmSB
7oikVpA88aAka/H27u3J8UUnd45TzVHIJrvnfLDFjXARs4PLhrKw9gvGrmdQTgjC
Hx9k1u3WgZCJQV/T6PPZJa/7wJkLIl+cdKKF+b+r6peiYiIMESkMOG66GUIGU80q
oWL6Odpa5vZRWw25g5vqwwAl0oiWDfdL72C45ZdHntDxCcEggiThgY0gXmSO6J2r
ewfNFnlx8sH24KyNc2HoXNNQAhnQKAvtvXRVIMpb06qmUS7YX3XwYrBo2zOAHhJk
FvU2NFrVKPQdCCE2MTT6UaACs4sOBB92tvW8xuXAMFcwq0z6f5B+zJBjvTjHaVCA
40pCxEZGVXKnk8By0Da2HccdiK9czYCemVU3Ubpj+4PZ9zWc2uSpOX48ba0xb/Vt
Qzz+9bUplQ8UrV+DPwaHYNL+I9LEuv1NDBGpwJH7pog5NvBBGxQYOls5vMTYS6e/
yUTwDLPVIbOZCouKGWRnu9xLVs4Sd5IF/zF/a6HjSbxzUU+T5PB8OKpGsFWwSCjp
EXEdOxA2of6MEGUztvXa5/7x7iSn8OYZYXRnSqL4/LggA+yQylEzo+DEEmTLc/k+
xf7+P3ne6nmcG7yc52WS/oL8aMZVLygDJmjA3jN3FSVvjKqhpzL5lmUrAVI5otsF
iy7vDY7EAtmgO0D+xzdd0vyujln3+lnjh1zCcaOvP7/xYUL2warfS4ahQLMEwose
AtuuphOqyS+CmeiSDBQ9o6+kGm3kCfU083Qi32D+FR4cYoTb4JQPxyKv3m0kyc7X
QaEnfLHDjw14wSeOuClIirerpUW3cUB9tUog49YuYojdiF21Wubwb5pGcLQKFnd4
HCKB8U3Qy8ysgzsd/abIQqqHYU914whqF1CeOLIO7AwSBgy4dxIE/BKyi22LCa04
D2lXk9iyrr0pVgB6vL84cjq83DW1waX2InRaYizf9Psg0XT9UFOndPcaD0S0aiOM
aWVlTF2p7In2zbSXT3OXSigxGGBLLojnzyYidC4shY1tK89tRzTzgb1UsabyzI07
LnZb6skWP93k9I9EQfuc90TpMpLvIsevHHkm18H2tZkJT2nqIK/Yyp2qi/blWZOv
ICGnimjeViFmwhsjbS8BW7r6cP0F9L4I/emXrHXSviPafVrk93Fn5Ma4yKx5B/V4
Z6NK+NPtY2QpeKJNQH67Mu+SgyopMdMas5A2ZmpJc6YSFilRDvjCGm6F5+M4WRQ4
RIzOYwNV3hWBhIp8iGXTnAlXcQ37PyGAapYOdToo4MA3kNQFNZFIOTbC+rwGD5Wx
aIC0lM6qdztP/edJ32O2N4vhiHSIU5PzhINVo11U9pRAhzhHJeT22qx0It2rN4xC
2eFlpwJ9A71Vq+xPEZLcz7ZD0MrnrMWP330lU8nMgJc2xWI4Patr5cfoVNUVLG8J
Za2rhIeXGrhpUj2ntRpjoqTb30CptchdPDQ+sJuTeh6R75tUT5EbkvYqQ+/hfQIE
dBeNNe1w6vgiCaYZVQfhlSmJA3+D37op3hE6UeKxtOBHUvXFDSRRVFU6qkBHOQW9
jEN89tPOXhRQ7kkfGlzD6HBidxbdbxuq5qNunu6g04fab3+nUEK95aYLZxz7TQou
sAfAOKZhYr/beFTHFiNTOnPfru8Xa0yKHZ61csPcusA1HvNTb2x+CsRI0NcQ+6Ar
Yf9gGxR9NbWJbrjWe4DOSzlKvkQy/voZ5K8emFY67hYLRx2O2bL76OjnN1lzK3DY
wUwlj36Q7ByYfr5170niJ8veyPRRv3QpX+ETFaATe5zdU/WWThui3i/b+IIdTJ4i
0CR0g3iJh/ZjDNqHn3iE7buuRdHdk4faUrYZpl4h7gjdumtUQ9nPfpZnVPp9jBvp
W8mP8G/JKxcdRUgS3bUW/ybiNBgM72oJB+5iP31baZvpPMf9FdX4yqD2W3exlnPI
5v3+bj2xoPuq/vfXqqhiD9F0QJtBDqwJFe1EeomrjDtVWlDcwSiWL+KU+PaVV8ye
Hzt3WfbshI0mvNKmuHbtrUy2M/z53Gt5cJXKay50c7teJtTl/ZEwB+Smvzfa17CL
c/wMr1ItxQlvG1DKx4x+dap6VwgkSsZTXrHaKB8NRP5W/a14NxygJhrEPNo9BBEP
hGZaZiarKSfiBiIDjbh3QO+6sX9uddeLePcruAEV0neKjf3ayCFRSk1n0AzihvKl
16SDaagBHw9CjNxKqwEyixFb65MmYy7yCgUP+278LWqNGe7RR1lP0J8t7I8ctPm4
SqbLadgCFpcIY0Abkv90EETZv6oUXc2/w8HFQycCQ7ln24B6OhMKB6WiO1HU4/jX
r8YTCFmyYsA6QASY0Z+bmXC0t8G45dnxjlNukgOphz+KpxVZ3tosOKXZahUSX9Pt
XGBTK1TYRrTNl3FUNPaxjiRAuhATnLs9FcwmjkMBC0b+4yfjxdr7WXyLrGHoqEwU
05sA7/HSBOszt2X2Uq89yeDLXmCvGX23PiBSf0vO8Rr60xcxGjjNBJL47qKoNrJ8
1NBNJmrAIGN0Ehz9m3UdEZ8QeJpkTOz0/VFmUiH+ERHhgFAokTSDyx2voMnSnxEP
2zwW2DsZQ/tulql3+PpTmwBQORlZ/N2IsJ6X8qamVe5rbeWiI8Ih2Tfg7mzuEjEc
/qbpXmLYqO/sabXcq93xW1VSGyyznLOHLZYuP7LRPrnexbsLvt3ImQdhkNC3rJo7
0gpIIpmeHOjIVV8Oz7sB9ISwp22ztU4RFPOAVRCe3rSBwRXoOYk5btt73kvF5uwS
rQkaawIUGFOI3r0r3caqVKLf9QT/ofI7WjZItCCM6BEr4vmcL4ZkKNf8I1dx6kfz
5M8kVYVsf3uvHyBPcXKGoodN+Q9KfX9uRs0IpyVqrU/Z4X5RHvnNrAM2C+1CaKtT
ShurnsQvivKVT/YMiiK/FqKNc7uGPrBDuzSWGs/uo5h8+mOizEL23hMOJxHjACAu
nVx4QbXGC1nMD9wpKcRu+iDWPnpkjkY+QPjQK9KLe+3Fjr270lzbToYxXZ5t1I9Q
sgecAtUF3PHPVwIi9SqikffCFfb0Wz5AtAQQ/N7PMNp/K6Tj3Vta3kuU6tKqsWrs
pwJK2VdRg2oZslUsgjlk841/LWPEhAtkp5g2Nmyk18PmF2RhUjZRwTSzPl6iV/jD
gKF/mD6M7Z1Mi0yYHM8+PFAlSsK2c0XDgL8tjFTMcHK88yYLt8nP3AfTmnBgXqE2
VVKLp4w/mKcBCpzFSYX4GyaNhPsFd5gfFJYtL6JciaKnkwpbKFDA6wF41445nDO6
2jn2TjBPvhTv2YGRxRPJB90MvAqUgNoAjDWCj4Dwr+1zSPkk9CXevnk2bC5XRNTQ
mwcGjPqTOOgCLdg9U3mt62P7y2Ov5jaE7VihvplzM2E4l2viFans0qssxJc71lI9
RiXyMu9WDnxdqctZh4ty524yKb4MzO+s7LgFVxIF63K4dzh/BiJ6v7+A4H8LRN74
cKwBwbD/V19Hv7JqYyOuCTXFZUGNSqQFK/kuijSdQZ6LtG4by4n1qgk7J0ijymVA
uK9KPWauYpo1MamfHXSnD8t1wa/xTBm9X9KscRJkbjxTC3jNuy+opgVDxbog/nNz
aXDpujA+gqZIVqq5BCAcKZigtxTlQvbfKPfKjJzOUQdI1Xp26kO3ikVQ81sEBYEY
HTwVunK5Yjejks9Wmm6XnNvLVYu08QxvyXEqbU0wbS4vV+q8QCzwaXyn46kKhFeg
aXXxefyEb/Odr2qiNGtOvRya3FOeBRWS0VzDiBE/hre3cGJ3xt0uEh7l5NOHkWNN
w2DiO8Wi0DiHv+rrq8ZxdFuWI5T50cXQ0RtQouhj5kIUdksk2OOFg+/m8DBi9DKX
i8u1N802CFL0nEpQ0YkAd5nGTEHludTT3kuHu020Gfk4IWjK0+/sb7CarTR8jGwS
Aq8Sh6RzEldPQ9XAHojpDd61eWlBhVGNku4jxDDR/xoHQoYRR5ldHAO5IyrBwlTX
08XkmfbZKZz70SRxwhGOxQzmkm8AZKfvsNaUB3rPeMqMfRi2DDgVT6fnC3Z4QmiQ
bl1svotXAjpFeXXaMJIWrZpWgUAZkW0aHEcsY/u8o2eWHdpRVKwsooycHdvtILl3
oslSY/5fepIJ35kPErCHdhScg5dSLztJWUmZ527AJE5T0eMXOEqcBxU4kXb1rjwF
UGGYu3JkGc7pV9Xmnt/Xoxbl3/Di6t7smJoU4b0XwSriel153QkJTvmSbZP/nqoY
MY/5h4c6r2EyCSquRjcKhC6QpUI5FtDQ6XC1Re1ki4Isn9eSGdsW+gslowNocX0W
Bf40RoeeBHai4Tfr74Uwg1U8ma4jwwg6EyWlhoF5ptGaoR+VDe+EjubkHF88UeP7
/aPeRgL4lO+oCLVDjJ5p31sYFU09IhjSvphtomUYT3ig29pJjMLWpQv1akdeaQ4s
ix248t+1uT8PcYhTy0Q8KOZmaUFDRzo48fSYq4e/4TR0FqucFMhdzSL2Y5v5V2qO
orHqa9bdzpVTwvx/CAd94NaufaFckDy7GEcI6sTxaF2k7H2BIn72MdnABKoWeqlm
U9lVoMuz98wujGEZ0L/3XLicR9NQKp77VRQXOKTzDZWp6u7OxAwenTj5ica00c1R
JUWhDetddpseRZPvsC/DOBG67cznq+XHi77K1ShATU0raaZUMbIfoTMY29HkKyoU
v2dTQ+bv4MbtxTgjbtZEpER9xl1Q/3aTwQtYtFoS2QWTQXhluyVzsqb/ZQXoiobm
CdiykgCipFkhboXH9xRV3LgX4M2Am9T1dIyvZy/tkbdXcPgUDu4B453EmNVHf+f/
A65Gv1XLVDLJ4Ym8hPOH2mfLGK1wE9kzrc99vKs0DGcycUyH89iM20nvm7w+7yFe
CrRJgBpeHWWilpbxTtyan/iGNI2sNvR019p4sGSSV/4o0dVkpklrOstLtzut9YMc
TZfIK8VPNx6b+BSyQYtqPnj5mMymIobf4CmPHr9MFEFKOiejZt2UjUkEKWV3Xyan
71h79ay+aciTRNfOOJj3NFX+Ra8W98fqskF9/Igyk/6ra2n7RcAWKT1VVtXeDTof
Wxe27tTRVoT7N+d56Ig9MDnVpQpWtIIG1N5QHxTeuamHxsDK8rcD9xnWsUbMumWs
VJkvWKriDAAKJEgcuZfvse/641cxUuICRjVwr7I8qNl++IH/MnmOWqn2bHNabVhn
Qxiyz30wMHseELNpCBSq58GuISU2dyl2y9CuOaFbggGuvN1RPMB0uG4sswqD6oiw
2ChgqPhuNQZhCGTBCXdPB70zQT1Ob57XCY1gth3Ai91w89+5xjCMb+6rbhsHr4Ux
+lDnK3zuRCB9bXHtypBsq/0jOHMLPNbGzxgvHq11RxUDScRWAoze5JoMAB7yzxmg
tyfAs0CGdOvcn7/RgU86Uk6BCZZhYdn9dNuGjDxCCCXLJMG6e6JcG36K2+HelVVP
jISZqLUHRDcVOcuMU3PXkYIDTEK/7SPaRu9gPcD033YfFnoNP919dnEGl/CxGNpo
+qZgVMGRkpoelnpLh2DAwKSXtXta+2+Ti5xjLiln74fFD3jBa0JgcAMwF1RKjFaP
Q13TyWqxarSRsi8512t7Zf729DILmwUIbsvrv6TjIsNIWxuLzZQbTH8HdVThklK8
Al0uMdS1sTHi7O6776FFB5sL7gYbn+iG+EQSfs5TGoBBtBcg1Rio1WAAuLqPRmGX
Inf3+wW/9Teei4VLkhyZie6tmJUEs64ixLjv8olk18we4cmudewMr6mnUdhRhTyu
4+0LC8tAgVbTCdUi0LUgZwnet1phaOvRqSwPX9oAktrC0i/b9BKkIq9kCtiqiQBe
ZeCr3UN1Z47Q9AMhpwJP9EN99fHWBnJkzq0IB9THIgwqZNdUCqehFkXkr4M/vLN3
XkBFHCUCrohGoQW+VCH/ENiZ7bNZNgIvptyWMofGaEyVugsT/xWDrmgb1YTAbB7Y
AmUKHGmbHe8SPIUUErpiq9mbMw82FG3W1cG/o65fVjR3D/3PnSM+pUnMr4wcu+fc
g1ew83gpTcbBxWQHPk6sqPephU3ZJbF48fPcX4Jxv6JTInMyuTiWaSDs2f84KNJU
K6nZn9G7DQ2lftJJgKVoUl3jg4bOq+t53+KpZlVxe8Ww4EPi4jdOK+9OP8d37uP6
KTpRA5oVn9OULy991y40ng3Uw8VImUKwIEaUrn+C/ZVmZaHpMbA8CXrK+uONauc0
OOV+o+NppxkLrecWB8Ju9CYBC6bmwVP64B8HERKJ6W9Z/J22dfbgsh81TKWrLAQ3
7YKpYJNRtPr6a+pe1YsD/ejmS84cv4st6eDectwM2kxzZ5ZfaxxfG/zvxvNc+ti+
vfz8io2rvBIurFatizsxfGyw+G9BGDy3J3E08oBE0AFs7P1UPXgFprEBU/oOovaS
GzrSvQTFIRzYvFWFt/JVMjedq2+cribLKWvDnJLq08PbIES6wAqBGynj3ergggw9
SCvvlF7T5ZGUCRGxslO2axeppZKahRIBlBlJgZRLXlfVCOrJtvadXpOOfRkkxXE/
2OqQJwMvKYJSzaZq1OkQ4dyqR/dVVDzjpmAEmAO70lcMUpy+u3DrOhJTNNM2IFTW
UDcocJli4lEMMYdKnRuDFZ/XOHmxyceg19Dv8O51EWNKeLaspUwdAwmjuf4i/KMj
cCAIauQqv3v7gXnPwsnT0hGbUyBtvQhjmzha1DJXNczqUrIVLVBRpFFzV3qJcHlJ
mAbiOOIGgFMxd+Ut8o8pqFnWoRAsymFAPt3NLtauusQA3VUDKMzivN6vZtRXX4Tk
WIYNm0q00RQjmV5FKeD+xqHVZZlqqIvsnutfLJnlDvspqdicpMBfNu3IjCmfRBMZ
UD4zv9nwNSHDD0yV3UiYcHZKlh4aGYUkR01pd2joOPpfGlEZlDJUFUIC6wxQWQ4P
UvZjfzprpb4JWQBs+98iUWXay1bMYc+GDcY4WmlFDoSpaysLEAGecA1/XkiZAGMg
uldJyZpJJCvRL6suY8t1xxXo8lZmMckbFOw/kBmFwsST6nDe9UZ2TXjQ5AYreRUW
r3ULF0mSt3kYJv43/Rv5TLI6I8Gwg+I3jAO+TzkAqqKnIfnqXWZC5wZ+8g8CKN3a
Udgyp7f2s51i+KdwAo9DTdfpYTjNHr3IFxS3BLBv6xM7Mw35uUJ/iGUJhS6YLj2N
+valURm+aaWZ1HOXyq84m4DqVVuuBzVcx8iZwJOs+0plbA/rDWBIog6aSgqzCidi
VBkjUCvNeibfyEF3xptfPpoRoedDYMJz8c27kBJJj/C/JcI8XQWE16oQdUQoREr7
wugiKRzs/QJc99/ZKofR10iAPGTIB3uxJ9xeu6DRFLOTDFVxa1YUrSTYqD0/5Pat
KBgQ18pdxBGdHYQ0lkyQKx/bERNbPn2uZMco3/lBqkV1ZC52obDXaCoOxXoL1ep4
r/IVujb7N+R1HNBZXQZUgGa0BGJTBL9UIsKBni6DHuT2HZBGGfB6JHPsclMA6MBu
p6eehvb5upQy61DIuwuLq+T+QopMyx6LYzWIK79XMO9svoXyu/OAAz+eYZpWbuiX
cMeRRWXRTi2V6jBXtoI8dUrROiWrdDuJhUZWhF13U1s2Js5V6zRCqxkEomHayIEa
FqPbiX29sv1xSPbah32GkOr2pO2ifZTgQkP/UTc9J2C/TaNDWqBaxLn0sDMB8vad
SZdhg0WB2Ax4uNHqS32UImOM/e2G6zT/sASgxJg2n2se/kvFYbLyIwpPVU9sU5fd
rivhoU2n+onjMquQK1+Dv9en7CP9QWSpTqsd0apLBLG2vqqi/Z+zULbdN76gh8SG
l/mlhnvgjbi34G0h9Aj6C8UVS/LReJSJbhAXApJykWyn1BDeSJdC8LP/l7ILGlxR
X3xt2pMcJpfpZxZcRK4exCpQ1GlBDwoCpCAJ/fQA2ekIDwfXavM/54E1yOCRYtAV
Q0O7xLyOwtcG2acywFonlPpc83Uju/sK39HOuCpzvbkR7Qkau64J4uOxy2Qhvz22
vgxjKUEtEh1kF93Hlys5s0e96o5NgZfQxdFfoXqkGUOyMYJuuv7cYL0uwX6P/mnT
bwa4/aGvGYaxmG7qiZH7gpgxWiOEAeQCUKwRLXkcyJM7eud7+3hz2bcOH64eWvu8
omYs8sMB2qahq2eylVOeKBx6SfKfNqg5phN88nbpybou0VyJT3LQBnZNPvtLciA7
62hSlIrMeOvjoy+DqAi9y1q4EKJfWbllMIBK1D2g77N3SWKg/t3SoIWoTEXo9Dzg
4yNRXKIVwq6gZ/oL3QOXAa1zYHwu7wRX5gJExLoX9f4+P3W5r1vHIgRG0yILwEgX
5YxdG6mh/2e8LAupZUZcVb3VGUNRyKves6tmDq1QSrTIK5nlIHzHGZour//3nyjL
dosLL/RL+6pxffcsH8i0LzPcQWJMRW8eW6S0eD9+84ja+CyD+9zki2dzro1OCGVa
Kq/7Y7O/ShdkwpfrAcN1BixX6ar4n/4n5YF+MVYdfySKhkH73Hu+PjlZbiqE0ZLX
shjyjvHOxic4MUtlhCf3T62qq7Gq6UhVFTK99kaeqoBhQoQhRBDVQE2jTxyPeIQQ
RGVba/byjQy1wtZnx5qE1Og+NRrJwlaIRbtBpYPKFiLSsXWoO5X3rocFJA7EyZO/
mYFm1IxPfsT/e9bkmwnDTkTilIG4Apc0HJ6FOcGgRYBtCaDfkphnBIdh6VHtjH6X
Pm4NJffLe0Qz/5N9Xa5n780T4KBFcHuSrsfeKyCw7oC5FBZenUAH2+0QmAa+zhMf
ZjVoERX9KmqSy7BAnPLQ9B8uIy849fC5s3/eU50j2Z3P/FKUFX1/e+/EJSUn4VR6
QGO5ijCJCwCGYpuDtU8n4dzUJIv7ns1VFIIx2h4WD0vgPnZ5AXKmvjpggtfTwDLU
cv/mbAzK2esVmIiUUVETdhi1RMj8mWIfUEauppXuw2An4XYOP/jp6qugct8pegRo
Z+P+2Nx2sevcOUwpvlDSjdut+y4whJThs12eiCEnMAcK5nX20Pnj0PM5+ARlDa4s
EA2k5HTExkwOTkkr2YyhBMZgrUlWDCuzZrOTryOejv2SXa1g3+9tnR4taNurvHC3
E7pqWsavLeMrRLYA19IyYSnpf+FHLaJUaG46l0dll0233O2E2nVuc/0N4febSnUr
xaHCAcuMbLxlwEARD1qILlxxLHha78hf6l5iN5pEaXEmFLUvk38vRlzS3Ti1sVgC
yHSWzlb2jITDe0N9twZddlmeiT1ZImsDQzbPNHGrOk1RuZY2Rk9/T59sx3dXESPj
l95uPQFXrpQX1te0e3xmNDMCG8wiUn3jgrKcf5eaxRDdfZ9klq3qguXXqtc1mRRF
UvTeHOOjhDyN+nB7D0uFsBnRiTrj+cYj73RURFOv2cIb2VCVjMH0bGW/RqbJILDG
BN71/dZzIzehZqx7BYffImhTeQ9+j8Av5EOgUb9E5poVf4My1OEfvGva80O8C8bI
qZNY8TPswUGuWGVVS1z+Kdjt/GgcqHuqO9r1hA+llc5bBPVB2sU8+LAVtkIO3tiz
yNKoGZPbStAbW1r9t0Wu7lRzMvk48UnvxDVHDWrhXAqjfqhtfmRgxJrDh6gpn+In
As3tth+lXBvv+rZLr17MDjb3lTku/TvGTZ+y31r/KKcipSS8ah2JmRERthI73GQV
uK+ZMOaTISIJEpEiBtHVjhoQI3MVvxpPwzJekXWbI5DPmiOSQo6GohjJoRc6CUWP
RUH/NHe35hRLJ+Adoy++zxTZ4qtvT7NvRQ81q4RviXAlCMVZsBCS7E45raMCoqXM
phXjs64M1BbvRtMgPFS4oGSQBfgRX4MhrLwkIQUX5YP6SZv7AXfOEbOHrEQwheCX
xZPO+n3Fb6Gxzr767mRhF+6LeugtJwQQ8u1TSesxykiC9cY9QtuWZ5Oj8XMLPjKe
Hlvw/Fkgx3g40rRoQk4MHUA9+aBaprLDuB9sbyOODPtLV9GnBrGrE8kCLKw6fpUT
2rSPXu+Ven1SsyiGE4bmY9qCBgAxkNZF5bh/M6ilpPelLqA0sceU2BdQx4T5RB3j
b/rfMviQoyMycoOH6VVTXrj78IkfHIlVNVyGjF73NKE2xq8yMMtYLUEz/A8c11hU
s6YuhydKsyWC26uHkMfNnJtWrV01ZSsanx5wgZ3IlrwZ+u5VI3C2XNODts3t6LB0
0ctjnI0/9p/KSJaZmUHuMJg7/0mjhnbn0qwui+Ux3I377Bi4ai2TFf9ar/C5+y9s
CuTVZBEfyvIi//6QIk4McVBiNgtQ3QvJnED4qSFrPnrgcSbgqXMdhmmZ0A9+CREQ
Fm7wRSg2BYFpnb9FELhVTNzFO2E7mpC0GP1VLK5JD/exy/jIKaVFLalFmER2xC8r
V4/oYX0Vcqs+n45ZdccrRMLj4+FK2D7asHe8r6UwfaLDpGEClNb9k3Fl11GoWihN
oRa7g33ATLrYggdyv5JpOkaGYuinFMfivyk9hB2lpA3iBfcLgJ4tY5u3oKxropt4
XpbQab927bNGf4dNzg3k8o2pI+oaTukrBe/Sw/UtZ0isElEsAsQ53d7CJO33zwmt
q4Axc15iXW1XnuEKbEI05FoI5vohLfwa0XR0eJM3hlI/YnVak1CznDHI0c17/Xow
NWdC5Eoajf5sd9T1Ifs+YsB5yUu7GG7qXpZRrnNs5D8QKFt1UsMSG5GGfPL+YL59
PSMmKBpdSgeos2afvdP5gnvkvsTrLdh0/rtKQONq4WNbOfOhCLSOPQo6WhaP6Fy/
d6V/XRfzAreZlKe54uOMDkXJbsKXXqMh3syhQdWbPole9ruhPNa8RBZ8mvY3aAgm
ODtSKBGDsKXjYRVQIe8n9BNGPxZ5O3mvXVaRSptEK76TW273eEF1jZGuvS8iKHjA
YC7z7VngjfHaLGCCCKMKOuHSSlKhqxJjlFuoNPK+x1rGu9rX5dLyKVsDmm3tAc8s
FLWIej0/BG+etDFJdRsgYiNpht22YUe2ccf4/JLTqKf0ByEjjGLYHl81/yVx+mbl
B1L+nMjwVSUlWLLfOCblbasw1ONAFhJKjxG7ujgHuEZ3nUS/3dX1TyfEkS0Wg0V6
VSO0R9XNY8c3lpXWLA8LLkY61BPKhRtiecTRorKNzuBUDr48mfEfdp/nOHvMkQvx
ih9CMu4b92fe4FgzZq/n9B4sX6o25UH6r77wdOwuUGQjGZYhg0RUqlsRWCPW7UkP
e7K+R7ynN3SbFH/LUi4hFsqq6wvuS5WLmnHy+m0+GpEAgxnb+CWg6xBtSfTioV7J
3mGazoollAq4Nk6NkPNq3108ZswOo3v7YhsrxpL/IxbgIx7Nx+6NQD1K0ulCuVJs
9vqC0uUpbWOmdrJ+0BgeYdtuoQ98q4yIHqtOf/Fx1XeLKcqtyK+0NGJAaicL4B0k
AaGp1kHDl1VmO3ypXf/H9qlBAtVNTRfCeq3z0z1xW2g4jDvHq0KKeqaTXNi+TeVV
A13B4bwqXLaleEZZ13Z4HJcYZza4KRCvmRW8a9wRp1xkXBYbdXZxetEdP1kfgd7w
OfpPq+EVnD2t/fIRak3sM2uBAgnhA6sBpXV0uRENbKGzuhZb5iBR3gmFlLnZKSXH
UD1kY2GYmRgfaGoFGQA02eqCkSWpYcSEsE4cbekbgkjpzuVzontg10CLX7WlQT8q
HD+u4Scxf9nTY4stjbVVtq1z/eSn6xpKGhCRXE0Akf0WM+1SAlyfW6KED9tzrwMT
/0756SsrQNkC5UrIISV0sZfFwYxKa7PiRnXshVRR+e6aQEweOXPINUJFJtwbWxtx
ULKklfkhDXHBcrT66kcCTNlWzrdgwB6a7BJ23yRZZm7+2tMssjizhviAlWIgb3r+
ik5G85l1fHzwiukI+2Ov2n1DCM8lGib0U+H5oNl+MRPrjKiaatM1K2ZtOorHC0te
2iF9eVUmO3HZpRmwjLtLLsT/R2THhyCrGFbMw1mta8tQgsEHtE9WSFjn1w4v0zSq
l2EUlpLncJl8+lUGZJ67LqFBLn0KIwRC2FFIPvfo+PZ0QQfo8htgoKIQP5CqbMlm
jFP/whFzd42ax4nD/Y1xwF/a6wkwWkWpzP/isnUq9ULbfRfI3EkAmGSwEZm55lVL
wPGlaqltwz7BYRwnilcXmfkC7lv05vQ0bF1ggGRngwzV7oVFzyouk8bTFYN7uiTj
TnNRkjrWJ0y2nISBcQ3RjThgsYf/dzWyfPHmglDJMLBu03a64jM3eOKxpFPghDbc
eBbT0K2GmYXQoDZafkVZE/YM+orCv1A917y+tJiXxKp+GIMpWl2rDSp0+KNa5nYN
q3v2xIaPrxOSIrtl3xHJ4F4vbF4Yr8ifgffskDxi6C+nbKzJHaoT8aFM5jEU2PT/
meEaendAnfAgANPClfRA3dCO9hVPL5xx+/8bZr9ct733wcFZNDKXp6ToNEEkmkvO
rDEqPPRp7WZV+eq/74Z7GYMyytaKZ/ubZ86ODtr8O63u4MbHv9CfxMD5AWCAAoMI
pJhrcrLJdP3SIWsn+Ep2J/eJ3F+ZUQFsFCvs8abXv8zbJVt2B2nvc+JuI5/mDNTH
l+T4nWA00eZCrDoVdR/cjSZDuNh4TQh/mTDtVxrIFtmrHrx1MT6eyNi9uEURxSys
uT4BzgR3s8nLMnHz1zzVFjemC/0A3mJJ7fqZfsfXzcsgTPuWC4LjUU8KxLDF4Wsj
U0WAhHCu+UcB7F5Q5NTI/p2kX7EeBME6eAcMs6xGJJwbbp8Cg3O307kUJE5AoQ7c
rTJQMoTAu1SR3WdWpSX74Z7wGFCYE2OaywOYxBjPZPmXJ+Wz0ki5hWKOx2Ljm8Ja
UP51CP+X+lJBsd3TZiWjEjs/egmtgWcqZpTSLJ9KDrtI825hPXUZZdhJSFSzm1TR
sktGKNvoK/tbq8JFaEHS0dmrXoNWjox1WeRvUL/L8V+ychDgY/u4m4MBaptdwcQw
l6RYJuSqP7H1b41U/CWDDIX/N4pEiQiD4TonuBbHUH8xV/yo4a14rb4isiisy/Kl
F+7XeLZHXTFsND/LIxhDhehI+XVYg9RDPPOKSnsKNqgfo44IDsL27KUHZgPiE7Cm
ST6iR+afWMwhqEcKR4iSSA963LYaJNr8+8JIvHlub716hyB7oBc5JgpgL5A+7Lq+
vj/Itsec+C9GStOMpI4F47Zmx0ZZU1/ySdt8AinMPEaraWyImCqMKd33eEUTM9ub
XsVHpae9n2/Ix7JrMn2bLzWBFYxSe6+36TZydDES+MlwfssnWGyUGVIi5GZtoBvp
NNt6aO8a2Ka7fI3NSWhUtQ9bIVRhXZTWqspjInzw1iENYyPrDANiacYxCO4r5ELL
MLrBHxJ9HbZjQ/7uxOkLeT2hKRu+kv1u/bHq/FPSCDAi6765X6e3lttrs84Kszvt
Xefud2cX8HG5rvZM2L4VZcp67HvhIWmFnXqE19QXPEOMFeA2Ag9xJqQoJ7GqdMl8
Hff1DrtxtU/7mDhy0rNq0YhD/BPp85MIayo3xD4JgFmGt6nS7dImuzCfrejI4pNo
bduiShZxIthOY1mOpWVthLTRW1Rc8a0aXfkM4H52PlkA/Tbx1jxkkK+MYHvHOPHm
cHxAVjW7qOg9wVfDPRv9dDwILsi2hWInF+65VN/KvdPn4GToVyTC+7mZncerwKac
pQi9zGxfQr+LcReO1arvf1TYM1u7aTVB5CpVvmdN798DVIgEAhqw3o6wv0aG/8v+
HUlUOUvSMpiRFB/aAmXDpU0I1ZVj3DzRw7baqXgw7lqfUKv8CH5DVL0cDvh/0I5s
dXVU6Ndvsc4JtTDgNx4LWBXvA9gWOzi0hlWTJYPCcsMZ0ADVqe70CSSuYZl1jGhl
fJtmQ2IrFvqCLFYGL4SKg3AGTIMQnV5zcispRj1vF2k2sLnWeikSp5Vuik+Qq83X
yR9ZmDqgbWo9xyBDj97ybHHE8+Grl4P7sKyAaW9/HkbAv0YQoMuV4t67rgVa/1ER
4RUy+pyzwOWOm3C1khqG3t99pNMNv4aDHWu/g5RD7G2HveZaOIGkOUEASno9FFCc
i2h9fin1m6Ho5knwGc+l77pa9EaahVNnWKErK197yc3vXsswJz4tyWdzS8Sw00UO
lTnYZzXJy49vxfxC0nQgQsD4hheNtxcIIk8Zix+fN4iVJzX7trZJJsMPwjMucLYq
BXBynxjbxkskpN7TOI0d8kM6vOruPK1QphltF6/2mTL5s/s8Jo6yqlKH0AsUNIE3
mUB1j7tfUAJ9bNoqL8TugrJGYLazracesKxvYr1AnoN7MRABqMKbrIOn8IUW/MoE
d+rWZCjcwHQYHh/L9RkDpIOrXNYkL9lB/rb4Fpc7x+Bn8kNtTr0cNdebXB4kEKOq
Z+X1bYRWHG4WS71IRuwCV2ztZ2E8/pGLGOdOyP+5SUX/jjDk3h9TrwIBv/nOx+Lm
ze7HY3lp21f15pd1atsWds9VsLw/Kx4PMquxlc4pe1ebFyCQ463q0GLvoqgIUXxm
4btunoikVNKE5urZ2qKzVWgsrfOCX8iwbpLDHcSPVHcc/7WR+JQj+FaO42wqFLQZ
J5mvTHULhMwGaRM4ftevejd5K+Q9lMm9fY63qWxDNUbRMovmXryQP2eJ0PDb272v
ln7ZD+Oh1RLf0oQRFlxhgPAYgvfskRA4S6BDztcp+0A+tAkl2xcly+St2t+HGTSY
AiZLnu8mGNh4Md290g1wKRJHT8363CJDBIu63V57HURKkkN24NhCIcSAOA3b8nDd
ZxbczSqHFSAxPg7j27lKDU1Wt9JNm4uSQAYiLoyJzXWtQ3IgyOZZSNijM86cHuHe
VwZV4AM+XmmfEMu8DCLVml7KE1xBiP+0p8TXs8QpXOkuT/KeuqZTEnHkicvF+/KW
TeXkdDmp/ZBDBT3BDw7bHn3b70OpUglaRFkG2NlzCgNuISo1rDkkcUvdf0VImiI2
QRL+cVfvQ9IXCdF41NDOQ+cl+Om92EOFi4ohSn//wxZ8SfWJVOjv814tH5hj+VEB
mT7dk+Cxfrm+HrBgwf71CP2D7GnVxmq+oaiMouaGPqgW7THde25Q/8OI02AQf8HX
okqlOFZhMkOIQb8rHXyLQxT+t/lkI6LVaAxMs0K+1fKgSb9pkZOJaicOHIhoKXH3
FVUQLSi55asKxPH19xbv7t0dxK+2vbEZw5P+vW6cUubCqYFBiiG3QAjF/iZrMv2R
hBlWhX9Cd68Ex4CCfIIGuNzAZhJvrtN3e9Cy507TC8CEsF6iamZL9/De3YD6eROM
G53YbKknPBQUsNeJblyvs+yIbMGGbTpZJ+6LO9G3IV3vy68bcHafTN+fVwXmG2RM
bJsv+XwCaNtVJTtx6YxUY2rAmOcG8a4Vw915D/TEqIWaIdN7ZfOHaebeWNoQPDKa
6dqf56jAuJ0/3lMJ105UVkmU2pM7GfpXTpFpmK52kYtJM0jLrf0ZdKRJRhXaAPli
qcavECyDnnOq480MQ9zRcDexoGHNDCYLRhCWECu/u65VVeiWx/w9XVLEXezpKe8n
dmQzGMvnisq/z7tIfST8GL5KdZTJ2DMXePWRVxe/njxzC3Hu0TmrVT7Hu8AXSVro
w9XD3S4vndNeLT8yawkCZ7GYmq6MZMUrR7oytHp6pjVFKHbBL/g/Km8HaZiEEYZN
RE9Q7fAK+f3dgDjAiht8QSlC3eze3RFpmG+dRN7iuhjysyLwr+Z4yo3aFT8B5jdY
NSg9Kdh+5em6oJHxCg4aXfe3KOG1wd9IkyPHh8XURUkC4T0FolwwB+NeM7/OJ521
bei/P6NeaS7dPv5XMPqvKlQFOpfcEr7wQhn3txUw/ilFKrVEEOGwMiQFelSoeQA/
oS3bCF4M68asRbPhnW7NBpf7887iXPRbPZf2tXGes5kgOOhQP02VgR4GcIN6V2at
aD3Q/OWMxxZsjz4/ZAe90VX383yH1y39OZrrtRliHabEWJPPshsWs0BMtx5nCxVS
74RcSCMpd/X6pIdpdV7gR//vbl2mJ3PJDjjgszR2MHunD+R5eEDjIppsg4YwAMgv
unqhPlcDSWDM1+MBuL7OLt+PP2cZTmGoE8+CIq95rCQ69NZ0cB4lPniomoPqNI9T
zAbySvIMCkvEdaQwQUEFsupl+7atWSgzE3sjb/IdLbPdkYEQgeTsZANLYqdhXara
IqYYxGveGBI38MIquNTYSKFCaZispebVJxzlDXLVpJZ6+OUI1U45ShMubUbTImwH
pmW2Gf4Yjz3HUSJ4wTWpZVtSSAz9qN1nMbZByhekjgvCvBkLadwS31qEGW/8Uvnz
i974HjnBo+rmsg+qKEliAudgRuGbNjRVBM0JrOIjdD2APn61w3QHnP6XD6V2eDv+
McljsS5rE94J2v8BwSOpmDX4DPrChBS1/RUBxhXq+eU+fyXbhSSt4LoAOIe3eBpg
C5l+NWMuf3g1GXUv2rLl6KQ6OTVLDuZ+dO3Fd87xe2ejTCSPUX8B4VsvRfmOsTeZ
tRg8ljEtgTWidaYMJf9G7H+KujXT5qK/7il7RSoLmXFHdsyhtqcEZiMHKWU9dE5d
s+S9J5A9Thq2WdD/klG95AxK/218XF8GI64TMk/mfna54AWnFMR5dkR7k62iP9nP
FpviufcynKA42Qn+zaH2X6lQtHIvltitJmsuyXncmtrcQlge9BIE+K4Lrz4z0N9B
Z1D/+5MJTWXVDHoWaA+gQVzXwMyFbL9LvVxBtWNJYvLu3fIPY3SWI2zYzvCwOHCH
w5IgbPqNTwlF5ilYIJVaRzRds1jqDueAyexbIu3oXtKA2elCAE4OY1jgAo3yftk9
McDmG4EPVdM74JVfdRtZOZS7y/dOYN/rfC8RaCKpO4rQGvG5VzYgtq9VXsQ7Q5Zk
nQthb3qIzlp+w4uK7tBQ+BxGb9SstT4fGiznEB5C+kl3F6h348cDLDpLqJLfVP/V
qAsAQBmv0XaFEKla7hE8hoML56CgGhvRu19mHO5K6WkKaUrAyBS6/CdLdTIaS83Q
6ElUfyAh6H8CWFxXdo68+K5Ia9PUFgk69jJNg1SNJ/xgvKMgKc6ETDdlk9c/WjE3
KDotW3FpXQvRgY0IIFY0OUNk/yFsht6r20j/Y25d+yakXbjhw/U1dg3JCgLdfbKS
7Q1e+fEDQxIJAneR3BRaGJ55GvO0gPISH3CacmYaR93q6XClpHf9WVznRB60zExI
eRQvWJ4kfczuA2yIudFUh5/G98mnNcld6J1t31hIDc7IYqYRLST/Q2/UZdLFLjQl
zCmXq/HGBlafw95Gu5KDxi1zWfoo7rwI6/hUbJ5sXsLoE5bnCPeIN3IMROnMxlUt
phAbPRdWrKKj/tU2egxAU8qj0HLaAbf7XI6sq9r7zqe+OqSESpEBSrJgO0Uqkdqq
REdxglDLBPRB/Iy5A2Z5Z3CSOz6OBi5QDJtNQ0KYBgg8XcqIZ794JTYVUqKNkShE
15KmJbkL2UQrf9D18fgH8tTvuuYoTluCuU6TiOR/4lEa4p7V3XwE2JFGtZ/+gzTZ
yhnMCY0nvnq8knB9EdfnYxmKW0mlOG2FgsbRKoV7WVDy5RjCSgc4exGblCrVIo+h
CWpNvZzFL2y5NgnPyzRSasWAhO3tSaorUnxbRQIwyraJx0HnQXKY9GsJB4x2i8QF
bDim1BvtuxYK5WippJJrKIiLW005lINS2CLGyL0Pdl9+x5zVZEgFC6zY0HLCCHcv
qTupeb5LGNdN0GRzDWTKKqAJ1C5OWA9fQZ6YsHGC9TqHGlIxKyOFj5wgZ4WGTQGq
JJ0dy/wtlXIewxM70wEw13hQUtjmQN+xlPmXvkwO5/PvTc/qZGuE7WYwcAWlBS1M
ITTIUYHzfrtbpVMcnObBSHswzUJS3W/GbqYusjWIoiV1D5iZ5/K4BvvXZJZCmoup
UMwbOt0t8KDlQ3VbwpTP0xzIico35nCsVkC4oyxEh1f1Zfz/NywR3ykA+Dc0G47g
jcq//oZgD/nZGBHbrLHfxYaVfZQ6hntOnJStrdEntiQAQtvDdNEbMKP8c1PiuOGj
kKLzOGvrG3XA+sluDLVGIKhKHD71AByFhTXIy9Hoz7VkFiqOA0rZgEmRE+SCcB36
BSz2U8Q5ESIlwr/nGwCWFWPQGezfHZibLmSaHZw+QGKh1vwNGwfYq71ByeeCfHsS
I4qvXIV08iduD/SrC/0AD6Bp4cB0Xq0B+lTUJZhPML9CcW3EHQm5S3QdlQARqzxS
tfgMkAnKy3EhDxjNXD2v8mikfbzk6uBKvYLoO77Q+w0WP5UHpW5gOOUcwrRs2WP2
X7W6KTXIOwx+dr/PYBIsCp/sumCotTuFaG7kSJCuFATg4ox6y0kx1PZkcCodPp+f
Sqs98j63a0nUqVwV+Gb9pr8v7dke5EGMNR6l5yYN1+yOfOY29u/F6YsIjpKwl8NS
ZEXm5xetQ9PV4+4EyVU8tByLKoT/Kyqc2qAzyScQ2Y3LBOW6SfSMQhvRZ1Ifs6Nq
9eqgfdHX3zP8d5NXnrJ44sbX4jBOE7rvzutq43mWGGczGVPSH3lt8i8qzjZ9eqIc
dY8tYUKkiyP1M492/k5gOv6WqZ5Ll9FVZox6a1aDaLUhXdmGjJrU/FajelgmwVCG
jkBFRUO7GhtE3Bxsgd+HnOYuZoO2qsxXEGhJ6Pr5pLjng8VMBR+WI7OFacUwEClb
sQnQWAfcw3cczOdu5+6WFYKLXAxY30fYkXnoqZzJanX3TxHGNbjwlShbxncqz+tu
X4KomlypTT2t/329UeiEh41nc6FfKTb68AwcyzW7Qt02y8+3NG4m2ya9QIwFdLVK
Vwstjas4GdV4vQycKEZoeQyDsJiihOXLNAgjyPJweUKhwTEipyP8mS0Gcs1BNO9W
k4OGCkOaC07w4GJ7qMth9jVvMfLUhBWqWntaYUrv4UUWJNLg6PDAEolS2HdB6J3U
iLK8leJW+uWgl+x9fIJFifmm9deViE9ImhRyNbQOUuVrrLbyKF7RNtgPEJDpXDHH
SNDwEN5CkwgXof0W3MtfnqpFNwi6K/qv2mMDg/3tjj1T+utZbpdZYUWWkFjjDtA/
Y6+dMg/WpkdtccnDKZxxoz8nX2/epDVB7PFRFhpkKPPyuBBodiz4KwCG6bs47Sjl
lpScOtXUqgJMh3rxV8KGpgGeyNUXbh3IjtujFxlpy1SQxETWv7OsuAMPpdwgWt2m
W45hLi+FLJ7AOc/P7FKX/j3wVhjQ2HtWXecBs7aKZTF/9eJDNPwXHAlzP91mwtLO
Y/KUBxPp7Sc3FzOAaLbUsDs4MbZKIH+ODnD5ow1CSN1LJuBo7ylMF7xwL/TfS0vN
yAMMJLkIzxgktyTEM4dkeqbM+VpRJyrsnHwokBFpoz0texx4Wq+EtntFK4c8Em+6
SBBg8cg28wvKTOtWtXj6iQwwdJlAHytC9+4uwq2ulXdbi/8QOmxSPsx9Q2BfnqZ7
IN8yhupygC5SkipcK79DV5Q2T4UHcJ5SnGsYZwwhdC7LzCbT39pb6eGyEYREaE3F
pOxC0SThn3gS2QE8/kNT/D+21noMioU5cx+QAJvHi4X0fwCG6vcT/HHhyblZza34
qbOWfy2PbmWNlvq+XPPWTiD9h2a0H1qBPq1VMQvtSJOJg6YE8UXwPvjHwUxD4ZUl
TbdXaIDk/Opbes9oiCgupqcnMsi23imP804Y0rVR97XcIDXgO08KQLhSynp/nMAU
G38CrEGG9oPbDQzS4mTw7rsioW1qGwaBl87kX0qWM1zcUqkqgNKzNwqNstR8J60n
02mRd0sMsaM92tX1Mj/OBQTL7H1NPmXT6L4kr4kPduRgLUyHHp/XXAKKVBQ6JhUh
F62TAw7Z4Fzp0JEKK7tlnyA7UpVO8rXof4H1TyT2AWQTaghCObCcckcdWTofAjyf
tO9DPh008cDYryjcT6y7a14CmwhNgfUxRoJRu6HANkesX+KYQhcJoG+sQIHpYnDi
Ysw3VoR7tlslHRdZ63B83JWsEahpRDdISxJX+Uuaw3c27caaqjFIcPVY05nE4VbB
cQG3SD4M9JNyMuUUDsJxdiaowVc+PxnqyyynmzEpmlaPVVHohytP7vnSZGj5PNHW
yMqxwtQb5aJFic9h0y4/S1QcSqmGcVKq0EpjRNKQ67CmQfWTpaX1GPMzO1peiAFV
DjzDIp7C28IE8NZNzQpeBRr0U12/HsLaZBSbNKeyUXoskO3cLFaa0efskmmODyFR
k9uRQIuwa9tCHjaiART9IMeDvsvG8OBeC8bQS58NROLWRtuuH0jQ02/zMx0xnQxg
vpmXdB9389YEvzyw8kIhwof7EOkHSDUmfTmgXdkwLZHBlfFLzGV8KoI+fNqGIpEf
wziliHK3K/+cD4MVgV37yoFea4L4vhWFHfKGy5rqS1NYkTq0xCBz29T2saXEx9aw
kOnNqFmsOW+J2eg4dHuEvIpIJ9c97dNK63qnye4HKDVF2UFFYwHkyi+++g+fRFdT
l/kA27UnvGcYv2mJ33JKVsJU9FAlWLt55XYBTfJtEFoxvPwKb3ehwRoAhCSsRX0S
U/fox+jz7isM8SJxTI19QcgtBeB1z4l3AhsxwF74MK0eJY77/UZzRNc1IHl5qRQv
Oj+e0G5NDf2uYcI+IoY03NTIDWVTmXe4dR+6FYLb5qjyQ0Jer674V287C9f2Ugko
Q/7hE6ByrWCnULLTHxsNrB/VZLlCg9UaJ6yOT0Z7E9XWlSjNphkQ63Ve2X5KlFcL
PTfJfwVeZN3zJIUFl/hdvP7yHhZIPg0m2VM76omSmLUYznVow6I2W0aFexykUqO4
1o+si7YeUzyiTAJEb4o/+vFBiXmFMvdrdq+nSnC6KG6+jgpEL4ah2ri/W1EC+/cO
KdiJmTXyKJEs78rEKruJptLwkxvkJU3mpVEir6Qtbjm1LErvidBqXiKQhlFa8z1a
F+R85uVAo3ytTO2pXP/tLoOyTTAtAOyx7cyCSF4p7cFjbQQQlrh0iXp9f2kToRck
U6p5E+qTIH5ejpebpvgmme319sUau6aHCtG8P7yujhUcw/IzL7HrFxGKngTmkA8q
86HIyI6jsXpoca/Y4CnXw6XtH6k4WuvbflZ97BvBPDqJSWa7wijWvuk45y535tTO
52JEG6rhYECAaITs5LJBtDPPZTKI2n5eHcjD81B0ehhW0gX3zpUuxmk7kO+32MmH
KgWZUIR6fh9vY7kZTmYKNOtZUKuaF1JdEopB214MjvXwau4tDdASj8L9NW/+LaKg
XZ4vZ0ghMrASUnXPwLzNnNM7e6f0h5RjIEznBV2SXL+RdWnNRrvduGQKqDvybTUT
aOOY3cxKyjUXlqjUSr6l/xFRvRvwz/uhJMaVZ2/NBSqYIKFIo6H1nlX7GC0EshBR
UHQG0bSQ+LNbDBDAyrBlgfjWTOKs8IeQX5Ka5rZFMwf2gWidylhZCH8ud8Swx48b
cFUYkHZ6PNxeDJd2txh//MhRTirk4G+xyqvayTg1g5psBh7vxvlfj1GoIFjUh8uZ
BE1KCB+zOJ/Ah1iekqRhTOdHleHQA0/5gIslMNel3bY2gg+lPRSWF8TloDHxf1NY
T/8EF4no+j4IrURPxo1qghcgxNGse5ywD8Aj39bhiFavWKiSB1XE/Pu8ZZSwQces
YqxxKqGuCZy0FJfjMy6VdwxmIHB6J3xoMEYVfTEQbU3Z2sGKEKgVVbSvgIW+F02H
PUxl+xI6unCJWzJ4wG5jsFLi8LJWV+53j+HnB/DMrXhzFrs6JKr0QLhU1bDC1FaW
RmD4rP/UIjbL5g4iz/K83DFNPtX2Q0MWb8iOf6gSURhp6toCgurJdQCoRYilD6Ir
9+B8hWaxqhzds/Az0tjDfFvurnIvzrjrcm+GFZxAhLo2F0VU/yGmbQI+cZD4PdVj
AZa87kMpbXs1zrCfLjFfnb8vrZu1lC+rseg2ypPMaFqtSoUbv9jm/CJWyu8Ifamh
5lCJ2YmC7xPVY1euMKEB6Q6COK//JNNlHoHxQADsWY+2vNXDNq+f1o2Xsgsa/rSt
smu4Ex+zgRdSZNYaV60mQFdEUzXApzlwCuTMXnLIGHK9o/FrXJS4Z+B+F0phjooz
dxgiYyTHX6V0diLSrajGBIhbtkFwaarIVox/5lajSXB9s2TBTN90lLRqG01bYttu
XPvML0eNsGXcbCUfufHwH5RWZRPN/H7MpPDKpI8OBCcht403Ls2AHMc+mH3KSp/+
ikf3gGRkw7C99EhPFeHqrJ4FgjKyJ/C7s7XQ/L5WvG9wS/ptTp1NH2rkpnRTqqVV
Dr3QRrrmGsZsEHu78AzdJh0HZmYUO2mn7sZ5s0Uz3nXqB2ekqve42zuBdg2i+o1Z
RFfhDJIYNA/VjlWFaQex1Fbd2cYiwB2Ohdg/4YIDwcbTG9ez6q9xLFWrLv7Tvn5y
Wt+QwgjE+h13FtkGG4gODjV8wBC3KeS5vOE0fLo8jmUYqmA4GeoJuRjEAmx7pRPq
KJ9HSVre2p8JBKW2cUAegYLk69f7Nz6PX8QtxxjYjxjwCbpDYrWzfG+txrSg1BZq
k2K6ElbSKz1Ne7ROmTE4Wqn9eb8uaTMFUoMpmy/qX3dLOqGPSHSDKtcOYW9hRe0R
i6nchiox0dQ8jw9iIBShkdD8d6xoDP78Y2ZOY9sEj5FEkx9W231Gzc21mZlTAARE
Bc624NPcbtulab/XAiYnX0GMY9hEEPo9E6kxykJHSgA/7TBQ0FCJ/zmp274tbHw8
DBlCL4sPZPXpNQ5nM2wQdgxLo3QpawiZV3YBajzFWti1RjHGzrrDw/gyVooRW9FZ
h3on7Xge4X+4HbZXDwnXTjjvq7XEUav8NzrsDzFZfFm7pxRkIahQt+4CD18tp5bv
+2rJSvHr4PZClNhDeN7pKEa9JCd2vc6lcJIHh2NQNqde8tY3fXj/jHWtDvMRmnvf
fWUSmRyahazJLJ+3YraLZq1WgrB0RQe0BN3jJwcb9bRtu5+/ZHVDPTCtcIwQoRMu
MmsQn3DwT3LLV0o4dUV4Yx8VD1DQJlyA8Cu1lcyZ9IV7QVKXZXW/BMSReo2JYz8j
RrSPjxcabs6veHbHqRt8y9ZISw4qZGDOfRAn3MQF9aUxl3pqYOp9wLxQUb3ZS/S1
65TxJxW4wSyOWOZlNdlrUzrOq3zkqEDaply/TzHlL6aoc95ewtQKK0cFMM63ixym
n5eBEJGf0NxU6qDDL/rZMORyz3rrMTBg4Vm8skYMeWPAZkiTgZHnDSN9VKMC9jDE
K+FYxnQswwMhNm7NeacaYdjXRkbMmfRsGaWSa3PrSUSrFf5h3W1wv//fEijA5bXm
GBf36qnXtGoyVLY/HTk8lM7by5698Kpp51KE+rcetfTFBrdYOWjzc7EoxgSsKckE
Du5WOhBE0T2tfzuJywK2auTYPVpHHb586DceimhCnaZyTQv7ibEahzyENybbuGsA
qhJowuRRu5ULiAS+Gx2ykpAxbMoNCIO1cs6dGQL/DzenT7O0OgzvNGR74QThInbb
ROmPcPXvnlL45jm8iPnwNf/1esRmojEn84x3j0BPjymR3mILvgpeklcAm+QP+tdy
I/YlYyjYuOm3aPWdQ5xjtop2DPE3e2zXzKqEQ1zXFwMo8qTvURiSPS8Me/8Kafn3
zmO33H6J/4ztB22307i/P1dbXiIxukdMAOp6N9q3hhcSfkGb/X1Z0yplaB4qnkjO
di4xDaw88BocqUWXeqrn1p+W0gMNQUcjcneg2AwZAls64nWQ8XYXq45PQagHj1PL
Tz0hTUaTeAOhwvPkENrLduyL6krAiM1rlSWksE4Sn/vJqyh0Dl5dzsFLaHouZXtM
NFFC5ilz0MTBetaaYGCWEJ3lFNNxI3QxQlor8K3hP3WdHsNXRIOTwBLrUzhCAvgB
YDhYO42e7M1M3YDXZHNm/swDFYvqqvhjdgDZbfQURUoU/JlxZAbCIWbXTFhMhBMx
XyU4iO2psFYPxJLnYuUkB4hZ3PtqEAV5I9GRpffKZg7ELE8ci+GxfDwdwY/yrIM0
51zdWa9lJa9uSwkTUl35lTcquJiHMSO5wuwXv/c8I1KPu5SsvlFsQ5yXQYoQoYFO
K3Ah/2lmnnHV/UkxZ+0j9jtSWlCF33kjVX29irLZp3uX/UFr3dUlYrRhtDiEGKg7
JjHD2uB3qHdyP33BZnGfln4eXnMVroa1wbVVYYyTPe/R9CVsRH+pTp1uxXMdCTO4
1lX3wJv2QwNd1qOo1aAD8I7beWjIZWqYL8oIoFuTFYnKKVS1ip7hdsQ/ZcLH1v8c
Jk7W3+saMD/ync2yORHzdIIhRJ3fQJaoC1IJAwgVEJySnXLbe8auRM2643hebLzp
AHVAs8rBsXQdwF3avvQAjmAprrNyzmQyidhjZX732JjqbWUg7YY6evyXb+e5ZLXa
5ezEwSLqyp9v1yQhsNE/TBYB0+YuJbwr7cELDKmyJn+hVCg45X9+BWYcTyG9SdL4
jkLqvVICjCtFqECHXsQnuLt3gI/ZmecNfpqp7WHfoHLfgoKj7oyDc/tiQp7zkTYp
KGROGBzaA9EY3UlTRa3fw78GoRgPGL/bP919nolndg4fHZOQ/5OA3JGH/An8CDfY
kmKMMEUGI4hSyupi8VROdtccIPF7aam6DQSVlA8CvX3vVpc0bMI3+1ES6RPl85ND
Yo4ceAXvrwRRVMcMNe5rOYyFnHb8mU/IHRQZK6upqusl1DC7OyZp0NblI0uBwgxH
JurcLXN5DhsKDK3iD9GWbtSoIz+/KnyghN5BdvZ9TjyBi6rQ1uQ/r+9PRJhR4B/e
Ow6BFErXzLnLVz7menZ15O0mj/ssER/TszsravdehXefZWLfwRiIzEX2Prm/W4pr
zwqVIdW4S4LveyTviv0BVdoYjHEKX3VFAyKkHSSC77cwdLRT9K6KY4XXQCKste0x
XGjzuk/+XJlh8tPdIwMV6N0V8d2MBMBd2w8ZnJ0yCazVMVCbPan7GtFHXzf6JuYf
xWiIl4JOdKviROJ8TJ5+t2L2Fq46qJ6sEAWDykRVcesDtmVqAbEgMMwMMtEcMUn+
UNXCS+eEphueo02ZK3F7rdpf2SN2htiQfSAYnD27QeHVOqQmu5B2byUlTcFL6Xms
ibPs5uOaxvtRKOY3Inc2GngI3tQxnvAAaREsA7Vy+tfnhP05l2mHG9UtS83knGL4
+9AN8M1paHD/yzYaZUkg29JenDJV9g7AK+969FkN5axTiu6nE+reyFphjwaHWRJN
JMreK7UCH4thZlT+R39i0sF14iZ7JwXH3m/nbGB4dwrl4Avkd0NotTdzvN0CY6vs
JkOtTr2b5eQfGwfHOFvBtZVC9h8BK8BlqeIlP+NTAkITB285QYt6lr6Aual0A586
aO1qJt2wrDPeTfBAkJJ4P4J6+pwsmUUF9YTOplBtD/0+wPNGe2TaFMjgWhvNwj+Y
IRmIAzqRTmb+sM6lo0fl9MEZdEMz4EDUfq4T8RhQuTEurgXnwnlIdivJ2hAP64V8
Y+CXsp0CrjdlsSnbwgTyyQSeSXplN5oF+SynKd877xXvgXNm2FTX2xgLwI57grNR
6X6LAtff9onAqbsR1GFoVliA1asXNJDKuvFu6jra31Ae/Bla3KjJ/tLOUHHZaUso
VyzzBzkxF5evAcCr96+ukz6e/Lef5bg3zp27lak5SB6c91ND3ubpy9NGooqXBOpw
EJIWFPxdlbWnS1wWefDw4JKtJOaZQsGS2mAaI17kqOPPK6k39ZnTvrE1m9UXfPgH
cDF0WYmJ2fGg0VBnQelE2ingGPV5OKAXuasZuiunUhTsEVu2PAp5XpdyBkzxbYFm
47XbFycZQX11wcVE1YguvsMqIxvncE1jygQK2NVPWTsYONxBZOVVUTfsSNpHVppg
dBwCmQSmc4ZT40qNEAPAnxk+McEVI6AKo9pNhaj11PczkVyCGgcPHOlmP7ofAYrv
1LT98dqVH75jsnLmCQiojmBz6UA8VyGxW1o9x9v6BjVexj95OoOHY7rNXvESm5JZ
e4EXpY3cM4fb1xe28hQtu0QxJay9BpgQWLRMcFiMd1t1UBTgLKpVQyZquptOZXrK
xZk3rVqrjiO7RdsBsq7Ba+eyOnyw/A5V3Q9isggQKDs+3qUR/6cfBGcocTMrBbxe
rFeNtWtJgbZmLUDCazzLakAnrxy9JXjrE2spqBcmX0lRtnM/HyTYAJfoXdyo5FGm
q/YAcQITe+0yQURUnzntPwN4zsLGdcnWyjZ/RwajWM7OqZhy8xt+/P3tLVgJOVsO
8pAG/EODo0QLnEy2obWh8xUX15Nl9owSjFKieliLDcEoazC5w2yFHjlSslnmwApP
M7Ybi+v2OHLFgUqvGK+xb5nGRJ5rlz94Abxrkt/TlLp+FvGJ0aNb0hV1cWwP50ig
fioP6QoX5BF1PaEHOs/9rXANaFMI2oH9fkG6JJrdnSatO+sgcxvzQVPd5jXcw9qb
ur+vL3UwyRsMu5bfOxUW/kduXgOfzSiBQJxZWnOAswJ6OHLUeo7FinQLPrV9gebm
k5nVTYv6TmmDI4l+Cb1Z8NN3ty6hHr9TVKcEW3HBPby4IuwrOrXPJRAfn+9zx/uW
pkmX1F+yHTTEKlg616iHgDxKxiTvlsbS0ZpeKWacW1VQosB5E1cOS7FDoKpx0Myb
SfSCsWQFhQ4kB9iu3RePzDj8WD6zgfpoLrjkm71pHnYQIO5UJynlk3TAf8pfZArS
VTNb9ChNEjJ+h597HRv/E31zOBGfu31HUQEcF4KXtYuTyzBN7IR+PJD686kT5qPu
4u7qK96lAxiWHgNEF9kr/VxE80/1et4Pkomb/VKk/oLFpOidc4y9sHD+aGVo2Fct
Bhh1Y+8bSu1LSLzaPqUZtR9Qy6L3KIdgadQEfdpxPkRddMk/Boa0dRv7qUz60Fxj
n/3RDPJcbDPJpoHWxSxtrn9kOI9PikdzUSa1Tiwz/87c3x7bJchlpUIGKwGYRDWI
GlZNabeAwFNHHvS/NBtpc53OwFCQRsOY6tkecXXsZ4Hoj49JeveEOAG3CT9s5T0X
LI1zMQkob766Lk/ZyBX2JxIHXyzRLcpY5RskDQwHYZNO+NTFa8Tn3HbXZ/q947Gu
Vb8sIiToUpVEqhwWke0a1kuZQ/uuj/Mt7H8lzhJJzq2UGwPycOLOxYZjecf5Mv9w
LgX8NyaizUQmAYXeaaLn0Cig04n6mi+OQRSbdTNLwagHtbXQ2w7J02pGCRg+/I+b
ekJeLG10i7svzRItzYIqA8fJZVVEl3T0LpBHd1ON10GB5TkWcOB+K32fU3UdknCW
X780hDQ9iMLJc1T/sRKS6/5oSGdCxZuDLwNHRqmXekym/asRbDxu5uDk+lKa2Ya0
whMHSAXoFRrp0+ET1LcddroGtGWOJS9GlbR6bAWafMGNx3O14A2NKPbm4L31liUV
1VPCgP7y+ayM3IjMh0rv84f9VpbJjYugAHxY4pgrck7kw3Jc7ETZQSJ18394WQLv
BW7ShDogwEzbQEjGYWw1XoVvKSfaJKw/rTw0dUtJceqX8etOoF8Vdo5P+ri5qinF
Bvp3ZO2OPvCyQTTwTGTrUkJOj/F4Zfe5hCC/PkU2HS1HBXVwUjg8PHl6rzcDIxWZ
ecwLZaeo75zZCbJfh3YjMlsyK0TyNtRfNEuv8XA6VnP8Nz0ATiWQOT7zG1jeekbP
0DVa3HjdAMCUdPDVK8JXWWPoeP+VLyF595H3Vv2xPEyNOLU2TF34WuLWlEHWkNPp
PeKKslDsSEPcgXgqRj0D9ZPzhefjVLlJ1nv974eosNT2O/gsTpqcr0EdUWNgI192
D2E+Zu3MrLaEIFKxEktcTJDXeP3XikVFoFIF6hPlMaj3ikikOlhgbPKOmNyCucwt
AsHBWDuSq0mPlCyUNrpp07PLF7oqFDsYHqtBvyyr3u3yZ6OK82udzIGdPkVO1FZg
CBySeAxB0CdbVltKsvQnWVrCYLOQwBxQoKGUl0pWYVyZKiIfruIHTgkr9tQnoXdY
+ZB08Tjehv3LWlc1qKOfLGOeIpl7qy69r33tVOMJfHtCigNyCX0TuAZEEIDteIOY
yKn1frTV9auS1OggmhabVaurDPfjgK3mhHi3w1xqfpcLA2X38h2CLEM8tTbq5HOf
diRX5VWfJJlF3KHD3tbtZ1oM9qsm0n20xv1biYmtPZ6wi6qCMBNJVDMJi2DyEJDa
TIJdpMt6HmxM/rGyAmzwLreuargAyeuRrUSxwoXq6mkH99MFUdXSOq4vrRA0Rxps
9cPoy0rVUn6HErg4yM7JsQuAR67lp/cLcktwfUwaEQG+YbWq5dSaiI6k33/EJqnj
0PcvcFvWtY5eALmoDwuQ5Q6MNuA/a2WngS1OCRRA+Ii1r+4TwLyI27qfnNqHZ1Qe
fwj38dJl2mpRYqVQ2zqTO0rnK6WK0I/Ug2Qdr7LNSM3dnTIkkglhlKHT2cxvizxu
i1wHkJTEzDfv7iuQu66/zRROHxKuIdYsPV22aVF9cZ3lPfai7vEYA2FGvfNgRK0q
MFydrMMPjmr2a+heoaregbSFypYJxjh7YyESHnGSBo9gTOoW1Rlc615pWlCypXKS
pG4qj11P7o151i3aeEY9EwFVbNfjisuuaVVOwMPBeQH8gD0HXXDo1v3vMwZ1A6CI
R6GqeKQhJyqAiZ4FaY3o4vf3iB18bmRgbpWM/c9oLaE1dzJ1b6INfYiCOobXRfJA
Gyv7t8La6X9neFIglJ3N3eBz/cLasNEHGTXhK/LwMoGcJtQq+tk0eJ0SQNoz3Eul
wty5EZyt/1YLJWkmab8YnIbzehf7AJeOqOheX6WNxC5ZYb52DQG8ofhPWZf7AZB8
7pTuREN0JFpeHUWJnmltoXWxvLXzdsJsZrC/K9bTreNVXzCpT3OEHf1J2PF1mm3C
3Z2q7OtVij6+/mPKMdtet+GZa0UvWt8Hhxfwvuj4HAKzyF+RvCBq360a3FI9NXKU
s+/FFfBg7SQb5tdKULPmKefrwrZ0NboKnmLb0K/k2ZPLvo78k7JD4AedpGYysqEp
yg0emW2qTdBRL9r+WW4K4j10yxmb/nutLfP3FZA40wR2OAORSEx60iejMFJNVeX9
W7KrAoikNllhp0vc/UTr6eEH83Ct7Ejo2DeSb8ArNIDrd7xkd226E+tODk8goGXj
ycRgDMHYawxC0iJoLbXsNlBGoN+kKlQ5V2WHk495OqzjanXHRUeb1dx3e5pjsPsK
zDcIoZ5NGKv3vAdgOMvIigv4v9SLC0avN52WETsDk49bwocrr910dLsPPuqzWRiu
8p3U6f12spfe/Z0QDHW7Wg0txPiVBqyieKm0as/yO3jJoZ3hQrdkBqNNlayTXf7X
0iIXmfeBGcginEZ/1VEkA0yAZxLcuHOrsKZ3jZT5JjQryI3jSYf1BodLyZuGxwfr
hfUrRceusFnLLwrX4TvCd5R/I8yGl/LxnjaqzdBH5F6XWc16YIjGvHNT2sU4CtNb
8psGtiY3pNg4m4mwqmMG6rVyBhMcsBWfGBmTJESBmm5wIDSQnjqGIulM4IbemIaY
a3XMKd7JbQM9y5RMvDx1ctUx7/HcTYILZGqKyumwAvta3UQg2nHnr7NP85N0TSHk
rA6JLCX7c1JrCm0ncxig28my3SKz0GoRPJjjYUcDJhjnuT/CPYrf26l/cMyOgRzZ
4X2H4opjuj61D42D3vl2UoUvi7bfNiyLd6VNzu0wm6je5I3GaMkBQizkez98HZT2
BaD4w7mKapFwd4HZq6I3t0GG3GXIZUZtR2PsqgznID99CigWeWf0srfFTPkraBA+
HzzIsuKaMuYCZqX7Xq4WO0/CUW312MR7b6ZMAJuxgPQv+7zlsHBw3HCmEEuBvZZi
h6FXeOR6l6DgeP2iUznT1MMlohpAT3LdiKpUPjbI9TZG6fGfyH99EUK8uBPPGP6r
SdoWLgTIoHlPnCyMCkRT1NTKkcjodNv0T4sS03Zjg4BlLnG9vz95l7ML3lf0oprd
mesPEIcA6H5HPhW4fOMtQoq87KyaCSsyvyHJ2hp0h65exnb6i1gG2gHB7RgK4dkW
MC3SHeE7uz9nMGjyHRe2BQu1Dz8eE8RHu8MmcwJLrgxvLSFQXkkM2siTD4HEjLjo
ulY+KHpUp3pd15Hm4YbXqLQXna8ZhTBgR5GKsEtmcm+bLL957hgEM1ZOrpb1pjlV
HVkHF7YI5UwWuhFqlgjkKx4Xlw/3ST8d8kcpk6TJu18lgU90uHwaR3/D2dROcZHo
YfqzM24cZbw7mWL9tZG3NJQAkIAhzjvxlje/1Elak3VCAXlRIb5Kzr8ZkmGwCvFE
mLrz6QaCIqCodT8coLhoxbSWafqAX7Vrs8poVmzmU+OFgTBO5Kx8zadtk1Io+Bjh
gx+Zs7ugyKYgZNBrl+t7ioIlFuY/cneCOQASlDsuaN1HweubFTZF42QrSG/sd2VY
cgwM3KChDZxOFb3fZtDqI8hpAojZARGlmehaFlo2DYEmbvDXxVTH2yw8XO9tD23+
WubH4W9bXMu78JDnRyjofT0ZAvuLl6Yj64kklNki8E6nHD/GMFgeggpRvsdBG0X2
GjMraZSIsejeyHEhepImBUpCk537Ry3gcuLJAiaXRsfzAT/nrglOD3kqFxCoCiP9
Qp8F6HY9r0GiTbgbVrFI+mB71nNJnHGUz2r2rcBdTGKmMsmK5Po8IgGXj/4UZANI
qAKTTaL/pOK0m05xv8Q/2Gw/l+fbXG/bY85mlUKCL2D1CgtWpgagnDGgM3oCcNHA
3ZZKHVzMzaWxAGUGiyWRAQQUa0u4HSbY+WljgHrzwYtSmZ5mSi1w0H7he+nkyjs+
NUCSg2fninQIE2WKZuWcYXrLF0LlGmpTh/ZsJAh2evfbh0xzoIpTPwFBzLVOySE+
EEqjP2I3UN8FXucnuhuwYLCkc08qcqTHPj9UspQ/orNriLrH+/LIsyRX28FLWHlk
Pe3v7aSunwxpJf1d38LLcdobZaTT+xD/G2Ezn5SgSWcZpJ3U2H9diFW5VReYbHOq
O37PCQZeL1l+IV5JkWGTk6r8UnFM5+yZbSc36ILlwdIUdB/Z70/yo79LO8/RuDDO
+22j1ee//JXJC7wztXfk+dbMgOpU4rqKfOOmybCD8oQuL0R7BnVVACmUnJlv8m3u
bshnkWciSPk1STtB7g+b6WhEQOPtKZ/KC5yKntc+IEXHuldH4kPFg+O/iZTGOzn0
gNeG3XvnEX9HW101n+SZs8b9fAyVQxNH24JyKt3ha52o5/QWYjT48Vz+oO+bk93K
dwuklPOEL8VZKrzFLslWx0/E8YWyRr/BBBLxUqmU0bPLFXoIoU2QNZ6QBOMCLCy7
7Cr3Y1EG7P3q74mYU4pGdXJ4njkWYUyxeGKbPwKJLPErurBiLW6F+GHZXQdFNC+g
a1q3an0gt2EN6If1pRIYRHHReNymUP2Ln8CMlHIM1t28St79ZYgXbkdvV9qMt2A2
+oeX7zXTNfaeiuTrifumhMI3WOR1zXIRBWmbutFtQzFq8B+k7g+HdD6X5sbRU3G4
zRFpNU6FAH5JW+EywqaOhe1avXeOmlW/thdlEVXK7F7L5muT7Bqvy8x5yboKKrjJ
RRLC/lb55qgPHyd+eTfLhJS3YydSN9ew8PiDzamT+wbGdUSAVSLzt6fc8MwbzvNi
Gf+SLry1rIViNJfkU47eV9r7qwSX+hP5Tzl7f2w+Dar1wecDxWzyxUzA4W3sTPJt
YGcseV3+y3KH/yxRV5dEM++9TpmFAYMA9QdjTOEnLcTOO01gVr9RDZEpXlfRDwO0
hi0lSnQvlZOOv+enneY6bqEmUowsNlfcq6an+hj5jtOuewaRd2nP5qw6881DfopI
TjnkUFBCFo7FczwCH3Dv4VIJWum8jzIOSt4LRolga9Hv5FVnjkCseuGBOIpdfkAH
Jbbwbl4wXVdH4aQ95YMfoEtp40X+NCziW/aLDmXvpoE3HsyUuz1rBQGZSO281BaV
Nfjv6LIFc1w6zoGsqbvFal5MWb4pSukrSQiRIO0do6/C5O4sNv7MAhn17qteugfc
9elTlVgTYw44C1QtJBN3z8DflLSo+f0IwAqLN4Cr50pXTXzmjEBvvpYARWEhzuWy
h1hiALdqLNCX3xmn50BhPEgXJ6xT3HYo4ENiAaj24a058lPn7cU4ZST+R7hUYuht
p4bDfrd7JcLpnUqkjOmsTf46FROmo6zPkYOgbMLHRwV5tEP8y8EY7iYDOnkHwydw
ad/3hLbHhU1jGiEomAFP54Cte5Z83UPPukAmQqElxUIXHs97MYiTsL+KmwRNS3MI
/ftZOQx7pYTiKHbiw8OMw61RLeRUU7f/5zUZH8H9JokuovOCOP3TEwv7jNN0lDav
xKCQtO/7SPuHhUIHk5ZXENvCF9xR5K5PndJ6ruR5XuW3KnzBcKqiHM2fhWfWs3PU
jw2nKdMdnQgpIhxF3HaMSuHB/phqtRGqFXsmF9KqW6fGWasY9PhK8HSO9aqta2B8
J6vpry1MHR0OHc2RrYj0rYQ0hzq0W5egSv0HpLiSqbAodqIVB/FZNqtIGwTTdH1m
iUp2zLTF9vjWUic90i68zXm/acdYmQm8emAyK2L2GfPSIy+3m7jbeczldRKty6pe
L3WpVgjOk+xMD2ptJ75GiXimSr+eegjGoz/dmDx/AcsBXTF8HRQUZyCBug9aRpyC
Ns0CdA8hSVNd4sTdqUEKJqlWeL5ANRXvzU2AEK277bBnAthsn5lonohu6N+BdGq3
Svu1F1ziNeDsptSDphw2xb+tEQ58kD8IKv27/m1iWI1X5UxI/arQ7sDzNP7BeXpB
E8w73iYB8GXzjKyI+D3fn3zV5tgqmkF5jd/iSDuHyaUs4ubRVc5FH+Jd+4WIcx9O
fS9xTc917DQ4SPf5SJ7bT7Yr5VEv2DKzEwaJUHmJmxNXIbBaAnOEq82JiYTN/FWg
lipb5GEpB71i1vxGolDV2HSt4X2RX+OKfJgx2e5l53k/SuabXUtZqB6HSMh4vHJw
6HWfxgkRNVDGDolB/mwg3srpo003VAKbqCD9U4XnIKGAwYg9awX2NEONcXUzCJAU
iBALy+s+ekjKSbzBW5EesV/MgivcTKC7NoqBTlL2sI2rYcH4eKWT+d3lhDQv/FNv
It7XgC/tIAIkz1TSF8XSYWtqGEIaIsuKG3DSF3x1otzSZ2G8drZzbGjWpkOeVvJ8
BwNZ+qLNr28FtWjdpaQZUPk6wrOZSgISoeqdvPvwmENJ93cO298AaAozm+RHfvXl
i0DDbSmOct0EpW6zz6bm3Oez8JczL6yoMyOQ2rQOApsQr+Y2EX3H/d7i5WBzgmO5
X2Y+tUjQGB/axtIFTZzQwYgh1PJVkky9kPCBELWBzx9cjT4mN+NB35Iu73CuPSkp
IsCJZNh+eUAYgOERV5a47stGr15KXCI7pXpkXAflsuGyF5DcQIyJ4dXpDP5sVK1x
mOnAVsn9iMav8pkB+9l/i/HGnPgUoizuwy0xOu+gAMBsG+Q7QrraPyODBxo0/VPI
lqQB1TTyw4q+t0AjV74GnUbJq4XiLfaFCdyP4R8aq3h5qsRg4qAzrjiWEpyS15Lr
skprswAG1QzvaK28zXCbDYpseHitYfJlYqwhgXKtZOg2Cx83miErMBhUD6lmv+Rk
oWUpEZPcu95lDKvzgr+Otz5sm8fFr32R1R32ooYXgGc7KhWETvPfKzZHolJYsipB
u9goRfV3tGMZ1fXSGy0AFyiO8r5AdEYzOXlpBhz+4AYIWuVLWo20KygxcDXBFHPy
Bhm80yi2wofpDMILFeM/iHRhNSc9lIyPb05Y31aBxdAvQ+EoZLwuzjB3ZCKTSlal
6GDobB1jSr2RH/H2ArQvZ70hm2hYcI2yrrqq5808BpoRsi4WSPVN5c6y6dOGoaD/
0DzlZD+viKSuF4mXQRTyfFljx4h0ytOOrFJFgh4PrwXew1KX+/xP9L7bvFjg87Xh
fIblYhhchRPWoKvu9J/a5ZRQTXwORt0iLY5ivhoJEdgR3wIeObyCueeIjHG/h9eW
hp+9uZtjAH+ijA4NVEnZKT9kQgn1TFuge68cPM4iPr81iwI/rpC3T7HQ4tMBFQUI
aODyZPluiCerMdYs1BssQgb7+V+qcfuJBKZbaAcZBs01dI4wBIOneb90yS4i5AbQ
u24KUGNcUSqUCe/SqoPRw8ylQXQMIl/eEYQ8unyuBh7nV7i0j4spndVdA/XRQMab
05QzyfSgntoBoCrW+FLlPoUs6sIJSY7X4YKD3opm/EDs3b8cdNALbxVPTbgKTFvi
wfHH6yUjrPgl8JmvEuL/veHtk265D8mO3OBD6PLElLZ2D47M8mFiwn6zEOyjPzA0
BiMq6iaihgpnFoqw1HVWvXrXTYOH0U1HFq2KVxPyrPw0dgqPdkszXbZvTk8hLuZW
7j34oCu4XRTG6i1LgGylqGRQyWrNY75AvlHRyFkzdB7p3g5m681pSlD5aRA0AgNm
1nipslG26DUDgmb9DWTy4v1pYPvhiWGU1QDziZi4PZ4PHtzurjBVRsEIcOiSLeB8
ajhW+GJ3dCjpvXzccf271GXYpS2Yd35BMj4WtdQYLrlkcduh+5W6UQf/bj3mvLTk
9yNhjbXyMvcQKWUOtZyZR86XELzdzx3PH8rcv2QSw8ASD9IlU/6xEW6112jc8+ZM
NKKMuuAgwrLhB0kE+R+oTqcTs3o0xZ46FOTqBAAkgNRNuqsPdWKeJFi3ijTLzpS2
EhAt2467wwsAlP4wH2xyveY+BAoMwQXo5xEfB4hAydu+FqdY4NRFZtojqHZmejoi
j605mVAB+tZsShXlrOC8YEozSCcWmzFifRbN3l806bLBOEnLWcWkzLK2kqq3Y3mt
vIPRcDI+LpMvjMTEu6GPtIVv9Iv/OeQDmi8sn2wv1rPJFZyLHV7wV2LGCXtdzAnG
GB5cIK1F95fiJE/Juzn0Uny6YIt10UaFpOwRKNKO9kHWz7FhDvv26vErcn7avYTf
IPcutvpwdWyl7bwE5pxr4uO8E+QDX8eFxq4QIkK1XISVKAo57cnvMUKuoDgr2rT8
60EbjZa2iXhGfQKX18eP1dZIu+zqQ4meOdGOYMG/WhcvGLbdE/Q/v8LK3DqP8lqc
VHq49tW2NhJ0NUdVf+GcBDGy/7ZhPXdSWkbTr6L6P0bjlMbiAGuLvfNGSK3uynYA
tF8VfAiz2qAXamW/hml+RJCmcoByaIe7MFHEof5ThUN2FXJ1shf5v5UDPPEeLm+6
y57fKDuJBqEXvHQaVTYqcS/yYZRKDx9dWUNgv5621LfS9SgAyyulgiQB9+xX86mu
jAZdbg+g7bwd6Glu0oU2IErq72ll59y0K7z0C8mVoM5yIPmnzUBmHzi4W5bw+Q/P
6stREmfk0RcHs4IWKB2cGVsGbzi0kVjELlYAXIZNDciPtNSVboAQiJhqMQlqnLjr
N3DZ9pipJN2So8oN+v8lyMpe7+dEu6TlXW1mYHTw4AzrL4uQeDrI21dz7kxIhmO7
pixbiR1cTAy6YWj4Y47W+FIJjGC9dctd09mEyJqmQiP7IRNGEz8j7pEZ1iuOEV5q
gMjk6TjnSh6pxCYQ1RAqdjqAThT8eEbDRPmRD54L6RGTwenTimSvCPGqnZJeyrvq
mlOfAuTLAVtXRaE2g9IOZViDqW3xPfOabkyvMJerPsvwBXW9PwBSdDGKNK1F1wxe
vygEKgat3QVto/1fK7zHOJzXY7WInS0ErbzJ8ijvCnDR20VSqZ2tBkVwOvPCneWb
ZiCvNm5H7jju4PpsyycHNwV/IgoZry7S5FyANWnV7d5xWjwnERviIPrHhMtYVI7N
9E3xgsaiZeBz2LHgIt4Nlc5CXNnH1WkMLXihjkYBwgmiVrCY4fRJJyYaSqJsFJv3
3bdoZu1EYhiS/uZQjcUu+2/4iwGdw4ZI7ED6gB9IV5NydNfqA6aKxdK9vX3JBM0z
aIwK7ovFedUbKwHyEBvfOr2ep9MzvgtdtNdN1F0qvdg33NQdcadVyKJd4iXmzauc
HimrAsKHIVFkWs+B0tHT/i8xIVOEgoo7OFLhOd5qnf0jp+4kfcYqR7xkUQHG4Pkk
1Pa1e4+xF/f3sye2ROfoifjJCWjxHhnn1UzkwhJaGXoNMrgHu3Kpg9CgLRJjbd17
tnq9Mcqiuh1Blo4ERaDFEsEpC2OjmF/b6R+kwxZLYwIQvNtabkVogK905h271tl6
J5COU6oSzsKPHIxh56F8HsGycfnmw7x3I5TL4D0+GC1kRuc/qO4Gty1F9qaZRCbt
goKc2ICTN0hL9KucRyEiGOVffov6eBFDdAPZCHvhk2zYCD3wyXlZyaAoRSOHMKlK
9g1SZ8HPS29puG4PsgENlGIZ1MmVjq1aDOv1DyiAKqZ/WN8K6ivOnc3sverJ7F8H
B9JSENSSUVZEc/SpBK0HDRm2EE4zx9uXj40MtDtgiydWQQfZtEXOVU0P04wOJUHo
K9R4Ncwv7tMA7kdAy168cRzHJEZ0Hr60UmnY7rXTOpr2h4oz13q9AI1VIHC7D+LN
g/TalKXqxA870kvxNBjqv3jAf6lbz9VFkBEpAzbicndx0fcJmhoLzw+qI5KHi5/r
z5zZyFreusmc3z43PnVSnXSzyEeqo3+3kRC2Knrtket591MMFTke81RGNJz2jHu7
ii6Ain6IW1vlJ7xklyub/dz79+MwinQtxHAnuDJxC0Qd99RiM9Wl8+foT+dF+sFc
G6iUuFpne/DERlix1cQ+6E3xJ13oa2a+8vyWxiv2PYRb6TO9/HHhL5Lyx8CjgKO9
3StmwZvXq6uSCUAcDGLiDdPxOcK9LKnkMFVHrdg/xG//OC20jDJ9dtu0Eye9dobZ
hUDnghBoT9YMG/Jw/0xf+J4uDsZF+wIfW5YsM1QT/7W9YwlSBkHw8g+FHg/CCTfP
NwZ+XbAPSizdheSfILVfqmE3qtOGRzRM/RIgn6yf/yqh7S1ELRnd9KPfibjPqlDs
fqvYgCGCLgTM3TZ/0FIYIL4drrGY2eK04mIM/PjnimZoWKqzTa5dSgnl9CBUIVQR
I+z/Jta/laHHZwfiV/b0B+IdKW3FbK6iTKzk5oayaAzGGOO5Pkpzq9WPb/tnz+Na
4vL6ufYrDIyi12KIAhb26DPsW51g7xU3T+o0wSSlvdpLC42sP3U2yFGNdafaf731
3Cedw7acQIzWFB2EKc/gsYjt3kqhZuu1Y00o7Wdkt8WWQvdxmApsualQroTbUqXk
RUYvGODleZZk/VZNO77RCZloz9Q0+SVvyfzAH8gIDdLbjj0aT26ciqNkPCgVP17d
x9h192mDp4GO2TIpY/uGk1Huli6VyYGiT46K7j4PztOyrijmARkqZnuhb4FlpGXb
B1UyjjXaWI+PplljyOgXTAqWmBxkeJ326c+LRYWQhaGtELJnhir6j7LFKTYeDb8A
X+Ce6jvRDv05+SFnrLKgYsg3bcoQpfTk49buYDZxHnEKGyj/r4PjBJnM2/QOL5N0
IQA6BTVD4ovNr6LnqE/eCnYVBCdLFNsU3OyjYoxpT2l9IOhGrFhStsLU7cQCPTNn
d2C1VMHmXSc1OzS/bPU0txAkbrrcVKZVIB5tyMK2rtONOxCKQtpApzbCIAZOscZM
Fn8qpl9AkR2xvkFZScYrCRLYZl8mCy4tS6ZFZXLuI0Y9t2bpEUqjvAvXR/3rVYI8
grGpub6kKrmzsT6HdrMWu4L00WL91mOOBczxkyLhUJNqIfWgOyQNSLskmVNAh9JE
LM+3TCs5Ln4VL39y2P3XpCiclKVpvp0jcgDlHQQvXofOHyhlOtcqNlZcqf5C7SY5
aTYf8Hd1+OALONdKmZwL0qlRj3NDNvtugsW4+HYRWTQpTxC0J3Cpdm/6+9U4m5Df
DEmzheatfLsjevVjKM/R02DRJFcC0DEcaxKs908oK0JCk0ZlH6yAjbUiNqeJrs4o
9TBKLb7lWj5/4tbhMlg4n804qy4enIRnjE1Ykl0vP6j95xdYkLogcTnUwcVE22oA
6bTy2AjTPsJYquP30vP5pR/cripY346zWlxqnDFssbLoMDIVcpY+Ir0J+2FbKG/M
VUpJgQ+n98IQGFoQ6kfvyNR3UIDGQXxT4vYjli6tchSKbqWzUJxTzMn/Dc+oEVzs
9MwWaVPodeyD3/V0+3hLXmsiQHURvUdSApoJiats/kfTWEBBLjQ5RXy6LQGZ/ZBn
buiQWnLkXyyYTnHm5nTjw6yeq0KQn1ghQ1obDTG+skfsYzT80CFY+x1+2g+sYcnT
iGWgQke/MlG9BM3B0fF1CAQePjIfzPl3Km1z4g9qv3eLrQtxeeBIKVHo35BETZXT
Rr/B2YYL0U/MVDl61scIeFrN1paiWf+rcywVHVDDohFBuEMe/j1Wd92Y2/pCcRC5
jsmV7Muab0zKn6L0qsYiTm5xRuJRjpQ9mgYCBoD547D91V8/XVwcxTGOG3mF0jL7
ys+epmDO5P2gXAav36de7yLn51P1I3rqb7GgIHxq0dnK7qytEmSDXHvMyvb9F6Vm
SPr4bO6+UL6QEhY40EIiArPsX0vbE5rujoQ9uTEPTn5c5pCwSoqJDkhEHdBXS6Js
1egJAMOZAGkMlSPgNxIbaM73KFJZsX5JH5XhmzfxGklgFNMik5Mpimk16Ay47pcu
zFvEAdvxLDDoavQFLseDn6+BvH2TkxAn6vsHOoBfRzVFiyNpSgEcPkoFgotGLSsL
b1Ecmn+AOUjdXlfJCSMGfBT4KX72SLmyNb3qgyFJBVOe2GaGr0TEj41pQ3rn+mO7
fKaeQuNszFLx3CtfNaHPSjvcen2m+aIbLSb06UMUkS1Pem/Q0IYW8swnQasWfsJz
i913Py47Q/mXbyqCdE5+2lqBEjoZmJAxUtjPTVLmTNo8oE5GaEQJvBSAD6LQeagj
R2KGnQGVrIxH56jsGZcAqn0Db5upyaknM9yuaaTi+996ZVc/PkR2KsC7EZ6yp2gh
obDeCbn992X6fgrpmKulGgLnnqHJrm27gI8wT3t2LNOM0h/gCj+oaNxMP0mJEKJW
FUCbjuccuMPBAX5KKEsdOdSPRB2L92g+u8Kg9TYiBJe4RnTQwP7JdbhBjQ5Ke+IC
vzNWbZpvuBO9YaCu/JADft8+fJeL1tmArySTk/8Vdd5QLUlOQ+Stz7D7fs1direF
ljKkAaWCm2RPO91krtzqSKl2569H63OEFcaY9CXAkaUiZ/T4QEfR2kPTu9AqjvN7
9JrBirhuyO6CUxY1EFnoclnU2cjqamLPXB/VB947urTw4AQdQtTc5fXOC+sX5vog
aBT6FmGrzrHh56yER3fII9A3vSaJWbu8ColaKbtdkmxXYdBmZliJlHvM28cV1m+5
1YXcTZ/LHMeixTIIc38IMHcAGUw6eUlSt8crUt0bPopTOEIh0tHbc5YtMd0qB+M/
0Hlcpbdwgr2BAlkKbxPLlh0wx7uIPDAiZ8cu3K/ghZ1HXfKTNWzrhDs7ewrYDOac
wGWkGRWp/0tsslU2HDVY1t6tT01YONtTJOStyjxUlM1xfU3aAN8DiaFQEMiHRYu+
55k3y39eQB8otP2Lx28og+KCntoXTX+0c6XNR8A3gyST5bHPIGS2tBhin0Zj07Ln
EbdrTxkArANxHaKzn80b8q45469V0QPdviunqTJqpM6Fxhci6yWH1KZ2JXq9FLLf
D9n3I0JEvNWCm1xFrKK1QhMPc2BqP4dTDiHTO4tQWAUSQs+YK0OVTPV1q29Fsw6D
l5Iv3UiG/3p1Lre/9kV/Am8FGKFQwTqcpqgB4Zje/7Ad6ZU3Co1gBP28Dh7N1Auw
P79QIb/EPCNmvJue7gDvqrVmk0HRJGtb3uf+T6+y3NUHCgKw9SULuPC+0JcmIYAQ
cXiuHH0ORTlKrUW5cuWnTVmPbPAR4sIXFVCeY1g115QouAC7te56MjbAlRtSGZ0x
oFXSKzMTSlCWMmEoEBJARM6aR5FnZKehsEcPqTT4Sh4spSdSNrksF0NLaq5xVELB
xRdMDKtpPC+6gWP20mS54QUYkOIxKmqtw9NDoWXGXGDGbHMDcG9hfd3BZsKuF9RP
S+svc6qlWCWydcTRhycLj2yA4VYa7OdxqbviTasCD7VfEP6lM9C9TKnGXddav28J
hhEzZsikBIVaG4arNu4TN/1n//7P1lJFVFrlnRfeHEhA69D97NmiVrjCNw47WUte
XWEj2VuFpmH5QKt/3Lt6n2edt2VVojG65KDqaEySo2KUgV2D0/3Y3+buZ94ox9fo
Oa/A0HzWbuq7VVZPsTxAsV/c/AZ4uFa/eHM72LY8CnIM/NZmXXEVqOCtRulNIfCM
mHhBLI+gmbkBNDlmsIKdaHvGrQvR4Ahk8gQlbAq8jTohVaSDf/Uljy9lmnCyHvUD
g60a6Clps750UMubarhv6BB3fsbLe7RgZzFbtOLTHFickqXHnvFddrvECxjMasAf
VP6fFH7r9Y5Qoc4SfVqnGy405YIKkX1dLtRSh/njZYQeWwAQ0hzZHlBYASqbgoOa
rR18yB7EpCVn+GEYjPr/9YVk02ji+MI384oKjRlaJFxJj2YPIk4jaFdulCTMDMXe
8Imq4DXQ9HDEhBppHdde6ZkwNp615+S9tkHj8o+JOTDhOcOtAYJpgTIwqwdVLDqN
llImuK3N0GdUpZjwzkIE5G9FMYTbS8B3hYClmj1+K8Yh+lkI2FM4nEd401yqvnfy
uFJlX/GpCCsfPVW4N6Iu6g6aSks9POnsSMrj2MNDwkmy0RgAy8XrulJruI0c5pdX
pWkEPOhm3NEvubxc/qVw/WUgetGBXPgxZCmyvFAkVr1ZljqKs4DToSJfYJhfrIf0
ZnATWevIQiHCrJHptIrAWMVEDJGxngdHHT5ekufS+j6I+YyhajhcZqW0cyYf/iHY
uCKYbFcyyS08IGy2PF2Z2y4zZFh7tm9KRXyYCsgdxIg5FgVw1UplCeZA111y7KlL
re3mxxSykIM+CsB45R6EJzxvrZOWE+TTjl/uivbAauiLKw5Z+opS4iiygwO+p9JR
kFDeeEDa7Vj3uFQEWIfdl173aD0rZiDp7QDtdTVc2IOee7guZK8MkTBkTfsc9HSL
V3+QVg/jf81sSyDbiSEvNxlIraFbRBMWfNSZcawud3BXswfXNKWP5daCQNLoiOJI
7UBXCSw3aojk4glFc0GaLHnlUeOtv+feq1rUlNIoj62J40q+ZTlSaT5AkeJOPZfM
6zGVu9qJRb/sx6PlemfPhj2Sj+vSRMolkHa5SI4PTHmDl6qEJKMblKUf6+A7VHIO
ZWUu0j7b1R4aQb4fP8zV9qUewNRqYgFP2xv8YHHcFmelLU1jqb27A1w6xkMlfSFF
6w/cSaXqwbRbTOBiO663HsscRcY3H707b2m1L6QJ0Qufp/t0O0oRPer1PWfM3Sv1
lxbIXMBI+B20FWf8rHISvDedjGvEAYhfUPIqPU2WURFiEEHmrqPBZQyFsCV3Y8Jj
bgFLoKu3+PZDsq7FuwnZFWbywJyEI9/+WMxBubHw/HBsyO9jmtJiJ2h38eZpAObX
O/W9MEW6HG5C1tH0JOml4ytBHPbCFh4bn/d+gN1XbF7djWwfJFqvFFwF6ajvV07x
pc4IngjR/9A7i+Yb7jIN9v+iYS1ZIDXlrPqMuSD5KzZrHv0V7lfFpa14hc6wSOB9
WuU3uQQR9dqPQd6z5ROXislQbqZJ7oMMqzRSbcSmDAC420QI6Xy5FWWJkbOLmPHu
7sPC0P4K4AIO3isuhgBuLro2g+WPjLUYusUYyoeX9p8YHSKO+eOuZfFo7sdG0o/C
qv8gmYWFymYYocsM0PmQrxCkCWoPaCMAEmGniBo0xnWs7z1qCLQrDeJTS5ZLs2AQ
l/pRHJmrdobqMHhNBIKM+VpO2GdP7MsQ7A9gEr62gzr5hqAhfTnkzL5LkB5o5pyU
FMVVIiH4pl5ePe/le4lNK10E6U66R1OtlYLNEByh2UYjxhdx1HX/MmhGt0VSfc2p
vzt8jV1buD8Tt4cW3Z5sk4vfE4uNqn4JqcZ5NzBDPCcJCe8TrcvtxW7cCYCu9Z4r
JQtOr9g3uVQHtvG0df1hHoV4y6lDYS5imRgGo7HPg6TcB3B9adEYL0wjEGC8cVFg
HJGySPLshLUmi2xh58Zo/sY1CFEMf4lsymfU/Fjmz6tiXEyY/9rWVEKNP0iRfvYM
SkYRKRMypJee4CccEHNG5Sdgsk4tUcjyiJUFM7O4Nbz4kb69S+HrCQOSgrHsDvwh
bfyk7AXO4iGJrlwXfiVJicbn58zjz1HRGuLuUK/4HC4dW5CPEN/VF2Koe/cZ1tfd
gX5Qj9NNHjyCJQMMGiuc45uhxFURunAffecrprOi+7VIPFf5qOzv/3XP6C3Pfnsv
gExUZ96+PK3ehTl9I1cw1/IDWcCeaVlrjVL0X5o7It/+pdvBn1A4YcISqD32LXQl
YnCZKSMD6XE0hwZlFdEv4nwSNerFjBcHgiotkvZVi98zgejlZ3giGpHLB7halkje
YYjYSYBRwcduhPPXYUg1fpYPVmub0qlVKMyE51TlTrFPHHfAdNZSpuH/etljI+Yc
5eG+Nr1hkrNriA+IO52lkdcQ15KHT4J/GNHCCFaih9149Bu8hp+1fPJPhtNsBXY4
fXBzVS6M9FZj0nNAdE29VrkPffpPO4UOLNUkLbmLvcU6cnSpaVUKHWgfg1juArDn
ly4mYLrhqUiZGZsmQbi3HmugpFJ8+gCO0RHbbAHIOhNLmmepTd/GeWI4FS6JKqYC
G4g6ZV/e3yKoKfbRTcAK7p8yx1ANAJXRQq2NHOWuN0IeMLZxW1Q4uANjyl2UT44V
NrzyQBQAvH2U96j01xVohIJAW8kiD+p4FW2v23ZcfrE+nOYa7gnvZy6ogy4i7n0x
4NRrvQlenL1gFf8U9YBvYcQjW5tzTNEWzx328g4j/I5yFbrtd6h0yBvdzKt2SX89
VXry5xr00tbqH9ur63at+CNkyzNPhV62HB78TbwTvvgilWGDLsVEka1gnaJb28FX
LnAvP3lZz2knXdZkmt4WJs5CZw+HeFAU0+7JYZqqgLPy6quKZ79tZLl3TX8DH2TG
C0mKtL4OXAT0RKI+2+Cd6613KpE6w1GfaVjadbtFzU+vxErUwy0v7z7mrCiyisf4
hyZ+OdVPFKAQz40/o8CJRox9sK5EprQvO5oAm+IwhuuQSsIlVEDiJfhJWjT6+uwK
u9wguflfzZGH8mYVIOeWsHjZtFLRd7OfDtVKQkFu0WCncqUmo4TgHfuayLxSEYGk
L7sK07lEnb+MWnsuMixYIHDsLofsIqP5jha8wTCIhglUVC2m981pHry1ARpFUQHF
NaZTCMci8xczUXri3KccUAtVmQaESc9h6l6wZoHcc82qHOtsMHMYDfkX49TbTZtL
dw9ArGD1FHglSNkJxvJFsEeuCAnAAZDMYgDnuAtddE4Yk8XhjfvTvgpa0V6/Aw/C
TaUCM/deC76XFtojftBwae/KNspH34p0hgD7N5DR5Ynl9KaPXltCMmcaTu2hW58G
7+4clhSzzi4SVzsy7yg3MZDNv5gL434qkRp4vve+ZKKr+97vk6hNLXZmktlkJqkp
OqGyV/uwoPOVaejJZM1S+3mjOTkelYeI5VfoaKv+zMwL0SlOBV4zIxZ6024+64p5
89bvrVU5jyT4oYrqMZR7UYT0JaZIRwPIB6KGh0wG2DTD3LCgf4At0cHAJBXJ8wlx
wHXrvkjhHmLMAFAc6yjUEllic1TgOr6HAmjLLJXquC4fnDRn9P3d1Soc0UF+QjkX
peu7EJ1Orr9OollqVVYDh7XqFM+beGANfouQiIuRKB5VxHhytQ3YnucD+oLYHBTa
E+Y+Ta5rmB3ZfbSjnH9JAGY+0zOVQs6FRY5BIKHhBcAE+Ryqj/87C6VKZQ/38iYb
fTJoSHhZSUETIg9vyDMB9RRd3hHVnIZWZtfZyH1nsWWathvT5ajcGmGWWUDRdS/n
ce64twwL7Wwo4K1dpixIfnsO0C4sCj2vs34wdb/3qvWPwACTs3MzJsDCAXdXHPrI
UyehyYeX5ecAdzKIDclK0ypkJT+MrPXOBPyDxLRUmScbAi/zsVlFm8ZccHhZ+lbR
yOhkAqWDIC0oSil7k7dF7BBQhTcrIupGUNS2Be5Q76BlAajH8q2gW8sP9i21LQH4
y+/rU53bIM0UmvPuSHj3aAO9Bz5+WuvvQN+dH7h7J63FBCcpCxoTsrUplhMrAT+L
9b+iSPPAFL8Tymo1mU6WB9Kdht43cer9GWIpU6mXGU3179MDHS2c1vPrXzYIajvf
RSSCX8DHtOpWcj43W5YEmDqLWFuMEJxF0/f9stN3YCKxLLMCq5BjpO28466nTykK
tA2YMsEUXHlrnZh/7N/vNC+XF+BuT1T8Qo84c4ejP8drVxockY6oG7QkM4sYfj4i
W6KsByjOT1c55sBva0T+cdwZnmv8aIpJTTZCs2fecTPLZE2cAGnpsRRM0EqqK/k4
tJvc4SwqVMOVjE9FPtdCQYiZMgd6tfvJDImyH27NbtZrz4/T2qZFV5MgmapHapac
LA9ZWdtQXpvVzuHkaBDw1U7+wl+crViZBaPTHQF8vygmYIFp21l4UWFkt8DfAD0s
ikBHx7f7Pl7sj7v6ukH207SfPaL+nG0H6FPcL1UnTrPIUsCTbTcQ+POslNDHkynD
69XvUgPs6lTweFW++Sfb/XdqwyzE9V0EKNKWrpLfOCT0HEjJi3u3ChWdB9mMhVjg
r7M13dmLI/CobQAaLBPCDc+a0nuFHiRr3yvooY/KIAJhQp6yxcGba1mDjzMZPQWx
fJ4JJFjwrvAzRp8OVOFuWZoYr497JYCJ93JKxLFAZHZJi6QAXxjC+SPBO7icYQc3
9kdvh1Gnz1q3XjjCWXmEpXqx3Svgs0fczL/7z2GzonQIpI2BdH4PqG3gKGMct15u
pRyosLbuQrXrj+3UluAjDXa5v+1CLuDas2Cqw2Mb0KfXs8rzUPYa+V8qjuzexf2Q
tvUXbbpkMuJ5QEvwTJjb6Ez+DjugXiX3yuKqtgLNTZCIDEoX4duRJy6NL1dhgGmI
PZb4G/f+qVCeFv46VJ663omDmhWlWGDwznT76e1XinPnbScFkhyE45uSZwmFKk3U
sLVnG+TxT0wbu7v41lcIOah2z6G5FWfbd+y1WEMCsrc9RXfyfpjWEprv2xDmkypm
8Sov2V/xW4uFXp9yWeemVVBG5lkxAXunQCeOo3AgJ9qEWaJ2PMu2UaQ3dP8lLRXO
doGdO13NW3wl2Bp7dkK4DCCqtbv6iKsAODvwn/HOH2zhNba0otDVGUZfRJy6aPiv
60+nEFaC+6yiV41a0uPIpswQNUWw2KcQsfRxNPZ6pBRpNQiTnaRODiezG4RoBRXS
/ZezpvraZYsYzNqKmXIZvGC+bQhVRcdRu70NSlTEy5jmjJtrlxRSHenSnCU0Ilbq
wjBVCkC5fp5MV9hQqSYU46S5e5nD23op4sOXh+wNaRWexjxX7gTI130Hh67Tqn2/
8bcdrssTzqYU7Y6CP3NNCSPcwMv1tt6NbS5UxOs80qzcXnu9aWN4Qq9brfTd8Ad9
QKvvfFgIvQn02xIJ3hgScH3u2GWZ1ZQiipLjF8XBn2XeAY4oGaN1qgDsqDdLVC0F
ks9Tc5KiqYGylDiUerG8cRPhyfwrxmh0LYQslBdm2R8xS2DAtJpdXa3Q8iYocLtC
BViQLAyura5PS/hsF9vaegIT/mYJjmwCZL9wI0oERmvjgD7PMuXk8A576Q4/p/ky
8x7q+/iyrArGRR5DVlZDD/Xx2S4pGtDx8a3p4DynVq2jvVXA9V0PoYGotr37dkoS
uJABdMXRClvvG5KKkTcaIgclz0XEFh2Qth1np8iOZdf/ptiLInyR4wUD8PnEKBnT
QGl2lK7CSM9kCF5iM5RF8RlzH3cfq6bDICu2kguba8/xBo1X6s6b/ZpoDnO8gh37
sla4djwdk+gcRFos4zHWjArLc8u/+XqO7p3nnS6MpCqb4kdACLtb8mVqXWgVBhtO
F30PlMhwohlU1e6oauKeCWmRtK0ld+cxJ+VcT70SM5047OnR1A2CvONc08irrRoA
O9/F5gGesWmScWwNDmSrWGkxR+VbVqg+xQIZmFXBFQjD/HcRSZ3/LexDwGaYkRhQ
4cnNC11ndZax+byRt9pF9zO489t2tzYrq88PITW8QWrq/ugx1urobS/vMDTqfvQq
umG3JG+U2I8CMZyLl/Gs8pGJKQ/ulQkiPtu8TkIf9urSS0QmtY4kFhqYBKaGSshl
h+NsXJ1HgP0soTxzmqOsieAjNENOFulVaGlHN25z4pGOuenlAXFL2i7CB0gSsk9/
c4MENlzgaQfo1gvC3oEB5gqZYPDXR8FXBQC5YIJ5Sx2FNKt9SLxZ90O60aktubDQ
QkryFZnD+FZQvkuO+7V05gGl7kQHArFDeh/caLVXqB2bIdxXKMUpkX9JlcIP2ZZR
7nkmAgJtTybHx/dp4/C7hGaTRL75kNnR+LiXs0gK37Gn3zWnxhV1cSN+sJjbogM8
V42uYLQH7UUc1KIpB89RYXJLNKzOyghLRWmBRwyMD+ekZ8/kOz4wcDi7P9R96ehH
ohJRBjgDSIorqWjFGDDZBVbiiW9ht4NRBPHAp8WjlfkrkZkHVO2mF1wygofK4nWC
SStK6NJQLsiyCgPXrEypPhFU/YHTuv0nqKyaYrPg4JKdq6wbUYHcXE5AS8I7/LbU
+XDe/OXD64k4RE/VNEGRLuVaD5ODnhlRwVBf/B6yOAbi7Dg4GKCBr2ZqjIl3vydu
Fpn9dXyTUd96o5XFWX+L4R/NvhBQlGog0Vj4NJxORu/3g/Wpn9Nxjd8ejyKZ+eFA
RA+aShwN47Esn9d43gjHBa8PRppKexvRmNjXl/15j428VdjhwYNIjcfniqRkXHvT
PLZAESGsd3bYCcGHncwxo/WoE7/P/lVRyn4+hLIlnbu2vSHe4+B35povjMarSJ5I
UIsdNJNbyebey/G5dNHZ4iD1yEwIeJd2f4HcArN0b6iV6r+qUzwmqXt3b1Gp0mlS
fIHPHrHysu8Bf0/OoAjhKn6a2acMxSi0WhErxECT1GBfRGhlYAmQvY07MRJZHbpO
JPVSbPY44qlwYu3kyUuofGhGHGZhDwUuZ52YROTRZvqVTiuq+QwgfvsLnrPHvW23
kBFtD/WjxXvUGnvcqcO85QrW/J16EnG+G1C8PRJpap25LIsdDtm08+soyuWNBXF0
U8aza4wBcFumfldMdQOECuPwEXKOTWVqL4HTyV3poF4DkT7fAI/JkjnIB/3Vv7CW
W8sDKC7Eo1i7ParWN2k91MTr+l2UuyVkdUCk/rYuCxh3a1vBAHk/4xGadZlEWIOy
FS6EfCeaKqEAXeWLrArn8I9GgFsquRaEU9A79Qe9nu8/qNXI2EiJE8p10kU9DckJ
GtyGq4YC3Fu2N486qNewxrkWSs1Sx0AKUangtLrzrOSgNdazQA4oLkaGswATmfw0
tvJRP2Rdy9L+HzWGkJjDDSapoBkTYiII4vswZaDC+/IH1DSpL6KXXy6qlIsYwwXL
0WaLsR7qlAetsT97xTGP6dXpkwRm+PI4gxJNEqXREg4z8zBULTOt7SfWgJO1SgJm
kraoYF3ED3YqtqRPpIrjbfAoljU2dBz23A2hJIbrIpdNpPZxZXjx1bHOQVpV93mR
2dnhF/TL9IsHya//ALyvLeNXeCK/KWiWZZxfPVfxGT6c20u+hbzJTzdGNRvp4DrN
eqxn77SqhfLLyFJZ7MmR7m4OewVn3X7BqrBBqvYRCGzGiJiwI5OiJPIhFHQMS4cN
k5gu+7BX3DcUswjAGOfUB5gbTAfjBeENfgBGWjuq2eDApR6i3qXO3R2G8jkC666z
lhGfnajOwKfk79yDoTozLVJVasuT7pqwACfn19WLCsDSRqUAoIMoVLSkn9w/X8LF
19+vC5ou1AiCA8GS9DzmGu+y1aUdWPewgO0pSV+ceUftQ3bJvyDvFTuCPCKAhR1I
Bxye1VJGhrP6JAd/M2imbF+9e4Tj5MZVf0FayCU2DXhZKo9oBPmXZ4y3N4IkzaYL
BAGzM0OgnkVs+M2E2Ij33m/5o7Tl/DVss4NPQKn2KJ/gRZwG2ZiVAGD8eQJhOVDg
rkBareaQqab/C2Zw5amWP9vmwdK2gssCu+PzJMHvaS3NOotg3zdsgWglAaOv0uo5
wm4L7fi/a92X2xb2jOX7pf0qsntXG68PRvW4RNG4JXQmaH1ZniBqSluOE9k54Nz0
dk9PcuRWXALNMuExxbhrXPtFFjPM65ydV8RRUoTVn9y8qgb42wvZIrWim93lO/6B
13RM44doyw8qLCzIqzl5yVYNXfr6TImzJFfkYMr+puOLS56a3wVEOGdtdNpbn6AP
OZRtn68iBp/1f7AQD+3w9p+GVwecLEJsGoZgp94rl37C+FIyt1IYeIVPJf+j8xrO
kseueKBbnlF+Gv/t0TXq1LueLMzecFJI1Ct0B09PVUPR8FFymGSs7y+lHzeRRvso
MgRC3pWBPA9h8OOu1bWIW9q2VveH0vAilmWlNG8RiZ3GKoAYT6seyjyt/lcHLs25
10XBNEhU34rJkbYzWPJg13dg61tmv4i9lH/iqCWI9JKcxdh5DI1QfNMDocczfspS
saM9nwidvLEXXILCjS+XJ+xgU2hID6gVhOXXZaNJzwvV3rxAsehYA+w9/YZ4tZ2c
vayvkhDpR6Q15ZYNbcI6Ak8/WnC1VTIVoBgSFesGlDC3Yp9LLj/HyNjbyUWbgmH0
kLxfzxXEW+gzJIvMh+sxRDOoDFSSCZc7jMt9xmmbagqNkmvr/x1gQdAwgjRUY6Cz
H9RgwPdMuvG6fJrj3LafRcHFHQsd4TToEl99xZ56tlpXGzMPJfQWY0Em1Z0/NK2k
Vd2pExYxVGrxhq/T22KocN4RaYyJzCvChqB+RH7bZH7lDyIvu8lCQaspQIshOYz8
YuJFY3uKCyYaONREYR6ms18tSn7O9sNddxhDbtBpxeYqDC6pS6B1EljwkU6fA2Av
TicHLCwY0aKyE7tp5+B7CvVuNymlSWiKiEMCIDn+LGC4jypg8VpD84v7+himkS9U
Od6X/2ljOsyNRuG+5jUgb3k6swnFEHrzFSugR5WMEmr79urUpvupE/i+QmS/99kx
XVMHCRMxRPLEfd5xis5wBRMWiQJTuHE3kGGu+EErMVuUiUtMPXmaVUsx43RDX2Jn
dKlIT9vqfYC0HTCgjzzQjR+78ZmLhyPFKU79iTWjtN3VdwcYEONR7F04w27uRCDm
rXT9gFlvJo0LbzZBqY+dF/TQ+JivhArzXAFp2DO93CZiU2WQeBCHFYNKeCBuXxUS
H1pWIqwikct73U8/RLpCBp6LjYOQPGJ+FCOUcis0IG+hYrBIDWynGwLWQIzBhd3J
QZfZRfaP0S8gH/K5mA1veL32lBjm/xhgyQZOiQar0tYm+3UCPBIIp7ePdM70AGXC
aTrU1VM3IuxWHc7StOJvpcGQAS3XPr7o5e55JQ+eAvaL5HZubxpmxgT3Nj0qp3b8
5oD6UaA9oSSaiOKDnflMOvbyPk4nyeRN4RyYjEMQ6m/iGqeFCRXiLOEXBgmIpvKS
Jk4/iCEqM6tn3X5G7KEmz7mJDcfauZr/a6rJSQZFdtlPFHXFnJUK+dNzJrPL5pOf
zl1tYHXhMUUQAhUu+wBu2u8fyUCg4JerlUULKCEBEgt8ommQ6KnBSWtOkM2bYXej
kvRGpFFIm8CCDpLJ2LbJAB4wiBf7zTWVWBq13SZKNXQAWupEY0IBfPJ2f/luelUR
O2vQ50+JGyLF15hpNCSELMoXXLKxPNM//YozP3a2rGpvZQ19JM9nrB8zpqFSdsQw
PmDvm95XY0hhNnw+7+69l9DUaaTlCCuaiMYxoeXe1DpJMWTCv80EiWjWp5Rjzlz0
HQTEGo0sIRrQCJtprNXS29vNLJtNibFd3SmCKoj3NohlgeJR9VNOTXSkR6SR0KNR
F+UTvAIKDcB473jzNkU//fLKO/sJ4O5rGgH4j5jyrGMtPNEZWmP0WVVOqyUOpZ9b
BufsY4y3m6u1bT+tVqJVuiqJWbsi5yJBTznc2SFi/JPPzg6/BZM8r1jCC77kTk7q
N4n1gEfrn7Vx4iYuBXNgvcOGxuyoaVU/ky2oF5dn+n+wL4jcRNiB460cZFEOcsAf
zKdbiPKaaaBwOrb5xXTno7PXTmcQmaHWsuotwNTd/7HhwOfR4Skb9D3rZHPMpPXh
/xJStM/Jw+2JtJIAXXSEaea9G5qO5eIs4mCPm8x82FnxCHSHtQvbDCLfTQrvNYfQ
Ly2YANTfpk9MPKC3HX/gIyl/naLoTpYa6rBKQ3Ts4dWvMybPCl5PmZFjzT11vQBP
UzPKVu4j3uoUMFgjslVhHmf9LcK2qEtE2/nCpPX0ndo0T4/Ckrfi366m8wajtLiB
u0lEBiHKWor1CGOdcj/PK+w1vCXgYRV5KESWyJY0OSLcH2pJCzwQVme21/ooaxyb
5WiAIjLHeyPYEV997Pk2Xrxp4MXf/1xrkc4fhAnsEJwxMPLkQXjeY2+4K1HKUZ1y
h1wj5sAjx2+ZionSk+6hR07DJVXtxrStYZsnlOJw2waI7bFL2h3VfRQG2QqG4maF
ruQv9R/flWDfQXpVpbcSZSMyeBzRoZJ72SLzX+OUF3FjrOvwBPz1odnmiH/H/+4M
xCJCDpn6T0s8c6ru02b75ytwdrFyerIWDa51HBGsOnvWA5meW9VqRKBi50XETMnP
vV/i9EBRepMdv6Y9CKlEC/bZbg2ffeDLPYZUG6fe7Lp0Cg9IYYtdo7CHu1HSB5Ap
JLj3q2OJYs8GsldhIwfbzSGQBWcRQcKVHQu++/zOLk3l8O9ar0LZl+LWTZJvK4jF
JdSiEUpGZhMLJW7MbkSVAKOWx2cvK8fw9nvJAl+G+oEmPe5tBBPpaN+BtE4TO9nI
U/hgh2DmmmO9JF7reiLS4/blIgDppkjYOQt7sqUbBkDwkN713onVLjF6fbeJWieQ
eSisnFlrywJJUyVu6MMkZp3Cgg2fmwMRQ9AFZ/edQS/LaWywLvBX7EG+e8knwj3y
kd+fis7aYFtM+o1pE+JTy8D7Kzk0KpnIPmA+QDXgvH64dDugWi7BWkk2mE2jov5+
tn63NcqeDAIWMjpUF4M0K/157i1ji6J25ByBefnq7YXpXntvC9FMvNK7RdG6UyPB
0v/4Q8a1sdE+XxZzBN1b3ix9Vw0b6qcfmgmDBHQ+Coilss6o7/UOsYFDREfm02At
acNeo7yOg2QxEKG7aqQlzMnhtw0gR6YNYxEOdNwkoaz8sZ/FboDZ/eAbNGeVOmRK
VH8KmLN1VX9gzex2psjEwEjMjXbhXZgdU/XvkUa0obH5xtlvsGeIo/EHARQ9Gv2l
4rad6EExvw25dM0tSEF51qQrXlIXiMdaf5yti1ctDpQNZpgFkBZcux+hyXtdIi+0
voa2jMcvHMwPqPBVMKj3EBBsY/lx4BgzsuAGhqopYx73E6i6biHV0r3J7/QAR5Tl
M43wLQrNewbi6Kz3/NVUwhdsVeZpjUgfszNDBGrgW2LNwxbDnFRFs1S36cNS9ZMj
TW6wsHoASZHpd9BBkNTbkf4v84dTs2QpQLDFYuWMQzwq1EMXE3/5eL0C57UMHlxe
5Wtsa25d+PILZamsuSXm8DEXjZ1E+ouSXdYAVwgjqthb9pCZpTofY4sr5ljKCOz5
V3g2j/x5oDyjLn8AakyxOvk28NlbL+EF4udpqhJClGLPoMo9igNYmJhD60RSWWh9
qGEZ8POveDnYcExrUK9x9y7H1PfOxht8ZUX6TemhCvHDSWsN/oHWOr6tLOly01QR
j8tWZUbcQ2CfXFhM9n17i91e/L5572La46d5D4tKrYiqixdYuMfGO27wALr4keMX
cMMoPu1INaJaJf68nyqpMadZ+tg6U8255XfJhE05KLgU1Z6XYhOc8FFYdIpIF88K
GbOhMn+TnMX9hG8XUf0gac5b1Gd5X3yVTpylbQ1sI53G9h7D9G1EEEOG4M8h29GJ
R57X2GSkheHBwZi08zxedAGw537p3DDFdkLe0CAs5RF1M5x9UZxpeh85SUr0vB5J
9m8moVLFT+oECafPHqiCh3tMMehKjIy7Hu+L2H/9Pxa30qjx8zFNIw1XRwDnPYYS
JJDSudVcXs/kRA/mYI/9STBshHvMb16v94VMPBlF0WKvP6rJBxtlmQSP1aaTvP7k
um/Aw2+sdY3C0wnpXeVz24mPrGwd9bdC+SgruPVCTXui9SHRQOGfEJnu/C8IbFx5
R7/iyEHTxHlPxsRiZj+b7FZBiTGNZ2ltcE4KH+mA8gbr1HeZRHowt8WMV3zDfYct
mKHkPj1c3f//7syZZgY1CGBzWbjWw+nC3K+lqrrxUkkNYrV4f8IcKZNozpxS6AmC
GW/lDbHWBJCZMJBc3M8ucJUJ4jovN9KVyps9RIokco93QPnuy2AYU8hcJQxZ09Pi
Z92KHgwQxPcLx9B31wsD1Gi/C4T/On+sLzGmX+Vd5YneIg2FpsZd4KrE1dynVejg
ZeIQyhUXmNiHsxAAh8jfkGirJJg9ApnARMUy6vVJ052REDKzzb62MqsNv6yDHJnk
Bjs2zWLVJKASK69MTEi+qD9sFbqNOF66ZvdkNlxY/tUzv1UGrD2kO+4FrBAcPEwQ
JDsXN/ZdRMI4lF+uww1tor121kVC0eRtCrAy1/ruCGDBE+ddQG63xMbFlBkKrI7n
wTmXcFC8gTHPlfzzbQcQE+fwI1kieOvtek913hRtpw+yjDDlPYKElCFuv1r0N3zh
ICO/sMBHOFpLfE6tKAyLWYObG1Ix7AKewCXmeLd1bD+CU9zJdAJMNXts0PjnI5km
nR/y3gQcbONR4RkcBwgOkJSkU5qi6sJAgPTblSv9Qn6Rk0hEN/7UH7xtUTxOkMeN
Ta5CsfznAcLkm3Y4IpO16f4Euo8FzjgHvdtYk4PMH3yZXYIGWnBRnObnD87bbluK
lWBE7JD7BZG5+dFYFkCKcFTfiN3JQXAnIlnmKM5hUXZXkvYpAtWUng3nbEPvKUCF
Ownm2c2U+4NPLOdqJJSxpaf9gNjrp+gHKhnq1BgWtrKOJZKztznYg4ym97e5419M
2ZBitgSxWWCl1Bc8M0PbqVLEvpbGG7WWMr7siNed6oTIzeaRI7CB0YkhpepmgCXZ
dn2YUyrGO0ZsYLk301APi0YpndeztGdW2Aoj4nvBxyRekXt6lJHxmP0i5NR/leam
AkDdeVyEzFkjE1NW9SU85rsDEktk8b0b1/zGT9wxG+ykxy2aER2ZXc6mMDHYwD1a
jojh6coilEJlCu2hpJTPgAPphOKXSrkkVQFhQUNsbMfTRrB6Wi7VWH0pyaO/Pjxu
h05hAIYyAaRwUi2MLNDqae2FL1o43YWV+asnv0ZtcGVUd/w8BTJTmqDWa97L/jzP
8pNXzrUSZwyFaWdiLXk9inHVLIsSsNJs6RvNf1vzIS9wMCRBXysorGXBRggbvJsC
9wUbg7I2RP6ygmBl5CnkPeKFqNOEq/kAyvZ8crI/blP2PrdEg1j7eyyU2ECsgp5d
STUMTgCiXW5f4mquxX0j6VHmuZKexLObXOyiG6f+sXNdlUd3/mhOAAvZ7qPbqbci
/mQkjHzdsgGaD/Zh7561CCxpRuXU1UedlX1Ppt7tU3XyTluJPw4QPtwKp1g4z+mj
zfbGI5lUVz0YQR/O2RLWBQg0alPimwwyiPFZKyaSrr/X/CJUwKmoJd5D+/S+Tlje
XhuqmWylT4LTaAjvQ7EN8DHeNekYAxhnhaZYdkTcqnOBPCpzOwhzq2y02Sn7S0TL
szX2cx7vRPCTP0PPYIg2vgsNJ73+ysfZrg5mbq2XxnbBGwc7VA4heSfArVs40z8I
b/skNfNmFq/RsTa2AxBp5qP1v5rUSJ/pZ/YFSVbrHMLEcJWri4cpQR+qcBoLE5do
B+gLVMC53hxMNtS6GVQvV/HVV+dUtmNS5QkFhe8GNRcnWkQl6xKqAUzZ8ioamtM3
Hudul0w4FyejKpAMrQvKVFZN7qZ72SlifmsIPCn4vV8+HauGlxM99Cf6jARlLygO
w2ncElpsiF84wAmnyJCXwOFSJZEUdQRvIGm6sIdkyG2mvwmmrhl8O2d1wDXf7WZK
u8RHDeQaUMUb2YjYwdt8XTSQ6P6/VMdFzKX8kIZVSVC2VmNewl/4uVHXpFQT81EI
C564eCrq9D0au2WOAPBnxoxap7MvhnpNb5L7A2JkD2o6wPCwi4vNZj3ddwhv4oYl
fEETZgVX9EB/vsWuksyoQyfUZAFdcAuawn1y/GyQax8G+l4XlmGehWf8kFlnKcJ4
5fe+ZXZ6VkeqgSHK+S+UK3ikMR9KVXKETza1VO7auSHYzYWkHKU5PHyEHFP43NIs
XZqRnWcXRAUx5r/7EUUwKzHYvdmu7c8ke6ibPT6jcbK2I2w0aIRxnhgLJwx0wLhs
SVjAfz1ydWddly2De3hxDlJvVoTBdPyY1o3phkWlAIQAswbojVa0E+E6s3coQiIP
xY2TtwCrrJAOFVgZLl7BxSfewRzybYOjKFM9rJlQsTQtapNqyWaKRA1mCpKQ6B65
MsNS5RkoC9bsPJS+s9+xrjhU9h9zkdFdj+pc2xpraSs9WCjxwGLiRRhGM+8e0Q9d
AnN7IY6n8s/wCqbqqFf/5QX27vrt86K/noprvhUyiOei0c4CqKvMCThtKeAcMTZy
fq0ZMR8u9FZhVJB46J4J/3J9eZPD6SEW/KOvXZKD75y2bqynJkA793smXb3hHgou
ik0MiyxAxWbl5a7HKLe5bKNxPBhcIyOaGTqBcVnKCUfiqOcQUdNYLi1l0ErOuGbf
+ugf78jQwuadd9MKW0/ms6828AVvO74Ov+SPA2TkHywbOvoFwfkHoPe8dHCM/k5G
Uxy3kk+CENiR3xg1zwmT9yjeEagecplfevXjzK1n6asHxRGsO5trJyfeb+zAjZco
85xQCDJ4lmMIvwLatHgbZ2/V6XkASuyrMuZYEPA5n+vXGn7bi1kqrF6ujLM8uYZj
b+QHO9aITF2Dy8R/72dyngLJFCvhDI41fV1sX8PIjylqn118RqVvf017EIJhYJPe
+z6vpu+0CySPQ27iz9uGNY30iDd2Oo4hK1Z4c4nhXxOeVzY3L4lsIsTErQ3/1GDI
rrfAU7Mn9CqJGuAiXWmKhKQAxxOquFDLLI5/kQaPjR8t4ppGi3Ab4nMtZcc6JqXB
FE65SqiycOVtWPA5KgdCjXlgYI373kIOLge84SB7sl1yDbk+ZwxPIqyQ2HrJG5Rp
SqKd3J3u5U5MzXSJLGMpDc3m9xRaHKJWb30fwQRaYO6Trq5mK3J7Us9B74/tSlTz
p6qQYEL+8IC/1F+4ubZSTYw5dB2VPe4QN6i/11O8Fm0PP3eIDvEBVwCAJPmxih4R
XV0DRuMV+ue02ZLzMdR74zKj+dqbDJaWX+/tp/hEEqKb421NaZG7C4PMWAgSh6In
ICHNY12vfXiqY+ENNWpRFCawqh7yWdJvh+WSC5RltMiUZhfRf6xzkW1rE1vC3Qoy
H12DKimcxi7Vtllr4OHc89bkC7UPODCVNegIIX4wTewuSYp7JFLLam+tHgiXe44N
VlcyQ0B9Sd/NAZiA7eulrim8oNTBVwQlw9ktXrPpHC+agYAUPH4eOI5fhz5YkHAf
r2/9r4tvVULBFaLJy6vVayipy2clAIh5j8pCRctk4wzgEZbPGDMgFMWIfhJ9wGLb
bF4V/5rOJl0hzLaZyxADzevnxiTBbFj/609kXCyCrohMdG5mueaR0UaamorHAGho
R9X6GLS+evLAO8FRXoOtBynd3FnupBj9hBYSoUoCKG7P4CbfnWQvjODMqX5fe7OO
/hOzjNAkzQ2GanhKyVA18dmuW/JOybzVJENgNEpLmaPu3qD/6pANdlSRU8QV7vbn
EKGS/fkllcQ/Cj87t7JD3oc+Luo2+8C3EWJljoDMWFn4Qu+g2Ns8yNSIpaL9VDYi
L9PyvUjgMaTIKjq008nP+qjfZ2l7A8uDPst1Yk/2ndZHe2+CEYKsNOVneHrjygBT
SCsiTrjHuIghX/s8S/+FGYoKQaYVc4CT+4WOfh9LkJug0+zj3Qj2bFoXklZOi0oq
ACVcZCTvWm2QO1G+mHOIMUX/CUzKvGXJt0v5ZdyT+mRwbCYSN+WohF6Dm6tPv6uL
kFDd1qDn5atr6BlRZzRyakzoOtf5yDD6rakUd+NvPtnFSslTJqA1qsNt0Q0VLC4p
fULc3LoQRJMN8uTVlHMbZ6Uyj+XjrvUETe9QELdSerPwOz9HDNEQzz2sKHd4ohzB
taVxZSg3+gncuRn26LgFsBkc2QzK/G2np1wIlptfYPNNlNS1YFrLk5NreaFavrl9
JawzQFAyoBpFhjZAXsAQP2HE1h7EgvdEMjkyLJWdvApChH1rcbCk1HnA3KcSckgJ
`pragma protect end_protected
