// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:48 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
euHQ5xqyp9xs4n9eoIymEYPGFvvDCL+Ad4tWxZVEJdOxXGHcqhv9Re9v1f4wtSrI
PkJrG25F1gLtuWRTTUK3728ncivmcCkXuRyloFA17Eqf5m9CsR1mKOXWwZB9NbuA
mssFl1xZgRTxyRIwIXkxZexVfOIS6WclzE85LwDkpZ0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11024)
9B2hOaEc6895YBISxDPyMW1sUfKl7j+GGppLWsaShotrEtU08CVtSKKNNxmGER08
U5Rm2bKYqz7L73XMW8rW1HwN8YBLw3bc1p6/qxinN8Y2QGbIRtTBEpGMAsPvy31+
1INvNcQlvUvD7Zd6nJqAfZHud5zRqQ1NXTFLfzzDmDoG+V3K32TX0QC7daN0D10e
5ijLB1FR1K5/BO0ZH1/83JJAPfkGEBXzhrbS2BAw6cNysgO1uckXsvRHr/ft8g+E
nWc1SBZl6OAix2Z+IExenBItYnNmiz+fjWruQJ1yFByXDF62u5sJK2JfAke1X6kl
U/bRGKJkgnX+dKb/M66IymSKmFG6gMQpZ0ZFCVpal4UuncjYGtQKBo9wzILcvVGZ
5ICDBV/nJm8Uf+4GnnLsupJl5Ysetf9FR+Y2t6/PcxNe5U+4kMyXyDgvHY+E2KaG
vn507+8xrW8pWnBq3I70Xp2kMrpjMR6hWSLAOR4iu9r4UCjVnqfj2MJVTjcGVa0E
669y7F4TJ90kjRWQp8qaV1rl3Fk8CWNg3l3hMRqncgfYeMcJV2+GUZjT2Ezz/OOM
nP+qxKnnWvZv4MRL6A+/XRWDKnrus9MV/ntVIGjaKzQQxC9Uj6rULjnq+7eOSCwC
/OHc5jlfs4IpnMwxvz4x5ei7vju196u9EnvdepZAm0dSCpx8m72nr8ezkxipA0im
H/IJxEdaVX2pJaVlt+7x97ijiJ88Z65jNXCkW+ezKBUlHIb2jaGdL7ahqHKRJGrg
M6q4W0H9tRZCTADNu6XvyOf6uHg8FYmYxUewcBzCgjZ2djzLBpIGCQH4Sjme0/hX
WPJwFCUWz701uJWDFRRGqnbKIp8goxXefcaLUb7nlO4qbEpuWAyDsLbiKy+OFsWw
Hd7HUDMvHqlggVkG346tD6H0bu+rB5Aiw6NfdUwQaGosMK7Q+iDCOuQksmb0EA7K
pwOmUbJED8/BYO4n9b36iMA3nSUwEWgI9LNJwK5I8BqHBF4PXlUKNYlWgHuE6yeh
LKsy8mhiXsrbc7JESn+8rprl0ZpRLCpfSFZKU+wisJlY1o527TnnuLr41/yidXBP
z0TRi74rplLyQSrLV153jGm0ejeYvjEKHQst30ECp7gUBDItls2zOqhXryDf/CUN
oD02+CIZOwo/xis877PYYcEcBgopgq/5MXW5r4ybsD1Sa/zkMpDZwHPSevZv09mq
ICsXQCknXIlvhXzXD6CR9zryS+6CujYZTA7HNS+1B/h7cGeV92yfX9jwVE9Lneup
a7cpiTF9eUGzPnrYLZ+fp/Abtai9DLnrrdPLWYajb6/zHQ5uztjpAKZ35IKu1Eik
FCfzkqeQ3l5kUBRKreKsXdMtsDBbSLI6mdhCWgE3R/knJXM0Q4Syc+OPrM8HaRuR
Xc0thKCOB5J81wjKn2RJLWZmdW+VoGagt/mwXcPnyxF0dtmJiSPzxZi7VLVf0RID
QSL3CsfvONteSFaEdeuL6V05C7gGQMYiJRufFWLgRjjmyIYCBZAaDqM/Cvgn1S4e
HnXJ/ZxVF5cjUtJ0LpLKnWYgZ2fo9XIlc5C269Ge0ZeW5mUvgbSlUE0p7I46eneI
X7ePI1mT3TCfSnyAJRWBHRDyU8NCdwAevm7+EOzbkoHQ24Iv0lmoy3qMgn4AkxNn
qb4cKO/BzJ5fAt3EjNeC8QIkdcottdD9m5img/JjCQPRK9QYz999b9kevTVejVJE
V45JVFfvVXHwEPTyJ97BmNZFt6DFlg1WaaLIdIfoIx5+xQdHQZL/h3Jeifa1MBZp
EtBzi4q+wgWPC7Sq88Y4GeEzOoIoAtwMB6mKBJZr1HZCyMHmnGFQI5kdBjlVLR8z
1ThZrJkzYfHwiGg8XImRi38yBWIXbw57Bhm1BqV0GwA8sqKlFDlh9rAsk7T6Biba
U6I8MFQDGnlK61EtQjOJGD/bIbd0NblMBYEsmoEG8EqaP4locLhXn8l6dZm5UDDq
r7mEKKAq2o2YyuSVuw3kVsoDZjMQFXCmYmBwMclYf+SqZ6ek/7aXJHiuhPhEf6Fz
00QNTmlSGhRECLntfO99emk84ca5TYpC998t43wxTYO9ERp/SwLILdhMusDabigK
qk/7NMpF1AVyC7eKOQM0uEEbW/w2T+qT2w1ejGgDJah2D6EUwZSHU2w1Y3Nj08uN
QYSTIT6Ag/vK+pDTNYOex2ikpAzpCTeB0J75XVenIJhSFG89QEvWZ01HsIqyXCdd
CACLsuhOBiTq+8TweJdjoONek7TpxRdvU0KndATjs+BFtwGserHcgTyFVIJR+b5/
yko0/ty9fwCC6ePkgBIgugUrcH+qsiyh1ldBpNDDwJ71NST+qRta6KHG/zBs4hwe
DHAYa7cuz5e4oe3m+Y+BTFlv4Z3p1kNAq2k3KOwG49B+xRBL5XVzqnwxLbFL4M/b
BGtedrkeeinjX0CeQaCvbDWp13Ph9gcByZs3nbpIC6cKFN6cF+RtvRzlQJ/NCMuh
AnhqC75E/Zd5EPVDNWPM4XSTkiBHoHOaLAlHHF2Et3IsGbMRggNmXLJQ3Gl70epy
lbMwWpoibWyr0pZA4A+vfX38NqHx6bauEBEHueq7RPP4Ecpwxk90YRmfv0cdzRR0
CtanVDzORIkAwIwTSOTzxP+l+B6VseVDTVLthinOKRzxnJjfYun+5nPLtOywiXvq
jysoSgx7AiI8Gu0SfCfUVRchnDZl0jmpnEKTc7pRpCQpNQC6PkMh6CCXxMHle+aC
AhWDiDMCakU93OaGX7TDm6FK7+XOsy8wERzt8M2lYukDgUBbBnAphHDzr1d26oVn
2EFKVcAo8PrFlD0q7ADPsgwoBzj65U39HLZngr9bYBgcrcBrARkTKPjoo3J4brx8
KR/QkYKZitBUTjP1sSdgxqCfcGeZrIgGblsLokAnjU66qUsJaSM63vgh8VRgB98D
PyNfAyl0lXUYFjVTj7AMTlgOS5lF7ilfMh0A3gPZosKWR0OPpCAp2JLl/XkRGVQn
rOvyhQgjsPmmP06Y3EBsudO+5LLjIhgYXaSapiSVx69IN1U+0m7chaoznLUDf3iP
QKKxTV8DO/lje2x48qd+ejXGS5yGWqBXfAmm99GwalDqg2LIcbtr8MOgHMiMyF5r
TAPVEWy+ke+QFWVOQOTjHR5xzsvtPTE7j4YPGLYoxXAIl1QG/06Ah7f1Y58yLgqW
1gbjDHzmqCxL0JZ1EqfEFIulWWwrBXpy8WoRJPh/yvH1OlO6SBXicSeBhvgLeWkD
qxyq6qQTR84O4ts+Qp+81OnxOnn/UG7NOt7QUglkI1hHnkdL7PKxmMM7PMbP/Gnu
/d77F7zxy0cG0K8/3LS3iat/EsF96qfmoTKw3Dg4YW5SoEJYkh54zj1dQ3BD/eAU
yUIhgum9L/vTlU0vWgl9KeQ5i1qQaaDYArelYk4xrpEzDsZHc+ngC7hnjR/4OLsb
ghCqBTxYrfMnGRHRlVY7uvO5K6sTCbLjLxauNjLNHTOGKFV8eKhSLw2WTSim6lFK
n9lWgltPHY8d6wkp4O0qgF/XdrxWkh25gwh7Dedoq03/XHVmHnqnDL8SyMyAS8wB
/+z0zM736IdPpX9TA/XEZEN6ckIAAmKRnZWoH03ezbOVwjsS+5QoZ06HD0FsQyFQ
NNnuhm9gaJaKBH1Ybs0nVqFL8YGv1YKnuzQqviwIDjlqird6J0gjRxeTWfTJ6z2s
mkinzG/o0zlpJEESIGdg3zSlykx9pFe0i6HRXCKjplv3KN8JTXmm+bjk0w4WomU6
8Ntu0A7jQRaz0FEqzj8RSdLy6NBGHx0vTWaCvaXYDuhvbrlELxrRJxghMJojptF2
Id+WQT/T/sfPusJDlWVx7g+HSU+ThAn3fJTknYQhLLzUlmWmQR7pzSTGZj+Mjla+
NYVjcj1Ga/4B6nb+sLxGxET4NJEMbzmv+vP5y5Vt7C3Cm92lu4uC9UNM6tZg6m7b
uFITh1WPhR35PmKq6cVkDdgW9JewV0K2fZqiRbR+hLfXAVURnQRtKahaOIr+HO95
QWj+XDV9UeeVNEyGDFwBrlArqV23agFvSH6cOrcB4urjmLLy8RH1cvimHf752eEh
35CSyds4WILQtaxsyI9i8jpFvE70dYCO/MDRXdDA8Vpiol9QBlNJUUIpDzztucpS
fzdDLXfnXInntHmjS9smcmCmMdZh4bzKTwyJ2ihEj4T/DaN9dzoNns2ORtnh/f+a
yhyjFAhilBneY7Da04C7hDrS+NdXYo/ylHFbfmVxIGmG20AUd3G6Oj7ekK2SirXl
0e3q6HoM8zbvIeVBDF8vbQc0ARp6nOwgy3dUN+DJPZqLgn+wPLzEH0HwQjvKP7vD
uV0uAANtD8qpPNUk9MWOBEToiYAKiOHvk/gvfwhc3tS1ofIEKQ3UWlQiNzT8pynf
P2RwHV/voS5youBrkFXuQ1B5q/Y4qbxvGiObs/4yQAML/A6MGmjg7FQAuaTVOYJ5
00LkDmSESEcs3NNPC/ewXTXIMfiMgFGR1B40JVTOFSG/Wv8k8lvcPJpDce0ZifaS
jWff858Vm4pJfc8PE8WDbLYvuF89qADl2td5AuY0mbcpYGb1SmqeX6jugLxaRQKZ
+wImf4rk2JGSR2qwtCQzhqHkEX8Ct7AQXbL4M6kGCyhP1KYvmO/DY82Za/a9bRm7
tnH93NmnWVgF/B6/qLzX6SgG77zrSnTYcPMcoHrqkNVqxp6400Fl+xg71E0Vq+oT
SLqWzvOLCmiOe83v4DIEny2oWQK/4m7A9iJZGHKUq5p8c28xgxJT364H8kFCSpKn
ltVgQdXSGBeX5z9uW+DLOlXwBSo7p06DUlQROfWpaMcaBARQcpGeAKEEt2ZAomxG
LUIARkZXpJgHtb8YQ5prWTD34Cip1egti0NiJ+eS8+t5ALH3K8keJvS+I6DYB5ic
VlEVSrQu+/obFzLfsicJUSWhXoeH4rvQIVVE56uLFRWOfBzkPqXlLw7OVXn0YowW
7GIBQPqQOQKEkFiVtq5qBvAcQ1BGJqsLoNMZBS7n0D8EMyz8lVNbsfPHA+0zE7MW
6Q/IY2fZvfRipduuLIL503a3fzhrMusiIitsQszWeduiMs2+v6fZ8sHxJnDektwI
9UiC+XNqLH5qhdX7UZ45b3VfdQ6Dh1TaAkUxHwm3E3x8fb55yzu+3rn3wQv4YPl1
cvd1X+xtSDGqi3N1LaiT0kraFcM5wYkFmv3igHW+s3jtsccXR2mVRyxf6kBtqdf5
y6wIi4RbMR4OHU6xxNrXBsBAWSRgRgZ328MevrnSdBkzXKpTiOq6qqOljkDtOVp4
KGzzqJOyBJmcH2xXsrUywBoCZ74BQaGs4nHScK1I5IFsU+Djk/4dfYcKR4Jp4UIT
dvBWQUXakxW8vmvq3FAj2uhCD7USzxNOdPKH+s6W0Ujlxfdau2lDjNJ4ViaoSpGR
p1NzF22zC868Jhi+x3CnJ9d8uBTN4yc0klHmLWUxAYIaVBYS5ABUEXr/06jHNHwe
QLtplP4Nry156oqo4hWRo+bTgtJH/dwgCZOeol52f2Rep1/zWKSJn9HptYTVHYno
duY1UAO52pe+sL199rAzPKFwpcBMy84kTdCS2zsWFa6ZDpINlJ4l18wLTL9+l9ej
AmOr8eQFTi9V4kdFYBLS78C+fZU2u+ivBkFe3NZgbZ2bv1cx8xIrU5MZ2XfKyYti
pGhkfRPST8IZnyraKTgGkqjFUhZF8XDE5WFr9sq8IcH4jV3JGrmAo9GGJggplBOz
RaFBOgyl7m9MPPaycqjm7hxd1Dst6mYrLl4XzSXXDW3zhlv92qooVxXrB5iUAl5h
YZCVtQEnGPPb0TVuZdpbjL6AAgT26/Vpil7xslcQxTUUovr1CGjKuCDEPb24W+YO
lB8edgeFm4tpoqsJXflYBnZk5o8ZtS5FeeE8aZOlwAzDgWWmKI53ryMzKlsHsLWN
KuaBm2DfXzsVzdybwQ89DUDmlEn+mXBBAhRpc2IzURzHI64YxpdGCXS4HO8GdZRD
C1F0/SoQAvrW5d0dBS/awtC5Od5hXa6tq4NBS0getWtCtxMw2DIkZgZoPlYql/2t
hjiykC1EMBabXTaN0FYcOzxX7dZ7EeTebtaAyJIfMYi1jVmTmz67UVqqWCpB4GG9
SWcCJv18ABFU5Wi2HwTPHGrOskWU/g2TFe2tJvQLHbSpDZgckINoXuy1cWBDZzFj
+hbV3yjqwNwxxE5r6R8r+7VYlqa4rHj8L9GEBR0b5rVtab1pk19ASTAVQwGnhnob
TJ+7m7RsfhfyOCEE62qUVi25z/qfkuWY6YMrKNkDSvOn9U8yNMElMsLK9wVrIlJN
XQdmkjaNaHEPG2GnyiLC+UNoxj3Kf58/vdGDOhTrUtwj0DGpn8n4QxfohibG4nbZ
yr4ojk/zEAVHLL9+0+ICEKQcYEoqzod4QnhyOz7xJ/0wThfC52A5qT/qQ/hyQh7J
gIhdaidXyamz8JN8gSXQTYAgxh7ZquXGw6M8QZqFnBl/7295JMV7vKscWOTu2YEL
amXyNfvBoQ2zJiimIfwgvH1/sG9HnxxWykhui50Y/FkW0gaJX5ZM7rtWopa3jvQt
N2vQIds+Tb+4c+FQqPBC93ddprOuba9U/S70VBy/eRq+8oMtflm6mIQ97rRVFZ1b
6AZJ36QGHn9Mr972yObFsOZu+MLWzEJNdtsLLaQ+UleZ97YRtgdLkcqUvQ89IE42
HxAYwOpH+0TwXorSpSTDfxYm2WHayFrsjPUd9rvQ26mrU+W2Ou+BQwrHjfh8RrgE
ML8r30npy3dHOwxZGo7R+22WLaN1YokCe39nU3Axd9szKPegaiZFHitAnZHTTVfv
VE7yY4lTnxXY3tZk3Xmfn3agGh7u8SNohlF+nJzBJPslHV41zC03cPjsIRBiqusE
EsNqWEAI8pTCL0626blLxPTl0ejGf0lBKxQyiJSWNFosAcdH4tapjZ3RCTHl4cuu
EXN+muYdIC990lZ9doWHObLek/J0XMuQTH/If94PeehFLUPp3AwOMrqqEQfesQSm
fPTCd/zMcvV02eWxKj7BlVjJbPnIysTWMCwtD1yCOMS6GCwycP5q6qtyvc5luLdL
byBxDVhheLQ7orqi3dQC13kMp8Qa7X9UPo9ySWzUitBwdMJpNRLVLViGz2SfqNr4
HT3RnW7LSAqGh61V0dFYZ4sfBQxABqwBgeW6R2afjf18BiusisgbqkxVMCll6apE
iMvpoGGY9v6lWFksKRG12d6/12fHiTvS4wi9Hwm6ay4dgpK0wuLc0kg2bFqe1+e6
BVFMGP5dyIcPR0/WkKXsFG0IOg1WKdUQGvKE1f9qqJo01xRV4ZZlKG9Opt+k9vTt
YtVAhWfTEiskGiZ5mLx1dSnPySramSswAw/ktWp419NwU5XsWQXas6G9Pio2qgT5
tNnM3DSLnrdBArRTSPw6oFDd4kXqPQVLETvdllgHtsPk0LkpgqixIbHak4jk/ngn
EbogUENnUflG8t/SbqsyMaNZKkFjrrR2cX6U3j9X8+BFHT6AkbtAXfCVkqd1KxmJ
Oj7JHgdusMvvHLTaHcqDqpnFMHXNoGYKkXJpuEg1ZEi/JGDzXTKFpgQlEBkWp7+f
KdT2LWGJ1UQEwZs0VaSdlrVLx5/QRlMGaxydRvbc1rIu3rvH5La5Uu+PzDT2jJ+l
AoExSqadAYgg2ULiZqZDF22U3D0aGGPljaAQvzrCLHRS4RUCiLx+RjcBLRTvDabb
kKgVF/Jzf7QBG8CLTusx+MTameo16o7jeMx1HdXVtKQ79lpPBDrX4peA1tfWRF1Q
QxFjVxDQsyB+luYrVuLgOenU1QB3PQZR2cREX+ilgMunfpgt+9Xv9sktUFoxcVNX
MMRLz66blt2zq4yXQiA3vLgzNjz9ebODE5aqjSQxeN5DZNH6uOovlJFzBJkNqJls
p+KoceWBu6mGG0LRozI95oR6hsxDLgudZLjMuAQ8wXbdN60EmY1sDuxfTW6DRUQ0
xnmyNpm60uARqXANSPv6PY0nDFhqm2utvUXrz0XafK6j0o5qubvk+RX+Bgek36gc
tTDeq9H9sS6odCTX0Q3Xvep+21t4GL2oEPubY8p0ebYgHNuuQUXeDqxP1r3BoyKj
lUUAB0mlzsIow9Fbv73DG2QPOTYUKHxN3qQFMAXQzREQKsaOmlqsqOXFpNc9XxVl
TmDWk2NaHz+fTWL9eNheNdXlHK0rbP9mA+q4kN0eBn403NlpWlipnSASp13hlLmr
9DaqShru9QwQTq0FL2Jjm70+Ue+7g57+YcVPy6CPh/yTqgh2UwdWnHcbNt93c046
yEGJ6m4DdMNaUA86JscoVCpyS1cN9DA1txvA/HUkbTgOPOhMGwN0TDVor9Rmh4CH
49YouQh16GDn1KQrWG7/jGouQB9wQrj6Bqq9mZyWCquM/Wgywi+vxQQXj/iEss1X
u/saZ9+CqUyODKRbmivwXBA3lCydVgpnSNFpe+ZpJC+qH8fVlwJoAdmGQvS7eSEs
EcFYxOaL8ZoorDKd6CN6buJYHNgJ0yw/vHETs85W46hI+qCo5BE+ciYLjQst2yTJ
OopQBoQogPqfzN+V4tPQBKlXFB7M91pHGqMzICOqshG7rqBMoWc3kKfeREQlRm1+
aXjavlYDDLv1evyhKSanRSxVvdbI8oVXktzbZwyRin7Ci7SShfodAFJk5RfZI/dG
cw1Zl7XUinMzTmR6qzAWNAB0ODLmftCzyi2ypOf845SJFGl2vgzsBS/A4A6B6Co+
xLpmli2/ZYwsxJfSSb0So8UYLeAs79v9KQ7LqRkdIM/R18Bce4dZrliVSGKLZxDT
MurJd6x81KJl1T/XwA7RGd64cJEUv5OqK7Buoxg9KH6MoGkSq1U3JpW/lMIFxESY
p5sjnl0cdnqo/Z1TU7DNqQLS5jUBJSd1nhk3IDyRoL152KLifXunJT2QyCMzP5w+
ZixrtCTNiFHIwTqkqNl1IceQ7ZqoDtIUu5QxUtGVq6A2dJJjq8jyIqpl7PzDBQSL
+oakPRQPdyRvyrwsyd+EU5D59P+emgK9pW+gXxHyurQVe5ze3qcw7N/P/T1AwQtM
xbEhAemECLrxuQnbmRUpT+Rmn3DSf4Cz/dnWsqQXQ3U+jrY0PS6NBch4HFXwA8HU
wRJw9uzKWUDKt8uzx3GpBKLUawjuAzy/DSnEuiTbRYeuvWYddifKxCLSSS59nxm/
4k8BC18iPRPh022e84iyMJM4ZAVWPzQ65rMu4kmpMjd4RIJ2Qf3sHFD1ujMvPwht
oiFcB+yPwqlfjGY7h5dTWGUEAsQ4B990E4TAK0NcIbpG4vjS/9+2Ln4BPnP4flmf
mopvzkBL+4tqSutFxT8gTuyFQ2J7FHwyFmSugW8yP/Koeh6wcFLyyYivBIkZSfnL
ZjVoyec2SgoaldBYMbu8Zbgt/ldGRQsZQd2G8MazsIoN3j3CYFYjyut9af0W2gvN
ZXKs4fMUF7eIQWuTZU94CXRQjRJ6ADHoIpADJ98t+3MQCJrupd8SBG3jn1DHqiaR
Qi0EIS69Esx/Boci60galmEPA5ZWR99B0OFAHwLu32OCVISmkA/MQQsJrimog/gK
8PA9J8j3TESlkZJCrOkF7r3qrDOvFtBQQJ5y6cnM4b7IG4Q+aPeXE33/G0UuDL4v
B+1tBIT//mPA8zh3ZbHQYptL6Mlj/zjslnmAV2QuIYp86Z1MgKwZLBJtL5Agrcj7
hLhTOOm5VwAHKLC6ctGs2SvEJtFc1+VJ4EMTx5ByRC2uE4An3zSM41kvS61XuBwx
7jLlj1JtbzaRA/75WMP2nCYarXpqc7L97fEtKS1/lYu0tIzy/R4UDJbHSrx39b03
x0cFd+sceHikLsJ5M1qPTxYJm/btbkAl+A4WnW5MefBeVkIHIP3ADbZnTXTpZxJ6
wt9uEa5Gh5UDM50X4n84WJsvBUiT2PPtiEws5xrGhaVQMu0IBZtt6gQWn9d6MQMq
9zW+hzEbo1sJrlP4EL/m0CB0ZSgWyNxd0EAZrUabq2yddpWiuNjAWfhSAZtK2EOY
1SF2I4RVWA2EonpqAP132WtkmHbR+nOB3i5i8OG6D1hu3OlN1o0Xn5f4Nre2GC8T
CPQ7PiNzTEHwYpYNctsADTc2ywXZGkcmyNIYw3/hhKV5vLs5jhEOsQgrOvRtMlhB
MaWu0EiZL/KYZOjLDqMTKb/Hve0GUbaVT7iTlKSxI7knR6dGfVn1XsJN7Fscrmtr
QdIVbSbkR/vEhnEGnyWiKdY983pDgV3UGJ9yVjrheR9DfZq/6j7xIZIyNXl4ibQc
wAQkD9/aIkbn/sMBflMhIW9NICS8iDPo0QFGXnayxcdsoC3VLjuOhZ9CGQib+8Nf
NSICbUeg1mg5SbTS4pkbEiELnrHcj6T89INYrhW1MazQ4AQ00u2CHVFg5rAySWpt
yuhTxBUoKDawDOAuRAy1EPsl672o9AHBrwcJFZPx57ZM4j974sgn3B7k85khprQ5
mjf8mg8knfUk36GaMR53MKzaEGnCDZp3pmYf+kKyoFdUwCzABZyXJPlX+dj7KJ4f
/0WrLt5Gsak8e0YkDh8Fg9Z6uTodRHQgwd6c+eYiYWMHZqTJvmNhipiLPheaTNdo
qs4kzc0zXjv183hQjWbVPAIRRGUySzjKL7l/8KRb7FnXqBVj0J4Gvlh7TVbuJ5dI
9ooGc7ZaqFLBB1ynBeHO2tPnUFw17f8vwadvXsMWoaKVEl9L2kTYSbEk+4EYV+x3
x8iQmrj8XjdyOfR9FueP0JrQXJjtOee3gUwRK7+iFetnfi19crck8aRxXoZ61nPF
XiuByKWY/mWMjn6k1jpyjRy8th7/RK46t5tSw8xXjshgUUhrMq2P/T8mPbnPo4jh
K4YKqEIe2NcQfnxA9hPDVTXv4qUgZ+qMDyrfAhCJZs9L99lpNTLcGza/xbMXw8F5
sm/I2ZcgiXWI6D4Pn6sOCavQqpXjze0iiyjNYIV91iTWBRfqctjAeh1QfLmndSPM
630uwU7jkriMva91k/s3U9bsM4jImtzd6JIrugvgxiun07a+1ECgBOcpRzqZvq+m
hUheC8c/4H5UcTFWCOiBK6KEbgNN2zsClM6UF8jG6BuEip38XpGmQ1DfUQHHCmvg
xciRtJeCfskCS4K/9Wwu5tt9zutlsWxXEpnPRTEh3U4obx4OTTquSuYgPAI6QbHL
5IKXOZAfDR2EP1jnxOJTMDdaSIjdyAUlAZnml5dnDGDKOizAoQtZo7SyogMBhGYr
l6QF0b9pfjwEh3q5Juv9ufc2hI/qCP9pePkhur6RPKBnuqfZ2iq/EF13BMWMf6Qh
nP7KvwCGvZk/sNJejJhYmpQQSiNSoLFtZ9mqKrMl9RorADvlYLNHJw6JWotWkx86
1gBVDoo33oSzShO90gIA66esKIZnHBlpAn5oTVJtQu7zfdWHWA4/rddek3y0RrGx
4OFKargftFXmRTmusYUOVEgazshMwA2eUmJAtTq22rZT9Jn6sTM7QMNjzFzZit3I
uBnuRQsw2Do0CxBwUi88CJqFqHzH+9tEh9Re/tfT1YqF7AT0LKGKPP09o12IRrTV
EnuoXv8mUZlq7E31J72JUG9sGjip31338rj6XJLYRaq/kvLwE6lcO2Z7ol61uXCO
pu9IsD6iZWdOAUXXeHWuy34qZkbU7gUJH5vAzEk8zNmiwDMs7zSiE6xEOH5r+umS
iSUdc3rb6QXnY57Z/Rz+hlFgJgtSzOLU/upp7I7Vo2rO0fncJZzRDtt0pwyLQ+8J
koju7pQZNM9pSXVi2U+Wpwc2jfCX1URznPBqUc/FKgaE/0RayrUI3JDxoNy8vYYX
ZaruG8xh6lnICjwbw2MXfkceXTXuSbokorOhuvB0fvCiFjea3Pqntrsp1FYde/4R
9hI6yjKjBRqsi/7FfyJEY4VRMEkUymhaUV4AC/U/hZRM2JXiDbxADmxgwblZLygP
4o2urPtRV/y/UUdlpoUVgEzfiEmkNGfwGUx8quu61vSrZmT0x3dgrBCd/EBBSCnr
bI+emMKZW1CANMmf0SycY2o2YuJqQmsWjUY9nTpDuCsqGRXHiqXo+/sMqdi2krdm
3XdiLOMKHn0iPu7Got3Nn5ktB2Chly5EhAcCjm1VYyfYsZAGjYV14/B1c7nrL7nJ
TRIzoz8JbNH40lX4bc79pdiYez1V+4Yi1/8yLPikR93zUWcBdDmep7nfXaEt3D55
k1vSZdLi3AOMND0AQXPUPBzZcX3wj//j4ocCnWObSCq0FyLG7LL/8i9Xo+veXhFh
WzlP0Ahz2D5ZgB3LU0mY0mA9hIdeRiQgfNkBRkKCXMLEj1LEMB91433vmLz0/N4w
h5nEXHdA2y7jvrjM+6GPh1AO7jYh7hqF6+b3NwbX4W5MZEmcZPfI4ElfE6YzrrfC
NqnpSC7OfOM7Bp9x9txXNx/H7sh0ChpnH5vABqV6MzCc0vTfHNJJAev3olGG0lqD
gJxdLbkQDCG6n730YiZKS0E+UUH95VGjiwp4k4IEx5XmvxCuJXO8AxZGk12jlIJI
xtH1R3/dbq886MUo8j3EAinWw0Frog5WUXXW6h58wAS+g+M0jaVILT+lwGN24Ydz
3VK58tl5x+TdQ9xumsVs5FmKC1OWh5lv4FdwY+mMEvWnLHKZU5ucaKWjeYMj/5wV
4fwvufHMXYu57d3yIkFWHixnCX8RjIT7kps9oTyVDRPFOWdXQczzf8E1Q2Hz92lb
hll4m+eM9WBHmhYwcvGAAfeK7OB4TYUtnLlv/p0oqQDXhMAz6oFwXRToaUb1LHMC
5/JuS7/hn70COIvgNgiuWtQGoFVXb7vVOXaN2DRuzrEKO5Pbd/QiR8H62xPTmAfC
E0kpFOG9pWXvD7CaNv40vQBFAAgvfcNg1eP1pGBkjKyEZ+zMoZ/OiSUuww2xr00U
0jzHE3lgqyVHeTtX8gRnSn8l8hBmolCl5lKrCCwWaK4VYUoxBltNq9XaNsGszuB9
OEPehTklRCRkYkoJlye53nMSBBuAwBGcVxJRVu1C6gUi+zsXPhQnyvwV2Z7EynDo
l12OEfdvgbsVhXELLfLPrOePTFvFGkCBiKN1JhNAFGcrxRjsZn6uQWXCjzY1tRmG
Gf+cZ0PEz5Pnj3Gsm15Nzc4JIWJBbAnZvmaqYVR2leSxZbDbPZOYZKlIh/jiofEU
yQj76Xtt8Sq5+al5Q+R/19PLE0960gYs7+NbhG3bR8KNDJ5iI0osmQR4LObnjcUu
LWGg3ZJKerkcOVwkx9ZKmf+bDAK4BikpOELLK5sc9oqtpLMrEV5BriC9f4QR+oRw
yGene8y+Pih4CoYkZSKr+qF5ugMMfgAOkoYJjicmf8/7HpNgvgxSgabpMFl8kajx
bvVz0jn0Sn1hZ1TV+pl5PExG4v2Tv534jhvZxN4ALLbVJL2s4cQW/76cnv29M972
MsBCK6BhPnBV/QX0DWZso4NzA1OIB1LGgYlsDeWBE3nLWApL1IWV1oC8xLRRb3ea
rnepms0E3clXm3yRvGNWhM5qzf+ghZkyzZz5aT7n4H85nHcU4281rAE4JxVymhcN
nZQ2pvNNqep1iIGfWu0nsTNFO+xH7GkfN+OVqDKIA881J6q2GzyOZ7pwebk5RvSk
lIOdMb4jh4cCxV0C5s10DyfqmTjPwiNJkMtUMAE0VWm51xA/xcPvxa9qdG764dzA
24vXliVGhVD9csOakfis/GXKPDbj10nBWIvyPQkhf3BjzTcmNgn2QOZ11eZ9EOJk
asJwep3m4vsnlrRyNFRPkBVI761ttQ+jOqmX+m7wnGUKprSLYhytCCU+tw7rduFy
wfHGZ8anfHuzjKRoK4zebxYU8lsphkzN/kdMFPo4xGWc9mPZMe5ma+mvhyh0d+wT
tXE/FDUCYH1G6Dhlj+zNaMfgNOWBa61VqsClybJH2f5LqD+6tDZr4Blx/K3VQn2S
Rdt1tqbkaYc8RS0vD3pNP2nZoIn5pd17cQ0E+RnLyfWM2UBl/Qs20AFhzgZMWEkG
D+N4ga3QjrIn/A3tpRABCSEZ5gQzFFHucwybU/rJG88oujiH9KNKsuzfSxFPRR4X
i5ogVTqgwpFQQl38EG1E6GhAH7CSf6qkwEOBnP7SNlkkH3Dnh9xQgylD2mN3dBD0
9oB6vOCK6CNdaPtmloaW8hY8T7iVPCHAUzTEUAnYYpk5j5LAV74oixOW5wHRE5bc
A65WmDlvKn8iI8eoDFmyS4WoP9bSUvBCmvGmQDUD+q0iiTBEqPMvrZ6VRoxWvXBz
2t6uDMsPSc9ihzp76kd25S07dvMeIRLAyAkanb8L9r1k6w5hKuzVIZJO/zemz4Ag
LmD8Gw5VY8e39WCtMZ2GttbdSdte+0wuOCpV7QBqvdfxPvEg/Dt11vFAJOpYIx+l
oKKOsjB7Xk+zpH04K80+9NPyB3k62MdJZgdxKdnxmiXkQsUeHHa/xXfcSPdHG+4J
EJJ2ToQcoV798iHPuRnICIyBFSH4WpdnUfvWVnBNRapwU9fCtCSKMWczTPfLR3yH
SsJCXYFqoi/7IB/oNGhIJOMGRAVc5l1uuPBZehpJcCJLOQ7yZS7d+YhrvxoDW1n8
DFPKhA/OrrKSvebMfUuCiJv2q3uz2g5dCHN7LBIU2F6/JyEpY0KVmTNlgfaudnSN
Y3wFntJLTCNaDRzxnJUUVrBUC7nC2ax71tFMYrkd5Bg=
`pragma protect end_protected
