// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
BpVn+lWheepqy7zqlqGO7tQn5VkKZo5Mmy8HTuYE86l3rcfshUWU/3CUDzPBTx+lAGpX5MoqapnC
iCQRHvnN2jcdY+/LfgqsZ2RiEVNpI0Rq9icKdAObBFTd3Zyud2GeeF1zrOykZCXTm+oM8uWw/B7f
AwBD2dGW0VT14o74vpIj+kb9vmfkKkAzH6kNrUi+Zi8De6opUf5phAlnQ4lgBKOwf9z/78SqtgZ9
I8DXelx5mOahyGH+lVG8l+U88Z98qMqbcLVXjZriXtKvuzEUiJrk5dbXTwYFjzPRYM9GgwRe0qXB
g2zSzFhLaApojW/cz2un0s7Yi045k8qXPxHwAg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
BMm3GwCPKWT2azQHaZVB83KpqnpdqCBaptGFNECRjyIxQOeGVZGFkN2kugxf5V4LZ7m42PtplFI+
4jh/BMTUJFllBXoghJBDnFyYkn4HXyfwdTnbexgWX3N/z5TrDAylaRymqW29lDIJir0FDp8h82jm
LoZXh7gZoNMxP6R5E5dpHg7gm/X8Mvu2DBHeYrNiWWgEhD53Ow5FQnorC7K91kPwyOqE3rGpPWW+
CoeM9BwbJyAHUl/cwftUeB0ToOODxot3rfwYH7v7dNzDyWDbfmn0fgZq7Qtp4KE83G9q2/t6Gr1h
5g11ccS4ynPGe7/PcFIeSa36a3fXHOFX9r1dwEJOWX7LUfDVORTCDW7yqyA8AEe+lmI1X9VS2PlK
czhkc1ZVj242phwg4sW7C41J4n81s/jAppeALCTT4o7fVYUY6vT0+cIQMP03qNKASI7fWKN1FDF2
dDuyjMG/srM2+SZP7/MA/KW3pMauPHZv5vdQ05PKNII4c7OCRGrXdHC27HWdX3Wkh4fysucTVCVY
sso4wgo1+4s17JhXj2pkvkI4lPnTUGCtAauPcOdT9l3ZuDccFMOYhY9K62fiyZs+9vM4/nC5Nv4o
5OdKJ9KjNzVi3zeBzThbUVl6lAWHjZqYEtHga5huK3hRYIwNxvP22/577Bxt1t78RkASbmAE6wsE
cLIxQdtX/biCt3+OMDIMugH+29D09Zi2/0YzdAMZtFZMesvydXnWV0fMxg6bkh0QlXG+LmmgG95a
OGxaOtDx3DkaqFF3jgsyRq05hzmJQ2ubIam6OK/fBIkTsebeInLHZBYNCWlOgJ1tcU1N3pb8xTB3
ielY60AbnRGHv8WHnrax5NhpamOOj3wy9REKFodhu65PySvm1B2+hbMiWx1Qk3cQiZjfodxYOf89
CfXmDvwB6kx8Dt7u2Onyn18kiq2pOdJS3Ie0k+N3a1d3TSAhu821hRuFkMNriBfIRqP2qxHUC/lY
Tj5/aUdZvHc+6D+epFtLG/qBxSG5hULoioN3FW9eRbNoOvvpEOkVeCaRr8tInq4RrGvgeW6AL8KZ
s6M3/34GpWS0q3daH/qYdH5cYVMzwkfsw6ENmjjhUQD+9Y0fhabvGs0hkuDo3rR6gaGBJ2V2tkqn
wZ/K4Ap5gzv9KbAU9v8+EFBOxIVS3qXAx6x0kCpZ9MVL/GTElX/9rDicT5B9VeDRFzkDAPHeLitD
HKZzs00s4jdQs9AWkV96LMGXyuz1StaYfi0YLYPlk42AFgskE7fJDlGptE8KnnS6ODLob9eTnUHP
Q7jyf0ZJZJIphuCKki0dAzewGyQo2XjAJQoAhGObKptxT01FE4tqHDb3PsjDqcCgREQVFyX53y+3
OYnElJa4GvMNtvpmhff1WaVSEJFbXOnjYpXig8FpBs3r1Vpsf46zNfBK9DF7556nSN1+1/pIpudv
+nW0tdPTK2qetLHg9Ozmyy8DQdQnorDEvFaatuwhrGzi/nAun1F1m4mKEroThgkd5u3wF6dAAU8m
/eI6scEqn9bhUwFHv8G1UMMoKrvN0bP6GOziAoj8lwEnqYA3AtH1SOdJ2pYhYGHHh9M2BfCOz0k3
P4saZ//gj5+S/Kbl0dFK0xC+v/Ax/iRmpputxjppryxnXApIWkA8EbCkI9LqJFHAv7e3HMwPIaRi
mDj3QDKc2Ma8hYeesdTyk0SzAnA6wh466ENPTC1LVvY5USW/LGLFNyy6F6YnN8Gfqj8/fYOAIy+n
/f7LPyg+G8C0UOselmRMgDz9KYhHix/u84arj9NTl8rYrm/BQx5YfM3ymXn2rDFbtcIdjjfcQzcJ
gExGduSbKAc+CMiPme1FicaSRPenvn1rmdLM7fLqzOSKHjkuS++dNHo46CmsT4EtSZdF5CboMege
NNkq5Is5m9iQ6C41SdiPi2iAM/xILKuMhMVl80fUML4l9XTD+bUToKNTOJ3U5HL+XdPR7HPHbD8V
D6QU62ltV9FJd3KYrbpk6ScHj6Iqf8EZG+eCYJIFS+sPJOXrOQs6twuXMZLWcrWV7eCEqruwq9WE
OIrlVcxDb2QMd/bSSm1rBZCBrFBFXUmCb002XS58/Ow6+orhxxrjvlLKcw6Iqfuvj6z9RoozyA0+
MRU/35V4uN9qH+831azrHWDSVlZr3R+stvpgaAKc+t+QIHVy3nt1aJoqWBTJaSekg6iTdz8g0zs9
jd7PQLdJNQ4UIzNEOWWl+FHrFjBz86eKACB8QWDqYtkj49fIoAKSoT71DdxhC3TKGkY4JECegQRK
ZA9bO3Ss9z81IPpRXV2ry2GEz1fBq6vYy9LFIq/xKUdDbiNRF88pkyNPKHsDFrs6hgASiL9wbZUB
U1wQgvFoXnYIwtfpR6j/ri6s00W13qsUKdEMpGlmwCaVDn7cxfrHjLo6JU0dlDHzEhqWldVh6t0G
Es/amy9SxEnPcL1Gq94c4wGE1e4Ha1kVHFkQ3GrElLlSCR/vsazG/P/lZ8YP2oiODhVviTnTaNgo
9O81RzbB2ldA0Cwwdmjde0pJyjgS0w+imKC3epKp1uBtEZNEZ5+HeqHDmpsj5h7hZlnxp2iIec3c
GGp6n2Uixow4wc1r4CwzF3pCVbZWHwWkNm68QkRcZYBhd0VxxLHj+fNbkg39rArOj4og6WmBXPsC
QkESssEwPiVrRBwf55QmkUwOOYiTN0CDrxJWqdUFxUa7dMlkpQTLftFd8FKgolPfIQ+kEVsU0O4g
xTXkmT3PyoMxCygz2voYa9YELPverumaUoNV0KOhEkhAEJHJXWQ8xkU7pJhze3QoQiVShqNFv7PV
f5EImL4+MCZEGZ+TFsvBMCoxsqjjW6uiLuWwTtIs3fzB4CVB1/iCrJ7LycB0mu5oLcZ2LASbg4sZ
EKJXA1xpevHFwXXL1VCi1PSVE2jp1iC1KcUn3TU2UWI7ziUh2gUWsl7eW/veEA9SBNChQKnCIY4g
PdHqmOyhMaSNhYq98HvcIlouW0+Yywk9Jn/MQzNWw91oOwNMSf4lACIsmyEkQqDV7DnXyHkwU6v7
TNJswCzvDslHFAX5s3JK7nJLr2N/iWoRwK29rV0ie/TlwJxqw5qNzaoi/Aj8gc3tgzoMUtYruS3Z
2gfjwNHMUN8W+p+/1XwyTz1OGQdmtUwPDzvLnV0NjyhlnRhaViwNa6Za+nRlWpjPldm+Lvo0YFNz
HujmsTq++YZZgTZfNgOu42QSSaKx+95xNTTQ/g9EED1ycxXUnT/pUs+8uEszEJVJnQaew/dURnll
nWYz3CDR2wfMmhSriOWdoyDbQjBoCMchS25qxfi4sbmNxIPQgs5HjBaYbn0TrU1wgEVS3Bq4WWm8
Tj4PaMmw8cUpN3ZADb7R4Tzivqh+dHfTPvt3UE5e/uR6nPAIYXW9by5zvoCQ7lfq8/xY2W1+YRMS
kZ2q/taPOo9lnznmxXxw6P/Y6nHz9fdoMlGH+iClMgx8s+1l1TeibOansQD8nTWoDnPkeCifg2N/
85qdkNhw+rh3oGtkPxfvE1YjajHyvWXWn4iSg/YCK/C4ZApZxCWLXY4Y9ndYmgzjvkvR3BDr2zhF
29RnimcbT//CYkhpqAbbRdSsLRLc6U8f1b/JdyjSpR+LhJi67un7QuGdq481tDuRNgOrGBZ0Csbk
9MD9DlVvNGwIc0OiXxNS8IW6/B4kPkt+gNd8aS/oK9URG75d9kp7nxlxjmnUb9d8WqWjQXjkOm11
Tmpha1SM3kKwCCtkkWWuaE4PSmXfLr24peVHKhT6usjwPZCOHGONiypP/+Q3FszcTNjHPYso6dD1
4uzPqlp+KN0T8d7gEtqlZd+Eq9BquqaJ6LdQOhjuEAOjAmt6APCJc6Xb5aDSuGc8/mCjiLalasBc
bhSMbE/y0q8hSZmIIM2ENkgK7GEUvUtE5PXpuLWlZuuBaWJaXUPrKiFs+KYIzW4gRiakK4s2OnPL
+gML1TfUIGxspBSfC5nly5WmRt28hUun1TsPaaYrTLU+U++qfqG0TPgcT/TOKGrUn72fP3rFIZ3n
xiNc0PkT7CxkooEESSILrX7g/b9qNab7ZR8QUtEwKM0giTXFn4O2/8eAJD1W3c3wbaqx+FyhTtec
CIKNJjaQ0PUMcTw68lvvDzHrDa/kHMidwkzJJFCBdlw5jLivqXsuFsUXktH0eL0AQQQyH4K+y5mQ
vhaqyYSIPv4oBjQzYKLM2ZxvDw1MjSVRD8GQkuFxl0Khyp1tNgXT/YCcw0dNXlfRjhbW4wMtCZ2D
fKysi91J1kHlPqGL3ardZkVbzMG6i4E2OkNxRRbqOUT7bWPTNrEp0cr3Ha7evOQfbeIkph4hXxGv
gtnUUgb3BujFie+DorvSB5EzJRwOavn2eERs+XF0bg0/Tom84gPVU8yDeIaWSOtfiK2u705uB8Ej
Ykj/aPb1C1x6Y+RYJDdz9UClXSBju3Xr9xLJCo1UXBPQvTnX1HhFml73QMAGSUxZCQfyZhEvx9y7
COJ2Tf6V3drehFMOJm3WuAoSxZotKqv6FCT8/5urgZbkxmiLvTdC7IrvG3i92Unpn1TLDrzk3tjs
Bcn0IDOtrIZOdXraxIj25WFMb0kRVKdGHa/V+qSb7tt9cBiFgNb4hyD3l6D6sUWbLt4BAMYftU6d
fDBuRh7Ldu8CBXKzVaqN1XK+6HyhPEODq2XDJvwYPMX+j6F9nrrwvbXP0Jttg9vk7ty91t7IWahR
U0bYDMcl+6eXmMxK8Q63aPB905Pk/ZobfLnGyd8BGPArvgH7wO8EXkq38vNIcJ2IXmAnjoXFIVZG
3zxntJmp+Rqwbv6+NfouBrlDROMZRel4NGdhgLsyCrJuoy4FLp65kn2Ae73tE+xawUFEmfzbLbtN
4MQc4scohPJebj9hbY/Rdbp3I2sQptXJ/cUtMlCCoJHlDlIAdr/M5R+XVymWzH1kSAHO7BAKTZ/W
FhU9LPiKq+qdI90nILQLuFVLBLI1Mmy7qYiNVohJ4QXMdAjS2ODIB2j+GQtMM3VQ5zNbKFinG8F2
YxoZtNABUFhtYXHOhdmTEbvguckJACJupCO5m4RKsJ+gN5hWKn6s77MPWSkguc39rlDypTr99sDa
MNT5nUdQENh/HqOxqrx0KL8JL3AJLcdDJeb79ZphuPEYR1RCHghLacgWkx2qXjzum8O8v4EVkdc6
6kT5UE1QZZIEhVZtqj8K+Ds1tm+IMThRGqAaIZowOQnwg0a/99fM/zHYZCOY+u2MDSzQpuEyiMIr
6HpIWy5kmolG6Zg96IY29RAhcIiadoCyiGURWUXtans0zDeEY3TWw99AuSqUNMwRwpbB11L6jdn1
12WPOXsC9iRmPzVRbHiMP9VGxNRO4npLUcpJM1+cqJmrOod6p/mIYKwTvoiQSxMcbwiQdPbfIsB3
UfjsFOj3N+FoJhBXD5yfma1tVr7Hc0HjBLSOICK7yvmGDFhx4+bnSAYjCM4Xtv45GdTGcl17reX1
DA9WdyIEMdrDpJTNfPUsiFPwxXN9uxLdMqNI+aV3hE13GgfqZtdaP2R0NCINix1LD/opsyne/1pS
xjCz6o7MgGRoHOCdXRwduYFmrF0O1IPd+zbpkc83Mfg1NZh6V3z/0ntHU4fDhHlksyKXqzKDWOOE
gL4InMmTV6vPxDghwJcWRlkeXbF1VVmLB/qmIUdECo1fjfeyucutBDdwINN3zpW2+wq+w6OD7biU
3KvNz7D6dMDu2tdAZeTKrWoi+52nVmESdEK7bLw9wx4syw+px1y1aXXr6RUMRUUhi6cDBOxMKgHR
FoJ9sTO7eA5CoUjcBgm6Jri8CJfNTepnepewsu0XCIV7w8JrbfySZ0us/OAyGxfyXJi2kHoj5ytn
ZsVpjbYeqMDmYKXvkQyCW4r+IfrjGg0K9YQEFZL06FrGz8xRqGdq3w/HKYuN/5GVBzwCcUcLkQBG
InSJWY0/KcKBT28k2elBbnGUGYXTDsaSb90c0Q1k/EoGaKWtQa332DS7hXAtMBlt80dZJcuQEIx8
lbjtT1XRseRYgODU+ynVzRGg8Zi4BHINlePzB7epBcwH1g/xgeJ9uSs+FW8HQzXPAJjf+1hO8Jk6
tIwKp83KXqbqoOluHruEaYvRSiVvF4pfFUibCKOndHH/R3v+gza/+X6NEidVuVkEEC8wtTaO1np8
o28K2bZsZ2NlP8SP1+ojbEd+31gcdMBftTg6sudf02IjsHLQG07ORwEiQuDH11Dn3447u99O844j
ncdwWqUFbbTbFGciKdyM2oyQaWgz7DBmDQ7ZxGUHi5E7QF0cvZrSmc7fVf9oeM7xX0jOBxnYewIQ
IwkxkduoJPvYkPC/BK1g12hn7RlKLFVtcBK4/KmrNXfC7sgeLZe95IV8t8GYSCCCTEMV82rOuqdg
zaTFT0X5iABJXqxtqhbXxufVqWoBmlxlA/Y5Tq+XEhDqGkflJ+EsbD38Ne0VpTiNFeA/h8N0QELK
jwivww8WqjnGZkTRQ7mBzuiTuaW6TL9pfAdBDf3QPZxrx8Qo5v0NaP+8t8ubWTzpszOAFtRgjqEO
NycvV0FkRGl5ScciK5J7MMPXHQ8V0D2pZZ90BXtPHyVSaOymS42W4RJeZQyIWhIh04o34C385xKH
z+JwTjDUwAWx1WZqGy841EMir8S10BkIjAK9LuHXeq2YIxAVqsVkLZn00jd9PEAdkZmTKlEazF6f
znMbMv4zwj/MuUyt6fqTJnQeL7LL+w4LxLQo4YBbYx0a0fsEEmHflJJ7L7SbJ1wheMXMo6Yd/liT
eICj+LHSSvkAxayZwxah3DpBeMsrTjqfEEnQMww3zu601X35Pm9Uy+u4DXa+tlz/M3HspSlds/j8
uqxpjxIvCI6QPUHJpfqoAWuauRqQmO8cP0IWaPfmMuFPvzEckKw/ZmmAdhwVaztI7BNG9Ou4oYye
0kBWyhy2bevRW/86ZZow4WoXWpmA+Q915wfa09K08kmQbfDzlM/TMeNZ+b2IDWi1YWVI3S0Mmo0o
/Kdgct8hHKsZUzGmfAgDZlS7NP/OY/6OmPKXhsFVMwXHcPKp+QXsadEuC8HW9K61X2pJfLzjrxkr
bqyeCHyiNsyHu9Ro88I/mmPtulolCoxiaD3hKcynDNI7pyGxYTibldKMXFujvmy272TTtVMNxiM1
dVEjGYKkNoSHVtfKyalvNwhSH4ss756TXFbOO85MTUuTcGcFcsP8tn4kLVZ22EZJuwSQ5EPNd4vx
RJfV2R9YIXP11DPKWC3vMCvBWBTLd33evI4Fb4uRa/mvRl/OM43n9G11b7t1Gh2qaHzoWBv552WQ
lFC8Gu6AQKq9ufxckuuFMqevkhBuMVRC23NXqEYYzalDoftPc1BzB0wuncMAyjieGvrfnsTrYYss
nPmG+YEJRa+dGuZdx3ousmtX0EtELrdKlLh/A/xKt4IrGyrpQHhHHK8D4dhR4i7AWAtAGe0go7Gc
RdDbJBhCNQ8E+RKeOXwbGF6IW2VMTLcwTNadUqH15/PgZhOYdAKkMai7DA8dZwn7crNCgDHssS6A
bad1FUdqh8Q0mvIdNYcKOHLSSJgVvE8+Z0EGkGtkCDerH/DcI8rLewi/NytMrCHFqvsq/dPWzSvz
VvYlsWXY04+V3JVkn3yYTBTQ2/Hk9Aw+l26nEopx7nRaXt7xgqYNM1UTidonv69JQqeQ401qGbbn
DKPW30CpWdSoZJqC3zzrcsPLKAqbOmDVyDZBeJFwN+1MZhu3cbSOCB+UlvnONewPg67wo/YJs8D9
44NqarPrLzz/wcZXuk5XUQGHEKkxS0Nv9YWOWv3yFY/+CURyAlZKBKC7ZkDove+O2bcVNdiOJv0X
NG7ZVMwlK++ddm6/s4J9Twly2+OZpeS0uHbLq1rZU6DZ/G39jKd7bNX07j5gAfUy2U2D2eM4IJSd
4mhjL5o47EpfXpmJMXbW80VJRX+HXpLL5ejhHdk6tgeGyRA4M9HJlm6Gv/B1Bi/MqMwbYfQovvk4
btydsi4GxBCP//SPW5a7JJ3wEBSCfPHb/OhmMCAngsPzbRZY8CSnz3vnPl8c6HURLGUflHMyv1u6
xI6NtdQrPAftr1RnIxpgEfj8bpRgow1KniKsT4KdiPg9w0Dagj5duyaxsuFVg9jRUXSTfXK3cQi0
uMqrOfxwk/8kJd3qc46EQpvdbLHcMX0hgSqZh6qBhwMrtwAR29uJzG5UkommeZxsbkoSxUvvPnEY
Ha35FW9eQzbuzh3ecyz0+5zW99xm7jUZoy/bR89CEAHqMJecuul5yecAlk2klnHCJynjw+cQlMWJ
v6gSwEYWmaaeKBUbje1dxENvorUcO9n42eByiaAtzfEq1cls5NpHOLyh1WW4BZXQy7mcnp2bZCJk
WhGRhLyWl4e8CMWHd7zBOZxl0jK/aAe5XrzK4Ep/A88hee1jh9YGqLH7JAINK1TtRAQHXHj/B+IH
Xv4MU7RX9pNrReqnLQP1p7dF/+V1nPyK60UOdSPchYze5EYFh9LLE0kiwd/4ziKSi59ORczLHZP5
gY0NkTgdPRo+reVIJ6fnFBByFOKAG4ze1ZfIJVioSuCKRekM8MCqVqPBikoBixckhPwHmn7dOJwm
CTENXkln5DPn0GbzlMEBSn4wckHmwH2nSyxECXFAwitlqqDqLHbSrBsNYfyKQwHUuROhIx270pPy
NOKCAr1Ss8NqMHJ3lDclZJgzVHIz2HHxxvLwRU7RmGThwQXYUAcWLgYahKYFYpCp5g/lI254NOHQ
Gg3jpURsHXLQdMTnfGfXIQ1KWsSrh2sO0MJQeq6ahanw77mDeDX9A4gTqdUgNSqzfV3iw3H+LwHe
A/NmjBxd+WknEG1t2JjxB0OidaNN4PwwMrCCD5GZHGv/S2EkPp83jy3JXSDo00DhcfsD/19fiahR
g8M2lDn/yTnG+XG7p/L4B0y4RRjzb7qSwqrm1UqFKNmeKNUu+lyTR6qR2V1eOlHqxWcepuQjyH7M
dUyzyq4kyXAPaGukDfi8x2az4SU4MBcwhgf5oHUApnalkmJO/ouVjnh4tpKPW7HGsNvR/njkxukF
MYoA5/FwQNx59q6dEsgg5z2iUKT+lljZolPIKLf9144iCfT+4/5Z+cQaL6Qp77XHtPFTE6SoVgAk
CVFqVjye6cZcPRxjpRvfawcpoDAr4wu3ViXCZDOkPp0KTg+ATZ2YSKtFXi0mrxYhMS7lLOOkmjF0
Q96QElirC5yhMdZ1XUJxtNbn31ju6aYZrnlGAIrH+OOMKp0YaxOEwPt5zah96TuuNBuW+fCZ5xl0
8HYRxhj4ebA5gY6aqK0zAQEJfROC5y5sWp6xJCA/CfspCxmY7Gz66bchLDNo2Z30g1Ndi4mnAJoS
J189RjWXl7pauQPIqn5YiXXfCFf8xDOuvp/wCnLYFvNpNF6cK2FcfnyO5emr+bkS2AQ1Vz2ZME0x
bCbwEgot7lDRrXulVikcREhT8yBlI9hqbCfyNbsztwqVQSRaRIMlGulcRjsh2kRMOdc6Z7LZ5u9H
LSnbGp3RxfnaW8TKIe/SrM9trzATEf3Q8MoHUqBFxRQDCLJjPx6EZtIphLGEOesQgXhWWUGnIQz3
SMV9mjXoKjhsIm91KppzIYKkfCT4qriSIzs7AZVOZDOCqVETsIqN924SnXlTybtPx6vwqhT6qaWF
0UB6F5KjcpjWwoKuwoAvM1aZq6leOwim79fqlNZ6Ssfj1rLNjbFQCJCSNB5oi6Sfqo0DNiTIceVo
jeLPAe93RjPqManSsb+Lqya/buZYjQrj2nGMSAT6FQAkRxXuJbOKSrsPgn7q2KzmH24iDlnRhNAA
Y3mpIVvmPArh6IjwBkAubeXcEi91HFp0HnjIlwFy2BnGAkHWwEn/VAQMkB5CvFPwgLZyTwgtXRh3
jiD4+fryxcp7nrsXr9xfcQB15eLld0uyZitivwIkpvFgmQD4iDw8xKyP+sbyo8SnRdWmhViju4l/
nDlWNAx9C8qByLtcPb5+26t2ILPqGhefHiiiMO5z1etojhAAnVe/gwQBZfIBf5TJG1UpBYSn931/
MUvRybIEGGc0P15+JYAFZMVu72ulm5TXm/LDOzpikdGo5lkou9BRihjFi7mz02Hd9l/tJd9joP1v
MRUrScwjuMgyhSbwfnUKzUF/XjysgqdUMXpyiJE5W5chSQ+X5ntU3UQWnQxv5d1PP/SJt1gVd+6I
04C3/tb7PVvx84jFDzW1w4oijFEZaGUPDho+KBn8LFdrr9rUNNKOO1ckUaiW+SH2vVNgpNuZFtOc
LwZhqxmLTqKA6W+GoWKdwhGR14/pEF4eSrZbjmaPbKZVOtIn0YKJD0NOi8o4sVbzQ8ApvQ2N4oz3
q8n68A8StOEwc7AA1l8Ma+W7g9liCNSXHPQy9fxopdZAAYE/pbnK0RWZtIkhK+Lazy6cEuFJ4IEa
fdxrnzzPhkg7EQ+wcaAq9SV2InD7PmzZSIWU6o3JQEWwqnANqf+7hwlAawS6ht5M6kJR0mwrzcZg
KsVoDjjzrBeugolsYttQJOlZ6uFRDMGxCFiitcqHkjvHH0yV8RRewFQYTu3/5LFnNK/gRHHNteZv
jdbZzevDO/kQln6tF0jYuPu5I1z9pbzaeQ7ZQZdz00CCstdX4qHV/cRI7Yw0XeKjJE9D4DGMc+cE
ojrbtj2EhUWAUgsp4kl7s+ZmwzSOZiaGJcXiqhVViJyn5W2aQ84KLwCavU7A5KckSsSQXnbzLuQF
BQvFkY+jACpnh3E6B9sb3dQBX/VDUIFkmcAP4daCCbW9vLoyQi/sid3UAETlnsJONxQ7MxfkBaag
436zKk4SDoBMyTcF4GQYM25Y03mpt97/e3k5MfOdpFlAw6CjZUdVYT10Dvraufl2RymxTW683ldd
KnMvN1eh5K0xiXVpvhvE0lMqgBx+ZWNx6MiRFMLo2bsucei37yggrpA8qONatHkt3O0dx9ZmYuGy
p9TQGlButQcKR0Arh7T6j7yIIXI35cDWJUKPf5QaG/NIotfnE7rdjm7H3DXMUEEfhhVUOKYt1Yfz
j4XkKjFLk2UxvSafOus7kLs1Tj0PN6s6eGsODiZhFSGZ4h2fcI6hbt95y6NL0PH9z3mS8i/YG0Cq
wNq1nYyZniP2g+8/I4s7EC/gBlp3m8npln8SuJKm9vEmUOzRnr3x5TgriDxa+Y03Ao2dtWPs/cuf
89WgjrMAAEu9sWU8YOTW1C1xsfH+Xr0DJ8xzmERXgY1Mznx7+szNz2o0CJfQnweLmPQpO2T1vrcu
7mGkaanSj+xfZEFBWYjt6+7X+Gv1ggVeP8fIEJsRI4+sTN7ZnuHrU1MZQqnvDmHO3W3qBShWpIDT
1awkNKBLfXSluXiFmfCwFOL26W4ZhCacWTmVrJAQP4QDSBFhSMeWaThXkhHpmMKrhDGRS/cwAcAz
noDgkCTQspy7sTM3nlTwFzsqVcBOALNv6+lkT9Q+W8Xf62fFU9/nWwCMeHXmbCGGt+bcgUlUFgHO
ZVqkJAaKuC9/QappeB7eCPBZt+eL6RDU/Eoe0a+oz/cg3TzZNh9OUduiJw58LEfvVDuGK7sldJn/
6aScG6drg1Nx8PkIN+Cl04j98ByvZTGUO3e745SkT1loFU42NpuOPOZPY19fqHmtUEUMfP9lhRg3
83aqLJJqiXnYvuQDv368fLDlFXJih++tGEhzoObkyYUdZwPVAJz0hjOQCYeo++Oa0rDzh2Kajeyz
QMAxR5VZnO1I57RVszLdnuSZTCCxD/xukRoxxLS3TsusU5vPyzgiXy/fk/crVnK/Sp/eXWGeskAV
wPV1/It+uEJxTXPrhZJsGjMBh+4qwigSUYBlXsvpUoubfNzVwgpjT9Ank0bNRN5t/Wd1kydEukpq
TDwO5tT9tDrePz0yvdyW/vBaxeRFa0Y+i+qL5iCTQPESz1UTOiPcOnFWLkbxeojG8XmmiYwiWQQu
x6L8h9ajbFHrVdJJWS2vZMhDUUNQK0qHHXOoKEoFmgHbSCLgN+MYJTfWNEYcCN8G6ePL3D8odJvu
RqHNIPOpX3b1/p6YapWyHJ0tnzks2EI4bLMYuswESr9Q+K1PWubb4xNT/9rs4RjsCA/JmLKDzO2E
NL2qh0uIDj19Lyl7KczL0AFmfpIh+AzFwU7hTMSkzZJHlGacjZ+VKyDt8o0y9OdQ4mtwuMgTV+6j
8WCoxj+3uTXSG5fHVWRLUE6decMCmLX0Z2+/hIWiCfixMJChdRAkeLzYo/GAgMW7HzNwozk2BiAE
eR19EKyK+LWrfaTvWrRvMKt+p5yxHOKFbIH2LpbCSQlELVjj7fQd5e6+6v4rU3bBFCA1dwuQgQSg
BRyGK8YzWBiU9cAIfVVKEUuorJXQuB5fXAkgTJEirebIof63iDcddyUTZV/yBFGizFZ2K5fdWlTd
yIMLryqyqPYdAvIflMwytcAoypuxAWuKFCflMlF/w+li+S1D+bA922/FlJ5OUsmW8uaiJ7r9X89s
asiiQNNKqlvDkByI0kgKKy9G4L35z+yNVvwv7ZstL82cwGEctDl9XuNYyY+GJ8cMx0ntXqiOPQcv
+eyZ5OJKG4A70bfbqFYaV3ViK2THtJ12a7tKhKfTVh9pjC9duY1tggPXXqTNC0Gd6OMYyP1/8hY8
guLslc4WdtVik687JTYVaI0uCi/9wXRt0sF8BZa5V9pgIfmIVXK+GKF5QkPalw5OJseCViYHAFjY
UyM8ctevtmm/3MY1YzUvweIT2SRoVMppd8y7843LVIaUyEZEVxPcTQFkMbX3qW1h66QectWb0sp5
FUlZuCJZZuw801P6Z27Md5gu1sOHt+eA7nRAnMWfpkdI4VDUgbw7rnyewCFcq/3xSTDPruZkdmHX
APveLAWJALDNL2oAlzEOPv2vWPMLkfiVNwbNBONOXZ7ZXLHw5EysBoEOn6/QRz2B8JhO8GJ6gm7C
gHmmBSTZorOpRkylmHg8wBL1TSll+BZuV9oL+rroVOLGCfp6zoryHuMDLtEjQ0vNKjVcRa8oA+3r
FFzjdJY+Rc/g9sZ+eG/zWceK6SR+LWBLLqZ4bJoZcm60zhZphadB5TWbUKXgfNckxVN4i+utMUMi
KNttnMiGlXOLihMESOGNiyP15RtNOi5a56megfisYtK0IZAssuBW+tG0tefO26OASS+38lJUZsAv
fULEbbGQoNzvRFwR89euzO5rKzLbZf5Buvt2m8cltgbi/QGFEm14X1I/0oFmX0wAJ3yycUcb4MJa
ccU7go9ere7JwW7z5WPx1dqnJL7guLe3LbN9DAbLPgHLUbgGy7kb6bjCREqJ70A5pP1grndSW6SA
1AvSCTa+2UobCojKxvQ3aIrqNOPmU6n/t6TM0m5akUUXqBK0iIC0cpWmfRyAIpxntemWdVd9qfZ+
oFiD1WZxgCf4TpY5jUBM6uhWAhilosU+OEjkd7HkcpjY8i2D5BfOjMqgDo2bFr6X85poG534U5wc
HNHxCKRx10FeFYOiNquhpg+iPG4PtyFZhw8M6GO273woaORH7ef1dwCDUY8Fpm0NTi/qjUX0iXks
p7zn+47JXMfzN+25yXaANGSnYTh/yr4vkjk7xkyF6kX2SHLvAAPOrc0Hdf8fa856vbMPxL7nLsp1
pafFOe8I9Ngb/UhMifhB2FRUv7V9LN9XfS5p+FI6VEmm7MvYa7T+lhJ0es26uaxXm7FXGEcKt+ZR
jpp0qtOp/vFBsvUUEW05DV7zDNbEhie85aHY+ezbXuC6G0N1pmTAagBl8Be2TY4JrR0Xhf6AnukC
tmXwjX/d9zEvX6mDocMA6veBvy6eZJ6z6/gbNcN4RhMynGwItViVQNPyJGW8t32eAGMjeSZMVOzJ
C9R2/TIhMhO1uhZqDa+Tel6VuIu4ycXQGDiXXnDIY/26gflJZH9mGuo6aimcBJLlrxtAfhUQHsgJ
3O4imanZ72S6irVDWVQslLpcRtpsn3bZ7XY+UewJPRjwIYCgtegwKkjQVa6A48VhOCdNrgTG2kB5
U8yMlBLAb7Dh6pnpW3bEcO/38dL/qrwdA6HHO4m4IbCEU2hKj17bioaCQZOUqDswe9yfdxI4mf1+
0vDS3FnZanekYnU3souSn4DEalD5uYyDB5HWibGv3breJ6tX1RMzzOm28VQhbrLxAYAtL+DsWJd+
tumUChEeolAXSHDgBQlV9bffhj6WNVAJKjpFxKjmeMpUbKj5Psi1PAEF640CUGb6Wvw36Tak/hjm
OU+4W1/BoDNQYk9fZv9Bslb5oxC8YwHJm6ccJvvVddIkYYgUIYCKPCYRdVUQXm8Zyb/fBquutXst
l6bTVcdc/Li9IQZcOIvUQ46shtOKMsjubacgaywISmUt60cFFJjXlEAAMEVdznibYFonlk8O5zWB
D50fMQpW0Iw8bc9q9oQR3LGtcVKxKj9Xe9lZ5OKKMK11anjAZwf5kD1gllpMPXoIEweNQ+FawdoN
jqV+LEKQXdUpOXNxR6nh6zztbNmu/dTHi+Kol/3nTtF/FpXG/kGBR9ZOfBdccgSD9QJ3pojzCwhf
+quq+oR57Q4drxAWalhLrUl0k4VdD344hOcnCnGDEDsMbrEsE8YFUvlZyQhR4kzu/kj+XR/sCE1l
QvV87LgX30b7cZ2tNcc71Z2RCCZBdYeYPfhtoA/iLH5Eu9PxIAiKWmMC48ed1YpBNsc6016PFI3k
M334R9N6j5QL9lP/f43YCV7I/uEvVEAaa96h0NA1Rpjsa73LWHvqguUxPB4kggBMFriXC7bze5KA
hu1Pjabk/oJxZICS2q7zkY4TAeMOk89PX9v8BNW5QNsg2veNcvplVx36+PDWZ32LY839vNpqFSAq
goNOV2caWRdfempkDHzTYlq/BlKdpY+DkfW2cXk4r7qMGSZeGeHWuLcy1iM/rwmjfeZA2PkDHlBn
WwLQajG42tf9dyA86R4ktqsZpMlVK7NfyxpsJKV4L9hZm3cVmi8tJ7u4Y9dCCbNx37iO4r7dE3uK
hyn02KYO+lcn4AHcThGoOusrCqdJIaQ2+udSJBwo7/lBWGRnqvryiBxy6FlagnVhFvD3/pH0vxrQ
egjdk0i+6tm9UPKUqu7CKYh9eyQk7v89Tto2apH29bb37updbIN/m2Q6Mvu3vZC0EAyKsN+y7uI8
NLMDritT3FxmF1VTSuwvqq+NnOVMxAI+eN+wLYYONrWe5ACYzZU+7Is/XOG6/lo70IZIoSL6Eepu
YrwA6RYMdXKTQxxkMxgxd+XSbSopBMwUTL/UkrYEU8zFuxbFily8Z2bZeTr3bC4km9GOlZG1gXPA
Uwd/Rfgbd8wOrPFhrrmaCoAnIJn1Wgh6y6Dr06Kx10tMJIknFMJ7AxUZ4A1AY04KLF0C//ofoKqy
ywy0upydOCJjfQBJiDLD1OQ/VZB8ogR34jPfCBBVfy0Glcb6kr7IVd55izvQSXu1SrJ45gxjtSCw
J0npkxiCYk9WmpXF705vdSfNBnC7KNF4PZgPnVF9EbqwUVhYxw5c9L0glPvuL81TCmXJD/T9dCku
LbsZ1KbuwdL2KPJcy/piBV+5JdSVAUgDp2ujR6d92/mi598mKJg3gXZTxU84b6ecPPsP1/AWFGel
QqWzuTWDZBHUfKgOg0xyTLiIQiCiBLrs+8B5U2KOc4XQrO7rgaZKrJlos3gRJ/qy4WF0hP9TYYfm
I9lqgaIeOjI5iQmeIOoKy0QNC+kQEljjD4wVIMQbUf1NOqo6okyvJBHDnBbUQvJQPUlkvGEwNZBN
FYNN+mLXOi3Ph49gI+G4nWlBTovPJ35uNY8TSfEndYE5iQyWs4OhgPkz97neP9xPjhABQnMPnFqL
ldu3n1rujd+yAdskPqimnCqV7evfMukbTJXpC6JtLWgdUYVDuuaCLT7xy4HwiJY7iPgrrNfAgdlN
WbUCzD2NWMsWoWk1Nm+kKKwmYGIECrXCA9PnMEGbLcuNUY4Vc1mdoPu0lQxCLiyDV9DnHDPpX3sb
Pp+lCHaAthJBanPrFtOU5vs/1dasuQks4Y7aPdCeFbMrO0lxzU/waubCT8JWCS9MR+S/aM5JGAlN
dfnejsAVYR39jv1oiTHcBFJabnXOwhRQDQKWYaPSpqVTJTmTNQsIRz3U05fOde+bsu3XQD2xbzXf
G82/V6JPmnuhkE1BeL/WzfV78bQi4ZmWxVBpVMkZkeTxYL06AN+owmyq9w6qB4p9o5zPwBmzDyZ4
/Cw7lggvUiS0Ql9vI8nsS97VGLAQYqk01NdNXKLVxp9gpQ6G1NzbVn/R3vdFk6wNzX1RlzoCVCyN
0kRJpjcPUeWXiU1KmZp+p7kvfiMbNEtiP7BKUCuQUfeaHHKfFK9l3boQkr4NEyPugy7AoRcUwdJX
wYyKv16XzVSa37OEIiyNWgDluey6FQUd0BqAWyu0FH7YnP0UBRcBarufvqEdtiPbLoVHx6K0vyr6
tPtMKYJZmVTZCZ/tQfpoEY0aTNNguUv/EZwUim1KeBOjzYMD2r8wHhdBTQWpdhgNJgX4fR3uIu+J
qhxn5Nmsqrr29HshunYE1JTHRPYUse7yzd+8MyQdxF7F32YoXuHk7FFMHk+WopF4yv5P03QPY4HM
45pqulKBMhhV+qp0oTzgO58yBSm3DVu6RfM4rI1CSjepTcwUoTCt1+sbeNxFgTPS7ygnVbZWU8hB
+qZbIvZ4hNAiPbzzh6dk3gG4rFOHTDg4tqR2Vl8iDmIR0FJI5nZOslruSArBi401+jdtZA20w6GQ
cLYsmmwUCGitWReRSJEASgdglycQDnSMekWW7cP5tLdMteVqSy1gVRUqbbzxVJQraQfMwu8yk0zm
bS1M5NdNFNdPQAfiwtyhJ9qqScqTNpCnS9Wo4Uiso/xVrgQJptvTcd3ErZNj/8HiDJk3rFE5cMKy
Gx4EHfi2yRRVsyN7XcbEtOCjdwB4aJw77zMAAzfbeyGWr+dn64/Ngm0S0P/SbOfzdUEdew9vCfxn
wElIzjKQqaQ2DvH8/NuZh6daYtvbITLnjdOsiNJC+DW1EaH7UklrhpGWGpeLdFJQHNsLmbY7rSl8
yXK6tCvUipBMVZ+NEpMTgc4XDZTIQ4+TwTU5KobdzBTJt6VNzoUK1vXie12M4imlOIFpMWSS8LTw
Hf5PjfTeUmYoAajWkj84JxgDJurqz9p1oYTvwmjp3nJGTEJZenH1t3FaCcAc2STWnq4aDD4wztTL
loLOhX88khD4CxWhyz1y8TLyd+YEMRlCLikxZ/W52y0OQKdT9Li3kyRfQ2mJgYhKjr9wStm8oAz1
diDcmPHCAi7gV3sfzssuPcpaZNH/QhKuFmIHWeQGnc7EfwjH6EHH0AcqQMxTOzbOdXNk8VyRjPQi
UsrKf1B8g7IHiNlwVRaYhMk3wW87YOeppL5YEZeQME6Mzl0539hZgkLz7GYjnAchWh0mEYbJIrs6
hltXxuvFIqIadCjlUalVX8BfYxtI2ipNcbF9Y+/9xK54CvoLh7xPuuxNS9nPi1ymGHH5kYzPoS7B
DHvh5Ip1kZpUJnHZe9pEpvBzhFjz8oWlWjWK6Q8ayeB/7DJ3i8+2GKIz9U3twFtvdlWfaL/5Waqy
WV+9j4jcE8Fwyn8O0A5B7NPimAfbdK/hn8dN0UfEhWA8jmYAa5XF13PhHwrjWfTUX5B78QDRmwSL
2CnaxmTDXzd6A2Z5j2Jv2oluFDUBxOeaKMUUGtUTb4CT88KGlx2X6/Ct+ofxp/5V1keh87JxL6tM
dtuaTP8gPZKrNA536MzIEnq+PF3sUeK7CGjfnzYEynCYRYJsIi6NE7m0rvynNRtGggPu2zL2yAHf
nniF0eymQi3Ui7FnqiAJP8YENYb8o3ylPyFTMPDiH8dh0t1FPIGR5xxSMkKwEZU9Sa4ZxpKdF9Q1
upK0KocbhaEaav9KuTqhuJiGzgpBVoskixNELLjaRy3te0nWoWkalowwQzJxPoe82VBtXkR1LkNV
Fley3SrhGJHcanzwWxvESnbwJpF9Xri+hOrXEIMn8UOOfty9ejQncrZODsh7HP+XTfGpqbEKqe9C
XC+oZrLzwd4f1xYwYEkPMOcCTdg6zTZGEhHAKz5qpPVQTAvRyYhp1eBTMlpNPWSUYBpNjfoOu7vT
SwCdBSy3hx0OQb+GUgrQichvQrfjGPvvvntU8yZvyob+vSB3bKwKXkAYPmmSDPekL24seNLAy9RB
rDOfQeGkAw+Th6UvHPdhOXLEqmXvIdpZN8c9Mx6VFC/CTq23he7sI2US51rK+YCm/vjZUYqL/paD
TbrzlgNip1kr0FDL6669M6ntnsuALd57mF5Kec2qozT34khiCPbcOXtc1SUFlzupwNKfbyGbrj/d
q7CZBtdHWczlfJYiCNev29ADL40kjoc=
`pragma protect end_protected
