// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:51 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
T9y9xtEIm9JU4YqYDgKEZAUNwNY98b6eR3KBCTD35LW+rgfPX4HVoSRxGjEOIfNo
3zet/cYgspReswBSxyA/3rqvL+UjaAFOdrP3ljtrnmPe4Te89AQxvzpRcb23adTB
QsUivvgO7lftgeXm6D1pxchLoGV4OfGyiFhfCtwUhkE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8224)
R4loQj+Fthtpht+ulCEMGnbOV5eeVXZmbqrg9fmwP2ZZ+W2kLrLx+/CDxA/brP+s
zqMP7zNvQkRNRokf81KGe7bsOxU9yhBH42sNmspHJ9GAz1dcgag1fKHJOOA3Qc0z
v4Qzs5AK96uAF3pFd4laCmfLzNo1xPZQV7OiJCQV+D2Wl16xWt2EDPV7JU6Saxuc
HrZk7KbD0XUkemM39sXpuJIYbv3XaB6e1u0tjh8hfbcikWEhd7k3FH5XoC8GJ3wL
QijeSf00IeAB/SjEAE0MdNJWjF+78iyg+wT3bKJNF5wITqG4WzcfnQAyC4NhiV+f
/Ra09KTctNmmD6t7DUUu9zrw5pAfRwn0yt0B46T4tTDqiNickQlkWKawsuXoFnRJ
msnfQXuJyh29SFK1yw+Xkp/p0vjRQDJP6K45M6B0PJbD52F4eHndiDHdfOact2DP
kJ+hb/tOfjQMut8afxWNKo2Cl7LO3t0vlT7xhi/beTEREH/ZWwewA3zhYwmH55E9
4pmmIrG8QA71dXN8ILTEfs7mNfXbRdXQYR6SVfV/uNVo9+9I/OXaU72Q6IDrIoHU
Xp1tvnjnyhnRJj06cIJmEjkcrKNRSvmjGrJ+zL5Dctn4OuR+WVp1ApX9uBeQCZXy
AvPsLns73DJFDfhsXbz8pEpqCKGnuyuFGBv6tr4/ZU8urbiGVhRd2iEpt32SLg0b
Grri64YLUHb1DLhJ+0kCNqLbZ3QsUlgz77sKwdzPdwLzA6LFsHj+uIcTilhv21O8
GxsUCmrJcPHOMZdjp2clL7/SDsmh9HzekiYbX0arbrKoRL/rmY6dXLBo9XMxgIWR
qoQS3SoZjFe+1+AgOhvaCtS4fSH3NVPgFbKl65MW/i1oUhOG1bsEpRtfIKpd143s
tbHe6rCSxvlft5J21V9iTUrH8fDUVK4FlWLSFH5/3vSYr2EwPVOt+fLJrLZzPLvH
YOQOkRy1R14kjhxSN0Kw1GP2AeuQ4u8yteB0wSZmzI5paRUM+myDYAcRyZikeelq
ZKjcmuEqwmxpY/r98wwbk72bycpGG148z6srhG57eDHV5kNHGaLtsLvqt1Fjl6f8
e2UeAyZlyyNDh4ua/FyZzF9XcOrGOXh7UvAJn06cxj1LLAeGBYTqH/vuK430aZ6W
y0FWhASk/vvRRQAE+oeT1h4o8qYTtHyXbYNAmzqkWD+cCLlDLNoxi29MeRIJIRIH
wCTpvo1uILbymFOKKnRNvOnltbqjnoj876S004lt9LQUfXsTR1g8rR17rDciZWZz
SjR63s4vjs7rUN0cwcx9liB/PRYBNdm+9g37BVChdIZsiwZm/7cKhZqOXMzBlrU5
ILaWrUZC06gBZ5YofFX8vX181/VZooRjNviWTdsLRO8x8z/oBfXGtKg4POoPyK6x
IAYD35NxmV+8tlbH2jAzitam7jFC6wbZ6/RrkeGR74DTm+K4XzfzuMUGlUhUXHY9
TMCegImrJygNOyT3tWY8w3fxIx7IwGVJiX+NnHR1Bdj2bcNjpPuVRR8ZybO23q7g
uuzgpCv51aODkZA7sFAR71kvlyceVEM6wYO0Sp38oYOSAmbHJg+Zb4uArkuzGs9e
ASOOj7Z/3lQyqmShpi3AeUW70IndIYWaEgKA+YWflhn5g6gVB85kMt3aC1jS1nXE
nd+LN5xMZXBzJeHMN+VN6PpK64MN7tVA8Ivpxg4rPQZ7oyDtMztR3ozdzJRqcs6L
52P0nBg3Uqvyw+wP/cf6fAY4WO1blKSe8m0GsJ2Xw4FBf1rWFQOjqtWPkYnTRzNQ
Jdq2SkYsuE0HmYP/JRqPr9YspX5edEPT2Ac4XngYdUiDMqVwaGCgK3lLvvp21fGn
p3BWB8tSrOUF1faLaZpzOdOktM1v7bzv0s1to7Bzds1+ugY9xWdgyCbVOwC4wC6x
4ir1YcIksG3i/bOfV9nfCjIbgjbnqnXhZ/17zGniONZqYXaw6hrBPI7vZJZwkg6c
9y8o9/sTmW9CLbfp8Ud302cS59i5XYgTAQ3IfvYxArM4eiOP7ZLWrAi72GV6pune
+EJRgnG9w3rhSJc5wittwUuwPcM1+Y0qbIo3Z1rcaf1QQ1hF7o2ZciYMQ9hUV1M/
HcSW4Z1D9unZpRVjuxk2/hMWwr0lrxS9nocz8MycMYqNrQI3o9ovxGunYFKM3BV1
o/foBfXlR28/1ucTpNRZdCY/Bwa7zylZ2sZTMHc31acgCFkORmsM5abyH88sGAkD
n2ScykBZJX/RzG5CpdZMFbTeeZrwkdkOkZPweHSNRwGcVc2rhoqdxQJymdmK6DID
fUUsmnAV9yj4lHqNaZbZqZB5fgw6DZSYjnacDpx59UPGgY0nnf16NLV1zX0QwMjw
C+APUyaP0TuO3yDwfRlxTtLS1xuqzDwfiETsPMPHsOsQmnPJjWpOFxcxNnOZvZ4s
ICmMOcAezH2Nxr/3rtErD/0+Z5Ph1/qNLpW0xBFDjxQF4MXkRiSYFufvo515MjlJ
cEd33a699Vp5eCTRDaRweHIxQJoFbZQ2riNAg5UBP/eKnee1en6/48U3tLoNRgY/
EIoitWHb01YlHPpJtlCnurCHQ2B5Xt5ePnSIuszvptS+gbm3aPnJODlJMgxJcD6q
OVYYnUOLvcx75OLA9onFAeaWq6lJplCqr/Zhmt9ZrvNbHAaAL/IJA3DysZAn4of5
+ZzTzSaVX1d3x69MzBhSxbnRupRMgz4xm/seDJrRwCUeg3yjNWjiiq8He9cGP3BQ
B8rAkKbSdJVx9o4WXwaC2T0OrRCruzaY1GRMBA3xJQmLDgWRJuEv0we1k4v1JzSg
7V4vEvX86ZtBoBxuVK0niFeJsXPIc9OZIQnT4GU+gDt0b2RI1vn94lQ8eidldc9x
jWMgeewxu/hnJghw+iHqcjJiTIOuxQdpfbU015GT3PLm9LSvPa4NtC+i8AQSezgs
LFz1jantt4uDnjnjy1EEB3LcSdGol8+vDf7zBmStO7a3mUMf892HBhDRxiw/1U7s
eVws0LpYTdRA/Tl8FE7sjTfcfkjBXL7pKYqoGiEyrd2mW7C/IuxC8KJ1nQUNV4jm
6dGge8ocpCTKMAaxcrk6xqmo2OGn02/TjdPv3hbL9ZwP12tyUELIVrr0V+kwz9UO
V2inrqfYcdB4O36biYJZZmtZwCmgw6YnByXyzQZ6Q1qP4nr/u3iB3qcnq3rxs2/g
IEum3pYc3DlrcO2zzfi60+y0FA5QXqkomfdf+9nP4IMaaT5ztcYukKj9Gqa+3N+s
0b1SR7UX3GULzbjNAPMdhBhPSVtryX7joly0NaVeZExTqrdTg/lDhfuoH8UnWTKW
JcZDTG9fFLMdfhk++5LHu7M6CsIR3VdBabY9GxA7EOO7rsmmNbEG3eWGIZJMaB2T
5NvAPz9hQubjGp0I9SSPsamwpbOs+OdGHdvpxRFyh2k47wSNmB1MHXlMMyFkmvo4
x/7BOhNhXYeZA8kTWHKJBXSmwheUQV+wiwbtpMLMk6hBVHx/gImzAW83nwBNfZqL
ZW08hOQTRBj0EtD5DbiRV0ajva2oxB3GlLNYeDTUkr5Vbzu4+TLsZmiPJefuElIS
9DlNszy+torJCaaUD3ZTGD2cmbYQBJCi7QfjduZxNgIcLJdCDksfDvjFYOPO7pAF
vkstelaOeCxAO9WXV/Dl9F9Tao3prI1a7YIFJMmzK5U1aq3tf2WW9TNJUQexyVYW
Xz6V2OA7lUbsN0mjhfHpMWLc1kbnoyX0nqx6oR+VtPjVyHDZFmWuBk6m2mULPUUz
8jGlqb61HAdjbJPzNyfb3K2+7CBDlyrBGQgOD1pzYVPpkn2XEhchLxPbmI9S0445
gj9a8F39ibaLREaTjrlnbCTSr4u14aOsUlFP90SGF0c3UxOxK8+6TX2qqzqbDOqA
1QIsi7xMzzqL/lzyb3bYf7jjnQChkzWoPorwqbkTlHUHRLMw+mbmlYSgw+TJKN/7
z6Xn4Ko1l43xXuldIpReJ6wUvZPwiudvdhgDqp9ZUxQmruj3TiMZbyggRXYALKux
GGdGpVmlTCaolG4bg61W6NROHT0obhvv5ZiAth0+oUgAXupFLoJf4r7ESF50sSa+
16wO7GcbMtyVPDe1ww1/aeNNE7wkKWM1zsmo4AwAvNAKVVzPtz8S9jYOri5QuZDr
Uz3QZk/cNzWCnCNW1WLhT4njBumwah5UOqQtnMD2218nCz38Mhy5Ld8boCKg8wHm
Aolj8Aq/g6ElAkB+uyLNvvjWmxzPiZyagUJ7K3bGbF9Z5F9r4K5NPtciay5YIF7X
Ta34OkBDcyDyYEOlPo6e0AvbNkHq4BvNt+PVFpG173DhsHsqAngVpH+T5+W2P4qF
k7eIMnzDaH+BXZvroDfn9IlIncNcPNzFC2UARGgAU6qY7zhziWPVRl0Dq0afGEq2
dLwZJd9GXlh8N724heO53l4MqgERjKhu/6VHbG2fVGuZDeQ4JOUwpz4YyPvc6fXF
zkc66R8QxGZrvjLx0sq2BSZbYTdFbW4eL9BbTshmLNPU8+g/KkVBGGNf1PyRmQJU
omL76R3gWmnbSPuNznVPSDnb/3kp1RLZMydzVvZPZZ6tpv+kxZ2DskToB1tG2123
RZGUq59nYoiqTBj5NepvwIEdijlfSdADhAkkLaya/spPjoIW6W6mRzEkAQf9Uut2
h+wqHVyooLvtE23BlXoGZHFixHK6znzukBGgw2GzvFdXcUqEqDNEa5yscwqLZhvh
qyrQGbii9FCtgf2VuMMM4l0qmhLhO0nFxQJwQUX5xt3YOv4Kly7XyfTRsKBYleAo
t4a7DdvWE1EWwvL7P1++rFFUaig2tv5Yeo93q7iKX146zwMgTJF4rG2U0IkuHkUV
KNTPcH0N5TfVmE03EE7bIo4uyG+7/ENdCFXbo4cFBjvlILmwF1EpDuaS6HGZDrrZ
vCjN13qoyahnlbe0EngwtiglM7Sbjhyu24g9IXsiipJu9sCjbHFVe4Qke17Z9qEL
5Lo3R4iC4I032DWz75PQseQJggrLxkSmS0fM9+WId0/P7a+ZGBCh84elRzTIGMWS
+/krTKLcW5Bk4aYPaOAEatYqbvLK2PQ/bjhaOU2vTQUqiDzYk7OnG4+YYx1Q5ctT
x7xBl5v6+Ss5WVp112OVwyEuivnhlga3HsCbsgfv6V05Q1JS6HCPXV+UdBh5kV5o
xg83kGFvQi0t/zjeYvDZ2LM5op0SxooErJkVeyX7KfUjb1/qtBchOuu8Bl1D/msS
xns5yzgEJCsQ7l2MahpjuioG2GduCkh8xb+HBtPWliGvaAAVC5WKVXdzeugr2nU3
YE2ne1hID4mSD8xbVhHZTB74wcUsGByUE6KAtkzWB44vJ7eyPSYqMRYtg0TF47ja
iso9adNuneEf57rSgkuOVfsofcQ6WMgr/dJqVTx3h4IBzJEWW8SE8871FE9d/Dyk
O42ANk76GjrKV7P/AXZbEhDt1DpKFrgq4/gSAcPWBbFzRikjWHsSYlDeX94nZMvj
jRu/urGvyjcUjbEkSDVcQvVfVqzKWVd9IbJUJMXGNrCHQRE5ImqxtWDyu3UKEOsU
hiSL0JmykKMqgPsATEWkujN9qN3cA54qlhjENtmDL7C33AQrnpbT88bT61HDc1ue
b3ed+UleasQUFtnJWNb2yDJCWNGZFuvjAJZlN5QpMv0qx7Ddv8xhOHFoVc21lJCu
yu87ueoYTaPv55kLl8IRGT8OiFwy7VPY3nUqRPLVNudl4yKeF1FDRL0IIkHGfjN4
LapPfeizswl7NCefIdGA4QOuIdR1ZW7UE6T53QCJ0ULBhHATiHs1Hhtg/gv+ypsp
rHC8hmrBKQiAh2sZkjkxoWOPs7d5TI2JKbBNWsVVkfqYL7lhRbXrcvwv/NpC5h/W
ZUu/DLa8gozeuC0A4XRMHzSGeLo3DzkWS+zbMeQpz1wUI/Lcrz273M2adSvVXHWl
Udd9RLUliehU9Wf7/gLOS3farRa67mNW4fvDTpdRQB+cKbk8s8gEzRGj3qASm4v0
DZuzUNrHvldFNuG8IuiraDuEskcCmDTRULz+T+zF3pE7gES45JWeLbekLQDvOppa
ut2oVNJsRsCj5R9YDYEHDS8MRb2iOodKJ9ty9uOfWjpVcjUFkh1X9XfsFrQsmZeq
uZ5SkDhtwo6ENs85WuQlncWGxHmH9Vlqy+7JXtWQLNoorbw50dcXke1tNMVKZ2m5
ti6cOfOBue86ZAKjGboDFI/xqhBkDLdYR2l2UKrcErrYl6LTZvtzW1msPScy9CF9
Mk07Gg3k7ELxkNxhHNenYjSwFdX1POm2JKOQ5F6DTYviIQ3SAH8VegkAJgJh/nep
T6jd09fsEj/fmM2HTY/8xzLf+ReFpYMcKanI4tFmoMUsckignt5IcJONHNFhZDZw
i3qmr96JQU9dolySEKI6S/EeoZoW/MYV2uzccd645Wag7k3rW2Eeekv//oot2lou
76sWWcRqp2gvP1MuRWpxpZasRbJlOQdlPo/vXFI6lwgshPCRjhhLeO93cM0lkmoR
dR2VZiftPwjaztCICowYs0F1lV7WLtZbtM4aval2b3EA7ZWyxs2r6SKl4w6GvRhR
WSVcEewvR5YcNnn1w+XXa/3Hzxi6YwDiO2Hbv9+76b7tx3qIw2BtRIg2+btQKnzT
XnbPJA7I0Z2Nlm/UclijE4IWanE73ZE7IcX/S2a1lFeRE7nuLuzBuAzSViDx/7v/
9KQb0YAMPOesMlrA5RR/6z7jYrhnszbP+zjyn8UbU3l5fx1Gnca+VCGKqOvdlcFL
+DO0bwmH8f55JrrqrO8AES/fB1GlJR9XhN+94pb9on+AGiXWqo1X31O+suAq/d/U
m4p3B1R64PDH0/oRS5UTSxuS68hQ+QvDSUPyJWoJh70Q7m/zONwoB//oCraZ8028
TLnaoy8ZH/InewSLnDwTVrnNNkniCszq0pb6//QMzsEVtDdBxClbMb9ZEsRIWE4s
ZAU1Hriraei9e8gWNpphChGV5uF3x/GIkVbFyqgNNT3+K62MyvkidVATAuTJKRPQ
VfeQIisK9s2CK31gXv3zhrpMPTeGYrIGSmbDheIUgJ8OH7ds8+09FMZBftgueana
A/jtiJuaDl7JdoJ4kH+gKQhgyoZnF5mMYxlLaBN1z7ZO2lvJolxCDMfXnmPPNnTk
aoAwXx9a7jwpdDiW/wtCyuVWuDJiCgrdY3bd7zQXvkoQWqo9zWrUmvtLvVl12eje
EcBHz4f6T3jza3LrdI4IEzgW6R2awHnZ1FJD6dKGd3pM7EDBDfaFITo5cwHpdHBi
IZlB8M7y/m67c6PkuJSbGvFEgDLJjkC7n/Kuzsx2WJO/QWmTDwpPabG+qr8pEzwB
5wVRPU2tv/towOvInLGvVG+rYNcoUXvvolUewtEfMLKBqE9n8+D2YD//s/NM8luu
1AHFKPGDFT3II1Cu3gJwkwbuCoMGIh5g2zVB+J1aKRblCc/wxjixxNiGs/Lc3bfa
jrDrFnxtROoKwH+yfnG+Ph4CVuTwDrnig4U6wZPIKmLWgx+R7NyEQXjCDBgEdzu5
fuCxohmJWjZlddTKfSvvZaTlllNhdp/XSJyOg1mid43A+Mqxs5kuUmBnAHt76v42
xTGDGeDNd+xaBzaT/Uttr63mWEebbgBTReBUuEKTAedChb+YIiyt9CVY69GiqMdQ
OrVJsUvLYFi+/BWFDTyKr1tnnEf/7X14dHseYKz54tU0sT2PojUziHV4zY2Hbqmj
75NLlvtcRWjKbOnGMMZB98BqWQkjJmbiUaOnDidw1raOEtPScvU2YnJszG1+CH/5
/SROebP13Z/lur+G9d5UUIMpVwATm5E3ZwBhF+xR7iKuF0K6rUi6OF35EoV34ZBZ
nQorAz8Vnand9UMbq0aI/4MKzFpuoyRF9rFuka05+Nd/EtATTIcLfgZHxBMhKWvC
E982LNej769aGa8C55ju+HD4sScPmTw+weoQN+LvUUtZjgapyrNBEbzu1gMvPJ+7
6qWaGFcObQIGvxb2eLdaGo/hhEzj1fRpIfvq0fxrX7Hs1d89/ck2fyj0C2jkqePX
4GYtTj03kFwqo60oEB21cqgwEzGie5JY7rUb5yQyC+4TZnjYPkvuTGtPKX4CCsdr
XFGJJWVS6AzOLWYu6QrJT4oQ7sQB/hXjJA97ceJuVLNf2dFvYUGh+Lw6gj3UNuIy
wVDIu017W8fkuGXPKkqdThXVvmC9wwdDuAMMloaNCVYmOp15enZyzVLcAYcFVphD
1AzrAxQaxsSTPwnBsJX6EYc/Bj8Nww40AgkakKWWcDX/SIIvA/79PRymh0tzr48X
XfTJNeMoP5B7iGXsVBu2R+JH2CNsJVFvuF1DAxJM69fqNB3KbQYp2XWZunaoruRa
F7YQwiq6vzqrJREAXYfUgscZj+8nTIHmIDYLit+JigTlZzYU9LQGh3rglY7Nf8TO
uq/74Glv92HTV4hdA/ixKy0K7r27EtBU17VfJ5E6COK+Slwhnqzq2LSUUP4B9U27
ZZXEf3gFz0ZmRhoXWogTImPHVqOcSwII8JtDJTc2Mkx4MGarTDJBmiBfMNKSc/mT
SOCA9qiq9PV00jeidmPuzkge0gLUQvj15Mfa90zBY32s6Al4oJ31zHPiy3TkGBJA
DoRWUGTsk8vRsmdEOnmrJRvL//cFdmEsDjDIGTUpyuKybSVUBosBshg2qMbPmMNA
3KnQClFQDAXdSN59RVpISFjRrp7PHTbKRtgwFB5v35TCbX/O4wfH8Ly6//4OlogN
3JrvdiF0ZZxej22MLURYZWx/Qzfzkl3YJyNKwcxK3xKHSPbZKWjnkf01FUeOG1Sj
Q/aeHLr69B9MfZpQSTf9vV91re6DdxkMuXYjkZSv1mg3vuAq402dUFq1qUSy2ziu
d9+oMx7oYxdcgDBI95Xlee69dmn+7OPGp6moKJmbB118o9ydqdwneajQURs5dKmh
NR9jPSaAZuAedR3YDQMltQLVkUUH9hCvuvvhP4MCX0PqiScKESQ9pA7ZakYnCkkb
t7xPYxhT8ZU19/rWDNjiPmZ8WGGUSYhfD8jeqOia2hDAHsNQab5zkqUHvGwZzpQb
Ssr5GXC2YofDBPjScEZD9CNh7D80Tq5EH3d0dyUL3ZuxSn7Z+xRSKJQqVb4mUIDF
ziphrPfxuqiBAi7dxZutmetTmEK6SviOt9r/t+czlejDYH/SwgtKtaWh+iDFAXUE
v9BhU5AfeHK+Y8GA/Znt5KBRKLYO2Ps+UBB3kLM4AivD/Us9V9q5meVaWxJcGUsn
wreR+9CZMiV113nA3yXH2qNs+kx2RV9MZaYmkeXv8EUpdXPYIIjuGAXYoujg/uZB
n2cxy8AU/P9j1mSSjl39vio8atxoRcadBz0quJhlM1QvrPsRhfv+KPXCUW12ssRw
sWwO51qDmoiLyQTd2fOZfM89IZE5ANZkhjkh0noSmk73L3US4PuYemla4uwIaHVS
Vu7MY4EbIVz+VIv46se9vJUR8Z8bFwqZCQv9ok67AgyCNq0xA1YW+r97VSid9Ldv
HAZbEZpYhKuN2vpK+b4f7I80WMY/S+j4F7WujfzhCtlsVLofwroJsmbhbnWVbT+3
33g6p0aEcQUk/LzS1Lpcca1cWQyHOPj43HmBKRI4vUXgUwnXRf+P64laZ9CwTE9S
OcIzW+gWNA6CjrHldTFr1hUO8BQMLiLolY34DLtMkbuSXoQEW+hXh/u+zuZwURVO
AkJzXKQTP8xySr2jIOlgsxIiyUPHK5jpLi+Os2ZEW1vU1xPXjE8D8VUB14FjoFzc
fRczhtfn0RQ01uueeRHjsCp8EaygWgUBDzm3M0EWPqR+CHV2PBKUHKK4HQUQHaLb
Gp702x3YMMObxjTz5v9oLRE4G20jstlahYx+4hLC3gOjLN9jvIvgl/VJT3eW0hpp
/INS2O8aRBWHCtn+v2TjEYpgVXsldCfzfoh2wBFAucY6nlk4rJAspbVyMZ/xpdN3
Bh2ugGd3h9vu/MSGoXd04jFl2iIhl1VHNteniv07SHQQIb3W8QQLYVgJvLTOt73w
pjMVfvyogs+OMfqD5crPIe3U7xSTsr2EliVyYEMZmlyuEI6+Oi5wKDLfskxGrWKv
uH+BbAHVPd0t9AXCE3AHix/IB+DmQAiaHabSp37+vTKRQTWjhNrrZ/lvYwPbSypr
XngJXibIXjzE0xGi2deze0TgyksP2S5/Tm//7W2U0z0z2E5Zm9iOXEgscsxjM0lD
iLfBL+TvjosupsIXvelIWqWm9Qvtd4ply7HV419kc74xlyWF/9X0z6YBXdN3+BNm
tGOCzMjTPOUeIZEzKrSTxA4Us4yftsUDU/9QZIH9gGEHt606qjOWlgJpl9vPYQKC
XjP25bbuZ82qsBDe92oZ5s1O1I0T2KXsjkvGrsxle76td53aZ7xxBJ/7rxQVhRcV
JLIwAOeGYtuDFEonfcfyAoZ6CSHUvL65W7CaRrxLhY0VtgaWSH/gEIQzXPnC2Rk2
ELHR+d87AbKng4AbZw3zioppJKXC3Ph1PQTSL00ER20xkyb2Qj8SP8eqNu/TvAxr
ykymMsb0OL94u/TvUntTIO8IZWZd7Cu2d9zJ/ulTdt8BYsR7KozVrTsG73h82oaY
HaDJUb+yBWHT1s8O4TVY3wmFFh+zN2eekzRs5LM6piooCE+QzhG5vKUUUdDvIa3R
ViuRRdARSwB69VuBBP4khcPoKYFg4VTDlzxmn2FoLxG+hkD/FHiBTLcqLApA9OGy
1q0fV5+f+YiUAMC1oh3dizW9RhEZ62rpCfjy8VOtwpG0rYjWeZXm+3F4LlJuOC+x
ZphH8RTY9aFjrNQOIyEehakQY1ih5MZ2MJSnTcR1n0QIq4e0qjLR3w82nAq108j8
TS3+k23vRZ74oEbIC1B8s+AQx9qnLHbNrLmuaqJCcZOPo0wxg19hvfItzdvWyydv
vzBZQ6kIYTFBZo9SMwDPdg==
`pragma protect end_protected
