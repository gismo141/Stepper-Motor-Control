// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
S5GTyUsbj52pICtvHH1i1dEog5ucOsBgc7rK7fkVIQSo4F/Di8pAF0FKxSho9PgAD8KyMOz3z8Et
yab+TMSdxijjVheNun3+8ERkahvZCOb13MGtJ0nSWYaDdT12mRkyH8i7Eq6TrU+Bi+uEMrAx76cH
fplPpQzX+o4EgJxciGvEUFCP8PwAIZ9Hy7hJCzWS2ue9QHbfWMR8sEWZLJmvqI3wjtn1j3ScQtRZ
qsiIH8PdlUcTcoF7IoXQtkL3rWAZ8CIZZ9h4hlJqBDlFq+fVc+bIWR1FWS4mGFcOnlq4qVGwTGpO
mlQM/cG+jM7Z8RVP2fk1OVc7bFXhk8U1s1pfaQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
HNnDkKsRNl3IWW+PdtxAFGBmrfwCkzG9Cwg8QQ+fUb66Yt7q9c8NEco5WiVYVejDlOKg/cZdkFct
JSnBydRxiAH9OUXeCQhvAnyokPiuYIQjLasx6lA8X2MB6iaND69ZCxuwUSlmOgsOv/SqqQJgvog1
tFVQP0h7Una1HpOwGalkcsqUU9rBOxW9zApT+B2p3Xaa08G/cSpGpPGuuWMW80L/hvuDPwjxxUqw
6IEUtctUoWc8whdgzYFZBq2beyriTV16ftl1LKw74XDl+pIBRF5uX8qQmXNNjvWhAAOL1QiqKAqv
SjhavmNJI5c3Ukxhy6Ai9tnWM1NxTxYxJi6uSrffKwKHPRtVTTaq0C57EWnXhFRuRaCGpFY5lZ05
bUJkP+vlX0rmbuLwp14cP5o2DIn9+htlf3/eu/5haVHvrL3PUqNsB6iIGP6U+/jxhvTvPcPaWTpC
jlIl8bah0aNGll5ZHn8KyfzDvdAm3D1lMr/t2qWdbSTUdrIBzkXyjJLRNEuuUaoeyeKG7Ax7XArb
RG7FsOGnxl5yO8pFh9UKLLDPINuov9Or6JBzmjeN4VrTC67WdJcDGDQCnkfyZokuRzZCdyc2/YfB
EpP2+I5MDRAJgjDDTGROHH0LeUbNbMi3gp0I4wgUkVhRJmlt+uOex0gtSF+ZAIYXcZdz1b2C87vC
vVoFXsdG3rZkdJ7wIKMBIr8z+HMAeP5bR5G7V2kLQdPGvsV171Rh3m08pUzlYcXFkvZ7EP8pu+dU
Z82kYOCq1rdwPPqkb+jFISy0Q/m5Hgmzny16k6UcE1H6mgZjDH90vCVCnB4d6+0G/2U0nVXzIiTh
8KNkO+q8Laz16qd+/0QS6wQ5Oh7oxrQ6sGrHgR9p/g0+Wrez6Hvk2HETtykRoNretk6mtzpNgvxL
Yicb1IfqMh6y85pTbzg2wyKN1S12daKcqYBL9G3SOhLdAWAeTbkFn/K9K7pzEQVXhSCTMXRAR9pI
HTmMBD6N/82Ry5YHV3iflXnWizdiXejwhNXHjX+aaMDVxxn9C0JCRoSSkUdBDIhQsCRg2mru2t4F
iC/Z90uz1JolruYP7GyLOQ4BOGDIVvHWyhedz8RBhxJzy7XwI9JVwEFHOPRQs42ZiSa2uM5tWjmK
DrND+R/pZVGB7j2DB5zYpncIPB+hak0f4FLAVDD4zG80xeUGEDjAqCscTWJysJmh49kwMszBxpPe
iSfusd9C08MBNbcn0YyrsWLugn2F2tu7B+QkX/NxR51iovoQkj24sVuP0ovw2suvaxhRyPzxnUp3
DrIcghXgQ5rQ7xUWflxUNCAKWq10sDEOgYhEl5g2t4CDK4ou4e8pnxbikneSW4HGK+qQZD7QM/Mk
FsCKOmsKN6ewMRS4JLn54U/nMCMLgjhQJoRNPuGqdGRecSiyxwjNTAGnuQ9xmHPEn+kTKh0uvOvb
IgJYfMMwKbYDg7Hdxe73ySLKn/KwBBo2TcOr0owdWdElbmp34rwB0ez6cAq1zr8BJ6pFaPv59KfE
WUhUdNASsA/PnDfqRyf055lfBoeke5scfnhi9No4O7DPBr+q+QHikjAIQ5FRKZPwrtWxqb3UGthc
pIoPfnIXfajfIUh5bJ99RSuEsWR1BzrfHGg7hD64sZmPxAwYIcyY09bQdcxVsR9459lGG4ITu9+t
KHX97Y7b+eZH57D3YqZjNlLD/Ach8rshWgjx9rd2JtmAwHgm2x8Kj1Teu1BNO/Km4tnDq/MPCAUu
TWumu8nXCvRlKznrmohJUwoVGb1wTSmVALoN57g3FCgSDaoJf5ri9llUUJZSZeyUc/Ih38JUVkWv
IsBfRI9a7MY4XfEFJo6dv8hlreEKJSwTrZO2bQoKNX6gJdR1lWWudxJwF8W5dvu9Bnnv7gsNcm/F
8Mj9/uq0RGs5reKuoEa9/5eKS+tXMvSJ1K1GBei/WbnPIIuvfoRYnScR40ynLQAswM1+1Iq7Y4qo
RESNRPznP8ns030vIU2NzIOZneYkdPCqGanYg4qtSE0+Z4/9ytA5RwyZuc5syhW4AGCx+GCH6Idw
TDaTim0Zj2+5fSO5kzdMFXE3JZtvbm+C39nqKs3tmxNSZcrANvrM6rTJ5ok32DRdoe5pnJ1BWPvp
sdyhpjEm4KXWPTt+VN3Jf1IXPxM+debswRAMZp+kZaSW3W31qwL5G+S3R+LEZyTTvEVej4zIMTHi
hazNlfQIs6WjFw13jasi4+we2xa15E2PiWAwwAXqAGwZPccfujLE6RSnjTReDGzdOw00yeU3yubr
q+MMk2hdd1rJfiENJSC8/PJjC1wCSfyiBFtXM/z3YN253tlNgabmdBAoWa500w+Zh9GKZWKnRHbQ
UObliQ5IR6peJ5CbC6ArRqDtXYGFrB3gNHfIB9S3g5AwMVfNm2Pe4KicMxW+6VM6RUNndph95lly
DtbkyGwlwil/qgL9DfoWI5OeoI4D2mNSYmNK7u7a2a5u0/TWfHU9cnun4OknbL0vw9vZ2U/9jCy8
KsAKmvKeBFBbmzd7uIvE4lrJHFWGLK+wK0m1HE9xp1xOvN0WWtmm7VDlq6CtaSteYtKc6Tm1yimm
ZjSkZ8TotEbts4cQ9NNSUs7xyvkpsqxy2yndig9wfIVTzNekfm9GSCFTO5N0/OmWn8ypB9VHY7pq
nlLXAyyIs68hjTBaTjT70CVeVjDGMdin0NyiByrqPRxN8SwcTHDTOETu7JNo3RXfR9B3/GbAxhaW
oo7bGJQkndASVHfbkKkCGJ9UXkPQAIq96lR5T06/B3TZIwoszfk3gReoFAyV/6dtC2mudGTZgQJE
Dyijf6DnkpZBeUAQMlcb3qTm1Ot4sAq2VoLwl9YDBaWpbncCFDgpqOewz7tBraRUTnvSrrpyV5l1
cwm3rJeJXSFQJshRHaM3dc5kYWA+X2xcKfVui4IH1rPm3wo1/tjd60YM0dJjcxzl1YuVEJTPv2qi
cJMfUW1uF5LeuBEUpicmVZzoXQqI1lrXO/Kn+hDNxDgf1O4nOMH1TU5p31hNiDGKHY/C/t31JoNi
sSpjITb2PA+9WV6GeIW8f8/qaHsfxb0BYQ6gh6yiqa0Zm0oTPPwmLEPAr49KfsOA+hbWvd5mzlCw
3HrZ4AGaqh89CCa7LR4KMR5aRkLR9Yue3gXAn/gl2zaiFOU6g/AE1yFjTPcLLZfzLJbdiZu0OQNT
GuOCviARt9aSH/vXfVjgBJ6u4fqk09iciohug/tHC/20Ms89J5WU062sX/MR9sVV7iw1qld/IcUb
GreJIkrl3IN7YkSpLMDELKSGXyBvrjrYqevclY5R2FAVUm9suEFO/QXN2uuaxx8l5vhBLIaus2uV
1a+aBiAV06R/cIV+r737eiBzvwOvP9OKjXTO2lb5gsZ1Jwn//M8pFramjVRu/fsn1zMAlr3s2fF4
Wz+jCSVhe/FNOXcuTdqd3hN+lUB8gYyOvvV7fh2oco5u/azBi4oBUmYLeDcSojefIDvUN/fxjX6/
T/tHxZNh0I3qfAPysV2vVpwHz/ur2yOcMASmg9pFHhLJyjAbCVTbgzfszFzfXKLTEFjvYzkcX6c7
/g/3chLJDT7zx7xLXVhc9ZRQs3ld1VIjieXOZPeV9a40J0SYLa5EkPwxOS0htSUUp5ZHEYztcy7R
EEZtQjUdgKF1JptJk1o0ikV4BHUIPMPIerTJn6hP2b3/92TzsGtPXn1VhAzzf68eu7FkyVDSeID6
QFR4C0m7KmoevYS4lOnZU2LMuRAgxufbfCLVujJKeP7r31EH0LhhEhrAVyBhlTS7aM+CvH+Y6FCW
5n+fqgFsbOkGrPzN5S+dsub+/GXnuMVMmTEz2pm/antqMvMn3VJu6nPp5fF3gJzOKq+78hpbnhTJ
84K99LDOaDy198viqhCoWLgvioDXmFjjRB9Isy4vZz5tV8cFlt9uLWG6Fphc506SwHrDuwdwU8eK
iu95hE1jb2kEcaMifbDmH+f+7XWwsDGW3RoBE+M5vvtmtt8xqJALjuSJ+gSsZKuTcAgI33XkPT2c
1yd/idLsLAaFzvyjwZ6Zm/W4pmzxFYkWgJMxSP6eJS7Y58bwBr1nXf/IugWGRO8SaB5c2suHGkIO
vPyvVz5nexnyIMqJT9GB5555XO9h2pqJC74L0UncUPwTaCmATgzWs8l/3T/UDxoU2uMcVVZ2Tb/Q
25wVUfEZoOEP8m7+lfi6m15hyfXn1LlwqoGj23gOGPJQxfK3aRjjPekb3SEU6BsD7M1ZpisySw25
4NvyQr7+V8lobpUgHDjWlRPaZyAxGhWX/lkDxWjnOv/VpOjh+0yTLVXhCxYJakX2mKW90Xa73zTt
fIQEMSOQNDoLuL49OrBH+MSKtYRTCBLjBh5YdUA/wZVD+NRy7h6cNFPC5mfO5yqwgv3vHbFcxD7n
rI8y/HHiSNtMN2PKPUbLibJim/3A5pN4BhjH0X9RPZ4QdYqBTVVp/TKM2Pc88/zsszzAQCZewIm7
hSUUh1NyfDQSaic37jHmXkHYIzy9P+CeNtgSusdI/F6u75c/dHAJE1SKr8IT8L+46E/EAsdjCG6F
gfKoKvZf5iYuTQuoND9+yWZoK8HJEm9UJimftPpUMXfDUojnMMuLu1o3uddCTzeLfTgGQmUZzVHD
v4PzBDc44G60JujmnW4RsxQoLyWp+eCdcgZQhm1H50+ZKu36yIS5P1nbva7hjriTZgSLCbZ3d3nL
QzkfSJXlzHvyC+xzNjlFBgkMl42JKBIEax6cwZMCSLIRbGpyFTQJgAQE7OGLtapO++NqgTJZ0xDb
AUxdHivl2VjeLUupe7aS/kUTNIFW4mxEJ6QYETXytpW0KIufHPE6G2MVKrbqkSQVu6qoVS8rgspr
3zfK2hOSJhUwfQeweA8UcWYNLby3PQy8VwW4nVLxC6iBYz1/RloF5cGP5n5TuFZDw+sFea37G6am
6aZZB0ZA8SgBhfAWSE3lIoO+DuJ6rxNsPQJT4fp9Bn6GwnViOyMqYL8UwFaleS07gRiJSe7GSa3A
TJsiPsp2SU15uqdzjnzzWX7RboZ8lJ3+6X/yb5Hf8y+mnq90xMyM5bP1sdHZTO5UNfI8pzbDm9dZ
WacGfEPi4mcKwJ+oAVu7ZyI5yy/7/zKUBtfQ5DSLd2CgsHtuygHrimekOB6J/OfFvSJGFCb9OxJ6
W6v1LPESKUvyAuv4aExNw50kNL7xdSnVoYkklBSMJ1z+LJTuJqJROp5orlM63tlCC+1pSagDZH/6
wJSC6Sd7LHJfdN/70gsiEDFFhspi229DPAnizNrU5H8WoyHomhmhkx0z91Pmofjs1a91eV0GNoXR
rRBq1J2iiRit73fi63RChcA5DGXWuEGwcach7/PtpcYBvAujJzrmQg70tS2FfJZn5NfMYBO754BF
xH6obsTowdXy7iNc5P1yQF4HU0B/pZKDOVErFFhF90mnd3383ymiUwRNwTVhIUj+QSzs8B8xCIVy
VXsnONczaX+xTHHxqMjfXEfaj/F/Uvna4Juye/N4hHU+G7JbzpHLqCjJsbBMLPTTqVqpypmS7IyD
ogXX86VsH5MNKbuNZS2YOoeBJedV0qUwbjucspe/hxctREA+66Hm5HybuGMuW++0I+xFZ5gtHGTB
Ez1GSSXCwEz+CC/xUxFQJjI5IyzlOPqZrGF5A49NrXSCYMMUKhnSvOI0N6wUiDShyw3Od667cYua
RLz1jCYnhCQRRSWbptpw3jsSjQKrdIoiCp+5mH32fkMssuNbAM8LR3dGoATMtIa5xpOxHsa7hFVj
Q/vp400V3z/cGT05drahHRZfd9roMMd5hrFMKs89mQjg9b5uw1oBna7htJvALuBU9BXNXhupqJuL
Fzo1fxooYkYuPowoIlKgwODMmzJwGNV1p0cW1x2XjLUGMuiGrfCJrPooqNJLsrKSoHpst40wzk4I
VJDTYDDJ+cJ4t2vsb+D/OVWPci7mT/9Z8wN2Mam7d+uKffZo5kpRAn1F+yoHrvJqc3ADca+xTZo0
HQUttSzVS/ZnXvK//9zOStA+63tzZGE1/tqSjiwpfAc9QG0ADB+xuEl870RSgy8ugD/YtdQ1oBU7
C0yNkWRMIQu/sy8mBmd0hfz3TPEVWUbFznl+XbnvQnGCzgt1w8auAKHLXzwl6FPwnnrrJ94OJSoO
q8Xt4ZBqNsNfMDJgF8GJiiOwcm+IYEmCqaKSK/0h+m2sW9WX+trl1SotYArf8m2rroCqdgu2DQrP
LoaepqhPeNTfU+Xm/qKLaXDH5gD3DM6+ziYuKuC3at0YtQ8Kadk/TFWJv68GGl3Ljp/91uth8t1/
itmQEwuRbmqcQVzRzTJggu6KmKL6ExGeb1MzGFq/1GIhRlRkZa2OZQUbamQwtR+kgE8QaeXWALJl
47OFnODh2S9oMrLtMfd3wWCu2v/ftfhMoMn9k+G8buDe/ab9+skDhHeDQwbciDVBQ01tSgEhpGuf
hYwZFufJOSfGrqpbHtN6WAQgDvpmFWbmlfQLOdUAWSXOYL1O8sErxAAb0kI/BQnyjrN7kirSqWBJ
K1tCTtvk1n5ZBugh67B5ybVDQZ03TNZvAd38RbxkPbkbicxD2zbN7cc3s7+WxrOIkNNgrfUNdgxe
/bgiM6+mkVWI/UX8PfJOYK4tKk4JcaWn7f5/thmDSHENVNlKE1PP6WZZl/Vp5zX5iQQz7yRtx1Mq
ru+TzegB3MYhFGRotFjVnZAQazCVG0UuXTLQbjuThQVFZcMGvAIJcX/4nuahCwOvXtxuOlvUdtee
XSqHg8rwrniTwLwh27hYw1EDl0BRrh1bivNcLgow4YWSFFRPWoGQ3FKX/H/1SNXi6ne5J5LYd03v
EN41wxMPq+/rWWwaVnvJH7Yb9gRKeix/bYN2ejhCthHRvknHyKXAC4mb3KxEY3e/eJQI1jVJdhng
IpzSvsr7jyVM9KVv2oigoH56u0tT+imSzr/1hUJ2HOQmciDVzH60duwMLwybhus3X5anE3s3/xO6
cq/7VtIu3GkKK9N/BcnO7cEH8wpFcjvfGcMJDExh9XMNbYwh8+jhDxTYvyg8f0bYy10w8usjzvKO
HcYDt54y8KRLfD9KBnbVklTNyVILEdI78CsuTPXKhmEnPDcKxXEZVjlcHmVENX9ITobCMA/C2khZ
ETBROwoaGGAm934HVaXT5o5uxSthxj9W/1wpskwTXLz0w8SseThr2fNgZ8AVyFmi/Jaugqrrxgjg
iDjKHVXHIgULeNTaX3z7fegMVh/UNEfo4Ft5P3mQIwfwhOkEnSTtPcRHWpmVpPl0bSl/PQ3IPIk4
CApjyfO9L9Ha6JrqLfhdbVxlqbhUR8qRHlLyI32Sp+C3AjdJeR5+8V0OwfOZSZWVXd610npC3+Kq
rQpiR6yof8UeaAGCFXgtv7dhxcKuAdNHR/YrwdYL/zIjmdzyydj9rgpHvjzaSDW3iP0B/kCUcRBD
BWUgohxmZS36vo6YdNj1+FeSWzeSvsMHVfJI6GdTYqxldqbttKFtCaZQwbEAPUgEHRZDqc0OFv6a
wcCxNTP7Lhvf0M0ncxcqjJTGfTcMaauF+VbbK9IVqetZ/Dx2ihR6oETfwWAUfPNnGFhWKj5KALWF
6kF3P2nuWdoaV7aFxSekcOczo+VabttXrI4s0sUTx0YMNZ6mWrdowSpsmNnd0YsI08SBrw6NDsrz
72C9kCNLrzzlBg5j3itxvc2XqeDke8XpBgkcmYd1N0uknnArtCYBuToTpsR3GLIG5DiKufTS3SJ8
mw7Tf33UOWg9p/XBPoVXmCGbNDDoLx3AUkJFf7eSxE34/gRbt5t69REXIHdksRVNnJtKWES36TDS
AVYbU7jiTguJulI0GGOiSasFoxDLIzTTaL6kXFU9t6KIMjRyvkmv/RQpN43BaBTx7uDvNChnoDRH
Z/+Ods6d1eQy029a2lHBPp/QYh7FYSby1x5/nADAyEO7G0xiylQ87inr9E5kfm71SbSrcsfenEh7
siXTfAbsm8eXUTZJ9JfGCyfOUn86P4UtU2CTV/boOBvDI/5hQ84Y1bgpHvnX8ERtDQv0HpfqHe7P
lcyvFFbb8hXN2MSuNsvJxYDueRfafmKpuGmlBHtnpDq+Xu2ElMwxsg6hXbz5AwlnnwTGZ3YSwHWJ
/p8ippbrdOsHe73wQnXz/rURAftVUwJANaUay4cYhawiM219fBpwjPQxktr/m/3pDP6gWYcqaHh4
fxdaZ3fkKPZ7YK7FDturIXu7JLFgapk4PH10Z2HlTKCRS4v3xDvWvuSt4UIrsZRe5lTlX32eRwDG
egjG1hFlD+vm6ObFQxStNpBjPVTz1U3E91GwJajqEEsbH9OfUZV/kkwaDlmLUoHqSN2knqnEgFZU
7tUApp8jkXlqTBehVFY60vUi7wENZwYZbyHuHVeHv1m4G2HF+u/fMDQtj0DKUE7w6IssfJu99eyQ
BiqWe1v/+nkSeKT4THk2TeJ5Ik4YCcn+8pSz9qI4jlzBfuw/R8hIKEw+ZOfTI3tKcYHHt75nFRCp
B1RAScOePzRngf1sZLtPH2fTKGa00M4gbFrKSbEzRlZjcixzQUelMRCsG3XT1tcRBkYGS9N2kVyv
UvG0OGun0rNTBHaCFrafBMxHlXpvDLVz4yiodOmvN8iEP4xA2Ib/COANg5oYaCErCuiXfKYGWihQ
3doHWaC+bv4dzR0vjd6dxmmKPT8xxO8/fa0rjMlCPcAVgjDdDFICjFzQdS9L4dFUKf8tkD51f7qD
MlMKx4gBGQpH4G42rYX40fanAu1ku8qr3qN6tLV9+Z0yuePEw0NLEAFF2Us5G+0sOE3p2d3s4gkB
Wj7Xy6v5rh2sdu0oidAXpJ5+EkmSh6IYlMqHSgghaDLGUnjWFrq6PcJskE4CPx0ia4YcQlZ35D+S
V3bdlbOuKFgewTIB22fAmkKu2TP/t3m4UKlbttkie9NWr8X5rrkmBPp+7fSWm1Q6JnW0DpMPs4dt
c/qGzu/2BeSsEGbcTve7gO3TvPS9CSUI1KoLH0CHKTZZql0tuN3wRdS8lCU1Yguvq4ajQtUTaoa6
Uj+TCHO4ul97d0P3044BU2wKRVekE2oE9lZVQprVGAg5uIgJXGyJORC63zPwhI5+QZnjn3UB9FUd
UXM5bhWmbqzM1ojMf7XcNt2Ry+8kfBdQu5vf0fDAuN2eRI5YShrGYf8cZVziwcg2GF3jEDQVCWfN
7WrzmL46SEGMQTWvEg9WEIk6rIQ+EzW+Bq4+ADMTEfUpnx4/ntAQN3VIzCAPHLGfb2byzFcnKLSU
L3vhftKF95UAN9VJqzn9jB+xfVkXSPatsy5ASoqXvC4MixWDJ7fWtJ0P5C0G+tn0QgIQwHEWcJlV
lWpZDVEb2yf5611gRT3FJgapW7eAnCRQxWl1YHM3Q9xo229l6AfysEkqg5VsCI8c/7HkIq5Ujm8f
Nbv9qfLu2Fknld+h655G4uKbC/tp/5qHG7pUs3ea5NlVTBhu0Lg0nZ8kme1tDZX9X8e9UuV1BUOV
Jv+zQpnsSFW1Y/toxCeNnME3IdnPJnS8X4Fk8hLCBn4bweIg8Jr58VsANzfL60J/5u/OmPL8NyZo
fzHsVLXkxuICwPsX5xGDk7mkm2LQ5JCwTClhly2MGaxrr+7113qTFMH40EXFd3PUdf/FKSkjPcqJ
E5M2WIZpy+ieFZ7jkcOL+nOYBcaaAOEuVO1qOgdoyOcW9XezFseK159WhsMeEa6P3AbpUB560okl
MtHbDjEDWWpGhOgQ5u2Kxuy5wCl1urcQ5c30NF1liHJAy3n6hUuqRPod34K6mKXzHDEzd8RyqmQR
EkCX+ps23UZdO1jf2g6XweNsFhoC3xD1ogxSTJHDYNJLW5kPuRz3hyr6J9i7qh74i+4N+WvDTSy9
XsNHHt+AXjZQtldjjOQ1AOGIGM8A5TkZ8h+ilTlWU965JMTpp2VZmLFJCXo1GYEnUXm0Lwo/4RUk
mOACqJp9xR1qkYAhjRyb1LCgTLQ2nUBgODrBzwDjrkdbnIW+mB1YeIVFS9ON2wPg56ySJAYks4mM
FBlrvhSkz7lgGhcOpKPKnSjvGWqw8kZa1TTW7Y+/0Joo/NsNdJQ1fxn2HETzbl7k5BSoQQLIbqxB
DS+567UGbmEJifsGvKA3KuSWEUE5HU407p7bdNk3Y9N9w3/h7fx1UXp6LY9bjlp2nssNKXuvd5Pv
h49bzkwipISidwdngQcVIH3CsVRvSQaCnNepRFZjXyBc1noY3FmXlYIsTIlrFd+ejK2sbdPUXgK2
6mLXnU/YBQ0e8KAaF5W6eiiaS7IqcHaT+npmGmQ1SQMp+CIe/xTs07X2Z6bRUOAnhS9Nrq2sRiOX
Pm1P/B6Ti+NI5pqokpoHhg34EuU/oBjHBeevpSZd6b35Q0DecQduxqKaXzCGehcx08mpsyyT3A7E
4/aBsSOTFNzlczzxRnA9NI2A6aH4WQL1AZOxooQY6sWrC9xWZ/SH+ISeEMNjLuYyZRzwND7nSQk/
duFf5DqQYrFac3sMhmMKJ5mv7Ql/9sVWAse+hmb8ji9nm8D5iw56ef5hMeExVTmabsd10P9htJw3
WpQS4bCpedhYbrbGqlXBmgsmndCkQ4m1VxATsleVFaizf02BBV8WUwPowqhepy6/NGlgqfRsdUEO
H/U/91YzgGZ5jlT3wxtQjEEwuN2eCaT/qsSORd9BjMCiXBvMKZpFg8vMFuuoFzUGdJuuWDz09xBM
jD4ck/rOyf4rpCcTkgYuwEf0tFuPqAshGQXav0jYPKm0HDJbd6Nn8/cV2hF+83qWvTXueyEeuxNT
swP7iVSLCMyucosoFWftPxpc7SF5sKg/FpXzCcNtopSnrEqAA1qqNsuEX0uqNFavtOrLjhVpZARu
cfgJz3pz1CBgLHTz6oqEFyZZ6K4WJeS9jx+jYUicNCvRH0krLF0Upepwz5NkeT6gx6Ze6fErPSnD
7Q6gE0gdES3T5BBKRmlsHmhkkghCkNkr8u2JK5ATxy86UdxRDQQTBiv/YdyF9Bvfwgv2jjsEh3VY
R+FdEeNVAwK9JwbfE4s+keCm3oRuUwT6iBECTj81j21MlHfD0+sFxCxVHTZrKsiB8+PaU6nQjccv
bPk8PNcLfjlVL8KB4AXc//3LVR+EOyEkCdKfW3UmTcfc16ErfoWTyYpJ+qZabiGKsMtpgGoDL7K2
WHLyqXSqTHO8+lJw6hc//93Op2Qy2N2nyBctPH/i0X9cqGVeobEUKBcdR3YnKoiIG0AV80geRVYp
rD+6hGm+46iSUmbXVi4YmgXv9uvUN+Hc3ijnRIQWd2a1j9mKUqvQ5dF7WX/QDD01NOG1HQkF7SCi
25uRx3STGUkNlQewZjzlXCLcSJd8YHxkNrr58gLzEGNTI6uITrK5WrMeC2w2gDumG7hDlslw86wj
ZMHiCq53OUEtSHZ92hlQ5221B65ibeasEuMq8TyGV9EHIZ+Krd/YpuxFdLqtCiUGeZHKCc6jH02E
7zY4u0bTYLc+6uV1+0co4ufIgP1/VRcIngKPWP+Su5EFdn0j4bYzPz/XydZVbi2zrMgqYeSqVRpx
ObLTzATHFrBe+o/2OIjAOXrt98+oMf18Co5Rhvh08bmUjIgqicNZ9x6jLnRjZTpbkOddFdWPzteM
fIvEV8YYpmF/hv/R7DvlaQNxuCo/X5P0NQ8syn8u80vtsN6yYB8ogasTFvSqJwLONja/U+ogHLqT
j/2Rvg+4orDctGi3K8hc6dXLVYoKoJmVg27Bg3AD8nHTItfEFPJGkZ2t1pQa44QHqEXhpDzSZlLr
zbVRT9AQGdykpPcWJb+ulmWBAD06IXEzC5TsQZKaFPvL4jr7pvuz5nfBbsmkaq0WoPLmh+jG75y0
2LXLSnV1+tqlsrxM4EGGoWNJBu1RzADJFjveMPhQ4UF1S/3pMq0XyhQ62GS0h0WgP18XUetXy5Aj
PN33vOAP/eALoCvRUL6bwHym8cNxrQqgcuEyoJ/c6zCt03uyHrtOTXj+DEglcrHNOm8r+ryoepIG
mT4VXXEeub1ZnKBRarDMtD9AgC6kyx2B6+uqB3ciEHyzaw6yEOjsBbwW+APw8w/tH24XAN4dvOhU
v80ld0nkfaVGCX6FAypi101+f27jRsBUTWMCPtvonuzpmT5I0m3j/jSm0jT3hcHerKuKaZvF5opT
PzwGw+9oelIHUEM31mMquF7+1dha+OyK1VLETsC36gcqFHxN54DzjjxWx2Ikzt2tRm0Z20DUADMx
xuNlJ7HpTVPr1daVV+K7M8jthgJoVTNlrK/hMLNoIvZvbN60zs+is85/8Dolx9fsSSjU66E6QtvD
sguCh6WZVB+qzidqzE5ainiwgDPJAV/jSDOfPKaqG3brjXaMNlVKZXh4l3mYzAdT9ihYuF6gqbJX
vb6yWZw0f0hMcBWR/y6JE+cZvk5re10fqGB6U6kwIrZ1gEtVOr01MmDYoPLP42osuPI+wjJ/4Yog
r5NCqIx5JMo1XJRUNFob137qiu4k6DSlgBDXwUwJXBvfP6X3ga4muHmP4vXTKMiYX0dV4EoJOdJJ
xOqxgtADAHAlWb98WVxNXrpjUFc/yBVgRNpIVJSufSo82NI4BRCh2ZjTDP9KLVKP76bwM4Sw+k5B
ZNB3wXS9nfzaP3yRLLHO5JS28ouB/3+TLyHbEBuToD+wj7dQX9AzLjXgCvRh4BhUoDMgR/gTOmY2
jjMzQ4DhzqQxDCnsD+4hy9YfhFE5vOKbB5s1pw+NhWTPEaoFoWMoMi9Us07qoq6GFAOdlOJMEqL3
3Kgwlb3BV2uDrvcIOD7w+Jxypy9GLVmx1oZmH8F15/9opDnIwUMyCOuHKRBnMvXGqpTfJJY1n0xC
V1dOecbmXMebDKLhPi+0nHIiZnoioCwuQJgGrkllBnRUCKWY979bZeBdMfvi9dpBswcFnBFempHc
APkGTVhMLjv5C6eb2z8jrd0yiHyjMKkDllfXaYGYlEKY0VlawvaSGA50Zim8KNH+7vGJDWR83Wkg
htm80J0IicV1qcorcN4oRFPaePeT59puHaoXrUD5caNILzTQitJzooX8BCa+EIcrgZbJCgodn9qS
G60jCyKtgb5I2cUpZABITJQfOg9oaQUDBjtvC2hTIMEkuilCJMER8nbOT3HOMSM1DVXU8LSvWWUC
NfakYn0VEl+k6O2yhXZIU1rPiY0coZ52nNCVcHiOHq4sM+EbcZYwXPEnyPQvqVoXCOtHlHKZSkXt
YSUdK+p6z6UFZFJTg/Kz90jFqo3FMkIaLABPWiZpwhUkM48FLZACiOTz03tsQBq8oyZ7S6JvisTP
6ON0DwjBQQ5+pboWHTxjNdkHMWGveXx0wRAUgzJaZ9b4nW2Mw6kJ2jBuyAhiWpmcqqjdcb7tuWqp
9D54QmB98gnRNF27slYONH57Wlq7kv7NFCCgZ34xiDDgjgcI02bEs88V2QJWCpjmChW2g6wWAoqU
r4oH0fssi4iRGgqPZrw3xEVmSzbGDLaJX4HkVWZR2d8djUbHjdtkp1yqiG1fgjB9gqSblD/9lBfq
JClTD3WrhIYzW/DBg0d+gVwxF/LMpcGrfXmuTq3FMaTTiFigAs7fkZ1iwkcyyEpUA5yCVqGtHZfZ
HKGIAI7XO5cdAe6wW2YzuKIw7HmjzLy8snmGgfNV7qRor36Dx6PxiGmw9+/lj95TRvhGLVZM1jmQ
xwPz+mIY7vy4hdMTphu/YMDbCxKbboOryOelCjxgp3gujzYfpoKqXu7R49JHQ/J4EwG9CGlsALfn
swY3L31ID4lutF3yHi7DNdfzbkDFH0YAFQO9yqpB4ksQZgRrzln/7gKkOnlfXJvyNgdNS3HyPRKh
lWKSK/iHBZvtLbHXKnHiH2L3ax2IS56N+qw8glDzIMMklvpRwBekQkDwrx+98TNfDfZSQb8Ypekv
lDnFQjF4ukkZkugvOCqDsMR/rvRfB0IffJS/MwAhUEI8+RqXMZMiQWqqCHv9WZAsJ70LnFxh0XTP
gIxJLPIBUOKlCXO+673vHtq0k951ya07PPu58p7b+647SVjKkD/HJLUGnqh1PGpSg+IlqGQRXuky
bF/tmTsVGE2eFmjaYc8SBFo0Lo4bMUmVgrwwZ2VvBNA4+FibGPZ2ZLNIsQdM7Ymh1khDa8oh6IBr
YL4JnvzHf9JGojHQm1nOArCEvVEzHsEbgiRy80rnt50dXtqxPyNx3N6m3c3U7/ClDYQAOmtzv5Ao
NKFNLkBE1peBnw4qRvsDQ+jIBwYextpfsFA0c+EhiBOUcRZ7ntwMZq8wo9MvaG4B4AWpElz3ATHf
IDhU0gSHJXdsMLY96e4dNFa1VnbH4wsSqnKsWQHO3S1jbXQ0GhoV0sRINDdQRpbzLGJZPJ9mI8rg
qIsSSlQPkaSFbEguntmK6pYTpaoyHrkKneUJ3QQCY3dbL6bNjT7bAYlzhoKFmU/owCz3qUKNmwR0
fcZB6nYKweqMXA6sJo19bcFL/uZk+zcDtZ7ubtn97oxpTmd7UPb7Qx9YI3PKjq4rAXkUyLCA523p
CZner370y56BLKREWdo6JZ/lK9pfejoreAC2TsKytSpWqF+29FkBblSCon5RGyhjBdjaLv3kQWHq
cKPqRtYojb1YakQAbe4WZc/RX2Rn40+levW5cvY++cTZ8mt0eY2V0v7l7wK8jKO7QBvTFySk1Jdp
L+/2whOR1R3sJTxHdTU4MTqmz1A7i/MNtu0vLRTz/r7PKfXd9gUbsQU2C0hvic4/tI7iV+8/sJD1
4GLJZ9udqPOoF5cZSjnH4bH37qDz92LMSVCqy2PC/9H5V8YvDfa7SAdravgRn4niIfRJHKgAhfbR
EOSH9UELlp4tyw78TWLHXoe8qREN8V5TV1NUnCEWiR7IZMkq2rSeQ8wcJWypUI52Iksdq2nyzHQx
NDZkB93nK6of/Atug1ovXYtE8AVaCQ5gxdTD95jbVw9xS8yEPBlEAMQXYUFFFMExN1VNlHO6jp7n
LgyDWTCtiHmeBoiggcYQKOCpk8NVjA4kWxqLTNYAugdenjKxtdUttwAvlefWqTv2BmaMQCQGcIuE
AioZLrHiWeZyVbUudArab/CePjZmuXct6YJuEqGl21sq+BJcBCay/Fj4Yfy5dLLSUXcC0uZfwnbY
+/qKA1Rj1mi0+BEnB1BSap/PEfCnxOrr8BfbZWrQxDvDmDpfffBpGr/hJXapV2z71MJSUdNgJMbJ
mojOk6egFMRtrgcsGXzdvkVDJDwxXwe9+3fB9QOfZ1LB8UqcfzC6+BcsPw7pH8aTKACFPAGjxcRK
lzNnGvQiMuGpHEj9bWoaxYz19z8yS3+86mlaoNdGzGKKoAlzL0be5zgLSGkNvhG4GWV4AOSk/py+
jrygWaP6zNFQq5605VRylsWSHMs0Ai1OvAqdOoeoJQpfa6uggJqnI/jtQfqbmCeodnyYpyveZ3Lc
U3rYz+uleMoOiLP3/LuGo2L4disLwzwnlzRnh1wWe6KNfPw2bXOSi6F2wU75KcsUxislDYyELQIM
zUNGbdRMTIgJIp4mERgMejmZwBLgLV2OjlBUBZyROYO1Faqnp5GJrdgXD1y9FSyb16Xkraqwma1m
vOVTY702lbGV5EUzns++K7bEeqnGxXp1wenjCWKbU0fHgcDVplV18ozWRYOjlYOFpryYu5o40qJy
P1Bj/coq+d9eBtvVsdlEKnmFLdwQASkZj/HSnwEroj5Kn8sji5m9Ntmn5uzNRXXK7LfEMsp2Xz/f
fBVeQRSExF31hSmqXpLMcpYNe2+D2U0QhJE6roU2Vxgbg9slg3miCU0AOqrsmCElZZ+UCtPX5LLr
`pragma protect end_protected
