// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ODgG4muf4C9wVk8ngE05IPWQquF8NOtDc55+0tIGU8AbCikCSt64WPhpPLFu6FWqJcoQdqhyAX5U
S4pqMA2x2srWnwgU0aA8CePxG2iSZTrNTdA4wUQNkeaktHPJzm7SMQhIhf0aN3PIkSphXAKkV+On
3XinGWdXjYVm5cKBVVQ7iP3VAGeHOHrMaDotnt6NetlOkFkvWll1fu6Ll68KBvpb3wJ9qfVeLuwY
ShhAn3sjch/9QTgmorGi6HHBWyiVMEE0tgq3XkM3yza37MYoCJLI8BAVfMUhvLARp+o2qLEHnWkI
w9j8b3XoMmyuPbAAx2z7x/y7dNUM40+IBHpe8A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
o3XI/KM4r+m71TSscDuFIt2OE6fQZezA0FyplGFFm0N/cFccGaZuLJGZdBki2cW/Uq8+NvSvUNcA
JbSifgt0FKfwfQ/L9/cfH3oZuw3S0/4D+vWcs6miWfoRKAR42ZH3+BA2oJyXVHtaUPllR22IZ2MU
qOWKnJPyxPeFzwMxL4JOtDiYS2ETCxpR6c6vlQYyVBhEfs4ZVD+jqmK7x9ZFxtKbHYvGbfthAwCX
6l4CaCAZnNVmhrPDAIHrtgFyPzCnR9HTxwmTCohjWZEz3J5zKgEeXTHy2nuCX32CvwAY1cgcW2Sr
tvpolKzLtpI1TQ1nRl9d6hd+NI8M/U9hs11E0Pnu6gNj/GFj686kKwiZPG67CDj2koEoyhp7gK3f
4Ov1RbWDN1EW3nGoyMsGIQ9LwQwJC8+CKwUyvX4ln1CoppYL16ZkGdiThJtf+slM9n4DvLWoqsZq
CTMgvX1HxQ0G8tlHBGm24z6Gik1PznMAfz4lfTgUCRTBwnjNsmKOOUHEON6dGnQ90UeGZJ8IRPv4
4OwJO9Q8Eht5XT3P2x/ugiIs032H5Nr+MPGEKnSv1pNFw+Ey1wQMUGh3aiuTtIunmeBa8Vu5wU1R
PwqXOM4ueea3oYfW88Bgsg4E6C1lz/IMiQwhrLShyLUe3JmOtS6VrkeiIcG/IHXtJbBWUpRjmM+w
try5jWFGhPidKJ3pICH4R7MoFNdv9923O4NYZropSXK7jMlO+K1CK2MlYc7mGq1dL5N2KdITPbvx
7cau2Svdr5TESZMbd5OAU0JT6mQCAlLaaghWjj8+/8UqyLEu5TB1q3vcKexM9QVHBpzhtZyRMAfO
B1SnPgwEDSX8SNsoaf8BeQe+qCwtPZ4mKraDONLP+Pz+05HxbmZBv+XwNeMsEHdu4hZ6wH7CbU8S
K3EzMeEVTiEttA9iwmKCH8g7C6XHV7S2HcAnAjVzqXdMJa2IWKOeMrCmbbZcKy0Fjp/uWQJB2fnD
fdm/wdsple9RybW6KGzBOdPdljSDcNTCgdJtFqk+yKHFEjEDGtikJqpVUQLBxpkkUiYg/SVF7haT
6yTkt2Z5/PbCg+WRCF0pHL4Dsg4eKm2HKFz0/NagpYgtcfNzPld+N1vZ1jutseOjG0QLp1bjSloN
3pn2WEc7B4m93+gphWMYdHhPaVRS4zNTNmNCUdeUucEzXeu8AP7H4rZEjKy19OJ9nmZXsMXNp0LA
kzW+vzlWEBjna7ZxZsbObQ2bf3o7dywDhDDnUW5WgqabtZI+fe0LBM4neCc6lzi6ABSSe1o11hHk
HmxvQib1aDKKpHZB3SeeBOGRg73feoPvbdlqZUhIVpyrLrhh5d3cJ7/7dEXpMl6sv9qjjEAJxQlM
2c0U81LAk4xriG0MkyiBuo2ow1l16MCwfyYAlpqikNSFPJAoTXt9dH8IeRCsICnvT7KLRc+4ByhM
dA+rQUePb39uZeXZEkBxU5s3AA3Smb/PrUMCTlGcKsx9hqen7GepoNcgFmd4QBR1ovLQn/ime1mE
mWZoMx2bQt2RV8oJyI38pTEP7/kPN+HNs0Z7rha4YWFY7CGRLat6YD0x2oaMy9ysUdIMlLyZxWLf
r4yQ/v1vF9DinmMDj1pn0uMJ9aDz7Ya0QVw6KvDWJcqTaUh2jyo+JtIucNlhTMx1dpUAdShw/j5/
5q8nTNnyRIhbJ8ylZ/EUpHT3RSn4p6jgb9N70TrAVshW7KUng4Ak5n//hgh/XIgGGAhNGCuIJ3ZN
j4pkQXr0ts6EKNFhVmfxvF0T2xI8heuvw5ndmP4XL6aadDDOT7RMB4/pKS2cyWvRW9J0aZWl4+tg
rkaug6wUQ1cTjLTodSJKB6epPAYA6elVN5a5J3OMm5mBM3C0ps8M3FWvtX5iaF+BBBR/v9JaOQVH
+5DkeH9M/FewiVwB8iz72H8tDjJg0vIuZJNQlk7C6GWvRS9/o0GGGN/r/cm4zbJGE362sjizJ4Iy
5Fivs28dma+CGMTXU3t9asv6mgCc0IuHWlQhB3FYPMdss93mPlEWDOdIOQMjGf0EjTdhyLKnP3Wl
lrlGk3zybZ/NpvahkXa+N3BCxl/8QWAwq5olOYxnD0XWVy55WUe94r6LfavCxGw9vwXu1Lag2GHD
q464rZo6iK6JJ4AV7rdKEi3hVPZ0VeY3erBhqzYCxDLq0AsUnMa152ufEv/u4inAT7n1ZrkPi4Fn
MiBeuPVWHnm6da0gew4J9WmA735BXC4f2mCCTQmjxKql6El5R/6Bh3ZgMtzDpYrnI5igzg4geDtw
g5idmGx5XiPT70KeQnukVod1o70hzaXpBDyzSpXDwAIkT3V/fivv1vXbr4p/LYcv+Tw9UehSxIVN
AG6UjwFI+grXt4VKERJKaMdxSQt8UQDkpLjrZ1IGlQWaae4GY25EDhPIsAYGir84hZlZyJPUwz55
aP/DteCE1A24kyJVKdK4PvEjXnYFYJcCJX2ZadSXvPX8PWEMUIjEph/9m59BSrHW4oU4MOq9KuNr
Ofn51adHnXTUzLEv4Tei4dAktXAx+GBb7ljqbJENP1TFBXqb3DGM+jPQ7E7bWSi7i2E12sUBKyId
BB8d/NGwDjqDBajs1WqQxwugCwzmHRcGgcx71XsiOQhxrXJIyEzkNybHG25T6hdDeO+oXenjDU0d
zfjrZrAIQwnU+Druzn3/1YW8lIP1uh1mhVuPddLK0WeB77QTWWda5P+sATTHUQwA1v6aK8wB4LRb
aQtfDbJpCqs1GYwGAOUNaFvZtlRLIA5i87oT7o+xkOpPj/6yQbUw0Upy3sR/X1vehl6tVXAMbKmR
2s9uFSQ1G7ldwjhvf+zPM5F4Rb08qVSW0wFZJmv9oUwyWO9f4BDvc/YTi1WJUhUo5uvBVLPIjBjz
Hj3aGIJMlm9eAzXu2bx+OhlGjOaLBvwiZCpjEeqm7+x1TEMzND5PyiFWwYn2huqoxJv2c+IXXmdz
FIaSGx5FexJ7+AGPB2x4EF76lSh8DfEx7kLqvCZHFvxMWUQ5QCPQRU/wUxGeCksRyD3gPYn4aI0A
EgsTgSZnkBSOx8eFL1wgUIq39Mz4pMx9lC/HWZCTKDDwpjQh95g5GqEDRkQo7xAaCaLBIhuVxuAv
Bys/HYKDy232iV7BUx2M7JOhnSfbMDhkD91cLCpiCuoiJMRLK/DCEUVuyGNMFHcwjmWzC+BImxh7
pftiyADHBoAPhvVynE6aLxbtPQgzxrW+XNoK+IuxZZK8r4CpUbhXNAeduvwVaiuQelYO43dzhJdt
EPX62hr/VLoiS25gl7KGNs94s4PQtit+1qPFPOn1SIKeocWkcGTocMWY5Tt4DpzI2zL90TYEbRmn
Enc0gICr1hyMt4KhZRIakX/URfuuet7iBZTlhuK1lNC3qFlLULKZzinONvHxFW2SUjQFwl4iO0aP
Z+P4BLLefH7MnAkeQZOJn8y6aHC5OWm2KBt0Cv9Pa2N/6b3yXS/Cu6URwUB7oyKPPS83z7GIkrP0
e+5bTmBydVVAgm481bAr7EIdo8vOcxXbaWrqzk5ZIj/VW8ykFmH+ZwGQNszOUFUu8tZXn5gCg2mA
5oDHZafnJykLVih1j4qr3HL0KT0eXhhA+nHl/x++Q74OooBzI3oBjHS8FsxxQStqt24QwEU5x7O2
qJgW3EE4NLZWmWg7F2aOfRCyzY0lHGhiKUENT94acPOCGLmuoTD63sTe1CIA2YIG4wZukvDLuBXh
v8aHb8nZc74asKHufvm1lkh5wjg99K+OhzEfT6ReGxgZ70ipPVYkncauojV6ZpYfzHjouGCpQN3w
iP7QoO7+6YihIHb3CNpvpK01OAF5bne43NffkXq7b+dMrMEuu/v+HaIMbJ2aAgFLGyOgy346SRgu
HVDyxkiJc/DyN5OO6BdRzxtVQ8qJL7k+XGiJyUuXifXCmeM9pJrh5tSlxT9aDeayG6CZtZUuPUWd
kLrlxgGZ8dK6Hn/SMGcT0fuhIGpbd1r8eSuwovpMXlPCWbMHf6ymzl61yFHPExrqreGUwO69Rzi0
tZszomze2AjaJ7XV97OjKAMDgrhvGfGl2AiNPYSj+gGMSGRsXOSB54AdQvu9GBY+gGOI1REoMilM
q4HdN3r8YIpUMLvrfDrZ/tESQkil4IlcbOWWk4xFAbVLuDwJXxyZZ+PN8ZdLxWxmQs9QZ2ACui7N
8eDPoFi4cOFgre4XzMx8N8mpU9NQTxX4lyWu0vjK4kCpNCtIIQzhJ1WoTvij7Sy0LwD6a317zaUN
kzPfRGbiOPX86Ymc2DOL6j6Su+U6TnuG3Yr+Hh5tNfbFj0tJRp1acEkwIkf+F0jkjN1Uwe8K0nbv
A7nTGIsIcl7OphxRQCRhuJxN2kFJ/BA3jMO/oLgStmUXOXjwXKx5h88rc2LT/zS+iu5A7b1eZZJx
9AZbGGwoHlxCmGbP3jF2dxiEHg7Oy+8J06Cg6SB/OVcSDYl9gKgFKHLpo01WIPrPrggJRbsAGPG6
fg+jl5IisVlvpxs0dC7JFgXRRX2vX+KMku2CifOKcw7XJ7Kpx2CLHuepVoKrBz9Vg5zYxX+YMkHH
13ZjjnMsB5Y77G+nVGM7lBob+jNKX02zbEzc8LJ7r65W4HuPMkRllGhhhJQv4jV4gbfngLZEUyQ9
qY7rtc0PENEDrhz8Mc7wxw/sHVeNpn/qyJUvvZrLe0um+elT0CsbLp36EFTiiMfLkfB/XMcDMZEY
rweP7u/tC38jbaOXw6N6ZCoe002qTPMrcHXZ8miYeJCrTXr38soSOPgaMKuy/SPVkpDkkxQAGef4
jDbNwrRHq4dpQcLO4nYTi3M7r/mBGmWYr9sOdju2wJ0AbK5S06oF5eMfiOmzY9d23GmU283mJvhq
7Szmyc9vzD/BDEZRiFrhGdZW36LWcCfPbs46JzorzyLFoJDP/+6vdxI66ELuG/IKozBNHihOHOzY
ZfTY7rq/VX+hsLO4n4WdEDUFYylUzUstwfaBSZ/7UB3vYIfQtxfJhhhziM0/rEjwT7ET/qCv1dzv
+PgzjfZA5uVVNTKwWMG88JbWSbYR9vEfgSUmoOe1Q/OIo/LMl26KDK6shvkinbyQFn8JDJGIRHlJ
OPmw/j2XyuwAFK2zw0bJTgPEtKJma81c0W3byWtjqHXj4uUbPyj9o6gNOjlGSi2OJqygGBQn0mj7
czd6jDZCo3rbV8GaEm/eRiuVTsy0IF8fskIUOkDiJag4Ohg8cnMhnSkzzzeknBjDZVwVn178PYKU
DJhbE4eUVW9g2/AVfWpGmPJIG1jOaeZxjfbsfZ/wjDShuPG2Jsk+opnBKgc5uaHrVOsWHbnTb7DE
lBHnd65it1yO9rQgaajgT/DKkLS5MkLvShD1XuZrftof4jT7BYvadKrARHV+c3W/PNR5K333hEGZ
KJ+0pdvBXjirvdma+9WMae6fscLe5CXkZAuvOq9Pm8XB0lwWOKZeaaZo7f4zuJac9D9B1g575Cim
TC0pyO+T2CKeIgPUCCMtzxcyjEPD7baVnTxo+xVag1oF7duNBOY4hzR5t5uwvgbn7Trxk3Q48yFu
h8Wrc2S3smRSsNDAgZEQ4CX9xhMqhEfbe6rR4dBVDoWhxZbJ4/0F84SBG2BgAjVs5/3bnLeLhqSL
N4JGNE5BW7a3aX43rkYBXkoNoWPR9RFLm0tuqKHvW8bPtH3RGe2NOFmKprRDWEr5/W6VfzRQftpL
ODbZOYdmjy2+j4nS8SNttyGhmdqfv4DNe9Uvr8jD6u/co3upe8OnaxQ2O7v+X7oRd96GHKFsAk6P
90D5d7WF23n30X/geIz0kcI6sbcmYMLKu6UGaTiUceIDw1NpBlWmBSgGPODMOonpBLF7WPZrmsa7
ORugRI9eqXnuPOwq9upM/iE4J+UYCyfcoQMcmhviuVoSYiIrVpI5HWU1GUkaL6pnN1D/PxcUvxDf
9RCjnPW49kONbVfCLC68xO5VO9o0zcUNeh25FLSpNrErVigFa9xFvX0ed13RpdT3/KJX7RfD3ToZ
w9FJukNDAyLCVKBU1DJKM9JaL+WEoZ2MJW9WyJDOsaf2Lu+hALfa4omeaqs6MD13xnEbW5Pih3Nl
BP8UV8cTQI1PJrXPPpxQz4VPXdt7Zdt1188RMKFB9R5ziW8TV7GXt2UGKgoN6QLyHTFjkuAEBKuP
APF/h1wB8UKA1jQCHIcVi7+M70zdECEM8QTAfL/DZdSX2DgRzwEZZ6YLWXnaVwhjWuMMt8EGQkm9
px0wl5Zx9iwyOYmpFkgEgaya5b+HoJmr4Ob8K7+Jr5xXp2+ycPi4gBtFVAVy+y8TXk/1Eq0F1u6A
nYHyLQ0zinSiBkFb9r7J98COIY06KaByu2jFrTRQfy74wbxRfO/dm7GDApoMtVmMsa4lIJi9Xnnz
AOKmqCAwE+mvVFrtBrTA0JrLdVLQMpoNyeR5pW19Bmxog/kG7wBT6sjQV3Tm+73Fg/88b2vKj/+M
BBQu62evpSdndQc+rp+Qol9rDaWXlcfhvgNZ9cnehCABS/raPsVOMuQpdeWv9bd4gBJPx7+UWF4k
1h7WHK0RYy8+StSHwBtSnQaq/876IBVmFbZSD4NCji6EQ0ZaikDUXHa6OfZLHAVafo+0Uh76nmb4
Km3hkyj/jmryQHRUaJvkXgZPPIgHzPlNUqW2HPBERuzg68RIs4RR9B88Vt1XPwkrBmISkFOFZjJd
ADTJCBI6H51344uXI5/caDiWCbopTMWul4B8rik/jEAEI5Guo5izgXwYoQQqWNTf155vFvr+Gp9G
Afmaqe96z5S8jYYDAOgEZaXPxFa/fA1SAEOGSqcPe3RoYJRof6jSb9FwGszwMqqSSk9CtoXiuTTH
5+2JS6YaoUJj/lGhb4+czyv6MVGqTnCTSYhtVUXxNyG+g28bT+x5noclzOxEpjAdIU59cHgOXAfl
PJW+v3DoJBDuU0LJO9eKa3Ygj8XgODtdR8xOtbEd+jx0Gmhl25g8eJFIz7EpkPCA/DoqM30/Z+Dk
0JZpF8RcxTJfc0j3RPe+FyGwN/+7sDMzgUeH5qcwKV5qSRNRgTk4L63RzcLJ6sXrz8RcslPcF+88
axfHsU5x1rEKoJdzNXlrJ2dMNIxAFD7ADdarDq8zw2quj4mt325yFu5xnE6/bs+6hL4wElFKhmuZ
0Q86ettUEMkQw4uFhjohboYQgPY9raTxvE/4KrkoYwN2J57abIARWuIKRPh9p4YhLfmIaLeTnQ6g
zRfDDSG5H0+seBQgaW3rhNIbeVqnHjdX0ThhmbM73oInDLDeVKmDCZxdx/9QK8jQ+QdBxX/LFpR3
8aIGs4QixgH760kpvetVL0Gha7Y08jRfazVE+fnfH0vS1AgX5ULFemDVOlvg/PxnIc2ye1WqWBqv
0/gy8PMnRWflOrF6yCGChyoVz8Q5o/XfQTzP7s4wMdxVn5b+L5wfIfJnv0W7T0KHpXTSfJ3AKqlG
Vkny5cG67ih3YmeVgChuY0+6gzEuSJFLWhoHvNKihQxcZO3gyTyhS0/Q2qMR5RPW5z662W9q6N9q
BfydXPHW3fxowgZ6gsALzEYG2UGeQWlv38c4Cu1xq5nXyN/fs2mXj6gAjLIjALo4J1/24T1baGao
Pf9Xx5igA/hoZEaIKQs9+oZQijVndjAd5Be09YT7bR/jqQ0QJbUQhl9qESsTVEeFWaWujsC0qKLm
2BWP4L9e8xRAgsghSKXluv2YDU2VgCbJyK0BpYAGiRP50S6IbyjstVL4l5vW28GamI7kFbDZWr1F
5UyVt6RkiIHz8OtjrMo4A+MHsfegDycTM+VhC3BUACE4pIaIF0OSZI53C5PHMLd8ZS7qss/9sMHX
kRJp6QYulF5kJCoV3UGmq1kqLwscchNc/qNuZDMIWLGx+hUBbK6sNJL9f4Ei6i3YeQwWqOD9YFDm
cRPTT1bEea//joIcinGGpAzPigKii88F5XZKhUJ/tdqvZhZVI20H1BoU+/aT1ZrVqEb647vla1m+
OJSCTn3MW3gpUrauLBLME2qWdSrxCOhKrARpLZjETeo6pp7pjCsrlA+GVj3pdt+Q3I3PHPnsIJzh
dDuwQARxoEGLCX+RUl4UEh3Sc26OKImJQiZeiZsmrrIAP8U7cTzROkf1zInGONiywsH5CbKSlpRz
28k97DzHLheU4KpgCyL6mwzLP+GSjQ0qQlkdtr7f/H5jand7S+K25VjoYlMn8MnsbB5v+OoG4674
oQwX2Ey3LKgKv2IbFT6jB7Q29VM4C7pTuOG7631Ycsmp3llYCA4tVOrOcq0Ssgj2DjwCskaWjGU1
3tdFh0XRuCdVXkW6tIHbrD313nGYoY4lzVB6KzdkjcObywOk9lNxhAY5qHXWUnoHoLmrnuRxna9l
LNAIHD/JgQTfO7CslWgMTv78cjAsUj3nBUy5cuAcwjBuVeo184SpWJc9Fuv6gc5bDisFrMyk4YZk
VhCWuTlysj6qo0NpH4z+btcgXKDzyT/ouxFVXASRCPbPMuDKlEiciBG39EkrRcqmEdlV0AwR3Lqv
wBavG5/E/V5NvO0nyay3iNnmfctDRqxaELZ8Y9tjtsx/KaMIH1U+3itodVQ8+nakalBX3s1uJMw0
I1BDD+zX/hn02yimrsQngXmqNlFfgejynnLAILWuFZksxGijwbQeRTsOPb2stGG/Fg7nyp8Jr6rS
msAHZ8nv5C+/mZwea5osmf/gvVr6lWJz/21yKoaLSTQ8qRfyDoLbpbS6uEb5Ug82djoZLNhgTZo1
yodCRist6ClwJABLVjEzcPUosXRGqFpQAwoLAdb+MLMLWoc2TlZriyDN76+T6Op4yIPopZiSzS3d
efpUoY14dwh53vs+nHTinQHViGKJ7uU87ak+evSeJDMlIOzN8K8eQ3Y0ueFWAYz84q+dsMSi2puZ
Nw9smgw00GWy8wkQtqftM3P2lhe76GQHzwDXtwFmLtioX3JX9yQCkUo7R/SNd0ewSARAdLXH2H1P
V2oyONY3yjUpkEIl4WA27gQnSM9tBlg59zQiGg22HCkqwImxaInOrN8WONBnSUwCNbBrVyygx1LY
Y3HZX521GEyjKyYylRpN3CK8Q0SXJOA+TwreBjNi4TZiHSvw5awBUWw3VvwBmzwxXEKlQtiXbm0O
ZIok6w75AP+sHs4636u32c+pFYn8mnfgoF7xZB9F7XxrnqkQd0XbkRx4fqyz1hxcclWH9feFhD8K
9qfNoJgV2xgAx63+16hvA2CjcWgPymfTVq0C+dnXGkknzS+wviP8Q4egYg+juPHfVqQuhBfm3GBr
qOUayAJPdqBk01la9pHtX8iJkXT1peXpKkPOZ3mhE18BbUVpajgB/J6kycDNERdP9T6RSb5QBXHp
i2jOdZALMcZAYXkhC2iPQEOQM/FaxJvHEQkG7tYppk7dBjfCZIE0acOB7qXC5WTadteRROj5VqVe
0ZLXDCLQlyraNP4Yua6gPPww7AeNQAkbpqlvyAJmNuOUOIskz0/vmwy3Ya+zSNJ89aZe/OEAnUhT
JJJn5b5Sah4/BOqqP35DqctzLzZx4yLIMxu3mF9HK1sRscgHHX4kvzcrJbjB8m0/IWudoKvG7nh0
PHBMhptOBuB3q1pyQ7xn7zfv7f7FScrGqZ9emQQitHCW/JZiNnknmVTVMw6kme6g8fcodgnHSYZk
kFHZ3PvtwTbtLwDD0bCS7pepfW8a9VK5IIqbtIm4pNamYDGWtef/VrEWKDz2CvWQDDGYH9pJz8yj
L4yGCNrYypXHHpZ7RTSygbZ/p1O7LU38wxOuaaBeznPE43pBBKL0jPxLyZYzKrZW9zATbNio6Zoj
5UUle/8xWtGP+RGZjiIqc2X1f3tsdoUvkUTyEelPNxgQbpDzha7AEZc+tQosf94Ppg5OdeGEVLSo
etlgSzFNRIuj/MM+h9tVWLJm4lLm7bQ7YB6iXdZKX1aH6xDmEsQu5yJJYl/V8LRAulCIFdRqsnrP
G15hKNyNJrkXumdElo4YLmCLKbQ1Xe3o+mP7AQ6NjuccyR3FMxBZgNGMXF1yNDTL6ZXvjVQFTyf8
xvuwv3ZBNEy9r3mwK13JKSVPniofqiOTNr6I8Ae+OCKpVSgXB9lwrzh3vZO0HZrg+Njq2gQkJ1rs
oFYQKf9TxvsA6nWDeNBAcx+RoeUOUyQr9QC2naTd5wIzA5tByHF3GDFuI8Py8UwBeYizN8UHKHTL
YT5aCpCT7QQIR1l5WKNfTXlpKNRwrNyNzzlFNBppOUFG4iVORf2YC7aQTkhzZ+r3RL6ZgNWsl7kO
JLXrScB5vKoBf7XFoIrTJNF7RhEqzZMF3S5hBoggDH670EkHwZX3FRnthEuDw+apgUc3L/IlDD6N
TUi6LQ2DpHQd9B3HXVrkOrXsIZvPpenxKa2/PHkqVL7Q0dSq5m11rGpeiGPD+8vARenNHAA8adHF
igzCNMVjV2Vjr68inLERxDhCmg5DnTdI9MeuEmE0wUNOSTRWcNQxERzwaD4hLU5KKuFJNxQmfuts
Tplkt2CH6v9pqWRbbtBjOjAbTeFZw81HTrlU2ZsgoOGJtyQV+RybT2z11nAoUpOGP73mxWy42y0v
K/xd6CvxG4ndYR1DFeTMjRPECv+xEvYgPUTB3sOOxCAGTZ7VSWkERxdF9x5rL3Sz6vRh7U186HDJ
ZzdXu8U+VdQ9OsrnR7MSE8x4KZdOqP2sO6QGjwl/oSDBXxxOjxncBUpfnU9lvS2BGkc5hig7TFde
ZB939KbWyi1TbD9nXTE3+Xnwgrwlf5eBqo8swvjFgNzMRjtuOfUlLftFSy5G8OpZnhKxKvjrkVN9
3c37iPGtgL13q9epAZZbab+bVOpM8/SZfpkR9OxTtYydKkhOyLHWgbGP0AlxYjBhOyQcFcvDum2J
nzAyJmu3wcZDsiHzaT6BCZBMJP0yT29kKbIpuTfDv5e6yrTHMzDQv/WSK2/5TSqORzlHXRApkF1v
Om5NmHPxXqvXcLMxeRepbNDZjNscmlLU72e30bsdMOX/lnDSKDh4qHtMVP6t/bwRp0EKuj8sdZUU
L7HYJl8ENqS5sK6dGVlXtKP4wZzgU1ZFfLQ0gwOcEXzspJ6bqn+iAqfko7Ae2yWv3sqhVfFosB+/
1bcS1XH0c+oAAUj5s2S8/S8TAMy7Lsm9cA7aRtcDKkFJzROEpwfAdhDluytyruGsdowtzLIMOiwM
zzUj/3D4noxDJTPOIFA/plcUzr+IsXrSo4FKh+PfgLZL+uyvWm7IzRpxVIAkjPU8vJpiGMnVDtSk
0Qo6YT7nIJmnF3PXq+ikuvGgHp6i0rhEEh51PE0oaQUbK3xa/F87o0Vi6n1+MPSoU8GdthqoomkA
FyKDiZMY8CTbud236m6TUkVJrY/mpcEhA7O5OtPQYuRnnc6NZou8vjEHEBQC6bBGDY9wkRpnF0Qy
PzXM7LI2PCibfvY0zppSQtG9avikbBUy9cEZcxoLahWW2lLARFZNVFBdwbtqRqwSgg8jV9bmsolH
KiILsTtWrGtUvBAPlzHvP+sruHqLV4vT8FG4UcwvEUBBkGCk6RrTghwlVgZvtt6ctg8CZ0lrA0SW
Q4XRSaESq4ucn9uk0bDIDj0e7+bixoDZiwe6KRTojwt4PRKNbjYrzwzB4VcBD5X3c+hhyE04tLna
RmEI0m2VtlX/vewlSaIboraMKtzrbxeh7cDQEX0vwFysUPZlQi735sqaSs7FxGhcvyJGV/IVJJ8r
HH86voZpLSpYSuLllWQ9cO1v6S1mh76MutFvvYNtUOt95fTHG0l4joZOzN0gnuRSFPKGAZYJ31dC
sSRSX74kdbfy2ATm1wdO9Whh/aGP0yyCq9G+7e+hgmlbFHwTOhNbyB/eZBlr/VomE9BXMgH3fwWt
7aD+sbIrHda+BsgZp8EF8PRCciFvC8fcSqYS8p02c6oluE/ydSKMesToePCGc934o1Req/fRJ2Ar
rLj82ULXkDHNgXE49JbbKyj4ieBNW4amDOeWQMyxTNjDePkm9T+9pAfzvy+yt2BeETF9CMriG3u/
Dtcjhgtue7GHvrQs6SzEcgOiCSJPtOMmsbSwyGGd0nuCVTyt/YbTdcyVTMdpESty7tQ0mjR2h4sL
ARjKLd7J9dDF1WI5NQaARYH+HyVAdjqDdrtntoPYjRn4EnISGAa2x6165te3EIKBcRBAiGV4M4Po
Zp27VimG7ME+NwjEA52tmU4s1FJNxdlcayE1rMcb7TXA15GbKbtVVACQpT01DLO2LZTUcMb5f59G
7FW821tSre+asxEUHI7lt2hbFHgvnhHvTJRyfBNKTvAaAPppzjUhz5Hf587O+YG6LoqYR1HOSAHH
01ULAJ/zAyzEOpkEuP2vq5VDiS9gNHP4RGgYjUCWjdt3xLFXJccIc2pcIH4YMGe7JW/ogF/Kyy7I
9DM4XVewHGnvJEwWlslXF3NN6X+IVLFAmjJmZR602WFz7mY5m1WzbMiJsHvF9N3k6mqe4W5W7gOJ
hAxvQuxEELcvILzLnWe8u/WiFqs9a56FEbzvPkWkZFBuWdgs7qcct66Ter0ZlSRsseTlIxLlfZje
Y0xT9UxC74sqQc+6VIxzSXktLt4BoNGrNTAUPIae1s0/DueXMWVprBZ4HKls8uaVAOEzLYK+hpoB
Q60wZu8kmpBCsnFSEK54BquqsyoEl/oLcKdla1bbDZcbVA68G6oo3zH8BEg3vfQNhuG4vfbks7vm
1RthxjoMmtPnm3iI9ty4mVYm/L0r1fheu3mN/JId0QMH++DSC6dECI4QuceBvaCd8UAP7Y104xjr
UnlNbvwWbCTN0mLnnyKzF/EXwY5J+16vaf3vRGuXazkYGgpp5KJ9Vmk1H9OwAKbX4yDTAx+DTU+d
Qqf73FCBYzli4WNlG9+hHVmAwivuBYwkAkFGynHV/XYcm6CXdfxPC6qZ2692EU1p2cJ27Q0rf3UC
fZ1DEJ/8YC9FLJYrfklRStzRQFe/2TdT+ahl5TmHHYtligBBjiV1UUwW660kS7neurd9mUp55ASZ
YlPI1eS/bnXIUvJ2R8nUPJ2KI38aiJzg93LSQcDjsnDJUmzP8joJvgDKBRAZixlrSpzEaJLmkODv
InfCFXapVpBpWZk6rogjvkSahfVt0btGsAnJepEo3iN90gdxcPc++tjaBfkBnyrRfVB0b3/OGWCp
YwcKMl7o4k7Bwpdfquvjy2ETK49fsmLboDzjA7hBUxk4myg3O2JB5qjmpyi9x7U4vVfW+P3B7rbx
beJ87pO0oau29jnt8pl4AadWVNNDBhkWiM40chG51WvhsJB9uv94EGSE3fzSeinn5hcUgE38Krvd
0xAsRI3wi9HqMAMp7X2cZK18p6ISjPl0TnT/YiPFZ9M0Ey9HMC/U4yxDeDfcxiuy6Kgd9zQJm3dT
b2HMYjFrJOokkYEBkx6qproBVkjAo7tp6uhRPxw3M+rnlxmrqlWEIHhHIEgtNcmEfJf5Mu059tY6
9qbYjBO02wke0dOrer4peg5IIQeNQA1Wd6yYDjILskKb6ewbqGTClYc2lCKLksAZGgz+WxiEbutx
y/k0IZlu6QcrpR9WI+abMlPQh1dHi5uAGKSTbORnW2Gw2NXNPslQbPsiwsD94//sAgfuABZoKRXI
hb5WnhV3w5UdSHdRD/s6SCa9kwnOQLTGQYDZD+o8FUsrxqlCRvnc7Z2gsfGqbSvvQsHWAVH9xh+i
dx9d5nLZTNLwB63bTXScRqPC/PbqQzcxR/qMHFkIvzcxsI6jYewRlM5DiPjqm9fLjYeyZw9LeBeX
TRSoJdUbHA/fsjeT64ZoGVfoBOnmUkG0um6IKJpH/b7iiZhj74MdXc0woK+2s5NAV+xFl9joKvHA
Eu9UyOagauGpxP9VOKJrqS8UoEyeHuKpJ2Xpw5LsuMroNM2fH536tIhuHKV2h7yjP6wnd34H1HNx
a920XPoqU5TPuHzdFtJagvu76VeMUr+Xm/r5If3JCNWnX9K0xvLCz0ozgzq5MaEs06kJ2ub3R3cu
azDtt1WKYhngBZV/m2Wvoswz14FOLFZSlTvxOA+vhmcE8xkkFsgvhnFhfwvXhFsKDiImakulVJTb
W9n38kt0fFzXdS7jGkomQo0P7xHX34qq9Ry3scqwkBTkPBCYPPzfS9Bye+CkrHgkMYq/qw5DdOvU
W+zOG4QUHcEd5Sar2DgsX4tFCY2WbaKXntA2s4gUzwuxu8dPQrM6yO2qwBfZruVYroFXKj+X4tBV
FkDSrsEaOYE/w+u7meRbWw8ezatTh+ynqDjlgCfJa2Pa6pn5h4LV6K4U4XdtF6b/uR8m0wJf6KLF
HMilcOxaaejDlOZfgnzW3fqzcTujV5fnnKtyiLdCZpaqKPgOzYs+htTA9C3trthyfeY9NihDQETi
fjBj1kuz9ow6XBUj8tMNHlBTZlIoyOoFkC7JZtiktGs11dQF7AB583GO1N5q4G8AmAtlbRlfkXzv
JW+jWC2rg8G79V1eSOcaDkDAYiRDsAF232IpGmUuP4QsHMaQterkKiK/zWyrjcuuznk1L53wbAgY
6wlWV2m4rAquMRo7Mqa69VhzwZlgxJhn7q4olARyAlPvctXbIT+IQyEqz6N3HChesd3oBZNDw0NL
QR1McW3gsbg67HE5yC87Tf/gJoIM4LxS83u4zeVajhIAsC3TTItTPp5dHyk6B/8N3KxGxd1WQEN5
/vcW7tmOOXqF47kWHLWa3/lRqIBEQdM7Z0rO7SKt3xQw+/Hz4w1bl36Ty3Epusa/4AK1AxgY2nuu
ZJ9SPttlkum67uyYyMZrKR0uGFFo6QJJsAwGdC3k7vV56k+3rVor+tRwP5WZsimXFDyZqjhpVSC/
pONr8y+a5iqEcdcl5yVCqXKZBBVM8JfRCJnZTn8IkhHtjb1XGhfdUiW634FeNlpFU3c8TSLHMk59
E07NEwK18+gQuri3Q4psdXXs40YcC3TUcbnybMgT+by8ErsKBm+4ey1sezcLtjB2UOjojga7CWYE
ZdEdsJ6PnqY3aPRuRzC2/L4nb6hNwGgZO8ValeCKoZHcAYzv5vWWV2TOJnvhssuID2opSU6zb/Qv
yr1C0/lqPC2CkT702WeLf11VbKPeFLf5ePv7gzcLAWA72dAXCw5wGO0je48yr2c+ycueJm5XKCYn
sO2Sk2rcNnN8q3kJz05PADeLQXiZaYgw4msuf+doKH1FSoMykJwsx56iGgoqXTVX8kIZkCRJgHpk
p+SVSoXwonvhqZJmj2mdxetCOYFtPlYNY1NdZmA/FCLMHuINCC7JHFG3EBN95eYznG8ukYKNsv81
Q9M+GXfb8RtgGKA+w9yodsY6Hh57iJ64ILrxCa42anaS4Zg/9n7oM8vH+6XmBp1f2l6n10LuteKh
rhATHXxBH1msmlV8cos8OH9BPi9YvXq9B61zCVybjB9l7muSXkuct1B4kVcYDmvAiVpUPntAx4J/
ayMmnumYVWPPK9VeSO4xG0CL2M65zStNWBLWY3PS6ph+k0wGeBlafly3xOIK2/G+bujPPWt49/HI
NHdxhSKDoo7OW31Ew9GUWqFCMCZtHeQU4YB3hDVN+wjp0tjAmKM/wi/E7apBd9wAl4GLq5SrFqMB
I7r/Y6FLQLpK2CCn/U226CbpTwMaOUlngGRdHv1XAcRUQ4OE6F5Shn2syTNuh8J0nMMwOnOXw9Gm
uBnqJmhsfQ/cE8UgWzv1KOkjt1eFIOxz82OXUgBUm/5wTbduKAhMi88H5fjEYksSH80S0H2iU230
4QhGBM6QwnUcJzDB/kXAgMpnTrQFDkckKKYvkCa963EkrrxaS4pscPYsSumndhc8p/Rpz06dd/0f
AAh48jTasE6ab+NFkIGOdt06/LMhcoRiLyqiXAzzhfwUwDVbJRai20Rhzbj5qCB4Ei7tZkAbUV27
M3hL7ErLwdYy0dkSo4SZ/I4eZzjsgfJ/hE2LW83QDkbT/bBmBNW2HjeSAmj/EXhBXjWkNA20R53G
fQnm1el/6rhZCanzCTPBo9x65tnh+MYNp4OSPCXfKbH/KiQGa9PPMHgoHwBern0a4hna/bEgtAct
3GRI8283gW+tpCfvGmMKkhH3OZVdveNri9wJvufjsfGU4QjD51JfOpZbnx75CNrssfR7phleJAyL
zKLWSg4rBkyp2IcwpJ0Uj0THfVzS9p8giJCWHUYllbObO1lGW+PTX1F7XGVVq+PD3WUT6j1BXUMA
JWxhN4Q1K7NIoTQmIf//9F5iH4/grSiwhUZh4TP75GPuFpiCXxYahoG+QFPdX7ycewLBdy7U3R2u
i6ilZHRUTVA1i49KWZDJOqUa7zjU86vjP9byxXfNlKWTB6fHhlBst8iep6iqV++q/KPxLbeiCY2u
Sm72uVuoAdlukUiNghuj/IncK7GtlzsRYMkg43Q80SQnVDTyNy4sxyhkFx6xbF3C3AhIqMg8YU98
PlyZweEj4taqY4JfC3KdtzPBVZZtygR6ZTlSPkFOMo9K40KXE9nc+jEya3h7oD/mAD2vreXSbubW
qEMT7lygDxTAruW/MrTpSAAnFfSHVEloeKxFusggV62o3gCHsJaOD+HxDUpe2lBBvabfe7pM4oZC
miQ8+cNOuG8XWxlp7/bP6ICl054RVvDPX+1WitNin6gxOVTTgKFx+lRBCrTqL/8xANUzxhYaBMrb
afd4FSULXsKM8dpHarjvA1v/0GlDlP71Wb9u7nUjboj8YIvV6B2bN1zY1Dty2ofZ7jsY1BaC8OGe
rU3rxKQRkexNtQHUIy+lJXg5YY44TIDKhJmfz3rqGjr0+gwy0bfgeuyc7s50rWNAnSZBqyn68juf
sOtvVeIiYzyot/+zO85I61gLQOqv9102qlkV+fKLeAyR+QXkOMv4FqPX4enfO2OA32IbffRM4aSV
Hx0COWlPtHQPZoAxOOpCYEbxsdNPC2QCzcvfXVNFcgcryvX3SfB8D/8mGXv3ynCLMhjXpe1JAesn
uSdY5ErCaYVkiW+n4ESFoweGXuXovX+WbImKE6AxifZFp1dMqTzkG0TgyRrbMwCEX105ZoowsgcK
ilY07BbP/lzUDNWyCMDZRgMj5Mr8wBzww54xCYwyWfL4d4FPZpP1cQ2YMXJ0Md+X3uVhttr1NEn0
smvUFhTpGlGxa1c9EguSutNlfFPT6Gx2ROr9qVyChhyX9VBWWOURfYtOGfRz0UcEUzGqS06lW2Tf
bowvOxt2lGo9reksjVlIFzcWQHtLNlF+HVp3kTvoNPLYgh+W+/m72CivMFyU5taCH4i2Ezpe1zfQ
XokdbWZ1/a/v/FnOPU+u+5mcsh13zpbnZStIyqEyX9Qg9jY5kJ26eFG2GM2X84z52s8sqNsgV+tN
+3WyR4QTnGcZBIYzijbNI8QBliKCqXfE0vzN+3bDgU9rXDf4F5lmJSBHRXDe9fNQamUJZu8k8Two
XBzFuf3iMjv8jjDbafrz/IrrKlBXwTSiO0lKWT0+IPurZjZpMibbp4bUeGUGH4+1o4SfEc/V3wM0
839jJnnbf3qGSpy+SqYMU+MNvCHKTpkNXxLfP4+vVoGOS/s8AAZCKYQXHfiuyGB97mcUXVJKOimG
gEy3YRi0O4WxyEwxUkr0j80D8OfEf01f7MygqVzS49EbTrEGN1rK87DbzlypWePecSr6ub+x/Y96
p+qa2LjcMEK17Bnn02eP8S0vjCGX0E0dQW8ciSSNkX3aiLEhJG+/mqjfghIu1l7us6vHT5Lxo9PX
NGDdvFZwW5SR6rpbECHYJz0DrdXnCoQiwEXV3IFCgKWZ3feUl+OAffsxN5R8WMJIIZUbvwpr8zdy
MgPz5+BbwkCvGlYd3zCtY8mS/Qh4wGBSstNwrddRut5330FfPyyDdbcU/nAc/f1eQzeU1gibblzh
aPRDR2IVAnNxn5yujWFyyKTvEai031Y45nlJd86sNR+Hf0OiKm2u7MEiTYP4QYGJAavOS1cIE1hL
Fih8SDTmJPY5AznkFBv3DQSCMYOd0uMArDUqBIFOxBNw3V5ZmDdmhd4NvWyeZ4EXmt+tL/MlFtLC
9f+9xVDJLJAOArlr3OGl/B5y+IdncGVHm8AcoIpp+cDJPU5BlvERiFe7IBm17M9asnT6tPEBhW7O
auZgKnqTpSr2aEw5tAIDW1mjaCLbosmz3T0RgptKdN0wpxnpnfoPKxukyKx3DntE7+rjqG2ffEjR
w78kVSuvMXnoq0o/u6nFQQ7LGKzKh4SLaJQ7jh9LBtHQVcZK9D0K/JC9P73q5DeRE7VCU36WC5L5
x0Gn/Sl3EiW18HuS6SS0qqRspbEaNIOc9kSLH6WLS99441s20R/Q+nmijC0wmrN/chobpVe5iLk2
dVr4V5tSLYBDSTgNp6dG9NlE53d03Rwq5pwk+EvP0+lJnEs3MYuLWWKIkr4ptvbTTanf9oGYxFC4
6zRcVKOnsfxnI6IE604Uh568Rv5dy4VixBnnsl6VTa8ephuVDchDpSIPwYVAnOWZV/duf+IX/YbW
YsHf4NCaruxWDkIJlx95IQKDyI4rnDy7rjNcpz4+o4EWo+SrHkKoZLcAkdlgOWHnopxjQFmT/76i
6tVuHr4Exqxq69QmUWqIJRewegXA3ZYQS1dQNsm/eBCFRyEMFJZw2D7p865QMe87lzE4kj8p8XNK
O5pYWSw4fx8jfJnWlvoPK7nL5ZKMg8H5lq7WsQXLzMYPXHrpPEwJcQ5aBMRcg4pSrprM2xJB9S3X
12ySQUTE5earTgebSbUPHjcT0DATgMivAXzym2iS+Edo3qrfuugvqQsWVZQa+D78Tkk10ID8Lf+y
1KVif7Twsl6bu9ttWmdGe/lGwKGcqpL5fw3XcOfTY4dGLRbjPSd8L8T6g/DCqsi/5fbxTIO0Z/2J
okhCjqqULUXoVPDCXXG1qa5aTSwOIn2FMcqRpuksIEyUpi5uqVRsyJ2/IgB1U2dg++KqnipTpY/q
iDykt2+ZamScF39pwOYhyROidFTeIdgG1EQdPIiByrWC+WaNaAzZm+Q0Pv03bFD7LcfnO2oMYuCE
aMUgf2Gi9ydI3tcTM3MgXmIU8vmfdkYdmu3MMLVNdLu7pYzBaqHMxxVZVS5ZGnM09VWuYqbO/R5I
9Oqsfuglbw7hRa9qgXr1MS4LfHlo0jD288iXJgzFnGAs0cOVjFKAoeMvt9uaLc/gpKBlsc9kgGdo
vr0ISgskNNjScSHxGxsMb4uwrwc7lNGxFEbRLROFezlBghFu9qK9W7UCnLD+g37jCQdlExqkUTcR
SQViFvubcBxXfSOgAQfrE9D+6R0nQnAJkIVJIX14uw/BVJh4rcVCnUzU2M3qb5mfoMGpHvXpT/pj
9n98ZTRUmR0kJE9SBesRzIK1AQC1iNRvAzNqr617ijox/1mzmEovQi+6OuTbPou6Emcmoa0p5q8y
h7pldTM3ME6K0/Bsyw6An2ITt4pXtcRDTjPZYkRsf/HxdRK+asGPt8WcCCa4XLScOznubJHvkkQG
x8jN9d7u4zSPTeIQHzsPrupW7zSmlrgbWZ3Yvd5BPFF25aZkZWsY0hVx2RTbt8QsYWYAcWoFLnhs
uN9lMOHwUicjwOQtAAEp+lLPeqB8nnbOmr41fYESUYq2NTEcpumQNfvQRkAYNNipPS+GjoSj7Jg7
qZfbgVxc2m8FcSlNyG9v9TA8n4n040q3Kv8eEsNRJRFOix9PppHpJfcBKYRgePNCl8adNrmMlkvK
sr1vJm/LE1cTdujqghwsZT0HzqwWbAakmPIrcpWhLokM1+aUyAeDXAvLrKj8D8evU2cYvHS9eVTY
9IoAedW1o9szUIFfDDkmr4FJRw1xubXOcjnr/CBrzxb4p0ZuuWskH+K5tfjOLZ2RcQAlp88VNd1K
NwMoJ5IoRaxAvYpLrcSt6oTgq3NXJR+HsLG92ZyWqenqGt1iOpe6PnuHyWq0grebvRViBUsCS/Rj
l08YGdvm6bksO5OigoesPjRuR7W+rqDsIrOdR9d9E0Ug6ZZdHVPq6csQ5Y0hUNCeEoTjrIumQLbt
gIkw0x+y66KY0pEgjWZ+ZKRWbjhJjKcYtKFF1RQxL+K5iqboooKrOR8TQkRwza4H3diHS2FKYwFD
wxKt4TnM6i2o+VCItNUhv4/qFYs9kRGDDyavB/hdQfWYAlgFSThfBm6Bur1qPQfFN6q598ZaqRBS
3wgvdBKcCOTHQXaj79+j/WoeEHKLdWR9pdT/w6bZ6uCEdsFBvb+OSvXFUPKJk2gTGsr2hmZdctYy
W9RzB3704g3Iy3umqDGvzy+tgub/DzM2/mbo5dbVQ3pgiaAN37rdTymhoAgrERiUYzgzmXAFWaIW
TYWllN7konR8O/jvau3YCbpXKnm6X6M7eOkzsnF/KHOftK+ywbqFMEDRgArIkQQjwt+Em0G29F1e
g+FXuAvqdKuG0bMGDnGLBpu0eMAKW5o7wzZGTs7quVSR6TW8+yR41JOvcP5bboNapS9WuUm9Q40p
f4L8WY8dS+mWUJ4x3YTum4W5OKzmjeXxphjptvHAP4qLagXX63kHKc5b2BmBka1MfwwBEn6ADIus
zPeqywp5SyAVl86PNmly3YwAxTvVFdNnUxVrQpi5jpSQHuIC6XYpCc8u6FDqefICai4fTW9Euhat
1QJ98r5Ml0AbwJfeycLhwuRui38wRjI68qGiI9b8IZ+OWwW4P3ivtchIfeMuPbXaYJhos7nlKA7A
I1Q9r8GpxgpAKXkgP+9prK3DdQzTLwzXdru5XYxhckiMlkgvTnzy2Z9f163I4s1SF77/eqoY+gTY
fFwFAtB+Rxi/ohAjVKoAAL/hpS5tlROi77W/SRvpWKQfeDv/odjoZh4OWAJcnBVYPIN5onpfOaXo
EBXBEJFvzNVIu3vgzbsJwjuAHZjzXt3R1JMeOBIVHgqFIptK+zx/oOl1AA825nmC5Wu26V/Y6RUa
HwzLSnrVm9060S4jKx5bE/0yETPH9vH12P5sRXHjHGwZu5IKV1hIsFU9gxTm2IO7h7wZLB43mwnY
4u2MMaL3LfKn7efaerAMB+K1iJJMG2UOFXKZ1Fpfj9vThKjl/ctj1/w4BcStI3E2b4fmC4kDxE2p
RnxS3zcm3CQwTjnEoSIkS4udq19JdvqP4cURUIM7frrB/EO2PrqmD1WNMDum8K9xDLHZePKDAhzX
c7Q7ZXeYp6tpGHtt3Gg0ROZH5S1PzaIH402aMPjn0jtkgWRYd5fSkYTTbh4v7x7twmCg8rzoDkIA
iArQSUvTHD9vB79uxQ54/m9X5iRIt1Nnvw1mEYUNDDD/elIhkjjrrZnxyvtU0Un8JsIcmcOLb7ol
jSzxdXiPfmhCxpxEeOupz2rjZ2gaXUOGtMOcHhY9QlDYkQgF7squrhY3bI+oFVk6cPhgelSCZ9Xk
5YTvPX3YglxujsOGRwLXKqmMC4FG17JkVTz1/iGFui7hQOdIlNaxVnTvslC25qcieHsOMjEVlejZ
3Uzqz/mQFrshjMEH/VQA/97dP9IJ2Nl4ZLYyFYSBZX7T7yLF8/XG6DkcMrt8OW0QzY6/WDgZ4WFc
pc9gK4x9esVO5YLAPkkiIWWnTrLxRdpd/CTvlOcDmZdmiMYtqlEgs4MBg+ml1KmDjGVg8rx7M1K8
TYk2WRs83MPo/BGi67SvkncXkABXykc7gz8F9l1A+BInfl9A8w86VN5Sa6ZGl9u4Deiy7LIfyDmK
yKf4cFSuWwFruk0HnX3yt4aCRUQzZ5Ym9GFQXsUHJhp2Ob74Zuy4c4h8KQo9nVKaJ/9wAT21HJqH
q2fYhM6d99YaTGeAgb4FpTHVQ6UrSNhAsdJTSXrGh0WNO3f/cHDjK5ltecIJ6qfz4gXbOaw/IgEy
XMugrFKbMgh1HSX/EB8J21f7udv7aGJrHL4HVhyO2fjbLSegqJql7X5SuS57uMgarxBx6MyQsbDn
vCXk8Lb/wxbzXfocmrZOiq+aIV7RCeMUQNXnADS71VA8TCGHAONoEoXVG+ZJlCmVpbjb0LcOdeYO
evTO5O+5NUP4DmF9F5Jz+Fg6xjF8ABXkKsIYvnSYrY6it7FT86tBBJTPcVmTyJ4d2ZGmTPykwpmX
lZ6Hr+y6Ki/cVcoRF3i0s5eO5yKrDgyVwkO9oWUiSPbLf2N4b4yo+zlSCACRpgXNy+uOnreYTokp
NqUL5+wkAnzAlRLqEnKNP3RJ0ERsOie0bORH3UFO6Sstfym8Y3fNeF8PLB4LqbwTVtr+sewm8mvG
T3Khd3YBgD18zsOiVPauEjsbVas7NugkupOlhRUsZ/e6/LnYAu0kYfQaNk+llJgRd6QWgLpv/EjP
+NhSFAHQi5BxL398JVT/ZDexkCOj6Rimc1q64/x6DiFPrFHFwD71M9Ma3OBKw4D5q77DYmGxyS69
jJKUVyMz5iEnQJfL7EgXDuqPu1YNDXnX5NDWKgXJB6cYJpf4EogHfI8J4XD00jkrPd+w4umnD6hw
rd98HZ4jLpM9y+kpsqeN88L6bzDQd+YuFTwKoRr4YJCb9Y8YBcyp+Ify4xmvuf0tkTEVHbXMGZZA
5F5j6YDp0k4kZmmzVrPYSCTUc+dByR/rGW+e9Yz7JN4e+Lu3cGuJZ9Wb8qQFLkJ1EuCJp7C/sFnA
Oh9ljDL8z/CdW2l2mfWM2aj7yuzlvq/fzV+sggboMTolyIzxFofydBlR0uPYVbImuXKR4S+OpQKi
Rb60RVgCCyuVyq8rSo9znwLPjoNXdCQuGkip53D7hfhoVooDQ214HwtAPr0VON6m3NXJTKs61SGi
cj81mRjgbG4iIj4AZ5VlJho640YpuCeyYqh07QwPqbacx8uym6L6U3m5MDjc72N1qQOHLboZZMf9
73/pE5Ecbok+zxb3XbVCXnwy5homdoGtXjX3Rn2aADuE5k8jnSMvR1aIyxpWke1ZjMt5SI65fcE8
FHYsTNRMGRtb/GaqIsiC/XiCZkWoPS8O4A026Y+ElFkbeIq+4HKNzyD9TQ0aRHpM64l5h/oOBNfS
FvQoay8vj2ROgdz4oSzXsJVkQzv5q8IOwDAy/hAtXJ1dbJMIQcWPPFg8YZeNyB/75O5r5VACUOEl
oGOdJhiNSuyhaZjy2AOBxObJUjYZhFoUpPfqvGR6rZ0P/7EjtylcOnJ2KgB2L8fG0z1s222gbn5q
vRlS8V9FQdLKkGko8/rCtd6dEGlsWkFN3yeO+6ixOq78n6Syn4ItQebq7c9lF5FUL44jdA1TpQBz
mrIe3V/FQpluNAsnj+RfVAWehGUYNDxK39vF8Lk4WmQw2uRJWAW8ojwhys5+0gRtZ+xrbrncabsb
2IIqXq1velWxywLjHXpUvKD2q0jZJuIatmQY5MHJObd8SWC9JEw/HrXyqaHJsTiH9+OUc7yGJGvz
LZjX8ouhDyYCdoNhIjvc65vKCHTLyzNTO4HqO/jaC6sTqepTQ2Fo9yeyADTWhFSwvmBu6MNzCNFm
0cPtfTbwZUoI/WCDrjYD5CCxE/hrR/Rvlus30oHRV0CLIsvUtgQOXBndn2RUl1asHqiPZsUPpjWD
qsHEbn8J/bjVbkL5jK+oDp/lDbMreFHbYES+QgG2Pnv/dkQirRRcZBg0Bv5kuGsUeFgVn857a5LZ
x5ZCflF+/6ZCZHEqOfsuytz5fBOZLMdc+QfR/YVtpEStb9KD+kHGGivRNzEI64ieJfIdmhr99luW
uYwcuNKXghJbNedSsf42MACHAFRmcfw6HHraU/9GIDJyZadqF6wnPaZlLuWskDGygLz6CF3Ahkkf
ftpTkwA86OGR3GkZf3Zd7ehWvyMisQLITYPUwg17erh+o947MvNvUrHG1fIOMyxbVu2iKi/3GHXn
3DDtummL1m8i790B1cML7xqsyHE2sEJrQ58WD+2+4BFk5f+JpY4u9IzFODQ+QKRWm2ZDPX0fsKJn
mifysihWXc1fMxo8+WKVnP4nRNMlC1JCp3R6e722Yic7v5zS1njBuYF76zANiAkdG3NjZvqiLwSy
jTS38aegFXaZ3yl+5Jmrjor4NHL5YqWEi/thWCN7SGje3pjot38YlBvoNHDoFFSIBmripo4USFxv
l+WZWcU90OEwzpY1566tECbCm49rq8zXovRCp/MQHoXxuubfwuBw2lyLyErORBf26oQELhzrwGaZ
9w5Xb9IDEGXUwD+j8iBVoi49D2M+OmS81XXJtuBPii7HTdrbDcxuA8pdMM9WLgz4OlXZiZ1Z7lZK
RI5ZP0DbP/ELoTk5r5QS3TNLL/g4CmZIAzafnnra/3nC0lCXy+QuB9iSG5XgtIdOAHkwJIgct9DB
VymGruYXg6N+R4TSofo2nDZP82sk9MYMxgymESJdUv+5rftESoD2a2TXRUduC5LKL7j91oOFj9Z9
oZAUyD/xQuH4OSwby5lPqCa1pzoP2xTjMd0WY9VZrctBK8qMpsqJjRxy+Ixsfr/hYpPw+VSJpZzL
pilecmW+KmC8IN4xjGVXPqalV5+v4bciTtpeuNGso0FUFAqCln4UpDqCDlxGKZn2/0Yrd6svB70Q
HjjqTLw9voQTEbWiNVK/SC2Fk7OJtvvGBd4fkjvQau+nLRyM8Gd29AbR/A8dQmfwFEvBMKCHuhKM
myEk3XkpY6pTqIGe2YTdG6AT8AYHkN93/6IXdkhYhF3tCb6iYvnDIRxWlzi3WmO3YyYRcGjAlc+A
+tWqdtGW6jU0YIqZVwxdkPklcisn6vpIoXpiYyAt+mvETFnTetpDc6GioJEmuhY0emqNotnFMLzY
NfwOHiF8DkCMv+7Pw7z3RnC79Tkx45/iNXIQwV4hF0GaZNHijG4yzcHvyHCbZsdSaxB1h3CPtZrB
mg4G1b5XJsQMbSlFeTsWCsSbJlqhUKUIEIkr0WWQtqLdsamq30SIHk0MTkGPtwcagMDpqKGpXLmr
SLER7ZFcGPtDDR+sdtoITOuO5qzcuJGggCbAO1d4pINqnoentWoxDyZvH29h50fs/QZxQoApI60E
JIVO7hoET78yC/DRMpK26KqWpGSCigfg7PupaGqwy/3/kyCZBZBfFXGsJ2a/1suN+kEV2/thtMS4
nwNtOB+ErTs2WpT6h3k+nEuPpXRpcvVJUW0KBudCZlgdn7zZiPEg0qEMdVIbarnszCeqPyFsTrUU
IEpIus7BQVHLSrNwazjKpKL0yOtqrTYJgv/1serGFyeg82huOHGsgBp68gpAirxxBjbFR+BvU5aY
0Rmwdyr6Rii5ssNn60thO6inOS7PQDr0YP0mDq8sMoXuLHzGZ6y0popwJ8NccsZi0i5a2e0YFfJ3
dwZEayZuuaHV5lUwjsiDK+e1aYs8akYAFediI5HBv2amSEQun/BZ9LfSVs5/0SuszZ3bDLcSie6O
P/GJMoGPXNPBH7x0U197jAuhnYd8jsEeCJEV+rN3w6ElM7r2BDLKEytm0mZhaTSsnB+X6JM/4w/y
FD04V1PpqQfPI+93V8fBQWGxy5xapbbea0dmViVYR8ysPGazxlto50VYeOsCC4Te/HtKAY72/Tlm
sJ+WHM9j9yNWvYRrhTJpImwTe9RFlMGxnLI5/WmEmlyDQ1hnYdFzobD3Aa0W0cQYwNW4Oh4yqPtp
M91nKDdus4Ynvu4qzFSe/HSrPbVlDQn/uTslhm7ywcXxbWLIujCD0t0IQERdiWm4tAXGhIbkNYMP
khLbBbjPwMt7y8bc16eBgl2Ht8CNJQAg6+GsPB2AJ8am8VWoJ2zXitengaaev/vgdUqOLCEyQtPo
7kX46EH3ix/sqYNOSVnCJHxhUcxRjqbovRtg9FHFlOMz2uwxIkflug0y0983Y4VyFxZDEFFXdvK0
LSiM9MASiQZMFMZG86B5El5N50KHyd7QscKFHuUYrv2nbRtQKiT5oWkNolNv4WLREW5pVaMK/q2d
pfkjjOhNoNr/FL8biqhrlFkIkUare9Sku++cUpPFfvhfm7/GnOjX2RAEsOxer2GPuzlUBgCwteQj
zzPIaupHjMk262UzargEMrA5q9VCCPFxl5wF9dGhnm78tG+JEr6UQGN2gwY7qE/zWqJOqftx2eLl
+TCBQhUnB95fSgJUuNJGAABZAh8R0UN0jpuoIcUmaflQKCCEOwhZs1Hlzj/GfdsBbBKaWZntKTV5
mtiyNIb95ckX739t0KBLwWct2ZA5aOvOHPHxhsiKBO8xlTpj9gLy3OQNYl7mHzVE7Ize2Sfw80OU
f9piFRSrWv+Ve4aJwwQB4Y7cCyJA6zXkzSHcBtldLQiKR1WOaxmdjaSQ7JJW9/stJNUnpIqT0q3I
PR4iPZfqRKie5AiQ17Xa8URDGpX05qxr1Mz0gSdByu1chw19bQ2bDXb/7U2n7M/Lqs94BotUOsh8
10DngpfnxyzlutQVvIB9KdKJ2Bk3XRoKg0fQFL8tU5iXKoq8lLxxgKyhpuw0G8VT6VPrHQWP8Ilq
f+9YZHoHWUbMwg/JMewyNp4a6BYU9Co2fdwMR8QqRvDKBRaYjd4cUSyldrITkMBpMBPDQjj0weQg
TQH55RPtPmN8Q5XrOFwFeNv3112EeXBhP3EDBP5fKzv1HzTwBa75vfcR+3ShXCX9k5lLAOp4WJJu
HSniF+EOL/CmluvG6foDi2YeFGeLzlEjf4qpH0yQ9ajnpgJ5C+Yy8h6Olk3RUwb0Xs/01LQc7Kwi
e7cZI/Fg7Q7Xhic3nFUKkq/Ahv6HlP4pwJwDs/O3sFDITWD3uCFz2uTmLsxkFZtaTD054a7Q1p2U
7C8C7ETqpVaupf26gP0V4xmdIbo9bXilMvFgN/WB9nSIUoF55WTt8jphcOp9SHDWojxt3yhdz1mp
1JnnNwwwW9Bp1Xm6T7aF+67iFpx481xodFbY1n1NnoOCPOv1GG1u9qmWgUn33w6t56QqKmFmcoPi
bOocIm2vA5M9VC+fJQ1MvHkg4kWMimVWM+Pd8E77PKrbZM0jmXvJZeVNdr1wyY94I6KNz4v+rSI0
9wLNjLRkkeMJV6OPgo1epTVlLVejm2k/QOw4eUM6ZESFw9YM6wTr7tvOESrvsj/dOK4KR0bCN1sp
viRSU69Tp6VMfPpQkYkzFg55Jx95DB6e+lOZLTouePEx7hxswrLDIm1Vjyeb2HinS+C5sIw5+Qkf
VJ4vluT3YVc5Te/dpkH8lHgSqycbHGtFic455kcNInXL9um05o5Lb4PAkBOTfzJp7PMLqPg6LMT6
QP7J7zwZz7k3FaXaiRAmqFzpKqm0v4+19LKdA3pmyJFRPCWmTChL5atSslORasfKtBaBgwUmbxwe
ppiT+QxSjwiA1htCRb1Y4iFpEQQOzmMoboCAd83iio0xfgmlg9D6a+z9EUxUyOL8fhoUn3sdrpg9
XRItl+7O/y9t4qjzjeWeYN7KWgRhF4bm9lVAVlgrw6OdOvX762bB/a4qoh4EmfsMhU9XaGc5o0+c
W3Mm6i2lKW79VW3DTxH23rtIFmqrY5rHICAyB9kBJs5hDJEa6q+MIt/P74uhLJRXHVb0KU389egB
xGfMj15ebjO9udo1Zv/zU/gN3m3YH8CRDmX2GApKOJRtfEx8N8RZSFpr9HqcPRUwpnfPw/J8FUaQ
vuQK8yUbB9SarAE5g2iVNxJM4fhgzFiTuQCRlzdsmtZjf+J2eh6x8ckp7xtl189DFGvCuaocG959
mn7vrv51RqEMrkXBWxWE5zapVoPHfr4zVdoMHmOueipTHdG3GqqsUIjXdZzZ0ypbmBRmKZp7CnTv
8GyQHcAWZ3kP8wofY9oxyoQlbBDju0QXhzli6qWmShC7NtGmjG261VQmJAgFJbfQsI0imrOeQmsK
1TJU3kCxuCDw2M2e7RmOwRrrpVEh1GDgjXoPsF+bH+KJqDyq4vpVbtu3U8OgXIlvldf1P6Ir+vdL
m8/4x2/Qo9MWwlS5h06TMixTz7mUz/rCK1ZnPqevV7yf1WjuPFrWs1BFIBDdu0EMgyam0NLAHvFe
y6F6TImo6aXgkQIP3wGD4LZs4GeT/BvXSTim3q3ccqWYwqCzrExQp1mU6m0GvLPVefQXABk/SpbV
gY267zKwY+z9CB1RamZYmXOXLChraYnTItdZ+/4Fs7TVMLgKO1rppW35CTDxqzmRNeEpeZIVSIcI
Axt0tRjkMz7/EvQywuWvVN+mkb8K/IXMzEHG9J/BbR0QQO58R8DFtTRB1XN8CwV1Drsqf4L64HrW
RkCMb+tEwuUO57YV/23sLx5vjMZffWfe9jj7RMV60nxu7Td9myNCk7QX/U203lL1mQl8RrLG7Ol3
sZYSBEYCFPJ72rOx2eDOw87zepx0Jxo8v1AQ3KnyQhbVG99pLCyQn5wpKrfr7RZtVKbTROFg06a8
8eVWY+IvFGJbsRykID4vIMx2xGygzAviSzrPRgw+aO6hnZvakd7etmM28ONiSduecOsjIUGVKu46
Kf85bNYjj4EzN03jqQ+kqQ1Nt8FuEjiTKRJrr2fEGd6J8DB/7MrxxKQeR0OKBOhM42OD/3F/OBjR
6mUK5v7FpFZ5mLzbYwYsU5VUhdAFXqxt9mQ55QzZyEloIlL+HxGymegqy3URobr5tiE40R4BF1EK
7MRiFTsM1wfBPqAeApMZ3FCuCYbsiZttBXri/LKgI50V0iIMnH2QxH3F9+qZj517C622ow1QI93h
fcP4rcYbUtMPhBjoNPABwksaczd3fSFAXnfJbHrAOLCxMk3UVIg7MuEvr6sDnPvw7QOq4zoOLmVm
sw/j7rkd/k5MNxyOGfTR17n95scDr0yi9RWY1eSK41XCAq7PEdxI5thofSw5o/GtySXZPWxrf6ud
VYF5GKXVyj4hDUUnRNcxwDkPKy59HuK6ETk53GUkCOZJANWbDHD9QzuaUYZRcqthpK0BUGTo6GCv
wlKA1shJAs/ouy/YMVNDVqGKpeQyja+J8md3EX0APR/WGtQBJ97+eapoooiyw/RFve0YrcJTy9Zx
BTA8CO1tqeMVGBaZK+lLjZJU5iUeICO4GbHFau9Q2yo7kp9OSgXmZJYtDK/KmjTL475CzxizRl/V
khQAdvHFv+Uno2kQnDNo2RtR2VuP5/8+3vrtZr2D7oXhHhCc88x7zyI/GPJo4TA36JOueyUtfyeE
61CxF5NQFPa7hCC5YscHHMkV6Fg/WCGtpr1mkF10T02WusrhC9AU64mdAEnb5dMwwhuqRurtcMAO
eb+5UnEFLiSOOf1adl1txv9+pmEGs5M+f6MdIMciz3Yr0Rhls7KCAV7jKkrlkfi8BgzT7hkHoc6W
8eryR3QE23879/tDJleD4OpAiOZFw5lYSrwW4OkaQoKbRJosL8nu8ILVYFsmEyygh8ney4FZdK65
yZ5K9KZa2rk9qqnjtxaq6xJs4b94QUcZGhqgcwhjU9T9jfBx83JMFKhpWUVClTrRMf4lO4PsTijM
G5jT9J0QOaM7L66chOaRGhNARSiM1rwaXMuk55Cn3F8HqhEM17BNh4B/rV9uRMi0hssEtr5ZdZGP
09PwDrArvIyIApfW1ZFXRN6L2aWkoYLeRqP7zrWWpO8x7J9yoEf6dMhIhQQY57lDHDNP4PE/jd1u
d83U+1s+2tQXrRpF5r1byhqGm3/qvw7VsuVWAmudO4xFHACkuenAiVsE9y5hO+0qmVU4tntoxLKn
8FLnq6OiQ5DOHIaYAGbFs5hVl0lao/8ATxRD6D92CY0h/nL8hdduQnXIe8dCF1AvXnLKxKiHuw1f
VPTJLeDvvw6HnMl+8S24+czE831l4p17Wr4Yv3adkZ9WZXTI1xWigfozwYh22qhCj3AH1Pn7oXms
EDilJvSzGI67zCQ27qO92pftcVwRANR8Ws/zGdLOqCRM6UjlH7Zt1wDaBoWRSBYKUfzBphIUlOmG
VOlwtA5GHS2rHHrxwAoSkVoDjbO4KVQGaendBHsSC3ol3o1WaUZpiv5kwk1p3ufSYdGp+BD50SJB
//wNu+19hnEaGLb4sslY9/aMjH4ZOAkqz3CMklyjCpBM9xAz99CUA9+D3b7Qmk6IyUdGXi1GA3kL
duLyvhUCUUdj8vDdbk7gHQ7snpkoRcYsvX7seRaLjSyV5uzhQf/Pp+uiv+tNhYZuMGc8YbBGYUCO
FRRDbL8eFyRmF8Zec9Cus6dmUZhAMLn3hfeSIQ1razdrsmw1b7eCMQUFqy6wy3t4QJ+wK7WimWNg
qndQBi+Hjl2BGSgdTDPmX0WaH+pfqf9TMtbqDzIMELNXUu+PgROKIKC9v/ZUiHeuN3gApHdxjdVE
GEmboF/sqiyGdldQI7RdM/258GAd26ojyLZpZV+Mx2KnPh3h/zzdY7UBZ5HmDXAC++i5F4VNMB4B
AAkYJKKg+9NCZxx225CTrKDZvmtJ401xYCYq/dycE1kfxPDagq7OYuIm6I33YGOBaYNaZUP6ZCmj
N+YSzPH3PphG4pcTElAUVLjg1WYIdE2Pguq3EFW5mtYzIr6OUwjRPx31vcyYlgKD+r83+iPjTcLQ
d7Yf4wo83Yl/BmkvfGBhWNUPhRNpdT8HDza5wxMddLwrGGrhit6IGxAoM97TESP3RLVG2onpz3sf
80Nrk52LY2R7LB5nRnAool5y8swJoy/GN7CZccnna46iynUTTr4x9JxmCCRv6pRB7MopXQhLt1k/
hUeScSR0tRzhHrn0n9q+K/iG3asJMvfxsPzmzMRq/eWgbh9XaE0PjS5JOOecKl4j9+Timv1kOhFo
Cvxmb2385A8to3IpxKqQD25uokFPCIOWZZ3NhtatiPeJ2wUCfE+xsCd3DlxUApd31j+xqj9wK45h
nsogczE+t6y5jg8BGl+SDlAsi8J35I/geUyGSlJiNxJQKiRXYOz6Pe5m5EpJnPi48O29t1RT3ys2
4U2m2rRWktAclI1iB29kxs8IrIjmc2sy3JGUOnHZ4Eb94QSUXW11J7p3fO0PhcK+knO2thFGNlHp
u89dA2d/HqauwUDHD2XskVTwdGR9kffmpUuqnZQbRHmv6SlXWWQLVWAIHg2pohg50fJ1Fy7np7CP
RG5MLZtebTniNyYWDo5mijv1rASF4cfEMeT+STjAfXSpOyZKWpxUDdWcoeZiq6wYGLLTjLJfk1GK
uwJDrgF5o4mhoMYo5wWAEH22mvoFRf7lMljQSYMij8pkz7J7h3rOdCP3qANiy0M41P6uQyPissAo
dhw1Vk+0IoG3Y38mS8yx5txaHymuXaWNs+wcko+jVw1HMcdmb+UnFCv8GH88oIV/+hrBweud52+i
dk8zolCxom8EExsapq6dyzPWuo8WvUfPQ0EFy2qL7VfK4txBb1UPywDyRsH7jUV1lhazy2Gz+bgP
+mYp230fNIT64Cibc2+L/erAWD8vEwPEgk6B4cInzIauWB+O/AiLskWwv2XqypQgVLbQCjoQbRxL
CVBAcVF9OxPxTXWs9UBhNbWRIQFmT8T0Tmou8B8yHcWErVC01IM0tYDpSglzLYB7ixjfdXJRwIhK
v5iDTlLh1ndFOSShiQlfTsP2fqKSp1+K1MDIKO8t6w5b82W5Bnq1jZDcuH+13znSy93HFMLtwTuJ
SvfSoexyMZTt0ikmXB9jPT4V01HrHF4i/t2hywiDEoOYWtfESK8l8xrxzO2s5wTE/Z4fcwxhDWWv
eFtCuoRWvXoF9QfstQM+8H07Es2Wt831GT2fY0bMVw7mntDT5FRfA4BVTNaRcLMvgODuU5/x0mbb
Bip54GhUNkcgO4PkRMgIbQpyAOAfCAiOhJTTzaB+xSAzBaW6/xlBRmyRREcTVRLsB0GuBBerpv4n
SAyVCGlTlg/bAjZ0YHSuKj1AeCKESicBNmr1pgItZTxmjwHfwUCmBx7RwkU6lZoOpkfK3drH3snx
yEHiI2G/bdBav/fBrnUHl9MuYXj8TRU/rXAgNZu3qtduoftsi1oWWMLtHMZhjXqAyky5LWHrFLds
WqMh7TGxuEF+2/LrXG0b16aTXLw78F379ZZe5DOxZcBirLfl+enMgriMvOVeT/U7C7lDR6cAX+NR
/GB+3CpoPGs6p1RNtW08x+fF8fj2mEpStCHRMB0zAaAiKkWgH2Fee/2hQ0FFp4Ho2wonSguaeWKD
Z+Bqcd7as4DlkAELTc/BLJcg5k/yhUpeLaGe+rBkdq+sILonDPXCrP6D7zrV+2dRRwdFbkDnkbiJ
oZC/zzzdrep6KFQvUeVu+wqOZser7RRd6CKvLQWIfKruQB2OrfXNjP+y4vvehG/eqP6MsfCviMYt
KorxIf3j0BYaFIgBfSstq+SxCvCbhnvTFdfySzlMic/neuH2AHpnFn8MBL/xEFFdx2gAX1ixJaMz
CNfk+mv4DO0SoBQVqXHj49EYGZkDbOObRNzR2vfqTDJhOV0Ry/jHaldOkGKUupf8PiGSGAuYawIX
qn8EbTHcUuKv4I4icmUP+VIRy/9Dwx+b/fjgkwvdjmLq/+4e9thtMWTLHIs2FMozzuQ+5w/x6jkn
qeNjjQjwW8M33a7RALVUj8TyTJYWuN4jxHkQFWulQyQHas5qhdUo7ld9hwBfRPP8ERVQgWJFloPZ
Rq/MQu/WSDgOpCrCNpsiSAwo1WU5KnWVLFhM91YUCvi/1dVIIU4TokfjYp50NS3gqzB7fvvCZ4l1
9cfb6+o2EMClnQ744YpochB7teNFLWXCnyoWeJXrjjx0uoTfgcF6dZJh0zfY5J/vB2E2xDAOTxNM
tbDMQhbGgejDbKzt09FOVJ9rCHP2yOzganJP/ylV830U4RyGzkWkO0B87JJJAOangDp9fxIPdQpN
5H6AxZFYZnnTUQDUE8zD+UIKiZ3rTLDqv2Z7MTm28DcreGU3uHJO5c7hFWGYp540BJ34xywzGq1w
9qbL8ZTJuJQhicAoNM6iwKbCorzE6hNO4P0EkEnGqcXwYyVGTZzrvQ/fimuAr7dgHujXSuw+GJkn
DLcO6gd1YNuQDjksYfskys2Sd1aIQU+BazzH6yWQ/PxAddtVH/BBQoq0dTKwuwzvzSj3LtEVceWy
ImMhdsLxchTsx6wHUW32IZT+C6RV6kMRl5+OWgPvCzjPNl8irxI+BMe2tPxR9BTxVL28dzOheFJC
dOf+E9W0NEOhDBZoGUXeImsSxvGVA5H1Yc4ahzav5RGL4/78GP4Qoq/+0s0FTkeMLfhylkVzG6yI
eZfuGjX9VUpcfgFa7Ctg9pbKzd+yV4fqx9uObt5sc701AEc8iLd525/nN5HlD2VvoHjLLWG8bdpD
U4s//P8Gljk79RANUH7fbV7/RP+n+vvigkq7HwoXMhYIz7+8FiiNml16/uUSqkwMrcU7j2mPmWxO
QUqCahrC4yajXhJ5uOd9+5DBcNfVIo2Gja1ea4o95/QCqu7KgOTFJo8/lZ2R/h5als6OU6JCrw5U
pHRbRoOgmP+oObVl2NOmQcQctB8atJ2349fFjARl/WIXU7aDOijNdeaNRyi4slyJSY0S7JR1jTAM
0KocY0whStgc8hGmA8YqOdn2JgqM5eyApvvJVpCan1ZsTEG7evXYcEPoSTIj9FdVGENfKbNMdVu5
LprnSgOJK3c2aNOFUYVMFB7+m3w2On/JqUImxEmx4BCzOV4XXhDIR9/RyLsRHUqQui+GvfGJCu3P
idb6b4PM8UOd+WV8M2dKMiVCtCjq4Eknd9sKZf0CGYuLeQH26N7QaR2ow8I9okNj5RSEY/n/KSVq
aSpWxSMOdFDb+30yRBpBVTA37hoOmk27RkY3HN6fQTBm4NXOTRNnWriGivzSpw72GvG6nfZDgUvE
1q6vnwUQst/lUx0SjECC9jKbYpl7O7qGPp+g4XIKhf6rDamuHIF5QRPRA2J/BBm1l2grVsQOBcLx
RTI4aYLO1xOj4eDBIxmhhFT25CFIRk+yhcvhY6M79pstGTN7bv6AB7kYjAIDYFv5N2X3nTDFp5vs
38iim0Fj4Ahv8J1Wn7iM9v+mNJORFvwLF7HZNLPS6vAFJNt1trNN/qfB0AnkkbH1+gdk+iAbJaRv
92P2zsNj+Xguv92QwQ3HUJPSHmwrDS5U8kuNdCLvyA7Yl4/el9WCinBwGYXh1pu9DmliVxuWSiBs
l373vXPaAobNQ1JmD4yRqyB24lZ1Hytrqvd5A0pGi3Gv8lsFUKwZKFd50IaPrB/rhJa1sANwEtTm
S16k/65+zRmsnq5EIRCUo2tc2N7soDRB3WhkSJXCUOnXeBmkMjHmSOvncNNOmnRqU13cm9wMVke0
QCMtOMZ58qRtx1yPPcAHXV/uvjFPwOCrPIdRxHV6P5zs7x6lSScP+/f7x+1LfmLyCReOS0uKekRD
DLphecV9rH+D+gdPx9xY04IgxjzUnk/c60MknR4z1fA9jQDsoQAhD8niGcTd7zC1od8RE2k3LGmO
Ar4RAK4DZ86YUydwC7JhX+06i1LO5v/C4NkggyE4eSCyUy29F3Wgsi2gR5YV1UEj4f/vRtGymKL+
5CGK1wx5IiCYgEA2Bh7mAsUzcQMWuBoPL5jestRz1kJr4MDCVvBUDen2qn8eRiWsy67aKjlBAnGm
pGzgXQ5u3SyKTI+jN1wLoWrUhfSDcNZL/RJo/q0gSE2AqIaX6bwwMP5tQcFTQ/UySatxuXY8qB5w
OxNHEwYijsnq1MRzw2nYzh0DRxTq8MK6Yz0k7K7TuSjSibei7kXLGITuGj2Ht3TuCxPyNgqRtI9A
B0aww3fm1A3YwpHnFzq7xbkBU5eUt59e1jJGv/zOCxr1ecdbWx9wyc5F7AYQ/S6/wiNQBye8YIfg
HDXJ2xK5NLBkRe1vbHu+u85PQe7yXoXFyDf74ZUTD6pXZx0zeqPs9GTh0VayykwNwokoCb1JJX4/
71gry03a45AqwtSIIHLg1snH50NszBGZIrDT8U3JcQe+ychPrP+Fq9IKpF+9AY/vsg2a9DBOhUaS
FKyRXxmnhRmWzAIE6LNLIJdpZkEu4ooawZz7EiI9ll35lAssNywC23QyjzbqVKqAjMkCkyzyafci
4bftoRHfN130LUn0m6YQW0U1lyWaqC9zXlmrcwaInGP7R6nsafPQv9RdlmYTlRiKUAHMANanJa09
KURHokkCaQhzVrDU3nyTgMYZobrz8flh1uR765L5Rq117lhvk8LaEtgnuPMwAS6IxgRQtuoaN9yE
LfhhCo5F5cSc4gORBEjTnbRBj2K+51goSRsCEsv4EVhHWOR+VNphMlvqiCBR91VFYT1v6wGAx+KF
A/d+qrI7gwpiBPWQlAyWS27Ut/Y3XSx566sQxsHAIo2dWbQQqOietbfqm6lg1J5NQx7wupS8y5Cw
gCm39v6lmqC+KJxCZFuH0jB7nsu2if8Ey1W0JaEJdZbbl4s3J0Xswz62ijwIZY9DQJiaVUFCXEB2
lS3pqhZEBfK+MYVU1mhGxkhaytlGbxzcJitzto9GFSFRnKtwJ0eLpn3JipMjkZ3NYjr6+ph6aZyU
rIuIFFczVT9xx4Qcua7MpR0nqjWCzvGizLRc5MMgX72ehenojm+cLWSXDpgb7KLhVZ6bJ/l8FuFL
PiRLtaCAEv+cH42Y6Y2SZxgdMXlvhAfG1MGaFTsXGVlEDv7bGIRly/4IVtIUI0+B+vUTY9ps9XIE
Spwk2n+xEjOJ94aVRACktQ2x5kXgRlkWixb/0oXIk/+0auOjmRuhL5UKdgzL5jXcTIf7MSeY2B0+
AHFzRh1U6/yaSHhQt9FRuFrHR8iUqLb0S8E31/XM8JXWyTga1gtWoV/32/6JSElcRX9vJV0oWAV/
49gUBWH1tft41JV4VZKnqzB5sWHn9EQIVMtZ6I+IbO3EkxNdqRikgdpErnzVJC1tnnwQGJwAFQwY
/etZPWxe0OI6W3JUlCYdf0YKy6I+Zucg1I8c7trXGt/7unXBPWtiCE6i64drt9jogyX5IViSDB8h
hinQ8WnPcYoRyQKEJDLLKz+8lilw8gxLNmSN8V0pLY0VRHg+vomssd8V6kikP+iwYGl04QL6O8aH
qkik9OppcmaM+0z8a0HWVmc9m0AmQiiWcxB0goV5VvP1Olp938zAZp5kMzzat7+RZ2Kt/jdZAl8+
cqvlT64BI2xq6b2a8zHTPOxgmG0qORog6irZYgsJ59oImwuS4ZHYAG2pk2Jha6Mfr60iNhY+WJz7
ODHskjE3H8Z+9L5NGxdSpR7imLVUr5QUWmtDwN6GNqTZ4J+1yL2Pu2lzdJkhpD+HHsr+CBBOZi1T
0ocqgEWUKop1Vk5gqdU1DNG2WBxWIAGoKgH7akCyjmoCHTqsCr71tNtYoJJvt0YYDxx+1h7j3wF2
89sI54nkwUaAX3BQKb0sSe6rCgGcGfTzjyyahCp9libsh5MYIe1n+oHkRE+Li4JNwYVY4xYXRhcY
OrbR5AhMQaTwvd99PTWIvrxMC0n5uPlJ9gcrcZX5MLdPEr12ocKwsueHrRfc195OM3KAT4MqtwDn
NJ4IGdgxWW+Mwkb+urCe5BjZimaCY8HDMSQsz7eQz3UxaX71JDN04U6CC4vC+JJSeQ1HVDMyqUgk
ZylNfQiZ9HV7U7EIQX+HMzInccBFkFLXbL2o1gfDYH5OB/0+PIgHgdfcJKCskqQNxXkPGCrAzerr
71/zdwAFeHzv6zf87jy/T1Vf6AehZd50yRv7/mEVQqBlrD2dWHDvamP19gUYdo93O3aiwVOni7Z/
MOWFNcxzibDosmpDIZvc5b+DF2dojr5YDX9yp+OCANTc7mHxYJwNA0Qj9h8+m4tIpAsILrXVpL2O
D0IWB3F4ogvVx/U3s7/V4TB2PN5czINGSWVFkDJOLfqKsFKu7ArEfJrdJpWUNmfoh184we3bHDN8
1PPCMU14E9pJzMaS8TgDOa74unCya8B+IDQTy3j7K0FU8tJPR6zYsYPC6PwLth/O58JfZdTQ60CF
O6jIjS9sau7H8ywdR8TIe3ZNdBWKCrFJBfBNCZqYcQAgjjJLxvzedlA/tT/cWlng/o2QoPKl0D/d
AvgTJCSHD4+XywnMB+7g+0Nljy2fP04kP+qhQVD+oLku3w+x1oIKnA4F0T2W9R7oT6wdlbVBLjpR
fDAlw4p6knkdlR8/weC8g8UEVUIll0g83Q/7yH62J2yctp+PP9tmKNaqdoBmVYjzOQ4xTy/JPOOz
2lbGJ6uEWw+rV8DpZWftCaQcEcGpHim1Xe5v8M7wOb0yPq+8y79a1Wcq9I3k3jmRHh8RXiylWAmL
oQIyFfDYeQR61Ha1aUFURLgHH+/2D1D3ohtH9gj/e6Hd7Fgf/iS1cWN62apypQtvcmYADKnNOSPa
/mVL6wXc93Dq3bBTHxRKHQ3BmHeXjtFmy2S88Ujzyl+8pPnag3icYdQC8S2CgYoEHziyaTehmaa3
PnBM2do0A6qZk69ojD+MbibRxrJreop2Y91yZpLxEjhjkdDqKwE6nZzgrwVPps2WLqgcE0aBmUUb
E6mJgTFgEIertM4EfYQQaFyIvRdDn0aGAR8wQnWuukNR8sdO3jXaY8msZ+TQcdpeIJYflE8nrjDY
UXY0+hwAxkPk29CJme7b0Y6WM63p+DIL8JdslhXG43DiuH/TCyLYcSIyB5W3CvPGLE4jZc1tiXLL
AwvRLGrmuWVX311LTK6WgTLj94Hi8gZGOefrP8B5axNbZxYuQCE39Ef+818SIX1PoAwgt4RYZ7Zx
1Qsh8QpAMF/nFmwMOOFH34zihAbG+4Ngv7yirbxt6gy90KRbQAHGVgC8p6yC5gnA7vBVO7WwqeQu
wM4xohZPXhnAMXVYtQ0yKG1jzYAgfPO+NVF5aWOR3psc20dVVLvZLHqCJwc4HtuNMVXAEGWYr874
Jf74DC6Rvf2Ro3isIk/9K+sCWHBa4wLyQgL9ufE4PIZ9J90jLaJtxiNKnFJRsCxwazp0SzsyTnM5
zwmgK33dUSpOAoIKBs2/WI55hpRZJsKWFcmrX0N9VCRRn6oMs1Fetiwg4QB6xPdZdPxtYnFdQGmr
15v/+/Y2pEzjSLLz1d7APfgmRIbR+A6Xi1b0tNCTNF5T49Et35FWu6ek1saI20LxCEMEOiMLFDYg
MYQpdoF82uKq85T1jE6eFOMDflX5BybvFOO/pdpve9NMW44WwtIfMe/lxLgUcJWLIl00XQ2av/TO
fSktThZcQ5yVckJ9rit2fgcoVeFXVUEkblwaTbvTyIj9rffyez67lAFQaStcZCW7H+Bcb2ZqAsA8
Ej7Pt1rU8fhF1tGy4nezJ7IZG6T08/YtHve9d2DvAiWVa1+52EslcVO23G1FfGLyw2ouO9qHWN9Z
vAfhNxlyJZeGLXpoC52aSkjIdeqQxuYFoJSxoZ0H0HQGA2FFyXOLadTZRf90qGKesht+fAjmrYxO
2iYrV0dwASC79RfYgtLn2SGOOpjl5ca6DmZrXH/7bZA9b/KT920gq2KoIHmq1fhXei9qj0ERvG8F
GIzA6MSvaOuRjiqhRnYnueD9ldjue66ft/BbmxpljsRapgpaaS1yb7Vli8AMo8u7T1kTI9vi3BR6
3dOqI0TpcZ2lhlz03/xYkjuRJban3eeuWojFxajP3Xd9X4n3vlAKFP3kwD4FNCY4Lg0BY7lrVhzT
dor4VOIngeGI/1nh+cImTulFIerO+8ksKXt/r0oiMp63hVvfFZt5eUIYDZ6iyNO/INudL6qpSVC9
wgP+UVo/2h67fK4yWwog0BBHU+nuxvJN3TeF5Ah8rl+n7SIXpKv/r0AeLmiwMtitYxenzZH7kid+
QvezQaVyXZA8g93Q14WI5LZYtTKZ1jHb1Lc9YK0CJLVCd+GY3qR/pufchn/SEpMoqgTUq74S7a18
AfLSzjIkJ+9FZtiJuqIf3sRQUtusmbSdJ/OMX4KEMiSZPYamiYLT/MGKV7PXTWQb8APe9m/EF1Np
wkpiQHRUsocldG84Ej8fwxVbHR0X/ZzDTQRDxD7M+SNxhK+bU4DcQmz98A07S63os6/HO5dCtcjg
AcvBQLUgst4xVx48SUtalYt2GnhXMDFOXxwTa6Sr7RgSrjeHXx9ig7jwJ9XTuNWjpHKOhQQTHHNd
pZlG3FkoQsfpAl9RxSliXD7YhTsav1LSPSFvtimM239ZE5AAiaNkw1HrYbrnGL6vYYBtBS6je1cp
/huy3LSjhh7Qp3yKnENI0DqsXluCzYOGZIY4KD7c9IXu5CvQsjkKx+oUO211WDiUV1xxPJMUwXpK
weej724PVG1+1WH+CMOcJKVwUPGu8/RrCZ+SAfjYiP3Kxpy8cLR07PogrnqRxDhb8sgKOYCqf9rO
vpCiDU2+8MWipKOJtzjdfH9c6A9kIHqdi06CnfOEtSFnooFfiZOcdB5FxcNugEyLNuMslbd6MLyj
JhY22dARycTgMr46WxdtCxbvo3/styflhunuOaESuyUowpPuskU8zMf1ARO9g9WFN1jNpfrA9WKg
+sU/3ATdLTqPa0rZ2BdU+QUJg6yKXe91IXUtDjMPZHrBKUbefIjXDxEQ16bym8+oSOma3xgeZ0Jx
jR0FQqtVfBgMTgz/8uGfA7c73yVeAkgpy9T7JA0CJ6u6s6vB3+wKewGwZ3xL42LbXZEyIcNU651N
yH257taAU9QtU3PqXGzMjdYwRS28WZ4M3JTlC7RLAPjqlCUVdf2Dn2Z2exNIx8FVqvpoCfgQ/5wX
rRwrvmlJE6+74SXiumHbZVUcLgs/6CEaU6mxdL0LrPmptsUAZ7xakoF5+PKCgzImpUG15KkqU9Tz
bnsOt3gwqp2YDZD2oO+Hznz3nMl+ISbRf0INOmZGJaar+VqHO2hp+FMR1bESPat7Fj2cqN3b9Wgy
GKn9x0lCstRl3DydAU/L8ZiAgNqlIn4eg9v6KrJcWXsxLG+3k+/SOSMjhUlbTk6mkXbJaZMuu9/0
d2Vc2SG8Kzl4J7Q9joItp2Wzej+XWTjuxMu/B1glurxLb0zmRRZqkaVcqMufTUNxUQDLaZPySF7k
IkNnW3tQpmLAwoGM8WBhNJBqdktJ3N/j2tGPdCbzSradbZtnD2bcFjuL2b0fcHqTTzADHWLpRulr
1Wea6aSM6IWhnHwwHpc3sLAzQQTgtHIpd4c726ou9PI0pIuE9roNXxv961IVPN963z72z9pPIdOw
XTJ/0GaLffAvITU7vtp8dBlgeP5YuN1ImRJTWimwXeWHiuBjrmNhWKguWYdqtzko9UiiIdrz43I5
ay8iKOXUSKGVL7z19V9u+5/UfjIdZm219hSUgGTN2ewhgIU68JFLjPSQ75GYxMIjf6G3yGylR2rx
qxipoOLNoD9AmYuJPPKeh0kxnn0qUIgpnfL0rVO3QdZlxdqLAtBhKkDyTMEGTAeikzWOpYhkHmrT
LxEBKapLb8TRrhUuz5KJ80dhOQyMA+F+hzRok/Raul3MGfMSbwMkkx57Dt9GOKdu6gZLk/yyki0h
4KjknW5svZQTK0E6eOC6C4DG8Fe2TRx/xak+rVGkMl12kwEtcUxtpmYh8XWmaE7iiaER2k6fN4KW
ZSQ87hGGjGRjmKJ4KbmiWVgduFwo/hrVPTS9GlByLwzqCizlsLRAEb2+V8IsIWAxPX7eZQgoZehj
8Iw5zWO5GWGnvZ/aqPugWI7y9EExj6XRyF/oFo+Il3roqE4youdb1+YSHSmrlFbfOovMIS/1iioU
UFlD+GENKLNtF/SMBsSzsgCR7Sa1GnQOo6Zk7JQeAU2ehziWs8fpacY1tZ7MF4ZJIcn6yxd5NvoX
SYp5JI+l+JT/DORBIVmgSzS4brD1qUJC49lussJZXoSR9GE2wdHgjBrPEHid2Bb4NBZ3+j6ZmgO4
9bdf5cxnBFY3t0xUrCialYWHb2lRA2VzQ1lpROcXKqGh7KxcQhWUUyMXlNrcw4lX4qU8hGYwOmyQ
7fyByChw519Nhng1CQj1PJ36WjBrqfrSjd+ZBeLFNVa7Kfdocs4gS+dSYX/FxWHzbhhZ6ElcKpZH
tEIR1irK35hUbRNwxgeFYuD4r9kL49G17uG5xtKDF/SX8JE84RVlyomk+DxS6cr68LRfetySKjPL
GPTdWix1QpBkFWCysZQr3eNENSwsbMEWMpBCGJP7OXHz/zeHvOp+nDA6lV9cQAun6hw8LBP8d2uy
3dVYSBTks9YHmbdmMB1ihwde+N9AlnLxeeIFMGsq5GDE95t/vTjrKvMPqeNx1zd4ktRzICjDoZ0D
djRfdLUGZA9fC6MsftmjytTrhhap9FzTUfAbS2zHbmaOa14Hr50lPuIQ0vLehplDjPBuFXUP3KNb
RJLIka3xKTdZJrcE0ODJ8FGAYCK4zB247sY2p0gZ91P/T48c5ty+8J/PVwgvOS1uHwy42kvwnozJ
MlxqK6ebfxIudjJP2S0fig88GPE2a730mcA1gfBFCoxx0cMl6gC/C2FhxLnBZOc3poKct62o/zcj
bixF47PIAyB6y8KJ1ELn5ITkg6xIiDpy6olIyXpa1LPQuIh5TeyMnJElSQXiSPQIhErWwlOg+hv6
IzYO9bxQbrua33WB01i7S5VnLVwt66TFip9woizrB4JPW1lDj1P19/+E7xyaukYC2k51sqq8Xr31
S3AqxU3NeCgJs6ObHMOgqUiXOIhAI/ItxN7k1yZDhjBeZoJE5GAAuVlejV7aZRVinQ0OJDOcC9Mj
HX5m06I0BqWvVYm5T/IIqhY1ZTzfFQ2tVmMkyXT7FMwccpLKtMxuT32iAr+qm4I8YDQ43l+ydFu2
7rD4Y/0UMbYdmaXE7GNlUJ3Sbtrm3jHALU76lX6IGxqDris4+t6RiRJGIgWqb4zNO3XfnsD8gJaJ
tIt6Saa1mUtHtHZhc4KiMDlhSZP72MKjmW3DK3ebAqWY+0iAOU8q5DYex7upKlt2XORXQbcA9zMy
E/OBA3FTYbJ3s6CGl5ymIOiIKbLKrApTaum32ubkivTvPVBbeE75xdmRQ5INJaFiG0PY7xoMvf3Y
C4fvkGTSAeFCF18yCtj1XXg2/+irMpEfbfzFA1k5G22a4LcpD5ysbwUVQS8MX5rX/xc3QEPnJJ5i
Au2qZyx4IydDPAxYJn4oQ3msbM/sY5cYZYUEUPycrEajSgjXWsQ9fF37kg/CyyURp0VmvGSk0Bsf
QrTUt1MsPn33X1EzCRHQDQraTL+tE6VtL6Ae2nxlQ8DRemadpVW6jozLE23MwlWCO7p4xkze6NL6
Ql0tdoAh2JHV7xPAfGZpb/z89zWSKnQmiV1b0zBVkKbtimwc8Wpfvxko4Ct04MiF+hWTxAgDRREu
YITs4F5Z6CwwyCrTZIQ4dum7PM5b98OA48W+k4+C3QiBn2kUE/y1eXS0mVMBO+YebvG7TStjQVqP
/8cFqy3tuAWEaYflxunSaaHH27NFTk0uXSKtLYo/HXZraeDcSawc1UuN3isQOmq0k2fwVFaC/FLl
vE25XdKZgpGvyMHQt8BqUgNGLHEJkPBuWW9EN5uEg63VtZh1Se5kzTrkoFa76rjdQoxFBDvZoEXX
hJ/kQTcEn3rusQ5vfsycO4FVnAWP7I+an8A7DxC7FHHwrxrDmjsQBsjKCMcKc+VMvnVzMIezO9jQ
hGxjF5xIbtcHaG5gjX2x3uHOMTDmpGcSYceMH3yw3t30bp6s8pkmAVYPRNWOPh9fSoGLuYJmNNyH
LszEijvjnVJUaSqC9gb9qZCzOAF4LZVt+2tPwqyPm/+PAabndQsRzgqFCm7iMSVy4wmKvk5W6CAB
1vNCc2wlTSTXmdv5T0KoAkVtltXi70vaXpqe0uu9c/9s4OmSq0MPbk+ClK14BBKotXiZ2688Q0w7
MMYE3oeAjTRprzLjCiXZ6zIQsAG4fibADCoEa603siK4AYMD1EFquiGu3A61mDSuWNRMhCxnH4nI
AtGD/8OC3W59Fkhbvs5uJHmOMD5Y4nOxh6XlZthnbPHokaFjlRES1Wvl21uoGxF8xoQRQfdKO6W/
deszWxeyP+BCelP4qeO2dUX88817uOiFubeB/8QTFxdgusbvDKsbtxcXS3iZSRjFLgSc3POiQSGX
qvtkO9XnrYZ0v5F2ODZzQUns1yaugLERO3u4AvJlFByokLM78daH3Kj8RnVfzdwSkp4uIcyj745b
szmaUlwH47xF8thkNfB1Wz5fFdQv+dm3SyZylEmrsAc/eL4HxFV7/XHDP2Z/CaZKN9SAaF60Ibn0
gj1xbmXMyJGTy16juf4MIbxEKbLsZwn9HI3JxI1LwXRMXnmkLZ/AYdjTWB9/Z+tVQDYHkiEQ6hzW
6ROg22wcDVCZAoVLLY3HPjFOsQ2ytSCbViuD8GOwsKNVzKMu5JqYpnQFMYvW2FbSgSqHqbSSz4Ln
VSGIK0JuZrOFKO36HKU16Lh/Nfz3ov5OutsSxM5VQHkaESVvF8hpUkXrcaKYfNCe7s9c6jEEEKKi
O+HoZrObAIty2mFc6cvth4xdbSAjMlAIsUS6kmOpgH1hvup5jVlKAhuJqGch/0rxNvxjM+w4xNGE
GDDpV6/NZ0vkGfBt3OCBXPtCCNiTto7nmvolcZu2ksN3e0cSR+qxgSMKbfwvaF+63sJ2BhPrK9Sb
c7gUoFmR653T84tsP3GmUyltOG2nBLJIOlGifzjzyRbdma5j96d3EJyMwPNp5/M2icsiM1fYQHn3
wxwASlSN18+zHCttU80VGnZDpnqFWNS9IeS4HJUGOyRBE03WM0vIcVCGdFYJuPV954pJORGK3/EZ
ZfXNG6QmpocFZ41EA9MsNVUWnkJZqoWgWWM0PIfe0wE4jg/x2w/LV+ud7HmccdR+3V1w3iTgZSK6
sUJr0urfTIuPMqoGH49uJPuBJb/YtnFkQDd44iAVjHeOurS5g41N1FK//TzlDLlCKAe+4pTQZx90
LMSCL6yc6/t4Asl9FaDZwv9DDFkAbksL2gbMFOAcVtAx/8R+STMOsI1XO8Wnej19b8MplNhx6vCj
DfwmRA2AjJtBs/GqJISFSAxku9F92JprrOhf6hC0iMtIPUsn8CjOXE5smd1p8zJVJ3tX3PIPlAhA
JWPBdGqOU/yN2XhEf902BBMpYuOvLTAWQlEgzW1acj55agUDMMNZGhNn/Lrkdm0BBwp7ecTc5tWH
jczDdYHR65gEzRSsCHGIspuxYyuI8TvY68UIw+HxjHiGBQcyf3s9fY/nxxNYTR2/Zd62zseVYBTe
ozNDIIg36K0j5PMfrow2echCqlfUOMjs0W5e18AGgKo/iEcjW1nswCUZEViG0cJcDuMh/eRftB9r
SG1AdWWkCaGIWOYHeoj2UlCAaRzDQ0we6CLaODpJprd7vC6+IBF2k8qREpvlQwu90ol/Y8hmMRM/
/RzCVYLXk9upugzT+O/UKOrnA/rYAJ1paz6PD45RXG7NC3Ry8TsfLO1+80a2p0uDq9ZSfDdSGbw1
4KNPXoFrTIoBSINY/Xpz1CYhS5GYAbEguUuvktRjHk0K4z0lIBl5TkIFFnXH7mWcpy1tMJs8IWQu
93Nup5KZcvj/8wMc+kIpuOx1VcpAEEW6pYeKlY7A1KQQrBlJB/SDq6bHgL7e+kxVdGy+aX9iRL1r
emS8etU22uQ2wlMpuiMdalwxEOpnKefC4ncNpF2+A9GGUS8vSk6L+jHUAXdeuTtPBit241H+yjk+
qdMmhxuziTopxjIDLNDUkP31SkwuDpIhg7sNP/HXPCY0BZQcpf6ZN3Cqv++JQJ1o9TNyOqgF5iPA
cNRjfccQGNGftWMTGBFqYJY5zItSqXn/oXD2gWIFrWGITaWrLApzfnAC/ihnf3131972z/mliBRR
MQ9mgBS+fogCS268ER5kLNnEnMMYUj4YMRY7fDe1s9ParvmGa+alHN3hJbidWOqXYwf58pO84iT0
Oly7i+unBqHvyMAyt3GD77iPBYE5GXa0xRrvSOBXMQ+T3Aw1jV/0uIkNuZOydGl64cHIG12UF2ku
O5PtfGBWqp+V11qRFTyPYsmR7p9V/6PNJKn3EU0K0V9Ul0FAvvuryY6dN0KaleSrvKm+sqfn7deK
wKRfftEZY2Qo7BAhilY672mvRi5SPk3hIlz+DxAmWu2NkPm7aj4g4A7xbAnlZ7piB3Z7m9hAAVlR
lbpUBhlNIVVFaugGWh3/lRcT9k7o3kCRleXFgTZdDw7lqAnhaFQ+wy7lj4Px1FDSfxL+xw8JhpfJ
g9CnozrH5L+D6LPtD3qZ+/R12ArRvHSvZ/pmaBMbJVFkj+vHEHNDyYcSJJ5ZwKIUX7eCoRecCith
VlyX3iR4UEcCzGqIrKOZA8mjFgyDXwm2YZ3jRmWT+B1uuHxFc3KKB4eALo4ZUyWsSugTfXVSh2MN
YKq4Ekq/fBVZF70I5+ZBZnYzyYSa6Kc0LM2Lul9erCRacD5mONI1kbh3Vh3AqhXsoiSLac72yglB
mK6TKenyQOlI6qiKvGNEmoTRZUR1Iv7pZUW0tHraZNqKAZPoIZDXOiJtquflOluzw/qeYBDjEkU/
LHM4OXUmLz7Lii2MqGH4N5y4B66Z4utRnQ0CQ0Ewgyot9AuybbnuQsWcgCArqH7SulfppN+KvJJ6
E6zukUM1q3XZL6OrMUECy0iqbOKcF/EoTzlxhJgvqA9kN/2MNqdKFFlqjjvCPhz3jUqCzNu8FCkX
IKySC2PA092XTX8Slo/kAu97UEUw8o29xacM2yD43smC6p0obQGt4BNqI4y61cBeiX38i5W5aTfx
3PNdhid/eGZ507ieI/vPHZ2u4udHqNuT+ocPnkQ+w+9yDU0u/JOUW6RHkgnTqbtPu6MbynY1cnJ8
GJgDBb89Fvw6oJtrFxMx7F4XIdy83uQazH7PFo9ovBYrAY8TLEPd0iky62q8vVK+ZTNjF1ieD3Zx
7Pzq4ySGcrftxuQbsQFeX5g5CKG1EtjCehcxzfnDGLet09giYJQSZgzgucFhaTwdjtCX6FohLZVl
W0nfTk6CvFAT5Il4cwd3Wlv1F5d4AEnuwC6xQ1my8bWtZRV4HjDFv3j4+l7iKEtqjuR88zCdOniZ
jMZD6JZ76FSbMS/la5/dI0Y1Pt53xYhhkrhAzC0twMrFqG5VS6SNvelFQtEfIYRf1FX2jnL/0Kee
OYgLyDHek3YJs/CbQgcPB0iFXNKtuXbxlSJKbg6UxkwTCLal0om1hHB6Z2qoPXxpzaXGJzW2O1lK
W1my2lB84ktaOGMJEnkVHMwFODHvyaIzzBN1ElsOmwNbEsJsSg4983QakZM3zyg4kru9e2Phnz49
6QCCwhgSq2+XEJ4abqbQJfcDatb3kxjVpxujRnQaBKZpkZErIzGhR5WlNJuT2L8t2K967y5aDAxr
MpmPunHLmAnW1ozS2GexQJlownW6mdaGaRmsHDgstG1BeP1MmYAyg1y0gvTz+4ZkAK8b6oUp3Reh
JWLmbla0+432FHe2KZYOQQUIPRA66eZDMgMjKJSU1LLU74uY5rSF/q6QaG8cUwUns5HmY1zG4hsD
evVCkTh2UyiZYi+UWuIew89ox45pKVHrWNCYz39f7Rv0GMWHajvYzHGtyz9Wtmxa7CM91Yvu8ojP
rkAVCeEgzk290Exyem1oYOuT5vOd6qEs2YL629amaDnuJpyhGCft5r+xYBfvTrrlsqXhldeNaLss
q3YgB20+I8UJH5KD7miedw9qmkfVS3z/ec2BUuSxfgttB/v1uoistEdcLwClz4CJwanO6xqPTB1Y
9suJMGoEeqiZ1La4Pmiu/Cf5IKBebVncHONhmUFtRbOCXZ6gD1bpzyrK5K6eUIgaEl5oxGR9h7HI
wNChUn5hMh88XltDim++zIDH/EQllUxIsO2hifXQNpUg8GheU+wvJKOisds1zdnD+a4yMSZyBx+s
rHwojDdC/bFoxXu1y2S2/XeAGcH6OvfCLKEVyKUCz1HJvZQWIrXAwIKQTQ2/vAgAxXzY1WILqsWJ
mA4QLRBKADn+vpBkOA6Dvsg+6KLyuk5wnn3vRb01nBQNDV6tnxxQlivuo9o6GkFPyWNVUPjLxJOI
y7S6dqkAhuHxzGqu/4iQZm1EMRBsklroNXB17UQD3+ADkoGC3Lbeg1xOyhsqlMZjgivzAmm0VFqV
c0pqf+Q1MkqU3QKpGWRWFmVcppO+H5Egfm0T24oityQwDDfvtwNcITq3B++ZeAMHzKwhjKSK9I8n
sQXqArxgUfO+NJuw1vL/0KMToU9v2+tQ5e8W8L7xUUeS3qO5PuE3pAjEZgpjA7PNMSP9OiHTI8go
r6+vVXKDVufsFafnbKxUFq+9luEI9SbUl9eBq27qfIix4pD48RbkySvcBOtgLM4cmc5rs4b8/GNU
2ljPbmNcW2Bo3g7iH/GYQUAQ9nfuGWJuz0L2vNNxZXlcEKZF0GWzZD/t8sSZ1b5yYdVhLsFf4xo+
isKPBNCtZkyBrhC+XKRJYPQ1a5jHOEKeS3+nBIhGb7Ri+cF57MGdKb6Z6sHb6SsAL8x44BmNfwKA
UEfoovnUWWYCuUGTua9yvpkituB090MGpLkeKBjWocInPL0hvnxz2iK5FQxrM1Wvqz/LMQlvSoEz
mvKoGDwJ2c6fRvzPix41Hmmnef3lsXwSLpgswEeHR79BbDT5wLrGLi6mAYzTXMwv/6sJ6HgYu52k
IbMpC/asJfUmwD+MmDuIh30e/LnK65Pg3ECC5PXLIfmDzzuJ2xB8+UGCx/y3Rc9M1hFdpZfz2ZRx
K92MNAfkmVDeByi609Ehm/1XlQwLuSd3XcEV4bRQ/v9SFMFn1yeWJcjKFWuSy2V56Jtz3+gXgUHy
n9Fc0eCesPTlc2nKC11QLnMRhUngiLWmqAyeh1ur26v045RLuXs6XAYv6iM+lPdwBcnSy2GBAjr5
z8nskGFGFiEv6LGJl6D5ui/6dQgaBiAMuomhDCfB/ejE7dkADD1H6IHUWgnKHgYN+ssAhAm8kqn6
YvdluiXxFZ7BMnaHu7l+wQ5MBvUGcisx3RqraW0A3TWyhauVYihfw6JeLCCHw4lWlkAccd8z1+7h
0str+bVVOSENF4D/0bC9Lw5H13ANj5lyHXhuOMidl+ldbyeSmWtaEQnH5EI8s8SbMeWDQLmDX660
c1luiXWcDLXDm6vuwXT5XOnp3iP8WWJvF8lYd2VNQ/z+bNeJZqGPn3jGgtX+zz2K8tKz98YDGAjv
TfJs76CH6xXr36NSO186mN8gCtZjnzAT8rKZdwT4HNUJcVhA+cxgcIDqgtb0cy5vSAeRAKx3mEzZ
VB81cmvCI0xLKuGu08wy+bYsUJ3XEFs096mm6lc+qHF+i5kdzRGfKdhox9MnajLaio3B/ocWeVDT
M4XMfmR0F5+52blh4tENr64rWOZ/pObRxnJ21CqPNxx1PHafUXP4sKDQij8r7bRX0g7mrrt0XNYA
1EQHI77wlKrnNBs0VCxGcezNrYjBvQgpfwkVQKf+9IzD6iy26bi5iAmcPCxx8LacY3ZNyv2t9Kpo
IOBiJ/Ll01pfkky+AP5F4CWqWxcACyK/GDTVTbVto/J4NA8UNKn2JWf/fnO91VvEMJPZSCNGth5o
KI7IMeLANz0/YboWwlPwlu/vISdIHny1xmbNMMujpmE2bZY7ZxcaIiyx/DtlF54Ndg/Fvfuv/Qd6
fK2yuH/rTspX/8XI0oZY/MeHbMNpJm70/VWrcD1Zc8xoIgkxx5dRUZcFFa5IlqDqtUCfP1gLOpiE
xU6xm7edbRez2Yj5OxGXEL0/E+fKJj3i7vA+ZMit4mFYZQ9T50u2TFSLRYawnfzy37RQFOCYU25b
hmkSczgZVVkMulgIiNHd2bt0mK7yks5hr/PexJxuhXVSGEPS4RbTJg1HeTSpn1BVsX+iDhj6uBRs
8RPmviOOOW5h5Cm5PKGEprs07s+J3kCeMjT54lINyECSZMcFMxiV3NEZyXRq9cp0rB/h4nPFRZBf
1LzysMj9eUfB87urVu2DWpHH4eo921THC66HVFD8gekhc41edkw6geXUyjuqC/mJuTneiPP6rriF
eLYans2KEmn8UAvZYU5QuO5mFcqaCZ+fQAZnuHBZyVdlTsqxdFXNtPoXnhvrNWACvhotSGIU0AeS
mycIZ+/4G6zUK9AGckVFhedJceSp3bgM1A2G5lYNKkDXJEfgitUIl5HkzMVa1vjtfU3oXsvu5Wfn
LjPUqPrx+xQkSUTtcB5ut4yWcpB2zaRRpoxINpqe4Flxx9yaf/6UAdLCngI0S/GoE8Y35cpXHghC
hzIr+5kOYIBnqHWxLuGtAan+0YyerI3WeV5Wkim7DYWqzoGPDMhF2SYAv92pjp7OLpLhCuM4GA2L
nOUEL6q4jha5njGdrML0oRb5UC6hQQdTBwF2viXAmG25SsNXvglk3Ilwojq6C/Taz/ThCUoBa48b
fXhr39OVACswbpq7q5Y3tAkD0NGckA9mRbUOJ3ClR5YtRX87DcyOpMuF75xef2f4GNv/ORX474B7
X5zP7ngo3CP27SSfU7Q29ffcki2jQiFZZjr0lEHRqInOszxp8K+sJlkdmTOwetC3+ABmH/W04yca
iRJxmfCIK4Ev4tvw42XSoZf4cR5vd0VBBi6a7KYu0DmffJxo0m5ibWenbmALtvxu9H5zYM/Qas+k
XQEJE6lxLJjHcVpZX3Bv0lH5y2QgkKpi8FOAMdsxJrnMXbskX88MZd6t0XQHSkEmLGs0X6ztjirn
TDfGiWjeDe1qH6a4d6mE8Uh4ikfi6SYbUM8DC+SXQ2jqGNgq3fbfgMHxYAwod31Ovr/Cn4rRRId1
DLv8w83d5+ynst+B69UN9ly8gnde3hUURK+vbKo2ShQFlcfU2jbCzxIrf+TRtp8oE1gRtH1icWSe
eUAl3xUUmmnWJeA3eIlHstdGu61J8Ll8ASnBcBY0AMSaDLQiP3TDKa8ysP9xq0AFNayEJsYDUMe6
kzGHse1BuWiq3V/rl4V9aebWw4Kd4aKxF/hik8/KTqWNpU5ldKuMJhug2Tn62GKKVI6NWqedafK2
xYi85iDKdkAUaUN44O13pUWNHM5RpYzhgxzTHadJi6FRLDjnepHC3Xgd5jFgnd/TIBvbi2mujCh/
qE3wtPikvNQ8MuBSDoo5GrUxg6uGCqEoVB35FqFadLuQVwHonxMCJYhVVAoJYGGZgtB5KHQvq9ZZ
3MOAmE4CtzJsQErGn4Kvkq/r1+YHSj8NxwkcmQOSpJRpGimp88outxu3b68PjlrhyOD0v5AMGXCM
aWuHsW2MLFx1gxK35LBOSMjhfW1/xYmK6OhhBhaakf8XKedpDXD/rxpNM/P6RD33j16yxDANWiAK
De4lopwZlgkfbklYW8l6Dq/ktWY1MA6BZOK9mAZTfeGkzki8stBbCQ/rL2J6y2EYlFiFtzrWh6ko
Y7pNygS2KS5NV/+iPow1CQq19k4KOclw4DXXoIWXtR/MBtRkNkrNU4CTSGRCH7jM8OBo9GlMIlw3
2i9XMt41zCjY5E/agZ6ecquFikWk2lpe6Dj4YMaIg1hZJVoB6IX/roSZMRepMr5fVpJGMTE1viqA
GI5Wrt+47JzbwW15Vh5BNRFOpqZZDoB6eMTdphdMmnuwxlYd76RPe4siLTh86ZDjiK6bRVzyDCqK
U/7f0ted3BuabzynSYzGSVEnWdCxtA/Ixx4nAI1O/OVwXcEPBbWlWHIdQoPBwALCs9gG1qKMuiIC
k6r+Iy9xq1AwxpcsUmXT6ilqjbbe1yEJ3hk7yWbya8hS8cVfqFXyJS8UQhIxWvvlS+IJTmPOWyud
J+T3pkG9bd5NZ03T3p4PVFES/qAMFDzUtwQZ4pOPzeyHnCr6zoWvG9UmpeqGrKKleGsej170kwUW
QiwPK55e3iwNFz/ns01MBXUKt+dpclFCqVAVqcfYOz0xVlzHv4bqwtLhU+OcT9ehUXXLVV9Dxq8a
Ra9R09Y/F7bASUhKfok4mnFCpIWkVaenA3BAQzxOFahh7yqaYTHK9k4b0NiK3m1VU57Gh3LWDk36
/IyWX0ytCc7xTh8ljsOBMMMyp/86xLRUAtDfD3ISiR2dlZl4dp22a0EP5VgxiLW130RWkYLXYfDN
avBOjwOWzpSvWur74QwhXujjwddDtd0i5TIFuK9X+FbPsHQ2kwNdAZ7i9yTcIOYVtJpObe4Iv7DB
25wu9dwR5DM93GfXTtOkKEGAZ41Hxay1EwGBBg6EaQKa5wMYYbjYIDHh/pbS5RCXdWWaOOD8P/Yq
5IwzucESNDfHYjyJi4M4T6zw37HMC/RZu+wWCa89saPdu0Khmz8QYm/vVSRIAtD0buxk8g+rbKU6
vwf73Dmkf0eMAZ5fKeRmFlNaw6Ut5o1umNd1+wdSWJ0789m2qp/XaqkpiwqJmPdNpOujoBpW6XHt
R2tAy4da6oa0xzBwdbL9RBTxA/cIGZd/9dRAwp/+jgXCrs7hmxTaYYCBNLGavrdmBHrtCjd9oVZP
CU9kHkUeY6bQcwKr5NuZ6pcwVH01WMZ9/6BHsojfpayWklbn4ER0NPgSboYprPI4854PIPpF9wJb
sLGUVCsWrvXhKQ8Us6HGC/X0oWUACgRbULZQhjU/qZ1rlxpCI5PK+0peXP3U/1TwauQ3bjicScYr
Ofi5OtEf9jkZgXmcFI7G91DGlrB9CZNj3ZIsB6BupyFwrE8srOx+6QJYygfRza86KkmqyzZ5Vlcy
1vUz2g8oxzaS53GhvF1hFHiMc7ZjfH9XZCmiqdWWyqCPrIzl6z+9/ueTOfgt1AsdCKo/9FjvltoZ
g+I0hKr6W9Wi8PMq1cVurAeDpO6bqDj+Q70f3TaCAgzS4vIrpVHg7OaeXjhpT/x3Rm2ssmnO8rsn
C9gKLOiuBq8UpIW7uraTAPtI4OZ0VHDDPUbNDLTSXAQYA1eiMDPPQKFir8jzNknU2ttoxGxZBH2o
BKyeYmVQtSN5kylf8g9W3E8WSO6N59Is0ZfRzKMihfB6vB8Vo0wLNnd5AdV4sZuhJx/GgwHqbfxg
p65wgpWfeuOqL84VqhgMJOvIMfprDjlpsjJqxV1SIk4BCisz+e/S4M7Z7HYXQ4BM4XEjUZYW8d10
Ome0vk1Q1QCvahfrWE53XaWznbJhvLuRwTylPdbsth6mnFCGcIQhZTzq1WRJAALeHqt8uX/sIfBd
CRDNVbRxCctOD7gLzpxpB9vGrqQqMIzfGRvU4jR2GTs/AtUipmdlA8/iF7Z7XM/KePRBQDEK05c5
rOCS4zNE9kXhuNJ35uz6vM2kbxMcd0O30/misYn93mHJHTuCrZuNfP/ojG0pQeyMS/kt6sBZVx4W
yta/r6xMm3W2SZT82Wmk51pVFd7h/LgaNS82EPI/p8VH23A5McO3eUwhlB9IBaORbjCFKE1ML72+
m1WWkTC7m88hBB78HrnIt+fGIhsce4DEK7x8Mscb+76wNzbNmYSofT7BxU6JrTnW9TOiHP94WxAJ
tX45ijNekQj73hs8tVaOz2SXoAZ8P3BBplXlX/SpfxoqiqCSHCbYsjq0MatWivSSX5X2ksesvuuT
bDA8Mhm4xMB/M54UQh386SGg8ko7kIaFGDN/lURF5j0C8fh1je2eL0oB6Afqg0sjlUYG3e/Y0Rnh
qqdeILQEewlxWO4nOqL1J+hSaDgx0iKXtWrLZN9yjTej7VA4X7rFXH90/ybpxvfI3p1WwISu4ehy
2oKwlSsqvHgKwV+VoQFrI/FjJRhrMM8YpllWJ6anOqr4rdYwX1W6bhGpZML2lMpVQT/TvumfEgES
C0q4TXYYiOBgJbrlMMYLaGkGRveyljCOszacdGBIN215p/027afc1mNhw1LT1Ip9MeO5OPMxCcUq
pNVpGqMRaWTSjgRUsXDTNJHB04/icOypEgbYijlVRk/uQMdLusFeHiq0Udb+EYXKAFppbLSOxDZJ
tFE6IvP4Sq0ef3SMuGBlg7MDKg/Q7uFTr4ulDDaM7/KiIbHj1iZrqjwC3PCbnPjP0oXtAYdVgr7l
i5QlgN0Cp0Q2FYsxD3d+1PXbCJT0Xq4MLL/y32h0jX6FYx8InycIk/269EVIRYCUSjkDLAilJOy5
tJzimpbelE1J9BX79TmrD3S4tHijwDEXyjr3IiBXrjV2FeBF5CYa7oy2k1rKvgP/BPz3QrN05ylJ
UQRp1oyGVtBI+mHRUHAJpxqIr4awkohkR9nRxw3Bolb49vn4t+srSc1sNj+tFKPnnz8XUEhqPvND
8TN/CBKiEa5G9OVszxdp/ubjjfTRLHJtO6Wq66BDUoBMCsc6Z6QWLwLtddHEMDWTyvLCQTiNoWhp
fANjw6zCDQvWFpcTFTRgwQTesVx8TkBAon3Otox0L2WcBTjOG9kisGIrMhmXzB4WFbXnnPOLG6Jd
BCCdiE1Lqp4W1wA6TMMDktgAgn4vQCOYsr3nECVUBhjAMoOEnQrGM0noWXlaZ7zY0SmEWIUV2vqy
uGNB1DEByOOWQb2KTa84aVLjqiI3rMfXy4exBKUsrVWXNhnL2KQy/aeaHsv/6xMkMcCTBy7IB525
TYVH7sWKj+bvxWOiVnZVtfQeavQnMOfDuNTsERUZ7HgGc/jTRaet5sIg+NGB2gitWN6HLnVfh+wl
1wAxankQdU3TUd3sIrRDD1mwcDzO1fapQTGh3kBD40++ioQ9QoQb2bxlw60lnqzi6bjTdLB3nggb
sfVCoJ9YKzKC19f3PUIC2Pcu5R7EDBgIpVGzBjcXFQpjluX2SyABfJZE5TL45zqQGvZUbXDBKAMz
rnczsTiMdAHu62H4aMNggi1Puizc/T4trk/8U7MUyODfNUMEs7bxpCwhpJ/2yodSxSp10emCUVLD
p3v6vnbMLXxfW8m3FjfF6pMiteI/jpbYBsrWCDj0GUhACtqeKAu21AzIi64P/UAMaVXm7b6a5tjJ
xRoA/9iu5GMP0HbpfGKrU5SQMwk5WbCSqFZEO3fHJM3CAyoklCSSdDvs5iqmLr4rZTLYUsUDuY3o
ELiVKtsH1Hlk/BfP9Y/fRM9mMd/XzgkVjGc9sdPwW6WNTsQkpnlHqbsugeZxhOZ3WlLhZO/rJCuA
fImlLPNl7IfM8CIJ83lEWGmWem0qq4y8AC2yvcO/cidjBPqInGj46kAiHvED72J8VXT7vQF+x4uv
4WVB21p6Bp50QB86dkALUfNItfS4uvEEBgxQrstduz1sVLUmKzbTGiIgSwniMcyNAzDMhAWnaZod
xTS6dP4a4RhyruBasALx5LuFrN1j25q9LUjB84KJdVTil60CYH0ImHiG/IaZysrkWoILCzzFlZ19
UX8YPn58YJlgGT16ZUq6ocDHkyD+wGb0VS4Zh4J4rfIX1Zk7NLL2bJWUlTTHBVlQtYegyCuZfQzk
y2zqQE6iPWzQfMTkP9uWfuEB0nmH1oXVfdxLo9WM/8cibjnvhKzFmZ5tU6ABk/sgASowWhAdIX7H
Ky6H9hoOv2ECd7vsXzARQ2a+kd1aY/ELjRn0Bfur5Z8yuATnfoaCbJKbBmx5DTxCERDlHgnVCKDG
2AEt7vSb7P60vnRvX1jB3Yw6HOFRd5NQXbivNGrPVyHF8wFk8W2mjmAFfP8PlA2LWZDuEJH2n8kY
HsoiYY4A5WyO54cUDf18QMhvzHhcJL9UIyhhxOV1keCjL2ApNbLwwzDCDmnEKqt6U9Uu9GgKSkT/
Rl7LzKVwd4OqlFHHE+pyyLH9/Qa7kR9RPVTD3/9eFJeSiaPNG3SiBVmGF+wdt7abUwjjhE/HNNfI
WKfXvYTKvRCby66YDWXjzCD/t0CwjvKyjtdyH6UxxCrVpxurOq1f5tUASLZT5+bTpkA4GLKufa3E
UWszz/3exVTGc3uNO2Oi0ip8bHJDAU55eF1I1bdVKuaVNlHuwRduJOO753mCps5j2P4ZXlhVDNGl
zC7NyvnVmmsrNhlDct/UJ0b6J8UZDTReekg2BheSFN3GcEQ6/NBcWkiP2bI31vCWh9vvkq0kJD0x
cg2c6reSuHf1h0VrWV/MRM1CBbsozI5QWUW5GywZ/Mc99cSnOxIBkaJk4l7Jv+jsnZ9oMH7xZgXP
u0CPtQoRexoP30kJs5+Y1kuO8LkvFrJVN7LV61LSt2pFQsd6OXBEFpGep2xt5WB9wJzS9bEXdstK
A//XpPQFnh+ulq8vCeeMH5cmr0OxONc9b+KdLIESzpZK2IZhrbJapykpoWR3f6wRcGXZ7qdH3iF1
6bsdgQ73UVQuxRl1T8UeQhoP5SMvUfNB7feqAb/hM16CfZuPJu3ZZWHg/32+h9wqhkbO5G+MIS20
V1TAXiy6kpqz0zmCJd76Jl5l+NGt5ejLmNgKcOLJJ7KehV5wmivc8VRpH4fN0BEXaGg5y9mC2Kcf
tDIbNwXvEdPRXS6HTEu2ldps5HqgBM/L2SQEQQ2NL0Aov7HOg9kCLYshLR84irBRk8G88qlDtd/F
csaD4NifYFtdDo+rKlwpu1rnExJCobcDErNv3lXaQRb0dH68uYX+VJJU+IrVx8Qu555qrZdslgkr
s7mDeKyqrz2ZDc6pZ4nIBMAfPYc+eAWCxlf5ZdqybcYuIVfUC+AQr+E4sDANnD2J/nOTtFJiNH41
Fkavz78IFKU5KjWelAm3956VXSjss6yI0tUdeXEiMyIrpg940nGQ6gCiie4tp9QRtGKwqCewe9/5
FKWLPxU1b2kwxxJ8/i+ankLOJPIbdT/b3+fTvaRppb1DpsLD2epDagqodXzmX4ylA70ySHe5G8KW
2T4mLh3qYz+rKtuh06NyoJDPD7NYkydCIdt80nd21QjjVzQq8eNkDuQUHgldmpg69/JqIFKjwbc0
x16j58bFMYgn2lKbo2WV+ej/fcQwIyjxp4NbxmqfaxFC8jPrLf7C2Ve8WLmZV74e6cGnMYJ5uiHt
+ttZ/xd3JGdtAHupxhm6MQ95XR77Lw7u6XkN3k4cBmDcM6G5Vxi+2y8GCttlnE27PWT8WqCcAEWg
snthgqkY+evZtcn9W++AFM3vI509AliwFYbdWdLF3FsREfK2nBDQWPKy+rtyOndKkQzOwIDBgyWg
y4Dc/o3547msUol6YctWiMzIIt+6uEc6e/ISdEAh0HAXQK10hBKMnm/itIZ8mWjb633QBR6zY6VX
wkMPjL29MsBjXXidUQwV0432otAdwrSSQ3qYarOEPunVcerDh1+wCFDWK+Nz97fthpfvabpsnyC0
TloG8QkUhl3QOYVUA80H4n4wcmPXSRgveU+kUZQXwW8rZrl6zEcYJfa2BkEiVA47WCt6uopD9z7s
p3xbdnRI3bR4UhzdEypj9YYrN/nwUDAryvwdIsOWJCzX1xhnGvQJPr0yhWz6ikS+R3HUO/YnK6td
aoDYVO1Z+LsfgjupPhp8ZR28k6jyIEspVBEklRKVub745BaafdgeofrIUOrjAUwLLfXCIgVJ7KU2
WaGkFBXnUGW+fcArTIwx1v5wROM/o6o3P7vGuQT1Q8wkbuIZw6K4qdr+yAEpJHFpmOgui7HzPVvU
w6b0/H4WxEPBq6uv/fmdWcsBzzanKuVQd2S6HzdzTOfkucpMNibS3ddqL0my+rnGhUWJRTvRqcQh
w2pBP8PW/0GG/oygPfEUNHpr03xJnk9kX1dwuYWAfniPc8g3Yv+rYZQRPUdapX3Y3Ajt2TBN808e
49FQyQe6a36HB9TMiKuxzcgVDw60A1Kk+AylJsCmPcKrU7nxu3iHInyxEpQr9GgZGjLb8zalCCen
IpT8Nqk8NdCSITc3sRA42Rx3T53bu7eWiUWi0qLWNS6LEb9lrFG5dwa/q/Brq4+8BqwtIQfWXPWi
mp+ddNUHTDNbxvlDXhK31xoWHzYvg3RMRuqfBArfCkHkPuXn2539bFIQVKk+ChQTmbCV7IgsJZhi
xZCyZGMX1BZQH9+2BXLSG7nPnM8C/y1WwgNrI1QuM0mbtvl9bus/aCN6EOhWEHNjrH7l3QItV/Ga
jc5aKT1wSuXCRsxjLkjlTXIgr6UwCJdwj4pbzyPlN/NLq5P+FpoehXwOnXCgJWSFGTSmg4i85u1l
wk4Erlpn6HST9FQHKpT3WAYbxcx3hQQnih0HwXptKibKER3IzrHdRY4PnocOYGLYgUpnQy1nD7Fl
Setzq/dcoBC09GvB/vzDufMWqIwmI3pZdvTt2PqkP/HOMaqokCGUs3VMXBaRQemHA7owR60YftiH
r3zbDFGYgHeTYqJqsppRlg7RqckLC1IQB4sl4L2EY/uV8sgQZvbCLQMIbiWEF7CxT7d4UcZSDDCV
n7nwBLnB9o2n5lyU7Uf3Os+N4STIKQRHp0wownObXuLtIVBXqTJ557wJaQ7wWPIVr/8QNihg4u/7
LcLYej0oLdt5NOVpcRSXfEUucwDQjcFmCpOJoLtgEXgnrpv3VuTZjqLshyj1lTqdL0RW2468T8OL
fa5GPCYaJc9gOvpn2oct6MuhMk7OyaVQGa2AwVAMWu2MqNJDU2JaOoh7pML+JFMkgazJhOMjd/cK
kqnVjLWncwrYWmpN6WP6GK0ayP3Q0Fh2RLatciJv8lEhpYyWlyvgyh4QiWmraU8M1i86pnd2AZYC
xNxH1bJeihabwB0J//cnLwhiqMcmp7wHGGbrHhCzJWpsCEs5YZ4v3TkJiV1+cTITZkKOGab/ij6h
TJbm1AQPTR9m+MC8N2tifdY3ys1stnF6zaHUw4Ou6PFV5JK7FNrkH9UBJ/r0rqs3M/eYb4DHroRJ
rqGIDEOEmS2VQfGfiFAa0fYmqB6KT9g8fKTwaqLzWTQY6CWXSPjo2c4M5n6JIu6vW1jkcxbyPurw
i+0UZWe7ElmpdYqg3RzLZHaEXFFKQgXYgFlSFxePMsx58z7VGrmwSLHA6zrh7EN/sfBIhF2SD5qX
oNTKO9AE0+/wYNVOXvorcyCMTIxFzoCEdy8PeZ8MbTq0EwEL8EWg85yIxtf0WyvOw66/YEb0w+vh
L8FAuq5xOE8kjwIAgbdb0lb19keNyd3ni8rdfE4A/nhK3pURqg816wzRDIY2lKhRHz/I3LY58ypL
Fv6yzeYhZiXc0VLoLa/gneHOcs5w0uEok5sbBmim6bUcT1MRmiIPF3GjPhOo6YtH3ztZeQrwlOZp
YZns3wrm+of03o5RdsNngUW9BibisuBzegvqR34v735WCQEeElkJvoJGW0r8BEnjqJxepfzw+OOE
cx8jAHiEIKpqmkWTqf4Uh0XWAW7YAPEVPyNz7pS2cDcVFZ2pvxre+7Xz/g3nS1pldQMjCEXG+ooH
sY0zgyNNJOdIQ33r/pX1NvQSNKzGhC9/3YezJY5vNVrZk+Cn3WOouQn4do4WHDgUxcwgmgtozrkB
pKydn5xAaosziDOgercITEyQ0IX4WePixW0Iu5t06B/en9N1eFl482JqgBf9GEgQIOLOoLEnUjV9
3q5bp5ur2FWO8b1jrs1mQLZZBuOZf/OtlsLOuegXj6xCQGpJtlC03E21pF5rwuCeYBMiKgubvqul
/Yuid1eKGC+/AlxogGNO1/CGIracqAvdgtLCWxyI3y2jwkbDC6wCTd0qLLCafeyJQFE7zVGy2Cbt
pmSgbhtmXv96ItERG0rxkh5xj9Gc7D2TbI4adoUvdhEn6HwEJY9GMgtSe2IcS5sl7STGanRj0KfP
4ElnFF+KpevW6jk9LZW2krRogYH5uV0bgozh/AytBeYVUSC+59JVrAql69GVLLjtXqguBI0qkiwy
3xg5w86381VVZpE8QXqWf2sYCBcZs/WkXybFbo0gG6C0Qq+v4tV6NNDJROaSiFHLZyArEEEXfSAl
0zyStiQS0bKUb1cpAjOmJkFZTqyG3DVkDKlbFnkmijKRBNg7XoJNCpR8AIDOku6YtDEKF6L+j8Eg
SXHuzurqsotZ+MN9k50jJI509ZfdrfYyMFKfCHrWWcrrwW5l0sSAbXismPqrOJS9Hn8KOB6eyAlv
MEe2H/OvX7Dw9Ujcnk4JP43nw2NrI0KxTrpg8UFBOntb5PpmCWpC/Rp4EpfS98vEv3Oxc0eO2Vs2
sW1yx/SHMkN2U20Xx8vS6usBoogfipd/sUmANDnh7eu0chneF9OJhi2UUYXwQGI8qHcSjrn6Bu0Q
xnDFtnSLrlKE1xrQbpz6MZhI9Q66v/J8/T2khie/JhbqUD1AdCz3CmzF4UrnFv3Op13rsx8x62yf
TbTIm6iQO90RU8UWwX+zagq7gmOv/vhoxNXnd0UtsQLpbaX+7474zQYA0dEFifq+5FUQ+AlaAfr4
VPssqOicOYMvHOQ7pbFJ0rS/q6uliEhYZkMKFam2LV4OZwSPIMaD3O3nYZQJwfSKgNFhUZ17OmMw
R9Q7SJpRWEKuWTSM2cdlQnGRZyVHEluhKOMkEdQZzapAByTZOH61SYW9wx3IV4UIkkWlj2/FMEl0
jjRSUZmbgOSnoCXxLiUQAZ4d7lJuPFgtHsnixN9SQa2e5jAABDCS3StyjW1hx91o6uRJAD1sV7k1
tRCJDxZamsx7avluCMHUf/OrY7PnJpCvOkeUMNyT8PXo1Eg7IVbspsMD2YksNu97NUaEyNfW0+WZ
b0zvob06nFzT9TclAu1882PWrkyX+4JE8i5hWlOX2HfioV2XpVZ711qCfNxxV9lLaY9LT8npnyS4
W/ybF/r8MtGbveIjOMKuRf/4PKQO6HFYV04CSSThelk/Pth8yC4SN0oZy7K4lq1mR8vLh2yF0QjJ
ZDuD3UCPJSTHTsF9G8VgQn8VAP4lBCCj75hfPdZq4vrivEW2VUrz5Dh/0ob0djqX4SyqKRKO4wQG
2f4EyS68QSCgLt8ekhL5SlW8FZmtMS+9BKRq5go1Bt4IXh1G68fB/TEgdFVMH99TvUkkDDQCrKUA
6iPuGvmuNVD85dbWxeZ6sjpSYe/PbgNorshcreHW9yWYluvRgwBFpf+M7Wan6uTHKbLigwB8hJ+W
lK+zylY6eRqcPpYY4U5PsaBYSy2iPe6olVaBNQlwAMLcOolTPk81Q2zqdjBqlvoEKPzdh6cxiRwX
b/HTdYhQGxvfhU9iyXpFNJ9QETD5LOEnt3aGAyyxwZ9wnRMBL9nBENu3JYql9dg0XR23rmE1v/H6
jckqr9+foVN1czaAHSvhhhQfezcfu/6bLnacYBdJgMn28nb3AuVMyA8P4uQjYeeLYfZKMLCTrB+f
dXgoLRCMbR7mOQKHrqBg7tB/y41WKA26hDxugwT4jKoUaYcVaijvA0vV2cHLUgYXHa/mB5Ov5202
rCinC8JA52T9itfEIBTo+4aDiuxPLJVaLxi+UEVeoAFQKwfJlwu5ynpTabCnC9/KomSWoHKb9i3y
zRPHO9gvv7o17zvS0VyBvlrIh/e4J+5HrY2QYkiHK0vxdaVxRVgYKZz4HXGawWMGGrAdlPnpJci9
HvmsLl/yr/qwb3/dmVJkftvMbbyqqrRQbJGeLHcZi+zqH/o9SJ9Hk3+b2Kl1pOYbWr8GcFUZQPXK
WdPk0BOyW1nb4qJi5+KmWvsHrbisfVkIJUKDTE0iMAQGyyWyA5trjbUxWQxD2blxb5oHsKcilRXJ
JA9VOV1lifMxddwEAwil5/ewjpRXRAFnUzwOcsyCldoTbABjK2Ry7KJx8w4hSyoY62RZDBae1dyi
KKzo+EAdajZgXdRlGZXgLaXyqRtpjRVAMmPMGM0K6IQRC9PKt5bLuMdpRYeolTY+n20HDHbgxsls
fn0YjiRaYOL/S+rCVAwHmKAT7JI0J5bIJyJIeya3LB9bEe6H5oPVcUauC1gOzopp8jsHagVaFWz6
d+UIPFe890eE7SSS6sACugsPGn+v4LuS6aro9O6bEQoUNZRjokVe84xSdgMOcX9smPc5GUEVFaRG
Yrg7R6kDwYx/JL3ROk+rCxryq3ubCty+veUehLQ1EusobXgBfh2W2ojkteMdeFQEL7OAsWcH1L1W
4S/JTTU63waLX5zubVzuZZuYECgLGZkwxz5oTYLAbeb6q1iPHcDfWX6dhrlwdom9fnXWIp0o5xDT
Vun724D0c/MfCksHDp+aRWA9AKHf4gvHxym2ca6UtQYZGEaWOPbweQyuy0CXO/g0in/9Cu4NYa1D
iX0Rjp1bQRyKV5VL+4NG6mGQjF36bNELuBZmau2VkyzFqAqMU2HZQBdMDZRuEd8QQOIBkasw90zu
k9cu626ZqM/CiQzpkGh4Qa0hvuPlPF8dg99LE8FY+4wPszEG3ZnGJBgzgxtL9B+mDFc9jpM/H5wo
l1xtzjVP50lAP5AkLUmTrDWlMWUFA5hN9Ov9rgFSUnq+rsl+NvPbsg8ckmviv4ArOQN+aYLKew1D
qxc332UI7PEBBs0DXdsLVZ4exVJVrhXukHDdZClYIMq997maxpC/a6gHz6AmxvEqsIUjUE2rON3v
w0XDkr0sHQbIwHJdvXvL5w4eUU+mEg0x0QGTiuG1Um8YCgrZ1a5JZclWIhqdtrLbQGnsMw8tS9rj
WJTKJDSOkY+HnW+v02cRN6Mg2aCFvr4nKIa53hhDTAuI4AOkUDQBCxoVxXs2zYx8o6CamcLamlmb
oOBVEuIUNNixnBaAMKTuOvY/A4bxS9tnTiSz8ll/XRx0jFF7kp+J5FRQsynpX+J5vQH57AjGEl36
3aGO0zBYpWEFITRCTzlpIvIt8xh90pLUBG/RmhzsYJr1K/TBlnhRFhKKi5nQ4EhsW0LUbOUrezO6
ZUgBRpcqddF7/xMJjAAPOtLsV5dUUT4vr2hBoqKxqp8YjJ/jOLgvAachSfgWOkXRN/BCvriLH6F7
JK1bU7muY2U8cqEpXFM/ATJJEiJ9uL6cxnS1IjUcZ/o0W8pM3ufxuYOZKy5u2tUEmzqMn78FEMTK
M6bFHQQd5trDjo4r3Zq/SG88gMLOSXGqRH+9AUG7rfy35lJuRBOR3uN13dMllHuGj8iXm5h6Aay4
VtABHYwX58p+Vxxdz0DzCYF0PZjhxihWUflEDVlmhDf/J+q0Se7WaUE9irWA8+EF2Ss8BxLFY49C
CeqzhcrkqKhgDIdQ2yMXUrhpp7ABBUdJwd4VpeRAIXKZNQZ5IbWDFKPQ1cDmh9hTTzREUFpNt4jb
rA5GGBq1keTM/ltmOtkPUl0Qysx00NFcbwgf6c1Kr7b3VZlA2XzcgbIsAHdJsti1sG73R7Ow6g7K
QUTm6pyHqBSonCyv8+Ejf2FdOSZ8VtA0AumXk79tpHjyxvcO6QdyQpL/gHNZOX6spEacmD9ODoLS
kfEL0gXRY7co5NTUnnjqsbMoWyWB9wDmHoSZWjQgC5sAFuUfzH3eBeyA376tHN1cSOpY/ivPsi3Y
XQuvNFqzy6na/2hpBAncxgeNOjYQtVkSDCaolEEELWJ8OcOP8SHy9LqR55moflpvFmoRcMcGPlrX
O91iTHuYXW+gxkxWPzIiFK344WUJ1FsboKhtTg4KFifypLaggjEv2orlyiHBbaEvWKATMxReXSM5
kFnrErn4SDzQcyjRbnKQ7UIoksKm54s2A/5Jptzlecx3LIrhltIUNCm3759Rg7BTYWOEOgyXZA1N
bTdJZgksGlTecgakFHTIaKCo7saE0RT+hP9Yk09fc6o14JUtCHpxSuaqIk2kAThr9PnYivf7Rg+A
KvveVNoh44ai80gTsV80ub1uP3CssZF96bd4bvDskqsepSglJTeeSnEgFnjk835pdnRt/jSa3bxP
3zC7XcxoeOp7Qj1iu8eGWy55L+0XqoDs+REHPEZbwTR8gbZvHN2SH2R7GKOJrwd7trS0v/oQZSXe
Z4bpqAM1Sr7+Y2HojLldqEcVNW1md2ZswADvUvxmdcnk8//TgPLMVxYm1/zFFat0OOXwyz72U5qN
Or08ebz+PvTnyWYF0EMJKWjxRbft6R2lUbQeD7me26o3+g1ExKSccXlQZSkYdJq1vumg9lEyNw2a
h/c1X6fPOYHAI0KBE2/wTsFhtKr6aDJt+g9P9B31K9MJhPeRZ60J5s+AfFefB3WKX+4j6lY1iMrp
yz8yOhAmnj6+iQfzGYLJULYywo4XToz1xA17nu7sjCeC6i14EBGr3nKcRxTCkeiC9X6gPzf17OxG
iU//9OQt+p/ToKTiLpKs5REdG2k56g16z0nccqeS16sVCrvioHkxtxi1gmpCfFJJIlBhmrm2rtP4
wvQ6+/cWnsv0718R5lrppREqMGdQ1f9ZfMpyKbL09pr5TlL/YCWRAw7SrxKSJzKHB0q21avWJBNq
wzhurgLz3pbsYCQZ7patepNtlV4Br0gFGdK2Niw8F6+fFF9PQxp0RWOefB7Y6Oo3vGDhTQc/I0lI
y1A55DYqQbV57dbmVQ3L2iwcZJcjakAcNfCaxjEdDaFiWyFxsA+znXnWdrChN3t60CEV6O0r7Ocj
PCXWl0I3feYHrVUKE80N4qaCTNdrfJwrHO8WME0K9iSdKswgiFIKGkPjHRIljc5DXBISJ97zHwWh
MwOfawGEHd16u8VJfklpIoOkgjTl+vqC5GESbkp6dNE/u6sJqEx1Ry05XtCOC6uCooKFksOzW92Q
dJJ18FwJug7fclNMNbaKUBVTKfPiCtw3WMyrsPohGHUlU+WhhjSno8ZsfWhAz9lzHeMV/2+Xcvcx
zjhXHTdQLgjwdvCGNqSWEjN2l2ZOPncZePRurrFZ8sCPMMdbqE273nfLDyWAOJwzyAIryd+aE2Te
+o1xbVLPoznT1gAkCcXkT/ldpnD38XNzE6JgqAGURZ7XnKi4Mz9YDTYo37nIwTZMCsGXlEOvGYvQ
mINfRojkcHQbscXksGQiRASkTsEKnFsueUYcQM3h25loGVm/ywwvgJiUL0qJhzqjPBaZOiTtEZJd
dpRX6zaqzqKUfWljNNbIzNRXQzznHK5Q5Z2KnKsaG4U67vJTvx8MM6sbAYDb3fJ8M+S4OzHxC1Jk
CsoUZBGmYIE2ICSwePmoKRXjwbTrkSzAAwUl24//ujknp5G3aH62eRMznAkOkigMj5k2ZRV0isaA
2PF0yD2H882MeFuXVvUuK4iP8xMkmycQXBeCFmg91oD2fcZDyWZO4KlTgCSz+iMFzE/s7OIEzfTl
nuMm2EFYDtXXlytpmZWaetQk0KEtCRbqK9zeYRprUBOFitWHe0+IyUxnKVuXw9K4U70v/tmzDWaf
GKsLNHvJz4kOz6agnoRxDQ1a3eRRJPrJoevZBTxBZfL23/7wkkoWCsq/zEbJ5OjilfVjAumPKFa0
VqNtfyp81XdDw/p1c6OOaBQO2NnUVDozoETrxo5Jsnv6JyWsAJz9Trff0UK6xL4+I4QLyE77QjOP
DAPuZJKQ+oIDwKQT1S8qTr2BH2FaKA+j8NY1D9XVxoA2GwKF2He9LHzWYYPqIbhrf+gHLMkULPQ9
/ilVFpKUDeqnOJNF7hWrclgkoFxwyXDF2I/7IQpA6vCGi/xs1dpge+SSoBakB7bxSFHpX/k6L8bv
wGJKP6fELQJfP7TL4aBf+O4koPUoO113lYAsmRcTFiFGf/i+dpkRnoNKvEvR1gxoQC/8YpMytenL
fK2FNo8WlKHgF3RqRvmPwv7Qs3uxiYrguJ4nXlQh1lr35SZEMZkM9o+yk5wAdiej1YAi5itJsBOs
eaCzppXbb8lo3Rl1vdI/k2JUYDluv1P7n2fBc4cNgjXXQ9a3CjHTCvSClPDwjBi3ufN6uE5JE/yt
K2B5Qzu6OnjPxdN5lDVlXJdHmnB/WIjAXX49YZVODensdK1ESnqsIzubhYaGPfy4t4aELRCMd4pu
cpICcaTCK4/h/SC3Wod6VRSN7tThIf7Fce8DLW/dPQj+8TG3ypetkqD+sEVFY55uWy+MpX+tP2fj
h47kIH08e1k7T2G2DSUbIY3iybNGG+hIhK0xfi2DX5cDeq2n5CrQHoWCu7/84wXZ+vwlOQAkPqV9
hRXb55xCKGRpiSksZdr/YGkCeraGT+1mGw4OjPNj7eIERmHMwRDwsLxtf3w/aEIlEun/hw0k+QPj
DL5c3NKXENjdBTlFntNYdyY9X+5y6RBa9WpTNXSsr/k1Pv61gLGOmi3Jb+vl3+vJcnfXtvg+s7xs
1H7F+OpbR4elpU5Vdo8KZgZjhZNWuBXJ84DSSY918/1g7+gwYQHDDbAwQd+GE2Y/R4nGA/lYW7iT
y3C89eaOeuxj5BOQ66PLUpJUcztaVYtwEBQe0KELXkbkzvKshgQ0zQ86DTC5W6/I+rlxkj5Pe2Sk
1eTSrQl6Q36VBGQ3JJIRJAGURcYLO0Z+Yh+UNz8NGh1BqPgo6KWXJ1GbzheNEsWiqP2BOUtso1Z4
bnt/JyXN37d/bptWjKZHfLvpJu4poDCgpGNksweTD8ofiG1Cu1S8ebWqqS9RI/9163ne5XlFemaZ
y4o97hLc4q4G2u2/BdwYGZon2/io3U6+K8AFgIHjRSoWGDt3dRWA9kBOj3SdXRbiKV8rxP6+eGzs
kSbtNjJoc+t/HmAmGxUapON/uK1CTjFqBeD/MPaQLUFj5AXuNJWiJOZbm7TFe2LwPPGvcmxecaN8
bc0gnP09F7DiiSKk1EwBNnxTZJwB6RijuJBI+gh0evKBhfuc4Jj76Z0OGOykK3ycg3REYCPiVgaf
RuswXhtUV/QKFA4CIIHqTg4T5SQv5TQsqqtio3IwHQurzmt5bnU+suTzprlt6dQCUTPmW1opZxQF
Fn2h27ZHjee7VnswDqDtnscC3Ok/1z4wTXB9jXZ1K5Sto8yg/Q/k2me7TqSE0mhrxMtRIzQ0G6Uv
vc/PX6thU4ZtGv6BKjpzY+eQxUpCP3wzltA/6mjH++2y891uAjeqWCvvvHfvl028AHjoUGB/1+C3
R0nBzrkFIvgQeOMlGK7czHHdVQOTgiWhWqFuk0+szjPLgmGcNhNo2H8vNx8GD7y3AZZzObvz1isK
5LTjBrK72Gx+EluMYwVmjX11XV9CmloANhfLiimCcEvw01ydw4p0HPInXcPiitPFCnvLmRuMpePT
sNMtnYLSqPTE8yQ2/C2dSmEf/kzEM5UTdqNTAi/1hWtpiBrgkO4edASnen2pOcGFgSI1VSen54zu
sGxPE2Ij8owKc5jNH4IN4o2FzGEAA3B1hBkTdSEp8uo9oYT7i7/DarJHDZrmh9hVqKLtiPFrbwX0
Lb0DilZsjBKJour0YGCPNUA+KI4zEJld7MzxgDKA+HRt9RsJUwlKckSNAynoFKlRIzWoms6+03c4
4SPu2rMBhdp8Fa9H+gLtB9xGCF6GXXOT7GWHJXAAmFhWBVJrvqTepoLsbKNnOG1hsGIn3Rl9xuyJ
C5Me1VAM5hsLHMJku2Um2CjEfCpzXZfhTio1XpyuuZeo5dTHwgMvulZVGS3gYcrDahF3o/MiDn+F
qDoEmbVE3zyyEnvM7QnlbYSQ3Kp+CRiAKXQ4Vqx8+IxaWaiXl72MhJmtlRR4Hn4mWA011qDHIg/B
rcLwy+CcAAi5NkMAsnb8iSNrOs8gABEupPbuWG5esVVSVGrdsl3Q+J+0QI0tvyq6yPbrIWiYjuT9
9WA1hfpR5wmc0YU39D6iE5CQ72oYqAgaBDF/xwpjyowXUKLSwC0Q//jPJ98qO8f2szKr/gTNmGpR
/Za4b2OrvprcGn+tXUsR5nZF8mtojheI7ENzZKiaTEseKFCRlh4Oq0Ik+8CFGSEhR3vd9tlN8Q5o
v8np/4aEB14266KJWYMkWag5GmLjoYhIQprLHfv0WQcWAIHNmVi/LbjlLrHVUqRuzlILSc/JeIb9
wMoxmFyAiaOHGYHxqVpty0nA7jnRjIm9nxPDU6Xkm9a4wrucXi32Q4dbr8LjKceoQkohkKU6hnb5
W5yOhf1ErYi8zoBI/BHXehsUVFKb9mXcpW9D5q1w/s7yv6Q0bgC6BuQpa+tRXHyyTZxIiACsbhA5
qImxDkgv7skMwwPl6rYoDe+tj1y2M5CVz8Mjl3IBDPEIKfdERkbGpUBQSk5RgrY0mY5jK/Gg5FpF
jHP7Buk5p7N5D8xZtHhFPYYkR9i6cBdY0IS7J8jSCEJPTbmGefY1xthS7N26ovYUGRVOJR6dHUBZ
uGEcyk3d8QQ6m32ExD7yjX0WUuWgbJxc0O1Eo2KVAmIVypK2h9mO391flt7PJ0p6UBLcBQlEs3s9
/dNCjtFezkwLGKN9BoWfIUDJQmSyctjjFKfXmv25aqHhkfzX218hPI2BJOkdQ40K0J5iAglcI7DB
LdzneiWBZohE2KGwqj9415OzmFvmZ+P7TihcEuAR9Fn2TuNbmygOAfQcVbKdjyaoFItEkIz6zj+9
Tz2BOr8fGrzczkgVSZDyJ2qhk6Exy0dLdx7R8f9Y5d2ExyewhkAhoKU+VzG9pz1fXWQyN/VpEgHT
zrtLFuMOe1QlAhJXfDcowGrSYFIEaJ8aUpvldzmpykeY8h+Bfk0wReJkiR9wloskb+KDsMgpmll9
a6pDQ4uOupF+Iz810DgvzvrpSWkxBMR3paH/bNMZB+CE0CniiDcCltQk7/O0Z/E2Lp7MKaFB8Ead
xyBfOrNqRGzAgfBeg59jw7kwv04VqT4mldrCrG1lRWtkNJgA72lSyVjfNpKTzlgEpBcT/iqogEZ5
q/+OSq9vn6SzXPOtRvBTh0tyGLYGUXu3x0vpFlxNSQDo9dHH/xwFMtW+TjIH1or5dT/kti12v9Dp
+YcX4KacWjfPtOU5D9p4+RBmMe0t3+wgXl0tAZ57qccgcfaq52DTMVzDrMCIODLScRWvwwiJ/p51
X+tlLgGAYDioidEJ2UxP0CoiJCiJqyxVcguov0OEvQLQ8/5MP1G2eyZ32/GtrBiYR6eMXLSDDReh
AY3rAHhCpswP8td5iVHh0b09z4ySz2V9yLIJ/3WuJJUdVmAIDDmv7pnLD5WmCzhLHypthzd94YSX
WoEU68hssIkXfzI8spKX/FWZBJ2802YXhHMmUUd/ws1aHq18pGDDTkwtrO9WcFRsduqL/QSyS+iu
XorhTg6nIqopfzWm27vQCiwlZrBEVyd8p9YNJ43xFLESEGP+6q2mScUlkDI+9fFXVZBU1wDj3boc
m3x9K/MKt5Wksxc98fDOkBax2r/5f6N99BriMX+UrKThyMx9AGKhNfBMKhZJZmbwvV2/cUKdyz9U
IaaDHhstJTXXsD6bFSK7EwPEJzH8zRq6hyMZgzOIOeRjr8AvcnW8JRp+Wzf5W2srJBp0ST9hmoSF
SGn8XJzU/Msz4ZlK+MEFmjUT8QWpYP3zFEYLPFJwyCJV/VgNhMAN0XoboQzRprIj2mCtOkxW/qu/
N5JASpyUo5OfK1uJjHSvgJbYd/r461Vroz/0/0/JWX5lIeus9TQizm/ea+i4uZRitoHmkYFOTHhZ
16pIFkefTRZ1Ap+7hKfmk2fKuw/mhLJKiBNKbSU6iDGflPFOhJTQ3HLpvqPQi+m16eN+0OIWaokM
ZAPB/0A1IlMVCYEKa7aJWWW2Eyu3v6BW2rMFuO656OLZuh43hyEkH9vtTnHscJ+baUOUBIVlESCD
fLP4Cu3cvhlqAf3SvM9n8XaMD36UIrkxiWAxTzFNmnKgRK/sXQQS8T9O6sjkw1MrMiOsHT56G3RU
QUUDgJYGOdIaTfAkG6/MnjUDpxv6MtGo5xz0vWQtTRAmSYEz73h8k9poG9A7QQCQ3/qd7nx0OSEP
v9rma9rjK/X31/E4hI7trvjJnrT1C+gUY6HkT0AOlh8YDjTbOnCpCK3fKZd0LPg7NKGN341m8PPP
ITCpj6QTksy3DT/GXWDvvxPCYiEqO5oHIpozJyRNhG6vWuFLkf2GSYLzWZBQHDiGv2aTzJCzIxCy
7k8EKyQd+TEUlyw9RAwziPO9BaAozb4oxga2mrUTcgvO9BfRqOElnTsIKiZCRGDckU54a0fbMPRp
HM6jdtfMFUiWKhnvp5jTPEo/AGwSZXLhs/hbFtSv+KApfR73rP03Apj7A1TdhdpPjmyG0TBdgS3x
IiqsQwwvcvo0kuprFLXAARdMfRVCVhf/Tr3ckjSXUqF43eUnfGB0PkxrKY1nccu17qMdwojB5fGD
Q0nuC9hgqtCy56A/NORS3WheP9YIR9YGxJH89sfOTgTcibf7JvAWLtlNcsrH37NoIy6nms+0gPOF
u88Kfw5jXj9QeKgVu+ma4zsHCX4sAger46R1grHXr0FzAS4rYvKbkIqhcA+gEP7IrJraKrYh1wIK
4q1K7NsAo+0Z79d85xKknLfiTUchX/kcVQmMp4eTkbTuoBigqmhYtDLF3jTFm8C5tjKwPeNy8cH1
E9/rV3teWprQ4G5lRhvGrikmeZxlUeh7LCoQDUN/t8p0xKBl/KQZZo186RTh3bDy90m5f5M5htvd
JGPbzLIMrnRWojwOjq1b6VNmp4yYDGHr+LRN4TA66GA/gK7E8qCeg8zECwCIFa5MNs0fyW8w2CR1
xkMgyVpYqUxfMaPSdgj2d/b0fzAUzWxZKEbSjI15uleHXy7SME+u8fHz6mgjTYA78ZvF0R+a4jWk
SBlS8x9Bcyfh086Zib9Ky1HQxf/+MqFM2qk56Vvog482hsbkWGKmjLSlX8qHuN8MlrfvRDi/TAEo
XTe6z0lofr+iofTdIYaiFI1mjDKYRmBVR2l42puOsevLqHS0xyokzBzo2lMSz4Hb1GbUUXOlp4ax
Sd4d3Yf3wNcN/eggCsjq5XLYm6qX6RLxwwSdbTECEbBvqDsp9s1LtFLQ8IW7RMnWUsm04XqY5Xsj
PtOajWiP2sfUGV0CcfyXuQuUwebE1x7Do2ObU6AxjwHZFLKOJoPQvWe0ZRJHbtBC1NUDuaKiHEo7
MSlwRh8IvGZLFmrA7PQuVW+oqU+hE8If5++MiwTMCRxGILgTVn0S3CrIRZMo9fkbkLoL45dD+tST
tk2AoMRSu/07IHpW9XiSet0l8Vz0/9M0xHqPeH+4gftePYnZeWlo8tGpXTHb7b1Nn4E23mhYBxqS
TOtmvznO91l0WfipqyozwRDDxbsoXWwR7sNlt9pEvfbPePXOBGCBhPXjv+R/8hCfokCUHNOYtEjG
tXJ2OHEFu5u1kK4wceu4/xGkSyn4tsmbczmUlJY3ZGQcCNEGwJAY9k+bNz0piTFDGbyn4PvU8kc2
etmdWB3jjDhuGZx753GVZsYAkCIubC+VwNGDbYU01mhdWulzoH+x6m9OzeSFfq0rgbWXW9nI1D/l
VKbfWfg8N6iZ/7BAtVCh9jio4j7BnfjjtTd1wW8/ePQy/Pl8kTzBijixpz5+Nx/8RwLIEH7h2OPm
wswOca8PUCvaw55OIr2S03PmhCIR7dyir5/kZWlT74Sa6dHd1DCDZfVLUuf5y8CqGqkqMfUT08A0
NLzViOGvuAK4MGyGfRdhe4ww2XRqzwpJQ0Ver90w8eMIZ6/U8jCHGMU3eUK6K18R/H82aQ+l8GWe
/VGdYfH+MaJjPvnLTP/I6Rqvj4D9NX579OS5NzuB2AD+itsFKCOlKrt45rSmkJXc5NKKnIhwDa4v
EexonfNDKduZ8qZgBshp5Gou2bXZd+s//IPNuGgP0x8zPsbBCwwPA/tlLIgEujDnKy1HQUmTuy4A
WhEcqUl6wAvnQl9zoHIx3FJkhGRrGbJbUpQy3UBnyfiUJuLx182XhGlCP9LNg+7AdnqxVoLUvIAf
9h4X4jsYo1kyG/kx/T56LQwpSFTJYL/w+JjUNLYes5KOtWLmQuKxRn1FMNekHabvB+FlTF0+qbnv
yvqmd7nhnxjlwU89Ce6OOFheE7vhVhfJGLQ//safqhdnQXV9gCwsQej6DwUF72jk/gwFHUlmARqx
5d/1G2vfMC5UnKXbw0VjGGN33myGgIpmAnCS9PGVKKl+KoWX0cFGEF8hdkOEbCgwDjc0ILYsqE8P
4m59OamxAI+khZslVGvqXHD9HPfmgcPUKnptaaCzUnK3bFTsv5k0vyM6CxcyMh+aFP0Au1LbwEBS
uBpnzV0lyjQahY+TGf14dKw6UEtuAXMKdz8k+gnoT/t9f8hKZfjyc0r5vPUumYD6y+47Og2i2Qzf
Ltp3L/EGs6gkfkV2BwptySwmh+qD9s5oUsMTzq3yPws464n8n+fK5+3vJuBWXP9frNqCcDj5x/CG
BDmSpMuJizXsqlNqsZUcJxfLngFHhzTgoBuEalobWfT+P5/OyWWALTnL3B1UOI1XBpOQwCbvPgs8
BbpbonAa6HeUGgWEeiWTEQvF0Kj9UvoxFxKBStAw22gNvRN0iRO/Dn26TERVIbLXsmv/vrheTdc7
qi79Z05TeL4ueRTncSrYzUBFb29eB5S2FUash5aq/Vc9Eu9bWrNy5qtqTdhyTmJImoUKDPw6/5f8
yn8j5rj/HfSHsaS9pfZjtjYn/qfQFtjchNsTLkRw6wSwmkd2/jBoy4uk/FfFMDTvNHCBfkV12SJu
w163Nn69hIDXZTrBWjU90dRo0SkxP9mJHpYqFqbTz4Uif4jatuR9eKNCOHm6c+rTk/Q8VnzUWoQ9
4mxp6Zt45k6yPqYkQ3LJNOHCoa3tXe7tSdqr1hEDmSVSJLuwP6rIPj3iz6TLQRcnesh6vjNRa/oH
AhWBr/Ebqti2oskKectEjb+HWSA5VzreesPY74OZqHN8jUX3VO8vb+OdJka+tangNi2LmvfWrZo6
Uc4rhD2q1iralwXcDcYKilD7xiXBMf9MLZ7zUy81D2Ch+M3bDdzqGl4CW4Z8qCZylEEFLemTaqkR
ll3KiQEdCrhCKp8dm8mVyKZbW+COdhOVForJDg9mOliQ8GDMew+pKT4PY8FIyG28NyGr+JppzqFM
YlqwbpB4rEBAUTUACfefGO44fLnH2bswWjexdl0SDkkR3ye9X5ufS5koLycJ2OAJmjIe0WVx36o3
m6k1/WlA9Beka1Inq5iEpXM0M3CoOURjPu0mTlRf60k6Vqdy7P/ZG9csOTuHYERivjSTTjQW0uYI
pd9XQhrSf7yGO9YQ863Mm7hNdKtkh53UktgY9S9lBGpceTa2N2Dqf07Pbl4lDrOKSMufueaGOMiK
Mo6OaY1xvT6/edyp3H+x6wK38HPcKBTHIx0/JNTU4+xwIPcA6AjKBO/PkOj38peP8tzGjAOAbQ3b
StSN2EB6jpWQCe6Od8HF+u2pS5/a/F9cM7WffbkUDPoRr0sEDEHTHfDY3RORR3KacW6VRRT9pDzN
6aaYlQhLvrtTSPQftfbDXPcO2VeF+8s5ghJOT7p0PBHXuFpBwESDZQpC6CK0EoHUxKHFiAOVjfW2
KzlGcqlDtw5+t05fwqB/uRKL1PlVnr92cB5i+NCUBiCmWKWE2Uuo5ZIRlhZTFlWfqXUj5pQ4rxJQ
Q/gXMCqtBIvMxHaX9jVol5AXUX7Ffds4GzSZZHhBir3caCXGzIzZrc94Kya5dbO4NO/5cOdE1Omn
fVd0Zg91dlUUhzUNTfdddq0x5i5MnV6IfZlEx4J9aGZ5VbFRETyhhnGrRS81lqfosSsLM9wlBEgV
/aZFiqFCKbPeZ8/wOvDjq20Vw6n6aDkWrEsCjRTJ7yRHJ9GMPzSZpwX6/5Si01luy59vQ/xAs8Pz
gKc5nd1fn/ixJmhzg7I5ujXhoW2ncPhczgywNpyo2H+eqfU4hVCdrKKrWvnD6fv68ACWXDu18gG7
HmCRAyZ+/AwNZxGtzZ8VEH1d/AJ0w1HAktDcViKm5/DYt2Lbn+aSB+CiamlS3Zgnstj0TYZBOKPY
yyVFVVNCFtoW34auMttu6HGxA0EM5h8am/ko5XzoUS3Hut3jbmjb0leGrgmc1gVgH5sfQJwM31HT
dl7n5Jj32E0Ly6H3CTUJbEhkjdMICVIn55gdQWh6vB2GJRiiK6tC/fwV35lmrPTPE3QyBkVTjiD8
0CtknBA3vAfK77l9UOuHAgW776Aw/sVluexZ6Z1MwZCLJwugxD8i1HVIROx2uMxfC0kPBMRxZ/yj
UMpcbgCke5zTwt15bjoYwv/5Y0yvLPX7/NLQ9yOfvmTUBGmFY3iF56O7rDrdR7p26whOkv9sji90
Wt/8xAIcunYw+IsqSw/AocqQuV+mg239u3UZYNZ2MVjvWLJlzK3KkOFRLaR7GVS0NNnJ0RRCm7Ir
uPTHg6ocR9QuIIbSl+qS3bN0QYh2d1zosMinfFuY6sapZfbfl3otgUrXrqP8/d/wXdimuou+zI+k
xcXegdEEe961kkrPJu/k0a7QHyatBCMd7fFp0bdYGxvuQioIC6OaJCHdpK/vtzBJQTEFoZ96m6BZ
nQJUiT1vmV8XLkO1QjJLCFbEIzf0MXWJnnHN72/bzk61nzGiT6/2qMvQuhCADx6/jyXhAN6xADMU
oq7IQXIGjpuu3J8bfGsbkr3BLXlRZvc4VVfHx9NKQDVxVXrqFHfgbSvXWJnppSvpdt1KfypAYzt2
m5WY0gPS23e/sKLahSj+Unl6yVQYVqZSwHRriEK1/ZSxsqhBGHvMzOExDUy7Mobkpp7f3UBTwAkI
4by/Ruf953gZn2uWGLBYTSC6BidX+RjVNKcrook+2B6V8McIRjavORuI1252GIjBIpjYqydG3VvX
WwujJza1Vpz04/nhS3Wo+7eEeOWS5UirFr7fLklGoMxBScmd8OXNQHTX5I6uw/BLy5eYRmGalSdV
pY9JpyhiTaCksfp7K0J6XlmlWOSAj9Ml/fev29NKGT7yrqo3hnn+WQvxjsR33gMHLdh7//WGxxdI
nglCoJOYvVcRwkzyqq/Rxhdw0JxC2wQ7xS1VPml3XxLAzV1NIpwg3QT0jZjZEJwSlpIUxDDwSV9O
eyt4Uemy8JsIHA86VtAsZChJNysLd0PanN8dDnM1TqwAIfTtnTA8IQFfV7KVxfylqmzYYaxB1mbX
+uPX+EAlgmH60XM4SdHY57I0PbPZxjzKP1+xscSe5xwK9MuJVVo9TWgT2V0KYOqZ0l4uyf4CxdCO
LFrMEGI6o5a32vsd+9jswE6usaKdm2WI1dTPEgXqVY+vHb60wBj0crpQy+aYaFcOxKTVFsC45O6y
6xWu0tio5So2E+UROl80nXxmo+6hATnnx5/0qeBOKAf62GivdW2+JmOFIxerPPpdeDnN+wkWWCHx
312DezgXUNLumoSJPw3jen70lx+gQq/F8KUzZASxjav/a+Rd879BuzVbqvVjKMHM8U/w6ydBSdYR
C2NhH5OSxDs7iWXEGIRD/x7zJmPJ7zvJHuC2sJSc0dJoW4+LI2pMbnrPRnmyNsbihFfUfzlujfW+
N/6ZsR2aH6HWF9k8/IGpIaNdSFLuK5lDFZ+51T1spBYbPWJ8Ny+eqY0ksCIgqRpXCfScdDWQgQdt
UIVtPfstwtBTqqRHFNxqo0a90cUNN+EdNYs5mpm8f723D1HjEMEky8OUeI9eiKZfUS9rMHJi6mVl
9DDEm1ikHZqr2RD3aoTK8qPFN/XzqUvz26RGxBbRpXX+s2K7/fXF4+UMCJsDqnxm72IKkkmCV35O
Z2sr8TIUGHHVnjD5jXO7PHZ+4xdTEmyAk4gvNObR42AZg9UiGXCgOaPZFe+bqeUKfPCcdX9CoL8F
dnSCqefAt3VkOXrYi8VLtRIE8NWImp4zk9IjDJQWggcIY1n3Uc1Zeh7bgLjwQg3nsW6MCVSZfRQr
H4nUng2kUP1sBtQh1mTSM049zKhPlkcf41yGN1+NhXrBvaHlEW4JRFrR9oneCF4CphaO+f/MTF0f
/LIiooqCfGbOz24sIgZjhzQGvkcR/VLbq19QugITWc+heY3u2ialasuxeZCHR6vxyWYhtzSl6/Gm
yNBIS0WVbe5DStW3z2U/QyasK/+HRvP5mLHxkIvIZU5gH4xXZrJ6RBVxVBwMSlEolu4Zpk+Pygk5
mHY8hEqD048TFtqGdjWm5JBSX2yKbPrB3RZ3fMct7LLs2o8l93BYIy0wPRPqdNMEe92IBkjqnzUM
QASi/5OgRctY4D6PoJK/Wl9VLHiQFQ0Tal1edPw2EkXJLyQ/2GlauoZiteM4bPimDrsE6OdO2Q3m
haBlMURRCluKsZ06Mbn30nYcD9TpFrdT5B6D+6QVtwRXgMMevGCkLZ9JFXtAY91aDE/iGfU3btss
JkJJkbDsyhDqPRmgIklocbwTwFaYHUX3rMuqQol/1T+dIqgC12yalO+JVlw0YRcffqPteAmRCQdf
z5WO78v2zdK7IRVcGek7o25VYdvZKwswPq9c/IgO+VqatLPQSGNXj3j23/QsbUTL8J0Ac4ko/Wyq
wcG/vdzFFoX6kHq1IyEfBNi6CSYpp8mOEmkB3aZSN/igfSwP0HMI9rslV8bYk51XWRuzWyB1eN8N
W4FYAOwHJ6C6Ce8yNq1oad/pkorS3hP4nR49ZXgqohZHFClBftz7acowU2zG9JFs4IiIPZ6EXwTE
HGGhiPKLQyQvw/0e59eolo4IaCiQYgG7NrzA+4leB2FhIyjLOQJVxl//4gSWwFnZUibgxVlrk2Yc
pPFlUEQyW5zaXvh25FB/0MCNqxoY419RXSHqHPf6Vqomq07N2GU+BL+Z/ZfJUh3+XukA07EznpNH
vr2wMbCt1FPDAgQpeOL5DDqiWoMspo2Q0qH8fJM1ZX18zjw/5Qjz2sFYDExI23+BZWt9nGe4gx0i
gexWmlv2yAX3AFR4qEcnbL2yMZCEkMLMafG+hYNK3B0Nu3lq3XUkA2isPPNfXXr2v9LNP3mDoMIs
CI+fR6f4oihScu7feQpZMIFCD1rWdwvlBP4UMnBr4jqTY1H56EXBaOUY2uELK6eS0oiHHvqbgw4V
4Jj6BSJCY7WXGT3w6xkYEQa/g1uvwKSEVudOlQDp/T4bPQI8C9qo+oZOn1hnT4zpHA583jQNgTXW
cfXM31avJc/wLtF5aOnTJ6UygVL/62lrvRrEU74Ihrhp53o3+6cbRgELJQB0+NsDa+xBvqm5L9qr
IjThaENXSOE75uHySwBGRWRW1dufI6OzCXlSgWd5l8Alepn/lh2lE3kSm+iImhJXCejH2/tRO2PL
MNdaKOq/QeupsRmFeAdeSji9IjLBNR2PPVu6hg1ovFdQYL0A8z4mXipmQj+zfo23AFc6UYLqJjhL
SEQ8Baec+2YqifdZ/bBcTlxZ40QIppwsTMB9liUI21GgAvHA9S63E9gQv0ntbOvk/uWdwMoEGtOX
kRcR7SZ0HAlDWKQJkez7wy3nAdQR3CZZuDkncipHS/JSTL29D8UwPNx0eo0VuOIQM63xNww+W6DY
q0c828dcN8YnU5DYQWcRbfGcxqilBiMzPXiEb5k+0jMyR6jmpxyFjBYU5O8j7LHa305ul6r/S2JI
NozYkvVMSGbVR4sBqoCoNtkhPtCp0ByhH00eVvJTtrPwavVFPasTZUY8VmLVYmGT802z3ajXFK4h
T30R9M5Yx3VcFcJrnAo3OpchixJfB/n+JiBk9ELKbggDztawOKBciW63DX2xceJ9jQ6oV9Lk6n5N
Ck1+XAU2gfELmN686yYfFXpnv9O5SDbKBeEmP64PmA7kI0RDkL0+l00c0oEofliaXVxFGBfZuLv0
CfjFwJ+Iy3GHX3gUWBFnXP40Icq18djl/Gr8OqetxcOJT2Sc3vIqbbWLlI08CYbIBJR48nm0Ct2Z
lrcdwRKWZjGhe6t4x20bL99w2z4F6xa426iYvpkdDN4TESYBSyybgfs/YC0r6HV5TxdOsW4CBNTO
9UPw04olyh0NMkiu73vOrzfAbsnRWPXHgJuxKhVW+FYTlKxLWWcmFvAivYaEVN6wzjnA3bpQCupj
iL0F+o0beea4RmeP0+vEkQKnADA2vr5e+8Jh5ije6t2x/FmNaT+FspVFfEthkIUPEBap/tm67bCP
HpdeXJWu8j6WTmKmH2Fkq7YdzGFIQSfXw9+X2zPHN2SloAD9sB7WlKgXd/72urCuXCbuPp45avJ5
gfpa+vD7ct85Joei+76gjSxZ5aFpJdnB1YpTx1MH/2bGRiCymfPUTOpBLtvLMtFarYjf0RYuPeCk
hY1K4i6y86eWV9yASQAPT4uK/p55dhWKN1Ioz+JMdVH9QOYPy01730tt8G/fkLr0hBLz+hj78NO9
CY/fHMLGTQefcOxIekss1NZ7/5/i29oAZgFuyNuVRWiNt32PoBvBamauv3oNgEjwSRneD1bCIrCr
iAjT+RdmMttTL5kcZQq1sdI7UI2szRyyTsy9APJZSsj7tqoYsqamwPN8f70MVBe4pkBhqiFyLLVc
0xhPzgzVhp6kkXc+PhFik+r7c5wpjS3ERCj9Pr4tO4qIRNDJRll6jza81JsHL/e3Buu/VoGJsFCG
P6z+DeYdpoKNnuZSQ3gvhZq9R6WtzNL6OeIUPheKo+zxFTLVdxAp1N+WkLFr1Tj54sPy+9b0Nzrc
UKdmGR0+Feo4tKNwOtnT+hX7Vk08WYj6RfYsCRHumMYinbVEtkbEAwWZMNXg+bFsQrnyzXCN4j3H
0heyiuQXsJU2/HiIAAYigNU35k81GKs6EsspYflkYiefOweTH3ZHgLftBBQOdIGNdMkBOPNS0BPS
Y63wJprOiNcjJN9XfoAeMqpyxsCZGTs2fGDrIqpuCBQ80uMpt/+1Udb9QHrmqrnEjg5zh2YzlFhe
UyIhnH6mdW5px33lC+p8NPe1H4JQ/w4lf2vMI6OgGWcuSSh6lrVrIouJ/PrIqkOM+d+S8V5km4po
M/7v7OzKvHwsonEcTeWGkp0u1pbf62mNsrdy+XssnNPW2kwI4BE+N5qTSv81Yof8AeZV8URYW3m7
87T5uibF+g/Obmtp6jOvg96+8r4QY7tq+2PKq0WmMRcZr6uQhP9mFQ+A8A22q2JN5nHY8y1bXnWV
Q2bX1NrE10ppWPwETDzvEHJoi98OWkmmV1rpCWPawaQUOgiogf/Ye4hhmAtHYslGB3CXUcSZQBX0
YXHFJvuyrclzFqUjfyemFhpz6J4=
`pragma protect end_protected
