// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:49 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
anlPtvWHjivrIyHQivvgUow3ivi1vT8JGgvFc2vF/WxpsG/wssEao4ZbBtyPUnVM
zeORHmG0tGxHZOVb6rTr4VCxS0fA2dqW7hYN7Gc9pBNxIuCVxWp8MO/XmZ2ME0qp
eBUj0LXMo4ykVVD4i+tggxTtswAKDEYwEsvjQPI8TtE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12768)
8QGCZP5aUPMpTqVf1mqeE6EdW4n3tK7Y3tdCByIHqNRF94lB07WXB5rctrhsHSdx
H/NNtOIyyQXsan/TATwg9UVgFQUvqp/jZpMmRUkQVlxJYc1cAA0XNg4zjP+aME5m
1RqUdY14D0CiaKr1epWKIQZnA4xvVH0n2p4HEPpmCWIqSvVKwa1tb/JAcZ6XcrGd
Wm6hQzm5viVmJ381tyG0R4Q+gdknHZ2COdXwhAt/n1rGy98zp2WsBFrBxVy45am8
awXm4eodEP59jHtPPSwdD0EZ7qBfbtpYXgsTmjpQYnZPU3/m1ZxFnPyXOJPyWNfw
A0bVjV5fMta6ygu2bfah5EJfo2KJBBtn147KXP22i4fHVoq0YxYJKlNMDtM1iQ4a
Z+Ho9L8/KhRIm2dGX70Qf+YfoPcF+VOnkBBamWqv/UtNZM/3x/kUbB5DquZpZYyj
YYiWyMHn4/IS8m9eB7CA0mW5Dr1bxVxGcATbHGGpzsf9GsDO6PI4boJRgTns+WVO
4IoUuAVndRb6tm2colWFQghD3jUutzjrHz0LaTDHzt9Fud7Ls4ThCv6mcNCRwfBg
FLoFi3KLXhtxw50tRN1ypm1scEkg6sbzXDavZxZC3jWBi6otdXecSSobNvnywzlL
NOU3cunhHAoAPHFhCLc+0ewsx4eZKBQlV6xra7vifyQMHQszbJS+IQifcUV0kiud
fQonwxXzNpT4ybcwVjzC+40LmRCcsdiv7ADXT0mTWkvcstb30R6E+Vd8HyZt2ovB
oAfBYoiR0P2+tT4xp62WWH5BkyewSvQJoppWfOs6HFLTsvvNmftsE5VbIPEN2+sO
YLcWIsB8jd0mEW7LAl5EZ7yiWntIOkqqz+B3Wu2wswvyrrwZJCZ2HdlSKjsqRlOO
nREl5mx3RnA5aLbx0aszy+8vimYvHJ6ucMIQsX6Cx3Ftjgy1EDX9ex+m56vlYbOG
PIYNJk8q+8IoG/wUmHWhFJmDZPDZ43v1LDgQyPQNRizfA9TGLVGS5ieN6zCmnNhg
pTdZDcZgthCPnzaTA/xJHtWFLstTjgGwlLY6IcttKVQs0KlZdbQiIdmkKLFfD5v1
NSz/Wp17t8HhOZCmFFLDFSV+L5+j6GaLMXy5h/ckqpCZq27N8jBuwpTXGndUKUFE
17pt8c45Bqe3iC3AoUQs2Wnoy0g8OmYQNQJkheCocPy/pYotqkQXY4RTSIa4mufY
Hf3/ns8l4SbOXDkCW929VGs8SFxyfABzisUpxqbSa86NgF6b3o1XuJ/B6pPlcXqI
otj91s3NW3lI4uAjHVTEVd/k+NwdmcWdydDsBAvFrlQKPBP0XmCw9//l3KYrnXq6
H2TX/b5DR6W4YFqQYcaJcEjcOG3gy28Nt4d/hrU7DG7KxkwL12hyeMMGjnsunK+R
k3qZUBALjqssmLP2JAyFelYqUhW38jG8htEUq07guQtxnOdU0mAvPZguSeeUQRjf
QzLX6oUKTaJRr9AiTd+4f2nCWIwyf4mzzcfweFYUyKCfdBsNmagj5kZZklTq9KrT
pyoTv1hDXKTUT2ycVyuUoUq9YBSkSYcLw3THfcMMFH8odO0e3e4H+pqGtIqRm/9S
wtmOmNl/SFA1PWgRRAbFhKXnHSbdpuyLuo1QIte9RhMRZr2ogBBC/K6taXc1b+Tm
xjk9AAal4RKyskmOQPrToSZEiZHAr4CjvD4DMc3cbNLA2XRPJh3HT/8dhv+RH/bo
BmMvmq6AQPG+M/idka4EeR7vI8DsmDXscJBpjIDX6VTb767BvMbalrYEvZITJXso
xzYICbj9kFkiNreR3pdlDDXmXNBZ4NupuUK5gwmE4jWG2ihxM5TUUv9FhfBnrJnP
rTd/AK0r7RyzdqmL1yeZQUWQaFHkHDUckHynMNuGKcOb+1XvG0moLHjS4g0Jf2SK
eDlQolSpq6D35H8N1HBFmxDm2CRUVS8GPaHhlxJ9HivaaHr8YeucTAqatpWOL4xh
g5qlcUBJ4rK5NRoOkRmBxKjlEBo2Ay5HJ8aPrnyGz48UblkCOByup5K/w3JjHfyu
j0Dk0OxOgDHRENbtUthlNxNQ9gszLiYBXYiWqWleohoQodSyfEaW5HPbIltABk3P
bVkTXXZ2bwxISMthVE3v/hOlCHrCw1z0KY8G/pQl/8inzbiWDgDwaW/NO4AX1NqG
dmozqjKJfoO/euwTJSZn4+N8F1o/da2Uzg5k5yq0QMEymCOtgTQieQoe2vwNDNLF
EaMCi/xRtIn+pWOa5hvqBiR3UwqyY1Sr3JHyOaGA6K3PTuZmM/FMzirKrKq5y/Zh
ZD3juX7tvgw9XBFF10TVEGQQtM5CU5KrRjDcWJCdavSk8up/SGJJJJXWEADxm9Bf
vDZF7eg1/LgPOie00brFlkQp7UTeWMo/M8vJYIrqK8QFoSYLmDjXqHh0/iWYu9UZ
rBHZadJmrgOwOOs6nuI8W+yL4NjwacmoOWPintu/E68gWDY+yJugLcgx86aRlfTk
gW8QHcmXgrelvCNB8w3203z9TQlpAtSJAhNhuH30E2d80mEQIM+ELkuPEAu6iA8c
ALQThXL35gaDwG6dQoy6x/14cdRT/rCqlyLA5kHBnerPCUiRGHJb8FFtDkz0sgjz
jUhC+JmegpJvfOoIK7qE3HIWe/vo7hD/VZJ1l4W5m+oYWSgV/auhHcZ9SQ4El6q0
+8Hq/YNhNAlRaEnHnJtbMfgClEPMPVn/VvAQd1sEvZ3iLG9seTMJ0voVwK69JjsA
70cXciY22sPFv+tAxzaurjQJW53FUvl9BpCvS+lLTMTkyutlXPg7rbtmvHIQR7ym
9Tst2WwLE/AoEFkSCbuil6ngTjB0y0V3OK9zfLDav66Fm3IyCZRGpZrAzcCYO/1X
e5bY4Dq9l5lOHJ7aHQygrrXuP1ZoQyIWjR5ZMKcR1x1R1GibjA7cV6Tnk1QJA65G
P0uUALZvF3OvX2ZpBVwuzUcO8KAvJ9fi3eUJaqV/tsGaBqT9VjEyYxd6a/j8SwA2
B9pYUeG8TPVn0BBIAzN835S5XNlJIxq3oNb1qFf9spmQ6j3rL+1M4V8RB506UxxD
0n7s+W33zccteliXnQJ1MGpRNel82asP6EofcjCaClZT7in44Tr4lfVVXSWRHs0E
8Rny/0roRLAfxRpodNW6w/EW0XzabDkgygkbDZ4iXWH/8dsSByj2NAdbqM/0ORmV
Nhye8hqdIRCL1pK/yFlVkhP9E86SMkaru9UCLze+X/Yy4uDfxWl6hmM30t2WhxUT
cvVd8C5JpbBUw+2ajBL155SkdKCIabo/EzkgzsXuYb/azYZci3VWXnXtP1R4rW+L
sSxY5rjlf6tl8/ZBN1uERr+675v7MuIzSx4qmD7gt3u76MQfCpuh/T9JDRNw1Q8C
hYgm/I9bByrNmXY1qYOhkg+UsdpGagw7FzP3GeHo8/Xfk7owogUQFPPs7+8IX79y
c31+pfkbv01XEZ0SM2XEG0WuZ3BbAujpjQYRrt68J4lYHmKVjT0QoPXD5WkYHJqM
uMBujlg5JSqPGArQXZ1t/G1s5xP1IFkFy6xHgG+W0jExBzv4EOfmSxlylyFK6kG7
fS3pv/VPp/VJuwNtBkEm7wiDLdxU7AuUfTMdZGKeH+sI2xe09xBRvaCZPfP9KKbo
dSnw5fsP002EOtELg+1ph/432Bt2ITvrSa7FoKoK/EM5Biyv4XfN1sLX/eq5whA4
R4awCIRrWYj+Nu3bc0TpNMSTwl+xCsQiZz9wHrMQE8LuYhrD41zQHTd3Q0OlwMYb
8AIxbCfOeOukLY5CT7pFGYGFj6Fe+T8vpieTVc6WeiLy3RdpEd9NfnyDuxDSEiAV
S2Iu1I75qB/wWCWkc0n3J8hx5yXJUBDUA63JTnVM52g24kYJsUx5ospURxP1GEMP
ny8/f8Af6ZNd+WJ+zQmfpd09xEe8akZfU8vKFuO8l0GSWeqfvuB7QDAnFECWBoQx
htneYDi+8wMtiQ5Aare8jcWNZm8qa4/83Y0/r5FCceTNQGv3+hB8ITuUSUjoyATI
LxmnxW7Uk3wfFhDsoQrfQu/VQPkqYGz/YlLSKXGwNlmqXyP8Gp1QmRaCK0f8gI2h
0jnZKByB1m/1QQDaCi+tI35luqLzuzr8bAMEKhT+PM4wt5iup1Vi7bJLbIkPmh1o
fhBA3g2cBof8eqJu1btT3sYuLvdODWOmzDBeVoqQqAj5tyBJYcjACmyVTJaMumXN
k6BHMmyGoeCv7U96GSJD77mzp1ySNN3msDmbZw3jFNGElkso31E4UfneyPTIR9oB
B/j1ZDjAI5TjLY4QiymjsMRTjBmUISFAofGuWJannaXvgAhBItY2J3z2fYn9vabT
zAAPHKsop3OASK7N4702Lopl3OM/s39dQToIfOrvkjZuQrGPVtBhRHZChNdDv4nf
rwJf1QBgO6Spk1Zfy9lNZ0BEa5tSTlzFldyt3oxwrlgbRn7pXhb9sNap3nYOVkXJ
3Uj/tzZHHtCC4zWIlAA2KXjNAqpDERY9Te4fU8tsncryF0i3BrK9dwugOajxET1F
TxCtpC0bn3C4iS2uOfSuNmNTDAC4mpFPZk4/O1Pl7KUqYbNwLmxReb44d/Dmmwrj
4S4m50F0KHmJVO3hk/Dpu2EertDBGWfwI8Vc4INBntNZ4o1iwdxc6NTe1JkAmcEN
yxwrhjbO/x3TLSL4lI3pZv0Srta/DS9Z95yOyfMW5MAL/ONO+s/jXW/DhG0w5XJw
S8IttPdbtlCE56PmIRmE8RYSJm3W6BqY643+SYJsX3MIWviXfzM0Zi6hl9vI4B3j
VJQ1rT9+EYI8+Hf/JLvR3DoUfRHbaN6v9S182klR+CTqqn2nDrG02NtJh9Bmy6+0
AVFL11y8XE1E8h5X6dWl8wd7tbdbRSNkqwLDE9jGDtijTEqZ9aANDd5cUyvy9tFW
JN1E3MRhbBCOWYSJ3s32SdgkbVDub/Eigjmw3PHD0bIejp/7NF5vd1oR4Ukd149K
vyzP+bMCc6BfAeOhfD9PbFl6Vb13ZsMxVZsGiqURQ+bGWyYl/76ksiUVjD0+2Ylw
OfDbJOChrlBqvhD8iNwPJbxYmLjR9bApUFeFN5ip2XSSJlbCghfnnHO7M6QM7ewc
emV17r5y/Lf1ZzMTzBYQZLbiKTjMJe1VEkqGM44+umwwHdLBkglE0bVALD4+9HsM
PJ2XgxrNq5gWbLKhcEtQCTqJKLA4OaxWx1s+lr9vpPATRwY/zYli0mKfnebRfGXh
T+plpowBO2FnVBxkkE9wssP6E/q8UO8CWAFtXf0RYnw7gJ6yYi1tv8yEsxrp/iPT
kpgkwW5HwaGCf9EdsFt+wSxchgK/q4SU9w7M4CJ5uAVCFgtGx4J0L9p+FXHx4YnZ
cceTnEhcCyH0ZSZPYJ3O16tjDcNiCdRtR+bS3NIJodtdlY3H/mrLpbZIebjG7tGm
60TtIba1bX2qBm1vqyPlWeLt/Aqg551WdWvcd2CfZlJBNfZxt+wsw5PEWWF2ILUj
lsYx7aulJysUulFDiL7EqiJCbRvjIcfheqeyiV2tTsWlAQ1tLh//6xtCW16Nfszn
bKc+8lz5zJbDJeK5p+YywHLAaS+pyUWwzYeBUzk4EzBmXkLC/HBgmpLVhBoNjdwg
7OoxXTuLzMgOae1AkB7d2QiH+HBDAQfnODUPukC3iiXJbMZJ8+QS0g1VVIH/azRO
AB90pTZGn4NyDHKc4fvLpIIPvfdlEmTSjus7EjIAK2TBsNnjiJR2pWwhjZPBI0T5
RAsx+v6H3EX6OqctmheHkJ2BqcHpYtTV4tLw/JYmFUuAQ7BlBCXhLAc5j7Bycayk
XwhgaCCFl8h53h7vJTkeizcKfEWZNvB+8+axJqAG7Ggevd2QCKB8uK7jhArVaVSu
NAyD6gHeS8DSPX0dLGZTTVnDCAzuLPexq6+5wegrcNZYAaH2Z7DKOddCrsnIQkh0
2XvKpdUvDQwCltHLiYU5abS8W71Ibt+dWV7qRIphNHgajpRDmrqzexwzLtBbXWHm
pf3g85RaeBBb7OQhL9COmwixYYoDORbMKct5kC23Fe4mLwKnfKjiTqRksybmVUiR
TEcoE3uLw8xT5PjxyuMQyR0E9dpklaCCrBVAWDeW7GZOfKWHZ5tJiNcjFRUuBL1b
tdf8+V2KL03dzPYBJ1gJnYCcryHu4OWLnJ0bjUi6ohQZhLkjghIkBXkAOV/VBezp
XeLe2ftX5vJYBfCPFXKzXSRI8brE3NRwFNNlpmWoN9DueGXhBII6fCtlqVVogsV9
XJPUVdjzzEZKYLReKPGWn/1/IWdaHqQVGV0eWyLSfqhBcw9/B8chqu4WuXZbZlwi
Nf5sYgBBlnjRv4MFMs11waTq4chGKvbYSeTdIcxPlz3KcxMfaiMosQJd/tbz26tj
yxL1Y2gG+NvtOecwuUNBZb0TJwxt+M10wMVM13WSVGHD0yhqV1xk8rKY9iJrb9t/
LYrGFaDuAu+zsyqODIJxmvm8pljFJb611vWiMOPGYLS9VrQbbEdD0oTH8+oWQK1V
aYbEiYuG9n4Hrf3nqvz6DKwdZGlmTi0uFU/WKe058Y6F0lhv7QHaA5i/b+YULIy5
+mkbpkpamJz/6oI2wWUkpvztarbtjgJ6etdujNJU5V+DeNLtU8DbZ+LbHf0khURa
BuZPI79q050PMe54UIls4FWH1a3rKV79tzd/xVNA6zVSsWpB01dKhLF4VuLnb0GD
LMFL6Mccb2w5fsF6YpKbHrDaKdufT02YTbxdfImlC+GBvqrDn+0wVGYaZBde84sj
F9e8ZpqMkD/0QqpkOJlx6FEqnxPtw2aZLZCn1XM1ReY3xxbVNIm+qCmVKoDNW1mm
Vk8u5D/WyuKRIz16OKQdIaGkdrPqKFX7C+56EwG+d/dz4SH2mgNdqnmcft4tqysU
G0OknVGJ1NEAyqB0tGg+UJ8uX2DagQaZ2HVor/RByG/n4T/CTYxLOjnivYEoYyyR
dYuWOtY/SNU2vgAcvWK1e/UjhxvnUF6llj497KHmxuBcmRtbgekU7//Lb4+l5qY3
6Xcf0PluSxKo+AgkRVs8F3qG2xVACrCM7Y6nfyiIIKuMWnF9kNcfYwnE2lbH1Bda
0IFD3LPBcZ0BlBexQF0N22TyjXV2oRT4yZKst2L/WTj68oJeGGNHFikgqi4b1O8w
uu0QjILsIgg4K+CvCCcENG5UGJyzcdk0wu5MZWctcR8kHizOzOL6ACny+kzizoVc
wKOJPfApzJ49GpIIqbGeTIIJhWx2fjrtOtzda9fJhFUsUs8885CF5c/8+gbn4FJI
IMfbk5pfx7FqoyTmwVNYJHyaeaUs0jMUjnUyk3kX6hD5QyEigoAXT0BZ+ho30bSX
nu9rkSXCNaLdrafg9Vt/7rODLjcG5teJzDj6bQuuvcrM21Uf/TD0Hlp5SqEl/axw
eEDfklPYb4eUjC6mw1ezYtKOned8aX0FHCagTWW7dhAwsDJ/d70jWsoXKzccw3JW
HO/2O9KpocEj3g8WsdiNAPQWEVgME5clU4S0siCAiAhVlnuM1jyNm40QI5dL7MDT
fSJf/33pCAo9Pd+WoctzGyvSLYB4MLy3TjfDzrpigbyxR/77TpGKgzplJJY9u6rL
IjOugpwz0bJG8NqLClVkhTzQV7rWGVbsLSUm3MUAohEfeIhuxxOA/CQky3ZtP5E7
OhBeXRVXyao4ovcLXxIVg+m8RQWPm189mxjPsOfMqXe0Z0qtImpIRYoHBzVZS6me
a8rePyox1thHaobcv1QY69VB3kP6TCxS9bOJ92qfvVql4A3ySomLjmEr08cBemrN
F2fJGCkafugmvcGRZ1OujvYNXYFasuffHfYxgrAYVVb4qLlSmOTudtdRLSl9g6eb
xXSDTxCuaXG8joQYkFESyA5XAjc2P0KinnMKxeAfDClbsXypTGqObnVksbmb45yX
iZTq1quLPSdh5GgICWBoZzRTB9VeMQJj22CXtWejzjuAZPHM6/harWdMa+/T7+9O
F2Q+YqUzXWvczBAqeRRClX03lZT2N3l1Dh7og6V5Tflm/IA5Mlhk8xeIuDd+eiAz
biHMSg2uWaKSMrB7THuZjX2njVczm6SiRBHT5bFYTz/oDmTfEXWkGqf2MUVXe3u4
mzl4LdzWgTl0TW2R8g0V7UhGWdEx3tfYvuECCzsBOGd8gLh+e+3aS35lN8Od6cYP
3tT1Jnl/Nl/g3yaLYmNFflpWK+S0U0+5vtNjN1yr0hKV8PEx5ZA0ZRymHXI1VY7Y
CA7vaoX1/N8QIjTjtkcT5Z2OyxLkHBhpunrlC1yvDzFZ++R44iMT3ZOv2EGE3W8s
CBI6j4f3lb9h3MqM09oKMK2DoRqgJCy0T694xJqIa/7V5Gvageyi+3vfiRPDa6vU
Nblgjy6rA9RO41q8QD4V5hXs0WKnzPt80fqo1jdqB/4V48RfFLUNAzGkAB70y3l1
6PDfOncSplDqHbtpn65zLY87Ap8+XRfMd+664o5541AP9b0LR6tO87Dq6UbjyfLp
EFuPgWie9v/H0Eyfn+uO3+8opjRTCCjQI8NnNSAn6jJnTyatEd/Y1vMN3/sYv38U
nX4WOgCqQkoSXB+/trK/oJJA/8Usgl6LLCAaY3EB75XwRPUtbKKhPZCmXeHbyV94
/b4WQP7lQXJu7H+9rnQ5Xv2nY3uAdeIqxgS3pQ85icJOql3zMoanHL5wpFvAuaNe
7ct3S1+P18CuSsZJ8vRfs7L2w4mDSCrfqVDdEApFzIs6HVDIjsmx1tPSOtWNOcOi
fEvyf7JlL/AX2rOit/cEkRmm68iRMFjcj3E0b2rsTMbKw2CIFWRBIVem4CGG0LWR
XXsjW37iNn823eMAQJd/M+fbYBHcU44va0gU4gs+E5oY/adKbDNMtZSaU9kj+ZDv
PWQ62zspxDkC6kHiPLwc7WW3CHbTm3VzvNf4O1TlbEHtgEsENjmOOzp0F5f2Ejnp
T9DSBy8bJtAw14vnENfa35WBdRpDkZgrOavvaPBbBzW/PEujFWlNR7laafL9sYQ4
F3LobHJTjRVOHSWRYUusJZDRZCSSM2rI5TNmqINCMjcnjW0teJaCW8lhKX+A5fic
L5HG7GgcJ3nf9ER021opG//qiduAJ1IIogw1hkyV8ctRIx3N70odF2Nmo3DgBBIn
4sQnVFaXLQblzpcF2NbDHSBmQODkZBG/wP4HePQLJSUBaC2A4PTzmdUxY3275Yw1
X6dqYQk/4xKSg7K6attXFElZPmdm12P2Nfuv0mvG7WKc1VnvSa8k0/WIMFali1TX
wEuXqC56EctbxUlOvjjDaYE6Zao5Uhj/EAhUxNakmcCY4wjZtfaRSDzyN8hSLVcY
A/XHplOIV9hhC1gsAgY8kty7vyAin7LD0XljdtK7InfnSa1BEMptbaYpoWCiNM+Z
NPM+aCybo+HnrXKrQIj/lG427/Nfr4kI107skqnY6A4VNSUD2rbN8kfo4gCuTGnt
/wlu5lCm6v9mge2YHlWYvArp0yOurymec9OD+pbde7HL2y5YTeUrncrka9Oi8tI3
ZW/fK9IYwVfn3c+rtmrc5/7u0sWgNnTUIpTdfoC/l7rIWSya7V4QF7vXUJbQ3tza
N4JT3kRi9uLKofNN46TPpV9Tu5vsprdHC9k6/3CGCwxuSYeDwFIvjHAS682Z/bPs
fXusjeI21Xy0n0cBn37SuMTNESy+tU2WCPb7x8HMRJibtUsTfKOItsE+L6wf2N0y
u0DRk3AhudtH8DP0PEwTmSac9k2RpCiaoPnXg3pMlE8xsASW37yeUJW3AJUGBVOd
ykjCIyElmsVxx0f3OrlcdGUNv108FMgyhOIon4lnk6PpSPu2yS5no9aJPrdtXl+f
WFlI3+IBFkHp3a0H3eJNG4r67teugx2nWSQtXz3X4xMZWVB74dX1KhRuu65QKr7h
/+W6o2HWs9/dcWFblz33vtm17r5V6TqAPMrivu96TCLdgt3V2cBQ0lbG4vtfGHC+
hahGH2xBiWcCsfn7rXQlx7rRCOmPhMyYwURf1jQR5T0WzuUEw8i+s8KxDe0pvM77
zhPNp4ALPcet1Sdrp4vnw8arxzeSuvXi3mz23omqQFdvlkf+ObMAvL0JIAIg4T1b
QxbDuS6hz+ldYlx7Ubo97gidGLuGM6+rY2+MJqfAxUDlKVR1BcgRjBP8aIO4GZ8t
LzWZc7qnJVkz2Y+e4JzAC6mUMS4e7gkciVY93bIAe2whp6QTKfpuQaouJ16LBHSc
lxUQPXULgDKPoresfZyxh+yOApxneCN4FdIlKqj9PmcQiMqF2O1XnJib3biXtkZj
j+8CVC7ieIGsbuBgkQOPiHIZYKlrZCbfzshq3SHpfAs/56YsyIlFrZ/itRXr4q+M
CzDXP2HqcXQuYkrUw0sRHRBk0Aa+IG/NgKMJ0H1T4EzjQiQWxsDE+w+PC3cabJMZ
ebses1YKahjfFnSAMVx8IsrWWpLZZYcCXVnTP1FKSYFwFIqaVgBpP90ano+KDvoY
VroCXWX9FG6lsXoGPd2J6wXOCjKni15s/mAcbOQDQU88vrK710Qv15xpgw0BqD09
lKB6673mAnJtKfqytWwBp+u3DcnJwksl1UKv0i4IRdBJ7lADAn9t+aFaSt1pVZa3
EjC/AfCKW+xkSyyjuxELlabaA2NR5TLDx6pE8ypOhcN8HutcE8Pef6eZleNdoAaW
1g5eTttlcui8RqywSsKlI3FpqSLRbYUp1deMV1kzyvgLBJXJuLY22v7vfHbhcc+x
gCY2KAx2FwyMWw9vktmpXF8vqqVjJwxlJQshCnWjGi8gLz85xpl0PF4giaNPLCpa
4FOfFyGCVwjrTUWvYMUsjeYLnUgsKj9iBO71C1nUsv42AwhWZIdCUyBOkuPvblr5
NZv/F0+svEjfacGO11aajz6o4uCFH5aFvOHiK9XeHN957J1PNtWArPp2USESToE1
1f/MfsDfm9Io3wg38aNSzciLpFyeZHnfhOeLUX+yn5gufwEHIg4Rt+0dqFGiKQZw
beksUqN5Ybf6LQNDj3KrFs+tS1J1NcsmaKiaWmgRYzWVFYoxNilueNX5gBJP5yUj
eQ1oeU04O9KgYgiKesIdKbWLRT0aiw2cpUE61DA07YqV8xjs/DGUV44Juy2qqfG/
+muFLCoPwrNb/N7De9lVyfN3/bbStqnzmrvcHiO3/tBoLy5SlgQt7vAUfz4UZU25
b/Xe+M/EybUmmlOLcCu0Sa7A/SOVatDPyS+zoH0PszuP0VIP4MYgOieG4ZY/TW5D
jDHhx8lUnslAEA+0vJSg1KlTj0rf55e/4s6I7gIJ6GjEfBUa6eCx412w7dQDEiiA
H3bz4huqN1H/+vOftb6Zzz6hRopbGsZUrsWE9xKsfJcayMRzb/SUHDv4Q7mpRha/
6ViTA0+VnVvJVrM9MmYOTCES42ee8NnYpJy3/SzUeLwiJgnS1Otq7EOMT2euD0YI
jPrRGNjjLIiai4xMfcPsh2sFxbA73sLFzCRcBJtP8BmrN0RW90q6n11p5ka+Jsq8
A970shzClIrpWfXSDNNB95c8mnhWxnmeFbot7SGtXtnS0kIxhoyBZO9yHU3ikLxB
2QEV+Ow68bBYdKD2eP24JqWDP3PmYTXWidzUUEQ0sigvCajA0dqPz2gFoMIR3HLY
ULjATAbiP6p/UdGyDTF7ZOB2oZcc8o6Q9YMgC9bJAtxu1rEo6X8yUfbSKsON4/Nl
y0QWgIRJVuVlBoaqlKYRrYHIImHa+slFJndvRQhw9h/940XuJx9kupB+thbSKbUZ
Lfgr91WVf/MduudyhXLT5nZBEK6xHVdATfshrn2wiFq97YREK3rpfeUQBT7X/ros
84MM39IEf5KpoQICjJH9vNs9EMbXw8bjpn20XG9x9WTQQUXvDFmyKjcHi3itGLAT
J1JFbU3Tb+FOBd4C9WUMgeJ0KbS48Y/RiTTmIPoTEqIa3k+ayFNGu6tHYRNn+S6L
RGrjybS48BaL4s4t7RBAl6uLLRxB34pVdVcwVPykD1ATcxFxXlnAqXJveXsFURu7
4H7oYA4I7spfnTW7B1/BN+Kxz6vRU2sHPB3uCNBxtZG6Tr8iEBkVOkvn2Po4vV37
BMUbvPCsTYiwyBdRk9pk8sRA49EH5yAG+AJzhksXaoG6TOO2LY3v7T+YK/TM4rHk
W0F6h7h3q2FP7/Y155P+LcWjIBkZQKQrIP/Ly1MI8ywb1EU2arrebBn4Kt0+YelQ
PfUNtYqDBOGd/scEz7+FfErux1aSJ9JNVM1U6GO1RLgiGEDsjMxs4q7Qa1ouVxeN
rEZEE/2t9E+kvwfviWhxnAVdvggLisPEW5gil/Vv6NxtdyV9W5XE3giRBOJ6DoyC
yfw8dmwxrX3pobzj5cBdysCXwheMzDjBccnyqrtlhMlfruVCEdVEVpttgaXfXxAZ
m4hAFsqNeYpEk0gXR+NHELNOsa6ZtYkCwErtC3g5c1x1/EAeDm4/1sDoQrSfkQtQ
EF0AVXLGMgjTk2Ri93PL6EaBTtKeUSH5+ysw98p0tmIyzP4UFbg15WoXVmR5S3tK
/ZESfFhMmKOspTjwdIZztX57ipZYn4fOUfZE9FUcdR0zxT+IwavOedUQDx+6DEjR
RBFkwRnDpqWmLNOcbR0HnJoxT8CZmvEn0VvT9MnzVLVFmC0w100RDmW1ukRz5Oi+
LheLKgD4hyLf1nXQVc69oUzzj9A/1++6Gc4uSyH2lRGIwuCcFrrh0ccyy4sJDuSC
BJGBYkgFnO2l/b2XYkt4wb9Ui+hzpKXAY+jmPIH5fCim2Mupwjk7jszg+nYrRb1n
8LkHeHF8MdOGiRM1DVya6/b4iUWwfw6Ok9ZqoN16qjE8agJ1I5neWXRPQwiemub1
FSndtHnd6jtCabg4G3HG/Lqk5BoPz4dasCRrMRhV7FwiH2CZi+DuVf3P8skQSvmb
4Nx0C8lYBNLzOwavv07mYIh2CE4JgQSPk4hbIylk2fLBu011evxnlCn70iAe4Tw0
K5USN/acrOavjU458Hi3z7fwBHVbnZRqgazVneT4kNyJcavD4yjHUhgMdT1sDpFG
vi5OQe8UEFIrdz6+GGc6riyg7pwSycSWBa9EpL1AMAlGeDF7TbFpwDYgZtvPj2IB
Fbi8ZTzi1HfEenHdy0EHoso52WY/AVm4qyR4KbaXmCJCD4+eJQ7QtM0qkL0oJ6jQ
MTQmMS9y1W9sWQCtFsKqTBEM0YFbL4MV/vTz5L+ghRgYiOxhrfIFOL/wiMxju/ik
528gIY3TeYJ5mJ8nNljpt5acrDqjuK6sLmMP0hL4NLtk33lNwvMPymy8gWxuZU9M
dEW5iYPsbDmB7hqMHz+5JO7LvAv+07chYSOylgV/e8mcm2eGuhZ4sJJwiE1+fc2o
1yt60Vwxr2aVQ6NkhRvVs9MImqLs6FevQo2jA6Pl5cfZ2zqacf9eIANRvFqzeE+0
8hbKddaIkH8elCMG/TAegzyszaAQLp/h/mkIeZK17AqdBO95a6M5dk2REKb6CnH3
Q7vMYs+GnhnXpf/lVNOuxrYEpU9eT0/nCRh/E9ZVuFCPM04zqPDDPwjd1rbWTDzx
7SjUcPKtsmVsKaGQqTQx8Tic9kTlCVzQLiDmwz99fOGu7CStTczmg5FFEUxgHJQc
YZbY+r0ksCf4bGHXin0eP72I0/jtELiwN+nlAOwkLculrP+ILp4rHaYwycbPv7bP
73oqY2OCqCXTf0IsQBMOqmE0gZwPB5PGjsDCRwQQpZxc8xP4WUmJsCUDtTt7jAUf
NjdoZ4pgl5tdkwaGSXXA77uiAc3UYNka8+LxZHoPIYPIZkuOGG1YKoUgkHjXLrDN
cXf8fZlgPLSjD+EmJYQ+NCv+mK/Hx+3Jjh9O6/Xh0y5+UDiyRRF1ofgzMELo7J6q
7SrKYuJZRm1l5G8Dzzq5CfJ01fV4KinCExKuGbrFpf7zmTu3Q0CHrlSPSSRIn2rq
70qwZ1TyIjtPXoIAtjKdEpQAwnfJmBOYADnmLva9q4RJxk/dJnh0bjrrX1knuidY
cwb9CaLu/tGPEjZqOFIiWgXBCk4eKm8ckxaldGYigrq5L7FGVL1Kb0BTRCV59ym+
y42uoxkjVYZQ/c3ov9Nk0CIqFPmbUfSY6QcAAaqw1v8CrdXy8vSCRxNWc28PPOfD
2lfU2QJgoct440UAZzr49E/izyPVMqn1MMNa4Ph4AK31sb8D6+cPLxRhs5LSErNz
YUymnjGNi/aoWm2i2lLAfM/qMYpOCTd8eC21jj1EBaLv4Q6JKFjAovq4Ps25/4/W
idPQQzgCwaQa9mEs1s3PK7vVA5M+zZP7Pzf4EHt17rOcED4dEFrtQnRu3EcDqHgr
LnQ3t4h9kvlRvWmSH0TeWoUTN5szcls2YwGE2ga61YyN4u/qM0kq3/RHKd2lAEdZ
7Bjaf+I8nY7GMDh5hLkxWaJZTt8rENH22YO5jMwpA/Ie3lf9FZ0Wk1qdn3JqsO4T
J1mnK/Q0wuyX4U6N4aoKsjmYiz+i/mixKNSDbPe4HSsY9OyLX8Xvj0uYUmOR6Htw
IPdv+ef3hsGY+NGiW1vG94Hioh44Ap5QGZ5slsqu6zPJfEFIm2xlKxVh5HdTGQFV
T5gt1Vi8dsjZ5s3KBwINi293qIxFtGw9/f4xynXp9R1Yl6b8bQkU+cG9roZ35aEu
b5+v4vEikYHnqQATFCm6odIGIEPWVbam4B7SHITmgNSRodG8mczGbP1Rjt4Dz7VZ
/puZEHrzCnzmopef6nYEODP1w0tB83M+qqtWvPBjNo+Lo+WhGsytPoFXXUpsMN4V
iCsHP9aAc6Obn96LqE1AJvg1AF1kIgB1QBwvMNRX+6q3DkhKOKV+S/z7sZYlkWJR
fxuZlUT1/8LJrdp7omh9G1t8aelYdtb7JkCBya6xFXqocB7zXsRlcqF30+ZBTBZ7
vJUzTRJ+EfzNywpmriu6VaE9dvY8ixCQjQ5oe9FtCZDOoUJWs/Gy+Eq0YooYHwOe
FALMypXcX3VSkOLpRec895/XHJ7gUJMRy9K+Lf7HOZjYWIVL1v4db7Ns0XSJnroJ
3onD905+HaLYx1IOE5z6VIo/wsa1cqIkz0LQ4LJpcJO8TQcnW1AKGcgPL2fyjtj+
IALQ2lfD5rJ4Fu4mu136HAzyhJM3ly2To1rbJJjeQ+NMoP9NJ6NyJUuJgSEPaZ4D
ucUF3NG29atk543mHEhrc7RPbSMHCQr/qpef8Ugi8ATp7PHBmmaiFpV52UCJMMK4
BomZM5fcj9Fg2LsOSh0U1sFQpktov2Q9NMPK/O/hPKBTq8aKnw5qAYcX3oP787ce
CkznVey1C7N9wFMKIQNv7M4eKIkmejz/4/cXt6TREdoBN1F233A2Dp001X2tBreh
HOXkWHG5HTezduM6rHI3ezmB0I8/sScJ8hv8vJDdvHWT63iy1/ovdyRIt9XtDY5A
y/Ma9UmyDLJzwgTdxEopmuRwtvcdQros3g6QI6svzS0k5Cug38lgrW9/pyupCqBc
i3sSnfJ5xf7Rt+DY40zbYJ2KBmTgIZirendTX3McTR7oMH1l14ngux8NbEZrGjJQ
uxaX9/6vmNvyaJq5cqfI9HzeAQav2lQyVqXKga2BwG8Qq3wydTju3fAzR3SzyUaU
UzEk1nhqBr1C0mY2ioJFHHWkELvgGTISY2CseIVoN5fKOIgQKjbfE5sYdcr1MnXw
saeWeWHRSy+KRzCKGbopVzjGFv0kvC0jJatMrqVBJcFdBSaEydy1gFt7w9mzm/Ku
2lWaL7FVU/9qi9hgYIy/IeX5jXs/NGC7bJUIisIID8w2rgGATYrbNDrmxt/4+gb8
Z+r3a2lM7F98pZh2iMFVXIa0So8DT4M0K5LgnmoR6+FL915nASezsYHkzbxJQv4J
7PcZsrgXSiE/HiSoFJlbQKEbI9eozuY5bLrVAoOaUe7uX1vlFbYhpWFE6sDjdiSr
j1s1gLu2iYVqf25VuvQvk3OKc/H+cb1gBMKJFQD1g5kwyxJu1eFlKVHO/Cd5+e7a
7nzRo7L4Ux5HhNgyF8fSeeozt1Z0fQAV2XJ/JH/t7oiLvL4WHJ+ocBCQQMyWkD7L
W7ezf0RZGDcGhaJRCPMtIa6WtfzfBY5BU3fkeFE2pNeCNGrRlvseW0KhyrNrDtTy
9yyvzAu+3I3Ndu94xpZr4qHZXedSdWyA06kKahrICM439BcNNgbEAgcxmqoRg00X
LxxrQL+bb/wjZD1fMHBoIdlzfCjY9GOcPAENEXgpyLeykP9QvQZTGtB/YVzbTgCq
n7b7P9WgqnhfXkRlMx0LWrNK6G00TsMNOB/LHKGOuSyJIf4eL3iCOK6m4FAaYo/N
ar3rILp6EO8CN1DTIccPHiqr2WAvPan2/i8pSH5/DXCvz73qonppE5N9LPEbX6z0
mr3I4uyVVq7iLqeFy/WxJNRXXV55laiRvSb08bWHQ+83ZsaTpa85gu1T6J7iVM7a
Dyu3zX7+WGkft8dmINAiQecPpN5ZBiANrpnopjS7MA8890QKIQxqAfTHfbWyTvDp
rTi+4E3h1MdxR9uFgQJMcqlejW83WHTXUCHWzqNlXD6Ca+9DyQTjubbu++aV7xKg
lOleCvYLkZbSZIO49TQL+vABqrYvfcc1lIkp0GBw7GGDE/0R5/qki+pHLDtGU5JL
zuoGKBTx/MbNsmNuDLEm/V56th+fUz4hxhrw/YzBt9QvLji5FYhOzS6g40sg/YB/
M3fgF3B9XIyG72awGnmuxJb0RjM6IdMpsohe/ZX/26o4Q8hVdmYp1T8QYI9CegYB
NoY4+czxLTjrbHeQdCAvC3eIEbI9GnWViEooDNbTjC0R+urS4n9RGU5WZYl1CrqD
gZ7WC2qXuCIK9jMdTT3gpQ0pgexCKea9fsAi/pCuZf2h0WpJVM7zN/+dp3mMFXaG
mxKIlhWK1vIdFllGLxUZjcHZQRBTr53RpFpCYCSLvBDbB4zTlZcHVEibDutRNhes
HL4B3Aig6sk0c8sxvLIXRcW2XGFv5sltQp3+eY97aIJo5VGjnAQqvMaPh/M0xFAH
`pragma protect end_protected
