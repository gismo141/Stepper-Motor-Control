// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:49 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c8QNFRXoxgeGiR0kGU84tfj3u3Ik2NS7dZYwhkwBPnEip+OAhmNdmOlpMWAtWlt5
UdcJgHeJC+gPT8uAHfttzLee2HVnra6zksxlGmDtl/KBxj2Khq+yECORfvrXtFb7
ZSmKT71dLakznsp2I2b4vvGgza3ohui1MVoVZz1CS8I=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29360)
9WbX3tbgENHwt9wcs7eBPDHCEGBDv47OVxsizf0/91QTCp0defBo/dprggaon9kL
MkqGXpSR3sjsWooVo1DJhYueKBbCzE3E6VOVUK2bsP0dYvUh0GXuhGy045AJNzif
wWtWv+Vsork/+kEdexESh5WenScdhVY0h3IxxkDvTcWDFL68CgSUzTIHzwVxJwiR
ETgErf+ZrzkH8b/cFlGCcIwykCVkVBl56ZSnyJpU+WR0U5u3Dn6jB1aL+4hi75Wv
HTL9I7nlZIPkwbpm7NkJ9y4ancpgkc8Xx78qAugF3lBKB4+aMNobY2x+WN/1f4nI
/FyHUQvJMqf/A0h17o5700JzeLPDLJnlD9asg5LpEj/3ZepqWXWRQ6XwOx07igjd
B1eQ2CzHRJxggEvbi5wseVQbZhaIQjHJnYKzSvxznAXZh9mjinr4EPq6dSjaS00i
zYzwzTt2t6KuwXnsuYLEyAzcn7gXWRm687GjZECt/fkm7dnLJOWLqxyqif0iO0k/
ZVy196ZUerJTjZarQbRHls1LZma68IM2vnEAiRwORyb37EyWZp7vzefVt4FS7EeT
CPXXspH4dM3H89IIhu384TuwW4ooOlx4qaCTVyub29+cDHdZ/PawFOIRwr3iQYC0
KKzQnRKnA1r4P4DqDEGnTpZcs8sRkKUNg6pz3zmwDRrskrn40L8JoEXpOjZ2S00O
5JGY0T55Dcrwabf151ditTf16I+uov2fA7feozC4Bej8pQudXk3USuo4NiFuN3R4
i9GFFiYEJWQk50GVCLZEbcxNRUvG6L5DDnwZupDN4Lwzc6aTYX9GGvVgX8eRK32K
yCKXciUmZGJTm2N3gN59KplXRpdfjHTlTrKtVVeL950loCVysFW5aU73NLqeJ2zA
ldwDdRskWwATtAvjJhxrlaGh/u/ggo9n9G+/g8aCGNKFxddloN+M5xKeiNLhiRlv
QyRqHicMhCd75J1hE0aLnlf1yx4TMhOu+DQ5rKCQTVRnSfBCJ6vIHC3aB15+Dxgk
96YXvHxpQOsHBQhKKZ04dDT5GvBtmKKL1+RjYF4IkgeqM7Vgdk1Yg7DVzc4e9+Wj
bRX8F4gFDX+fQk3d+yUg54O2aTWKtmmbMuELdHmlvg/LcfGYzTs/Lg4oKqvshzoQ
Q7/rfzsfm3jIK7lB+rqCs759W69kdFqzZKt+KOSD2p+DXhzsAjZEEjH+9AIk3/Bi
lodchBO2ad5kG7b5cDKQDbj0qfoWI6ekYQhexFyGo92A7jPGvGR++mkV70OF/ERI
tOQLJJXA+sIE/Pz7EO48Frq1GcKnSyECf6no7CAvCVelf3h71LKCuMeNib25JzGH
J+3JeHzI6FfdTzTlY1GsL8e/GM8PcmJ/ERXbxJp7KE2GSyww2BcNODe8ZV1cegdQ
dJUdPnkqCxSJL59FLh+D04KRy+qC6vBkL7Pjn7ynNYo0tj0fSWAT7YLqrdQ9Jtwb
494t7JY2hFKwiamZLwXtTKtDQuH34D+ThUg4SrKDpjxYmmuQ+sFlmR7Gp+XRQFPa
yr8VlXNgyDvb6gqcVe8rjskv5Zf//90rKiGIqMO1IEAiegU+SMO8OzU60bbg7FWZ
sBTs7DKvVZVSrU7EoVu5sI4WRCuHqeanwtiD9CLEQN81ESPpGkiTPB76D6LGIC++
so5Vml67Lt1IbECX0vNMylaZz/Id75aJT1GNGOXqOwbR6xQDO+W4B5d8Eq8gzT9B
hnbV0ckkj8W9RlYGwz98bfM0chS7E7w1ayElz02Uds+Zag1kCedUYfjoGWmiR0xQ
iUkM3CalEIsa+aKo/nI2G4blv2eOBirg9egna6GQhUMdTaDRqxeFsopHmonW06w3
J37qeheU2JVzySPql89fVzGa5ZGUIe2RGZomHkAQgJ+MJcxa8hl2NqGHR3elfBbh
n7w5fLbRsAaDhSjUTPUvWeqU2NAyTZPf9UzjeJGjv+MCnVB689dRNp/tph/02dej
TgEoW8JeskuQjrpUDV7s3ROmGcVJ7s5GbrJgqda9g59Dr8gyjuMJ0KDRq/FT9W01
WTK+CtAeANiE4BiZWbGbk9vQuGPlzuKvzyd1I9pDPeyL+iH3z5QR7cA1eaD9WSOk
cpprJp8/2gjYwaqggBxRvxFyom8ItcRTLvrqtUQAiZMmTtsuzMds1b+gEijdS8Ee
lmcKCbFk5kEaSheZlQ1kfqRy5ZtcObO7ejHYfFnpBmDBW7GJDefTTE4GiXARCD8M
X7Ug+hdpRo1WHdHZ5uO5vp0cuDsqTA+q06n41ipNc/jEwJDEn7wOp/ujX5RVnaqF
bixEaFkY5qQug5LN2AkiUK9d0BsN9w2kOUELq5wkZtbRNY7OhyXNtirnIqovlzet
5zagndxplNf0lccYETkT/pEfCrCokozKb0ypFXgpOCIMylaYmCJHLanMVerliqDq
OkxvtgImzOAEzhdRUQGM3MARpYyorV6NXF9zoZ8oMzMRq85oaoJ1Dh+PhK4ugiDs
aJ/ue2FJBfibstk0KnJs2Z2u3aaWlt4Q33GytrckS59sDYHAjtoy03jYjlJL3gqR
J7bJr29/Qq4+PCoNRZ9CgyOLAxJOLIjfbIorCBP43lws56UKhcSbcztdkk3aFWaG
zrnkT7a7h61f6urT4DwHwvwl/xspnnWbYGHgo9HXTsW3NMSt4NBIU5hTlSpSvGbu
3t52tumrzeDQ7cwkM8npUC401dbIlfX9ZbeeiTNswY65y93BNoUSwCSnL9vl974E
sRL8qfgAOw8i7bEq1hKFMoKN7lGfWOojGyQNyA9iLJX2oKivgAJzGtbrHfhWsj/o
3f7Oy79ws6VRkrOLcNY3tDVG/qHfqk3HXyH92J21SK16EeuuSl5TdAbD5pIo/2O0
CQOLrPv4oXpfURw0sCN3XO5g4jm6HxyCM9V3p7YQPaiZU8Ff873dI9f7HmP9JrwO
BsE93/dbRS/C833aP/DSdOItwvcdkIu93noUWPTg/3RH7pHOH4BOB//kGsxght2W
Ra//v6p/Iz8PhFn1zB3Jnd6LHShisBYwMnw4TdYlyZ5ci0K9Kcc7UIw4Q/BZOZLc
/9lvGePjkFhIXxr/CdjYccF6sbr5aC+1OGBaZ6CX7LZfi8Obr8ihB7ZUlUTHODRG
jrWAW3ChR7mdEbAkT5NI+Ga4vh6wbczlqPZRgthB2rQMPr/UDSjx8fM2c3d+iuaM
N3GSjT2M3Za8kA7QmhxXWM4couIgFH6zVa6Bff7mp470mfFuXzlLL+SKRxI4nu9x
lLXdfcbISUvbxtzHOxUQDA4yB0sg0+G81nGpjMJqG5xqKBaSTx5aa3sI0KO2ACmK
lasY6q9nl62zuykWgKOYfNXaFVDEOqGHZ+/6+aZ2qazD2D/OWL9ZXG+mdu2hHmEH
9BSEy13Wtlgw99PJ4YzlabJmJzhnp8TosAKI4wPRr5vMOBgYtoFPAdaY1SpYjWyJ
uNIU9S9PDo1N7/dJ4kty13OZCtTfQff38Iwhq42pwNWzYVMi1ZyS4BF3EYgQFWLE
fEoo41Pj2GlCHq7Jr5JSkq0ao4FVO5ksYiHGFDjFXwczdWsXve1bwE2yH6HqLim7
mV9LvdmgpWIW+WNf7rNqdM1PAjfLLvSR/PixkBb0NrTEB0epCFM9rIbj2sAEsJqA
3CwZXuP9i0fRC1AiaCUOR0oPGS7Z/T56ZfUvzxtl6NwMgnZD8YOyDUksDhpMRmPT
RrU6SIUSrBZHLeUx89nFQ5uF0+KndABgV6ksmrV3vNQVrb4/Nqli/w4f3E39BPEV
yeL/zPRwXTpOShlgfwP0WRn93Kii7ItUT9fxrGFvb2PhUrwLbmcvvMtQQeD6Agcg
wAc7VeEEd4l6EijtLJfw3CYDIhhrXOM8ziQcqV63sbLcNnfY+Yb+N2aCSeutz/xw
DrClq8h5PcJzvk5cd6PjXCy0X7obMIkhBGuGiyNILsrN7SxA/OvIu3e5Jia+wWek
FloxQL1qm6Cnq6rM4y0dBiWSZ11JzpC5nwX1hjUnpxXMe27V6KzOABTIxtsIe1Jl
zCo/yHl3p/MIYLe0pLG+arb3Pp8yq+gZ9gz58u3DLDRud72jfx+yrEodJOWD3dPj
gF4uP+CZjahh8Qccj4ZcYV38Z88ucV1PsLnTCl+O4py9czF2tPOq9/mF8EN2CNYK
q3vSwumWhA/i6VjG9wyg49ITIXUQUPifGHzPO7tuJ9Iu2uC+SNESDDaJx7scLeGA
K70qjU6td79ExUivx7u19r+UPM5JLCsLNB3kVF+NNsMvAcHjdV7m0NfzeuffisjE
QGmPfFo9mi//tFd7IvwcRQzcUNq8kvbuVxm3JRtu9Ml/R2qgg9TJnbByunXa389E
LVYBPdFnURtxQkfCCXsH19UZ6EydCRTQ64Duk7sj/I+hVJDEJGU4i/aEIhTcRjLF
uP9F066j3O/WhBni4Axx47IhnePOTxestbCaoGs9SrzOoN/JVsHPKX1wgcFPvqdH
nMooO6YAHVyAeB+pQ5LmGt0v3CxECgGLoXtPeql4DeLqz1j3Ho/gKRNLgrNIXoT7
pt4sy7D6jieOaHW/HK1NbNizhVKPlAadbUeRM/pGzOWfMmHjXxEnH2wefyKsJ4CP
PgyUWpqtGQ9iobKuBHTIU1lTMRtzdVJZn7F9sJfRL6UxAk7RozXeDQxMssMnioFJ
aOBQUhpqSX5ekeZpxQBWpooXQjGNwDRxqffKWMzJXFnbK1pg8yJa05ySHQPvrfHM
Zyj6mK+tkiMnrTOZHtRvCvk/uohQ5Hj2siHJyI1C43wFci8fO3HuUYBDXeazbG2d
cNszWJ2saLzeToz2SVJmO1A7O/NRL+jprLH8T4QxrCXJgtsaCUBV5CQf7xc7ee34
aBSXuWCLUn+5giBhak3EUmtvxXV9t6SuS/PLH6SChk4uqnGJJZ08vm1MJjycCtUC
hIJ4Q77LmXAfrVfo4/LDq0YtWKf/ucia9mOG0+aU0oc/tU56OnztdLcwPcGIpY/A
p1hu6yH59oFWUAXX5uZJxhn60KNKm0eFut7gAkHvi1+DBt9+bP57JGiloAAa9Faa
2970wYlZUdy9gE0Ecj8tBJJMtj6zeboOdbNFmiWRuqP9Xy1aF6cYNuS1uaBvoveQ
WLjwPPdOQO0QPieYYT6xlzbSk5nALQIRw+7oqYlxEHmaepGGwp/9G2ctvu50OTO9
FzC7IqeihQAT+hs3ySCY6nFw8U2pqWtGUqxI7rZAYcgIvhaBSVGwX43QyNi4qFHl
MEfmWjQPbp1I8Nmx2ApT2PkANzk+s3zSNT4iDxJiBmXByQYX6iW+JTbHpVk9y5p4
3HOQAdkElgTitkgR7UCCziBI7pGW4I/MO+oDpzTT8FYBTRlFL+XNmrw0NHUwSnEV
WSgMQGPzjsYQnVxBMcmBN9/uogSaG7YKeErno9VsKHaU0LERPGlZJqPZ5WhGDhxL
v9yOwga0D9afLmEfvichwTaVHa0ZUTxELGOpjA41k21sUqjCHU2avnoboUxgDdQO
pWWHEw36w9n1nH9kD3orHuFmZ8FC3R9vdXJbPo/5FuGesWUC5I4QDKVB3qf6j9Hv
K+ozqdl75/KT7vobVQMP7RQnaXL3HNcTz5mmWQ27pWlQJ/vQv5Jdn2JcBxeFwCxd
JlSKYPRYbpPTPr1b/Y7oNYx9NWU0qpfTDsdQxwvMVZch/H44CRWxvm5g9lwb5yoi
LVKUo1vokQcGU2NFp3LEgkyOxgPIxqkcaxcpdejtIH468xqkq6UpVrXLe5DWal4O
45qEmPV4iLys6Ip/0SJOadRWn6us+xMaPjWNaEduTc6ye0Oxe3PsP+i+FYWfMUzn
8VZxCPCTyhtlo+RdN0XfG3SMK5fWJLnlcmo0oumlIY9NZRlMMjJBne4FaycdnXyh
TbsJRi2mQbfDXoU9WGw8mKwFfLTFs2SZGErZ+7y0AH6+ycSGpSHiUKxFuJZ37Hd+
6A3uDBc19guVj8X6chZCd8S7JrklZ3C0aONVw4IvvYGwCT/6tgnKbi9qseWnbSd4
c1o70cIvGy38nQXZ0REw7hUXWzcYW8uv2mMI8Qqumc6ojlFH84CxcCKXdlnahNyG
7LshfPyxXUucE2HcMbhxH49njmBtYv6gYnnBEul42PEQI5+YXJioHHvSSoXgu9VR
QzptQAT3sAZxWPCKc9nFNEZ6QpBz1sLikLU3WmzHnsSo1uPkXNyHPdtJsbRxawsE
5pI7DgaoTPnMuZnnUhMzcWGkj7jo/0NaIX4Oux/rMoY7QjROh8sNBj5451bcH1GC
cwolADGQzMzY+Im/TWmZYQE6Zcg2z0860jA4BINtFdETesyvBAq2xxgI7zsuSAua
EF51WdZBpS0vdN2mgo+wHWvsfHIn+eEAPX8d9uvIQ3OEyBvp6saNCFFgCD3n3Tgb
VwwqDdQkkNIluHndN0MUoVBfl3qHp04RmGmSZlJrT1b8ZNZyoqFKmW5XNnJM8akU
PsSnOj+lScDLaL4OCMszIZ5AVr1ubMYPBRHfqQvc5zLdnJnOs3pGq1rC8XF1efGR
94r9l7K/+CKqiALJE2Yj6Nf/iCZBFefC1Y8Q+VbTQElh4tBECpP/0XT/f6FADoXF
CQR1Lala6Mtjx2JS6D1YVs2CP+6+Ke8tSCclR+RR9YEbd/pT+A3x47Er4rdVIbss
qGD7cfof6AjUPpF+DyykWfTNkoNzQCjY0qm0Vv4JFLRblq+LAGyt5JJ9896cUVYm
yn47ahaKoyDDEZxTk9WBLOoCk+jRr+EeC6fzly83JnPb495z6zhIIYtOw+7FNQa7
umAwEqcb74SiJFfD/fJPfC61QzsXAaWdqvWZ5KtLKdfh9OYRDMGflqWD1iJsyMBX
aGiWuGknQO0DAUe4uFGqA8PAeZqn2+6VccxtIWId9C1usqPWmjBDsMDJp9PuL8Us
5Bbll9ysQdtq8wpY7XeeeJShzY7zz4Thhzu16Tgjj+peJaK1rRDWY2wFK5ZuRYSt
8Z3JJXjztVyPz9JvTnbzWCuZlkf+i1EGi5lIvU18nWxaQNys0YUwb5zOG/ivQqOd
9dQ8Xf1CxKSgcLS1xSvFtq0xQ5D04Sj0cRPhA6OpZgz2nX0ihr6T1iJ/vnc9OTVG
hWPWjq7YT5veqSs/O9ObzI87osfSqg5Ghr1B3bl1LABPx2AGgitbaCpSMfkDM5hM
0i9wlEwqFGncy/iTT6C79A40VQOzx5YYA1bbVqlHNk13664Ov0D/+r9T52D71W7u
CidlAhUzHUqenRQHB3A4ADorxDp38MD+YiB72HqHCSX24Qq/Dj6eVPB+Qo5MPCN7
hyWQl08C0TUfzbLA1tYW5KYfqqrDc5ZCYRVTtrBJj4oJ2hpNgLxqXvbTMCjDLSLj
Z6LMs6+6HaFuX/7k0gEWiy7IMF/f4vlg0wK/dvpHDdmEgAeTYqRD8xDNXFvfOE5s
5V0052KTUZxDJ+AWbSlWorElfuMcTosBPkOY0qWg77+KwWiSVedGpcGLZZlBT9yQ
zCsbhNdBRUWaQ5z/rbyDZXO/t6qhTPF+vV/1GCb0skh+95L5p2GYEU5HkfC38RDy
gLcxzlLkjc8cd+WVNBH7DZZWX85LBrOsBTsXrOF/8C/jWKUCbCixOXu5ryVaoa1N
Gef3YyjHl1TL65j1psmNbz1AgCMHlgksZspffCAyTM9i6Rqd+QV8fJ1rbF/jMYF9
8dMHS3qFJ+zWyCTo7LiiJl3ixBuPyDAoieqxzOxMddgvMlE7LobteHMb4Rtlmle0
PvXT3/9IKxM+e0XEbT7z3UV8Qqt6akq2R9aeMhpVv7l8GEdt1VpgZwojKpPJmLLo
BCkR+lcM0q+y1LbctcQxA6/K6SsibvfbEI7OCNO5jMMkpKDGMIcVDRyzJWlXzAyd
EH/T+7Hi5ltf6iviXDy3a32NqFa7oSl8h18jXxm0OEBflr/3ekC3LZQe+viCkg4N
48kEqUg3v6vkwbzLNz5nQ8Mhqcx9tv5Jyit2t3g6BnkoT3OjR9QGtSmnZvSyf32R
01l1NiNJfitoOTARFhJeKvQJLbEzaQwAq0VyAvMx6uB/sGx6wOjFR6XBTaQqyNJ6
QY9arEwAWxdg1CvswJZokEZ5M41srGIJXbq2WzXbDifuzWLYBiHfmX7FpIarKQh4
tNCDJyP3RzJ/q18XB0kffUecdIkwMW4FHkjuTrV5Ma1IUX/8R7rrpcDVdsgJX0tb
bbMTAZl9JOxwYeG1G2IwcGub6FPijnQSrJMxmG4/Sg/J3f1YCQzCgRQcHz3XvNs9
tTp50ynoseHAZMlUH8937qZ5rMFeLMuCi0U5wmmQCwWvpjxYPqN4iSJA7EgbpsB8
AU2wHcGAQJMLUhlH/d6d4rwIwmfYZDUkZ7GCqtMSLkq9xgjrOLGoHslf+EErSYod
b7I2VZ8KKNDmh+kYm4af/dWH1p99cKXbBdAS3lqji2hMgpPb8MpEQOjn04PqmeoQ
qYNTHcFUAZlycugxws8OEXBtze6fnMg5IeNDnJyDDDembk6eIX9sztpI9SJvUpEp
P6scjw05cSF8nCSeOxRasuT9qbQXzsKG1ypXHmA6HEXJNpSiSsK8Dbb2LiGnungb
R1XYMGnlvUKdheq8urJrOYI/n77N9DmCryaY5Lau5uvIYIrIKj/lrWD9xd04g98c
D7vgUYNkm4ASj2ekCbnmB6bvyeeISWN3qfs2nlKx2nb+UyjRaGyErksZwcZ2MOG7
vE8nU89FVipKDR12v9FU95qqbRHdcTh4M9J+NKRcPAdYQy2HKTqQ+I8O7xhQGe/6
myxWCFvF4+7wyzA9dkJaYTWYTPWpeJpmWC67nAfPHzOm6ZOi+w7rV+BX5YkkmGfT
LZww2BQBSmCPHDUzimvZohMANPyNtesRadBIVuXfibJmVaIz7D5rspuQOhQbxZDF
JGPAMaD6CQRCRNLItIoIbKD5tbvKFoRNmxOx/UITidB7/K/+7VOqk3oJbwH7D99q
o2rOvHsUzKX7Zin/+I33fV3euHrEqwwCfEsmluaLCML+QdyTufC1tlx8R5OpMQsI
X8LKdEJtOdwof0dpvMuW5O12KKPRvyPeelJdpvcQGrMgtke7R/SqSBNJsto575g4
N2E7IdbdPcUVYevl6HcuChv+WUbGALD7H/U+i1lMfweUNAfvLvBZIulJ/qMkx8zw
yMCbXPdlJI7TcKcj6rqdKeDy8B3fmm3sROGrwqPuDDWuuhmiFDx+7XSJnRYzfhJN
tEEc2nzKeLEIKfZJ4wCP22fFak4xCVwZqdgUUQH7k/yBuD+0o4Cu3RxmNUwngi/W
1uSUJ3n4RWbEIt7qhEjVJwUkZ6FmyLgVYKyoOL/PVkK9rVbzz7/vzW9rltMqtUfw
B7TaUdVSysx1t60RfmV9E7P1sVcsJC4hwR5NTNkxn1iiQas9lWig5tutOKrYe56A
PsbXxI6blH7ypI2qTRs3jhVMuPzgI9VA6lr8Ew3DFklfYD1zqLRlIPS85MCgl7V3
NIWlPFU+oCWVgToNKp1hDTa19CbNm2DYJtWClxBJnaK1XcJOxqS09B+tvwuT+DWS
X3kYNASTdKOMgu1nOz09EOJdEvzj3dy9FXEYkT6K9S5DtVUK55XsV7GhNR8FaY4C
zlNXTx4mSXqRMtL7DyQZMlVTnHea+xFkjPmXRh22IANcvlT0cnp2elRd2kjzH69L
MwLebSCFhMO0NxmCFsssw4Gj3P+jVeRfN+JyeHzdpqpr+AcsEDu+y7bVyl76ilcy
VbY0XI901Rl0epwx6BVIZERJXipf8XLis0Te2OE2PsJfFGeP/kd5+iVu2K4jnuhS
fxaK+3OMqVCm9+WYkhehoWaip5Suy518KzZTSr2qk3yAZpBzo6Rzd9GBJj1jZKm0
GfNtZd5BhC+qi6OZFXg3fIyI38Ke1rlOmPtmc+7JS5JvTal3QUrChxjm1QiqUBDh
Rp13p/0WZzzANIF5STos1PbrdBKQ2k9QCRo5smrKwR/uD+jxSqZCAh/GAflzx3I6
bdN/jgSdCrakOIQlCmYUaDFLbjbl1Kot/NTNJx/AvJUc6PfsGnOLXc5sacp71U4/
TZgloGfEmGikVnX6XDoGqp96aD+Ytm72xQRodGkz7Gkwk+BhVD+zyTXaSXbselQE
LSUAqXgLLUiJaz1zBhZeT4m8qYXAwLrfIW6dQGScHBgkzEDO0ugSdvIGRcaLiDl6
AwJXzSWpNAwPLXbm1PQ8+fe1tOc9t2MraWO+h9EvCeXkrl1W9mdkNSNtGTnhGIDW
OMoe2JNKItf2/mEfzEQs5QVobrMAZLqjaomkzENDUiExhVxfwnUkv0YdhKsfmpTl
1mFfZ9BrO+9mMkO+ELcyiNQAl7DtXa//tktO9EAtJG0s/laJzXZ7e4fjXR7Lovrz
VwXE0yDBpo0IOhFZ3tn+pGZHG/wx/EfRA1p0xB4xql8j29sMwCYl0lvp1x03iczl
TMZ++wIS4sErZIC0lraLaRzeCu8Fi9C1J40CS1ZF1qqI2Yii5+TJyGBXCSUrU3SW
V+SBPkeIBDRBODS3m74NRdP9vwTeQw27wHlAHLH+SzmAUsoj1OiQsJvOQyGT/xXH
HUtAVjnmfTghQg+S6zBX/W+h9hIBcRkKpLTJSwLhG6lD9nTOQkyIrBdv2BcnHI+I
1tOYk9sPhNfZqUOdGEtYU8fp5Hleg0UGPTFZfNjpGgr4+H12wLj4J1n8pQxxHkES
bwnMlSP+7LR7aO+RsPS+BHB6GEy7ytn+AgkjtEpwL54gt8sfzZtfC2B+BJTUozSQ
q0KcnSLHrNJHRbkPyD0ToYFYtOhqzyRFBaYdqDdIC5dAvFJ0lw5FKxSGo/kKsCvN
ODpvp2KWitGO9bcB9BNwc/qmPri8jc8+YADEBVwQX98hBwJuB+TPIIGrPgdXd1at
x1cVCMIVcedFb2wkJbtslCRLKPm2HyJ4wxumO8efgL83DwaQ0zD6TeoCyjjcSRWr
w3lYw1f9e5PwDsmxgIg/KkcO9orm/at8o1B32OYHAbTnFux7E0Ke4/sM362l4K1C
srjqb0BQ4PYzVrYqbm/p0QSRKl8OndabeRp43zrhgTsHb7WI+LB+iAaJD+a6BBPA
CO24FVd4Gv1aYWlYJJxyaZGM8TA47wi/eV0vw7W16g7kpyjSoGsPdyhkZaNa2r40
rXvNgUOlWtf7K6Auve+kDPCwlV0po3I+dTPxRKJpGnlC2esRUFX+P3X5YiGnuEru
RPKKNYuBVpiUJz5zvK4NNHu8wTCUdTgY/ONz3dLRiWuFTmkwLXd61iGAVRivqp0s
nr9p1K7P1CxR/6mZhyoZ5C3jd+nDfwxkzcOk/dsdlyXpPnV2KjSQwnu0LSqjCQb+
HWpsPsyZcppXvkM3aMtzTUPazHclcvK1+IFaPHTFIixUVObds5wAfu1hLu6zZRKq
LBQtVmJ+Zz+QiDWSQepffZ7Z3jXF1mh8n24nmcI+VsCcqmICVyGVcjpPn2P46yCe
X3JXqReoeD7sGLlplRG06g6Jn183JKrxhFozAY/pjlKtwbnfzN2prs/b3y/C+Mt3
9IoxyiQLDBV47jzNUdgSonGKiU3ZCPuh9CsPEjaS+GQUVmu3xHtffv+I/rUJIVLR
BlXQIDGr6pI8S4VlCHBauoaqg1rxsmq0B91djEKSTbrbWk3jcGwAiQIoOVxHhyRg
H+JVQ6JEbv0gVbscTyG+wQ1/NJbjd30kBrJM5HwB6pL5DzhOtTClpfY1hKpF4X3n
I9wo64uIQn/yBvXdsV1p0p2teheNSXgmGzX49gTy1XruJiI5N5cwev/wdrr1WGmH
YM5TREHfUCrQRmjrHpG7xSdZ9IXF2K1wWINCu0dwobocB4Sv5l8Ttgq6KEgnvNoA
uPpEOzyfz9zkD8MvcQo8sR556pVimwnyjyAQI4EoMlt8GwQcdbkba7dWllnoHlJW
dzLChF33NVTkhMUxho+dAL8dJoFp7I9cQbjdqbLyxMB7xUdvh56QfkalzUhg0aP0
LoaqcaPUh00MFXqBiNL+4knnTaMIYyBVlFIwVZf3zje5LJyzVDuQ8ywsnWx7X6ma
u2+YB/82Dh43A5is0yK01tx4DUpPW9DiYpitlOPdFIIyDFe3Ab6LNAlfw6xHeUWz
cCw5b3wU9A0aosw9YYMtVrMtqnUFGIrsRlMAO2nm2ALYTueOBuvTcE1wGaO4Udc3
YTuD87sdAccB1A8o3nq7x321GZchkaXSTVH32R53op92thkJ5KAHcmkpc/byMSwa
oNubpEaym0YDtB7pwx3v3Udb2UWlPTq7FsAJocM6iexn+SMkh0FZENXOualrtSAb
+zmfB6eehei6mNfupC3rpDa0m4t4yQhWRiruuCziEx3hyqXHWyf+YzygTdD1lf+T
EZ+w0+/yEz9kj8srElL6FaunMCmOpJIyWJ8WlpdVwjpEB2tkLJMuk2dZF4Vd8PZT
V0OLe+GkqA6E4sduUgaFJKuXqYKvaxk1dDQHFTvJC/RUs+wtUo1MoivjU5Ymozo/
O+F89gbYdO9YWMKQ0TNBhBwU1eQpVEziX0rxyDTKd1X9kNT3pzbp2uBcT/vsKJD6
NnV/iuzGYbUczyeeufHdZ+6rD5knV1r4zIhCbMltkoK0TMRV6FXwam2ARFN5YXo3
s+ER+vXXJUXkRnz5hO8da+izXu/8+koK6qW7bRjpQ+Tr+9DcBKmzrrHccnv93t6A
cpwYZBa+piDCxzYpQ/s5tTlCpI0DiZqraDbHAQqpkodzoxogvauI1gXylmrCJfgb
wTff4Z/fOgueYmoLh5ir5DlcXli4oEiRYBbbmb6kSp9IegvzowvqmgoDuwoYngzr
i4sULIpq3XJqnLXyYBRIlqAdzbp7uPmTvwdC4j4OjJogxmgmEGSdLJXz5UakWAmz
V6UkblaIf8NAJSMGGgR3+teNcq5YDAtEcdPqKrxjBvtD16Jg0mTJJfF0YDm/fEms
7xKxdjrzoBWVGc4URIw7WDQci6FXRanKjTdVSpS65K9GpyEfV/BQXyIVLotiUV+E
/geBw1yzAdWSNLaEtH+Nj6KIHEguZk40G8FHb7FLMOvlG0YeNvnbbrXRpvZ+fp0N
GMgMP5LgjioHlb5R4WkYgcJSQ0x7Rx9pQq0dw2gVyQdxqUJsGAsA6bV2KUs1p4G8
qVqnYJN6xNTZcS9TpuokhaSVazTuJf1IjU6DMVmUb49aRGL1UMunow2YhMfaiPzE
hRbMoYiTLy4X7d+vVAqqDb5cWMaXVDp9+D35/dtuoRHDe3fsdAmaaY+fm3TIzRBE
krlHl+bKi16TmX8mSQR83VRm75yZF5ZU84WOYCuEA86xQGwaJBykArDdyfCJzwFh
csHpFhxEWLosG5P7l0VamuSuf/7nFtusrxzoBNmPoZDKQZ3Zjm8rBvW6Rf0bCQYO
yEfXSL8TH0uTUsM7mgkZeOzxKJihErnQFgnEZgsv44c0t9fdILcttmUqJumdFq5y
SriAhNM9yYD1DaFBR99GL+hM7hKFG1swshmVB/L6GXsYGsqcyq9Av16KWjOdl3zp
t7V9apkTR9ElsLLU18DdsF1kT/SAQWJuHvVA7XdES9w3OQKlaFMR6fNrWFBSyXfR
UBuE4l7V25TEUfBM/BqxSn+XKMXpcjp3PC7MiGvDFl1/FEMUE76FNtI5loamvJUE
6g0KNHWSHhJG1Jdp8AEeBv8ZU5Vc0qexi7Xu30ui7IoKhW16giZCoQB4Zcf9v8id
BjRhElCtyv64OD5+juKgzBcKAPJERHJrOhdNBEy77eCtmlpJYw0gJZERei9WNwe0
bKC9fLUcgXSnV51SMqihrPYSEieWJBjYGWuCh+IPmjoPHu9Ca51iRDPYR0TFvdy0
ABT2ss716GQUgEWnUa6WqkPRC41HP7iNZy/K86ZOztXcmQWQAlodg9AqshPrqoox
cyBBoiAFJYV4xBZOSVRsFZwUXiPl0cFzQON9+TDzk1CQ04hMSELV3mMyTr9oo5To
zmdwyPugusW+kKeqyRpZkAfUQDktfhm3YuOc6MyZTRp5KgbOcg+rfn1SBTIX8H8F
FcJXL6vexH9gi5nxF4toZ9DKhg2zyDupiqUTaOPM3YTDPx4XF6xVlM+ZQ8q/D2x5
s7jJLdaC54tvZ3jzV5np5GXsKpD5EMD65MgdPDfrmg+AsqVakgu7O9cl4xzyHYmc
eNc8YYhgdrtuIy+XVUCKO9ZrSbd+5f41tE1ZD5OJ8mK+yNJToEozabUNDJcKjjce
HHujRW3LyXHPXrv//DELgIU1dtXSNnHluLedhuoDhlvbnTd3BqxZ+e8XKYG8EIrF
yy9lf8UOfrm8MyOenxj1JFzRDmzXNPZYJtnfKqAINcnUdMBb0Dm7YbIqAqfnM+mj
KtpkFmu+UJr6eJejZiHZBxdcEWbpH57KlJzlJ777LcYKpkidkxUBcxBnWpKzLf4f
WwK1JB3qszzdz1pP76p8dOo0bpgWsxsHQkqQHWr8iBtVClMfxppAO1ewGUa99iXM
AaUY2R6Hpz4QuFuXwfAI2rKSSaHEfO2ii9XxdPIudyPapKWyYl/b/IT2OvfSVLz0
HebwCewaTZDFwgBiLtyeH7meuMTNBAhV8/HR5tCbJZqRosDIo7l889KNh99l8jRL
oW1p5s13h77R4nIXxjdzIQ4cYkLs1ld8JG4mZPsqzma2EF1LRnDcQthcu5Hr9R9F
5+25+SZxopw+yp10e9In8x0VFQWn+FLdKzvQi0iOFd2dM9l44bU08pTuozS8FvOy
WOvlXcfRLeB4/+NGoBgcHTSApAZTErOhuqUV+t3rPkBJjPbo2SuMHmntXYIjiIKR
SjjGKw3Hy95HaYIHIV5MAHNVBSdtfG2skBEcEBomXUzmy2hVXiQ5EtjLEimspnnu
IoFXHn89TGrxQT5qIE2e8ETX6gzMLcQmIGYAjG+KrlhaN86y6+RClNeu5tjyCUvE
75DMaSNNPo2I4NLgzcHVB8f3HGP22ifDl3bQhjFqV+EBx5gisJAGKxn0Yuy9o0oF
ppbJzwJhPHDP7h5t6lJqhr54I4hmRZ0GzVSYpd438YMteTFWLBTDOQqVGI1a5S7H
NzHDCeOT3zJiFoFDxNMo3NLJo3bb2iD436lvBu/3tMpJVdetUPb4dEwaQ3g6FRVd
7yfyuaLFUTKsqBpPpN15/8x8+SYW+1q0vH35LJzXkpyxv6hjseyPRgEINSMmnJa+
O/xnYJpHN9oUfcfcaH2EPgdM2DeYhDny8I/KGWawE92I7Cg0Q44loUCh9PrL3NMM
OJeBqOwGmIDGw0wTWsWjdwtmmncuEsnFcn9SvssJeDUHltjWIRrN3IHX2eWvM2ah
T7kPnR6JlRLUyzQEKmHR5CXrdnOPX79hij2f/ogu48gUinYZULI00Su0cOIUaInD
KkoJnoEbMq0ObHuRHo2n3e+WnmFGIF3sP7Rgb367Ofy8wHtDgQAFGv/03Tt60bvs
K11VDyNELuhf4BlToQp2iz+NcGf+dVp6gEL0HnU16+ev9ge6F3zX6N65V83b6elM
Y/OEzW7uqydNVbzHQPp3D+cWPwceYVcjRNA5sOBbK0HE7JXfRdDwPjXnbv7VJjeg
+5QrNQo9j3WELRc3cKLi/+9u9PfBys8La+rU3iFeqatpgGvrvKmYuFb+nlyTTmW8
kEd6MBPtqPWSQLHHuucoCgWVtyPKbqi6c4BzqCQi9Laaikc9sikIFIEnBu0Ao0qx
hL5R2VclHvwgEF8wc0C2y4EkE2OL/y05fTn31+THGPji3OXdI/KxFuqt77PUupWt
V0qxZ72Ja8aVKbxQWHGDn6ptW9XY67CNNfD2cf8ulrhOd++Li8JSDUInken52Z1r
yruHn9pjdNdUugONaUdMWHZeAAmuiqpZBJsSlb1H/nVNuGhLgAPea8hP8UEKrpvG
2FUDDzg1UOXAomcbI0dsJFeAcKAX+btCLBgTqZVKSmhfY3jXxot9X1z6IYeapCsJ
T5z9Qk1Vf2tz8Hew3GN+lkn8uckAZX8UIz7GkkxogOztXK1aht66RllsPZhj3EpG
ytibPhHDxPCmzpD28Tc0JvmlTccQNs1qhhldpHxKr//kylPkR/KSKQ0MvWWTeulw
SzHVv2U/pIgf0rUPhP9XZh3+CmADRS1fneYi4hCzV3b59wYhbbnIidq2AxTSdJw1
4YNoHv7AKgznTCyLyukvDKxXoUSrbAHyf1bim0qT+yFNeDap5Jl5pSEG5Bf9K3Oi
DLkrkgPtZ/La7942r8hxX73QVw9YxA3ifWkEBPPHZmbiur3aqcokjRsb23ALjTtL
CWqFlmURwfFEHfg66ae0Dn//prGbGoNscGYRdaRlfDmtc3x6LrwcDTgZ6NNn5IjR
9uHPiS3FMUUtRBg7F84Vx9AZVL22qUmebT/Bv/SQcERKM9ucHsUH9fEqMi0L2Qq3
wwT/YTM+H2MWJgpEgYy0wB/i99vBYjHf5ea/YEDvzWzMlyXAB/I8BHcl3zg2tXV4
eW2wa7x6uprkIuvotVdqzmUmUugFC569mvXSd5PyPDN/JfrH1uo34KA/6ab95JS7
gqBiA92cl3QBofpsmw5l6VeI6pyBX8yOrsW6L47tBTpFXU1GOCCm4EbPZYhEf0iW
ValQZA+eIJpJBggjov77PxD/F2h4GkLx02v0Hymyaq6pxmzS2YshfF+vhTaOEczY
+MWyQ2Opwd4NhIzObZsyZEY/PoNmdGgyGJdvtIoLAXYRtjUUJfSO4zVo+c9neupm
RBhBpR+MxtrID8Aa/sBwuxo9lr5gOLA3KZ3DEUid5yANaSA6/Emn3vVMx+tJO+Nx
vbjm04kOzSzsVpVxbOdl8CAWNb3vtVS0LiB4EsiAA2kgo/ZMhY2PcYjb6zhQD68p
3Ppb+2SUrataTJgxVWI4J5JCcDffvlPR5t4IhTcE3K0AEzHvUhSpibmIkgEcPnPh
AWU0/ptt6XWkpp7IZVzAYwUmTeoirBINs3SH8r8DdilLOtEAlfv4dXcBRsqfinKx
PLcRZd84eWiaZ+hmsbHvjBDxPQ+Zlh2lRaYgejiR0M5mGoRcmDxR0h19kpRfTteb
Ue09bzSSCBtEHZAVr7osHJR/BJyu5I+pK6FeXW09egtXT7ov1ETapXtXu+I83Voi
EcdaRy6VHhCeNPZLySxrFA5w9cKN0w1W6SbnYXVSLgV6evtMZCDmhRFc4DpbssEL
wZLowWVP/RwHNFSbrSK5sg0yuaQlq/Sc+SKYDOtMVEApkeZW5/ddom2VNiCPmHJl
kHzvhcVsJZt3BCK0ABJ0rpYf33QS7vuUX1WJtO2VGxXwKVgT8A1MR9gp02eJLUzW
cQAHgCqRBNJkH2W1ZeyEZPCDt1y2JXwd8PRZdjjm8SMyvwx3NKGZZChlNyemErA+
cs09w4bCgrKXv9cSE9bl+/QICKOJXtSyBPWrLOjqvSW8ZPmCTcq4iAWAMHyyN0Ln
YHXP0VLRuumwhBjGFuuDryTKUR/Yb18sDkjN3/DrdoH4aTs81DpLtABgIwYsl2Xq
xzctOcCac70sT7C0yq+xM/wQN7Wu4lqdpBva+XbRnIVWwRp08et3pTaEacf7cbQv
/7TOQ5vCdyXq4EH78m0F/I+iYm14J7LTwbMmK9ZdGW6d4Xmhvb2c2gDuWZlPIQC2
Jd8rtNzA0pmQXfnp7ytvQEuscI70dPu15RP9sc+2b0WJOW6nBbUBRDaIxQFsfC/C
qUzGKf6aghDCWbATlVjf9ZYQNm1oprR+S5DwMvTNrAVOfDY6uar4CWdQJJG6V7Fi
96nw2M+VsMHr2x1+bajSXPkGdCrfiWyO6L1zMb+oYyu3eoXhap8W0HJmHBgm/KN+
duwRznO42b5bQL/F8S+PQ6Xd7GICjfl92IIIYcwFiGhO28ghx2tkijGYTykvMyp5
AgY2DFm5gn1SGmpzoE6BelBLewG4l3ZH0gcXY3GrSirP2wfKWJX2zT/yAaMXyKJX
MARdcb8vdoG+DyopN1omiOmaFORfi1URlXAnfIU/8pW8lJFqSiR+Uo5UiYdCgfYs
G34o3oPNeRMJ9HkPOxctQfJNZF7dt9JHql9F9dx1gWjgqzMKnQ1AhuehQ9isIIzY
NaSqRyvawRTyYW5xdGzz/gZSzNOrcIOXSZpFUAJsvasi+AhkmK+f3NH2WSJuztAp
01xpPqQ5x4DCymFN8bRRa6wLR5D7SPMfIx1Q5E4vOtgs09IesxXj4vqh+tdPV+4A
sSVNy1ORj7wHuRpSCGI5e2omwks3rhAeBjB/G5eUP+9xNoVgADxQgCHGIQdb9h78
2dBx4897djjZsyx7IeDcYnsSA3mDohJHfhHpAr88a/8T002dsgv22H5Yc/iyPggY
RSHh8sgHrV2trHOHtN6OK9UzYv/o+NiSpsAXESrLoqygikBDEeYA+JgwcDmbnTIz
SO5RDLz1K4ESs8V6kokgtwrUo9PRcZpbvt6u8YrumTA4C3C2i1v+pnXWOxMnCr+6
jgXnQ3kIHAfEPEhkkkNG2BlSlzWbDnzzkw2B/kn5eM/CyQFKeaMOdvhfn4pYh09w
dRnPabAbhstHLYeJv77P9OHr+GNxYV/v7y0LurxdeKwKJxN0u5IcdNaHfOJ+pMPy
nLlxffnvh9SziCFAwnmUQUqUCgEpqhx6jofXOxWm2oGflGiEG0XKVQOWhnaHLfKi
xAgD9DRwEhDZT3ts6B4MDS8FIcPYt52tMk3N0UccTclovrIxNe5hJFhkSVx5q4mi
c1toJg6SXjtSU1xoxWMbvgZBpqzPZj3Z1SgE2mvtT8x9NE82ZzJe1DfblziIhZNp
0n/WgbpZKUL/U4hST7yrN3Iapcde6CTzTRfRdAfMPlDiqB01Uh3mvQyY9UDd892G
anAlViSh8yVo86ZmZNzzW5+giz5Cr0cO6YaYvLlGDxAGPC/RW4B+KcgaCwXwFUK/
ubHnL13GWNlSj99ww3wnqL2wsc2NK3ekEdEzuGcavZRaVHmCjcAezVHDMwq8vYal
bVQj46lhWt4vytC0lOWmL6b0MLKBmUuXz/VLxJrRU9mSIMFGXah5Dn0wUPD/OrkQ
giNotUawkvXfc/B3XGqjwdRxDmspueUWTdQyBXvX6vvMtwQncQh80w8SDD2osJVe
aIE3jSpUlAJxW8ud2bgPPYTAWXZdMBbpYXPv/BnkFcWFS41KGO74uAaq222WmRWt
yJffEg4kGQQ1JGQCo6e3+VdR/1JHT9RrQpP2wI7Kdd98eHnnsbrMYw9ZHCyKuL24
m9Zdo0YacQQRJq/k81aNfc7owaSGaUC7/t6EAO7KCpcR4DK8qp44Vu/5T6U+RcyC
fDkoKis2BfiURpr7Lvp0OKsbaN2QGKZYPPfO8jH8HCAKHI8kn4iMU3dNz1BlADCg
+brf1lsRAItvdGK8dbhRqADLGzFrVMjxspCfvNhAiDHWjkFaW2ISiLcWupffxBY5
+q7l6A2FeaPBgvz4G7QW1fagQpbYj72HhOhivRg3zowaZKCScgzb9tz75YCVuKJq
P6oDfJhHPSzmLBqE3ZjnMXOocVDR/mqcU5e/zq6zCALp6RSLTA678e3/53LJlW1B
i0WUk2zTEiJc/dKsBJUNPrcoOCy59ZyQ4TjIx6FjjO2tk1zHNYLK2OG12PMEh+63
zrf7WzGYn5EYvrs3SBl5vZQloJQLB+PHOabbR4VcmJbwEpVpfplU/+WeDabXRR2j
AKxiNBM7C4+eZgoCluvAjDEzZPqW04yF+RXCbg60Lw+h3RWHt5w7e0XN8y+9Ku4U
mcpA+iXVwnSin16TvyUJhXzF1LxQqtjmEBQSM+58DcgzGQYsI4d0WBfPaIp/A1gC
y2Z+OqZCfxNM7VGAv1uPKG2/AJyfWtaxECW6qU1ILbdlh7GHaSOSynAV2PCY596q
bU+e+RYQ/j1xwzyyScZHIuNqBBtYAhoejm3MDVyM2dOXfhGnSrdJaZjhkxIrWtfs
zK2k6uyhUkZPdms4Or/Wf4en7BbhSR3dYhFHWoxCWjBR6qP8yFte+1qhhTIx+i6I
m3LTKIxXCdtB/F6s+wwsQyKYFJH4cQJUcOMea6phLQUC/wC1Emk2EPxsKbuF2ywr
GOAaDUihZ1IxI9GVsHjOunYXy84oICywsbqx5obGXdIG7yA6sz7sjS0ZUFSa/kVk
4xR75d6Ne++9364HsA5nvg5C5QWBtrVnj12Yj8TVHMEfo0iZxOBgF3s1skQoBRM+
u8k8cY+bRLzA2UedZWfM43rFWW37eaCvA3p0yUZCbcklugngNl/4hoi2AOvesXVd
FCjpHlW4XxM/qz8a5/RThmhTC0TkqQnxaA1L2h1ISgPRUiuCVLEhtT9F78XKNZgB
xgIo/bS8g+fK0idBBt9zbMdcRmJKPw9NJ46XICo225TgEp08amkaSadaODnL9cGy
WZAV2YC8OvC/2onfwvP+hSCHHdvztT5aQWk2WtKz0tGvwA5cgZUq3BZ+yTRyvHxs
U0kQ7QR34D4lA6bVfdEa6KdWqFuGdNupxz2ejCgfYLkbB/yXir3p4HmF2iM+YGU6
zydR4MUk74cgGXCLonRCEMOSAvU3Pqys8ClmhQ05ttUpCSglr14vvuYVB5Flkv67
HOlFHkUpy/O06Lo135MBWDJtpC37qeQkLFbmDXHh9NLolWx639GU881tUrDKKiG+
gxSoglwvU/5nDFiODhjRG6QcyNFRiTb8H7ljmOQSbI+nkFyrj8uwGFaaH96U5qhF
Em4V10tuyUIjlKWeRABtM1kIaHtXSoS+E4eMBPrsanv1j+yjJQo6ffQ3rYyKnoaf
WGlh57kPcJksL7zSZzw7r3sw7EtrHJVQy3peA5avHh/quWUwwqBd2QFTleMGhNjn
fJrbzpx/Omp6UP7f8U7VVTJ0xXkgQTa83+eT+jnndYtMbPIJs3R0IrLHNTMsosvH
eJ8OHSd2rZa4p2EuLodRgLAmfTfbhOuI8DlszhtxCmgUyw/Az4TR60hXQ+QUjkHx
S3s4e0tO9GueM/ZUxv9J8gSS4++vErRXtgFOak0uwh3w/kc2PUGP2+K9UEuJcGLI
H2ZMQUCcnsTqimpdhE5/jS+TX0gGotKvtUXIpFedL5qGYSTgNZevMTDyNsWF7nUy
GUul5U57omZ9hkigmFE8Kc+Z94d4t+sZUZbpO76MzcL/c8sgGC+ojplTW5DkF/gy
ZxxH3OBQN906+c7rvmLvWnPWjUso2wV/5UNjXYdvM8LKVQEAdYwKQE29hHpJ6Tfq
Ep4zHK2LB0uH0dScA820pJYGlmfK9EovPwRm9/oKHzFdgGndSJDQtN0+mLcOg/Ft
KhWg4tNEcJY57079pBF3/RhiEYu5ZucLx2BgRutwNNznsrduf8HLGpZx1IFlpyHw
1CQYDUgXfSZ/jlUnHmaA/pxbZSdYkP0pf97LStHPp/3kjJRruJ1GQMq3sT9Jaq0V
aPCiXvVMuFUo5kxaXx/LXH44pytbdvveojg+LApYJmB9vJU5+dx7qqweIIoXlYDD
wRwB/GPXqE+JlTMwgUHGsPMeUVB1pFZYO3Qc9MAEtK9gjN0LB6YAdHLwohZKnXU5
ICU4PwMJU781wfubos6HeMqI5/LkcghJU6dia//XYBsdYkGoqAcAHwD1eP+RZqji
XiQQ54JJtdv4X+mMI+2u+9yEDhdERy7j7baNMXo6stw5K6xLy6HNbZYwweLotud5
x4dcaEZwsQwml/7n+/5WE3h5tog9JxAxz/jWr+fPxZySaTFJV3T2+w0Zo/703wct
htCabH9o/imXDyDkodYngZ3i1LFkzi6zzRTyZ1M7WkpfWID8qysSFFyuj2UYdgCB
ru9X4J68l+kRlxvk6RUBPNF022uhDP2jOxT8S+lkgROumZMfH6Tz7SPPRC5qqSnJ
9Z3Erpe+FzkeYurTUq3SIcYG3KvlwJbHJDFLs5E2uP8S00fn2gHDiSkEUvR3yDPI
xXIVTirlrRZEx/1lrZL8bUJv2zy4MQ1/JH4rFY/VOxxykH1d8C/N1SDU4X3BrINu
t+BvHliSfmpHOs3Iy6NgGqKlSZ2AMo+H48ugdU8RVtcddqJgl6bB3nSImzb6kTXd
ur8KHdcOcOl3AyH0agR8tsl1VmlH6/XfdWKA1KJDSgNLMTrqODXlJ/RIE6n0REmI
dd+oF6Y5gJ0E9vsxrKvbQ0HDIVgsl6shY+pxkLt7T24CZAQOadvIYATFoar91Ibh
QanPIrKy18uM+NvIzUnThppML3zibHivqmc6m/yMO2W6veFuiAoT70DRrrTjm/QT
D0ZRMx9UcUK7oDaObUsvtOcSu28BEA2RYxixvkOQZNsOIvTRVlxzdAp3nUT5e/tM
O+A0JZjScZk56q21JHtlZsVcDeBcU40sjvoT3jXr6d8SiEMbaNsfk7IIsMDRbK88
Qzgu28FS4KeSNz/e3x4YaUStN325dtFiT/Kc+4yOV1Ry9ko1fMwlZpPTQfdPc8qB
W+/kL3gcEGutF1gR2EuUubSskH+LdP4gkqfbrmDaLrz/y18Zq5M97hQld543LOXI
idB3BdyYTnXBE6YdBUX0PINx0eTpXjRcRsmSwAwwASh4a8W9K4JC3ep3vpn6XyFf
En5SHSyJfGzyPbD2IDrVmBzD13qriM4lV59bL0hnMhG+9eGSRaKuN27osAAMV2f7
4e8dfYNzqYO7fl2Bl+GbNYlqqByZGm7V/WTSqm6KMkqjeeCPXJ3KUuA/tLzsosn2
lnGLG3DYnB8gCZj18YDoy/l4Q2/NVaomeFdmIw+xnUJKh6X2966VxGwj96FNgvN5
urR7c/s0rMB8Pr0uiYPgeZQUG0cOHJ2+SAX9QiTb5J67s9MuhjTETHDFtbX8wnae
O/PkXg3qzeNuQ7SNa7jI7rluaZqNHL0QB5kiCZGk0mKlKSh6xvT5OlOh0qNAIFS3
qW3nzdWyBQzsGSeTt8E5SIa6S98YGQd0Fi7dNelgwDNFMc0iBAV2cAV28ia8uRlp
fOoTWyAkYKf0nPtQHBxeaN3d54zJcGCa+oIO1qwryUS/GYSAIi+fJg5DMAJ3c/Rb
IXkBgx49F/kQCuzNLuoTUNFaLiG8fVCkX155QqE6dpgi0YmdYTBOGUGD3SE3FC13
UX2dRdr7WNltFPaEPNaybIPONgnf9rwGAOAF16ku5CluMPcQIa25XBsvM+S8pIUO
T/ZoIoljRBcVzbaf7FH7jJNaXb1N2b4Vrzuon7DkYcE9kRxyXd4+Huig12+k5zEU
NoVTVkt9Wc/U6Rk2J/AJ1m+XE+Ab192XQW7Oi0L5DP9mINJdUntvBRTUf0vQFRD8
8p/obVEaW9IIGWTZKkBiSF5fTW/HMOUK84yFER79ND70Kxr6o+AUEe5xFXkwiuYI
rgXnP1swbDnQp3cLyziTaDx9Au9gxtUbbPAFmV64GGadoK5n+lMUPhSrg0u3rxSv
Ad+lckK/9E9BIKPQyLd24zlL+DUEiFtjzRaDv3VWIHsFIxGqMRD5f72LTG7SIu+U
fXfqdBmvWSVVKMOb2x60VSbNk2SlzAo/HsjYG0m79qpvPskgG6axZLnL2tQUKGdS
0f4CaNOQDLDZUUw1ALQA4K8n1TZ1Sye63sNH7y8YzGnb+nZ75xus3ZMz80TU2pea
nTL1tNzg5ZsedyJG0UwM6RPsSLJ+Are2loq/qSlMPYLIjqP2g+x3ONe3i5AzHT3R
anaov8DAGvTfA8jXbkhBJ+uI9bN49hqQchQKvTuPdXYzwxMe6ttaUZ0VJsSPFQ3J
D5DuSxcIYeKm+C0BJyymjugZEysDxsLrtVXz8zBjsWUC0Wk8G/fAXd+l+ljGJirG
A/oH+9vK6ehoEZLZnXbXFf2epkWPZVacY6x2yq3DBKoTxeu5+yn+gK68xe60ih0d
k3twjHrgIqW9XF3jdX2K/7eGCis4JAi4GVxOM2GfFjLR6EvWjf9L57Pamzdby7JK
NWw43RhzyhbbhRO4neSiM8KRsmZWzjs2FnJ6/s5TPjNUMdGZ9Jj65xIq497zIiKv
lLCNLcCP1oa626kJ3El65u+IYrM/m1FFsSt9SKIQGTamsD+i/gVKhFOfx5nQIsfe
aydA0nmmQayJN8Xja66lc+ew3LBTM3fLltSsIA2q6lwUTwz1g1g/fOV3AIw6O8DW
GqSZ1W+meHqDQSY+Pg4N1EmPFkhdqEwSxMKWyHSkoacmS7o+j5iRLX2nVB/6WEcH
7GaCm0uPv2x+kwEfTx67XoLJwUJzzzI89MCGy7+lycWF7SvMbbBEXD+jRq1ETsn2
V/amNanfhC065RnK+dJZesrQFq8MKymTh8ANPt9ZpM4FCoTLT1hbjUY7htIKU0KO
jh8YtQDW4L7EBfLQNjLNXLw8hilrNFlGkYi8b2+QWIu5gqf30NLLX3Cxr7gDnQjf
vn6ocwXaUZal23/UrpIBZEuKXRGUrZulMDFvUpqszvTbX7z14aQcDV0ys12LnTfQ
ZEcfU0hVJy4bm1Y/mVL41bblxOrcOPnwkUDiReFVaxUIRcMRzeIPOrTYE9W6r3RZ
5bDGCuyv7DX+6gRpiPFssn5rgfvb3nMN7dthPkIo8QvWUGg9y+k7mwoznF40ZU6l
M0qbPQ1zY7KrPZOExH/k+XPZTlOAaraSv3OF8nQter6IgzBsNtBGy7hCej8W7mKr
kb7xV+ZK4OJUd2kqOPUeRm1McdS54qP4EN0kQSsEofTvgwT2wPZYr88yfS+9Urrp
gVLgr4z0xU60xpjaoBd9+7ofJt9/iozceGgEpK3eEfaiSNtRjjnmbjyRPIyndkuI
+1YJoMiA2f3t8fjJQa1Iv/yT/R3doCP+2o3g+a4+MQgMsgn6NmUkbFr9MpH3X4Vr
w/YguEdDFnFYnpo2JCCmAwpYqfSi3hKG1MCwvdEja8i4YXeqhTlJ3ziuLAFsEA3F
JQipNI8MuaX0FwCof1dqL+HET3mC2TskxGMZSYH7+jJF3UBpPS7qgwh1vOJNaTKe
pnhUxULdhoO7AphqifpmgNzdrreQsO7CVpod01RMfdgOli3/RCa7rzy8Gb2gzMzr
DUfwuT5YFboDLrWv8cqVpV4jMRa9vSu/DDl5A9eVPCRSO3ynK0Ukwg/WZuIgqxPi
oxePnZC9zb3Rbm+z6W/5p/8ttcnTY2x0LX5wB8Dz5Xuf1+U20NlUMpjGwzKUBsf+
cWUzj7AI4q3ydRttQkU8vppdsDa3uEWSaKETUJw+h2X5ley2v9ascAy5kebAT5tU
ci85kcZskkoGr/R3ZpU5g9IlPoBJa1xpV25xFmFge6G8de/8e1CsCR+YFeFHYwGn
DWFV+nBHFDKKY+cKfKhVqq3Cewg/QLUiMKuSWkwiosQnKh0PoHtVZviqIsneGfn0
6NX9bWKhxlWMoKaXizniUj/RvCpPWqhBcoxqj9cp4azRzT6VHT7zNO9lOJEAMKZn
POeNTMk8jWOOWjysCZX/0j5DtBBZh2OuZg9WJUAM6bWk7Q/FmpK58n0b169CTfgX
q4lll6RwHh3DAxC7N3VunG3MF/iB0iScPy9GRCiVhqeKYjFRFvbwkVB/+/lyoZIj
vXvOFOJteOx628mpqTjM95Ia/Vro9spRQaEAPokYzbACIyfBTSJNIRCZ0zT5Oqhd
fZljLkGRiDaH5q5Q9R2fmDlnUHGhx3lYIVxPba+QOFr7QlECXl/GQwD0uPKd69i7
jWChEgHx3PkVgaX12oXLel50Bm/WwYXu5XQ2YYT7VWZBgVOZlXiVgEhtx4GoknsG
qgoKmvGseK7v08j4bIrrlimWSenrCyDS2e7AoqWLP9tiNhBrcp+f5HIho9UjkfwV
L2TlrOsz3eUogdvMpdWRu/vh2SV1O8+mfFs6sVVfOLHDM81fkf7wSFyZUMCHMh4O
WZZf8FE1+O2FgsTgza26/HRLtj/1YNbLCcogJircW/m2+aqAK+igOxEBoLj0iWez
4xYQUh5ATqMaCFXkPGA54SeCNZsuKbAVKpi7IED3u3oRk97kVf+5+OudnTDFrQdZ
ep2bqbVLpdCfiZRS5IAKXjvzKQ0eqQ2F1CoqHn/80w+pIbtbHl4iLjsnL3yR4YA4
/zlmiFmSwOI/kwngUVDENSiujmMWpFtLM2KIuLQqyjjZYPAWqot+Ok8B3u4kAhiy
hoyWlZlFIkbbUX2AkNDnG24FyIhpLSXA3Ye77ZLH6bUlm15JuRvHlP4rG+odDXBM
+EoUqjzLNyVLjDvhh8zeHY+10KDP2IzB3EcmSroOqilsAGch/UMkxAIH2h38MjPu
Q1PPXrexSYHo8dbX186EW08JXJYUqgJsPE+pHmujrUoPmOhofXMzb6vfGjLntaH4
Q0uKz3OAmUq/JbjG0b29AdbaGXBVcfD0KFXt+WZ0DO5NDfWqd+b9h2xwpqcazQTF
zS8YWePLnHYdFS/ufFCTjT5iiNfWFFrCnu6J06S3VQF4QQcUb3hBlKR+lO4EioLt
WS76jCBmjPcmZan2eF+oOx3fwoojTY/cVkK+o/EJaYmMtkysINuxBz1X6Vmo9axm
PSxSOaDaxMuuhZEjDxJvVJUJMwJlKPBL0HRY3p2hae7PwEeQv1IAXlcPU2qsPf7P
Ujs0INXcP0VxWN9WAGjmFhf8eIiNy8ZBPYHJWQl6lHSjVOpLZE0pieaFRVGO9myt
OKgUxKOOG5AXoYaJFy4PMTYWXPhPYfmUIHeuf8l71RPP+Wc24F+jyIFoR2JDgXXc
cKkzdSlsUJwIRAhm9o9pEOdN00YUKsjHLVFI8RYe5iy8AAQqOPnBFKJVzUgBkqrO
eoVFqo2j/zXFoiIXJybIUN/n66d6xxA0SayIJMF6ZI/NQJrB2O8S1VybMB9jj6nr
FqwiffkRinBgm++iEBIlIqS/i4y1trmO/z4uYZYqeKFNqSFWj0qkmF7Khw7uZZ/y
OGxAToWghCVPscQiaJoUu6SZuLoBCEmFOAoiA2LiIexgGA5TbuzLIrsjZtCpihJ0
09It5FmrEvfHoJDP9e6jrtlteYEXgU6DKP7msWoXQsflQnS9p72yMnPjnAdBhhRu
xeufLt23Yt1Nn4YRyb5Uh4RBPKQADDGJ4F+D+pGLfx+/iTR6I7oaB+Ah5X8zuAeZ
+dDtxiPDDMsmqsNhVPQMIuxX6u/KDvfyWM1TpBA0BlMsJ1x1OzRQEI8X5k5sm39D
k0cmBZfMMonyEMeDa+pCp4qF4walCebUbjTx1s6z7aJ1AvJdp/rkbkHvP/lcI5vf
J8fUmRB9F41d3QIhDHWW5RAgYS8ECko7AMSpQn5+V8ImUHC4KiYS459cVfAb0X1B
Zv37JWkEIzCjjSiv49HxEFoq7wcqR8bW1gkz0UHgTc/owevJi+404E+HRvEg4QL0
a4TOWV6DTqEYcZ4iRISJGz3k14Mz56U7JFPPu0a/xpdklc6XKldOgRhIzjBi/9Uh
X0tffMzJPkQt6UlD1TciPuOlLlmtcxv+a3AhOY8/0ElaZ9JrvM/F4nE+0RfmaZol
fhTDPuS+c8tR2yViYfUB1qF0oJiNwuDsSWG6Tszq5w1DCv3CMfeH10uXrqniuBWq
wBpNhgyklE9/w4lGJnEx5DwBHneyYt4zjk03nB5RrHYZ0i6l2JrVVHLHa9EMN4po
kqfo7HaCflLZlXl9dheDaDk41MncD7gUHk1F4zx3wCWvMp9dj3mmv+RWq6xrZsNC
DAhydSFHkrmGlOlYUjVA+SmOG1IsATOUU/A1JE6C/dwd6qrb17z6nh+8dZmYsIXl
0MnnM4OfgSAciG1W3l1dqotLLRGajWnoXyKuSvFA/i1p96JKw/31Nw5F9kovs6D5
6bk3YnKQhRioEqIhHxovpvJFhuPEAgpTTY5zRIXtxQUlRdoXE90DfjWaHjvLXkCx
KFlq9AHToCJqPV2KBST6mjufolTMWm7ZuEzGZA1qLTZ21npBgme45TBed1RKIJnC
mlaVMq/pWxXOtGxDYsHx2vPDPTYsqFF+G3KQUWn43O+CWhhGSeFFFj6qiZU9vL0S
OgyltKqrktIxP0xFQErLOyAew4GxhwXnCF2iqogH7cCo0fQs6Zi6gDiaOpmLc9be
mdvHBlD2kgMigpCQsjRlt2sDAuXf7Rr2AgZLKWbewmRNdUKSa3MO5uKk19++m65K
rU5irR5CwQHym8PdtP2giVTht7YLXEK9FCLLfS+MIyTwrZ6vjsA1wfTGKBqKnjmD
e6PL+bIxeyGDWiD1MMT04RbtZCBsyUgoFXgMf4DNm5rvXEKQeMInqwDrVjwX01vK
B7d3ai6RFbeIuJxmBoctyxnm5fGQZi0QvwlgzuZW02gCmQClXBxMOfhu9M2T2h+h
oEDulnj/8zV3H5o8TMkKk+oSLwX5wfDJUnV7FQJZniEes9Gk1rDvXp5MLwGgAu+E
XWKzd6MlZFa0wCJRwbB6PFKJ9CkkcmrRl4M2jh4bYvy2yUSFJ2hJS2nRtEf6P7Tr
AgRqb9EYpJ9UNAPirWjmpZhfow50ovUC0OzR4g9XJyQOr6S0Ii1aVLTASQmfYKED
grRpW9duCEls/tKU2UnSUN9BaAL6WRsTi551Ox8HXiyrtwxnngxEh4vD7KajVDHF
cfd9r7BTG+1r48VhWKzY7vQAwYfv98AQbbVpHH82tOzLqe5yhfGP+NshGNKXp9zK
iWhBGkQCyruvkC+Bq4M83/0TgMwb8x0ZDhR/CrfyqLuy0oVZflYR2YnD45o7nQfh
b0hPo015UYmmwkG6HsKqNnvJEK4Py3stnMYtUx2HGLz2SSG2S5YFx6X22+xnaZLB
qBwNjZJQnfoBZNrXTRRwyexui53YD33ZoqTSbf3nCK+KypHC4Ej4xHQW31NLN9Pa
/g4VDFWhXghYyTv4p34+/oM9eqS4bcjvDc0vFFnZ2GVwqyBMF0a1gOhPtB0WMlYy
9y9m2iBgjvpYMyA1EA+othzPykwcj7fZ4vFjHXb/3Bi+AMAbYKMVJwBVzzaWVbYl
Dwg+OHwLzOXAQmHByFDCcFaqRXeFoRcbxrriZcAXhe0A0ACfVEnEV6a4BAUCLR2w
jdIJNAVdDvXp7SpE0x2QPF5IXknxGXZT4mbyA7aXwDC9zdafRYqAFWHX/D4nWmi6
6x8yByXdPojx+9bitgHGcswVXWOslpfBzlohnXEbOXlbqd4H5b9zD9G0tlMYXs5I
wQW2rraIEm+W5meLVK2FcRCYBF23clfwychVhwAQ2QRN8IcP3gP6niGiGNXWGNv+
liPTr3FpXqIiUWUkdeqKdPqtbHJnnF/3AuJOjM1TBWFIcQgl7ji1IbBV6mYmm5jC
N3aQSYWmXfUKNrCWnA10gDOaQcQDLF8BX1nx0JVAmSDG4qpf3aWeEjjo/UxuT9Ll
yyc4tKz6KiAoDnuhK/0V4IW1PY+jhAYsRiOQelRGBEc+mZeMBCA7fe1ccDaulZ8g
Ov9BJGYCyCakinXQf/Ydhpp7N7HUXKdl7J0goXIUOTalkdbe3blpuKfXCZz+UEj0
JYtpK4Dqm/0ZUQk7nfrnK45pngug6MsQXBulu59S2gEPxziNy868LWvjPFAvABCA
4Npsq8GpUM290mVC2SVxcoPodGuxOc4RviHx3eTdBAaiiuH+BKvBWd5dt7gHbOXG
TRPZ9XDRJC+Tw6l4rXzkWFS3izO84AAqtnYnuevHHD2h2EQnc5kp1aYZSqu5LZ4m
19lNcxu6ConPNbyW4TTddH56ixzO0XD1TqvClfQgTqc+HVN8fk1ktRmRwyWT3/9t
s3rZ+HvtyWJtNoDpoeAZ9YnGqms+Sm2eCMclU/6NUuiqlRTc25vNXwBpzhG0kHxw
CYarWzn6M3oGWCMq3XUOlxDetmx41jsEVV6BpMRITNx6aK9VAocWgedgI7o6iz33
3HjaEo1rnHdkTR+ZMyqGbDZhLspR0y2WtiXpGbSUpH9VbY1nbFZLRV9ghDZZeRT6
1IRQhA2uTNuxMvFlL9BiBtAVBBiO9sOch8ybKsbYI6fOqV+l9vvEzPvnE1VxROP8
0/FYnQqwdCkpHzVTP4X3D07o6Ysfpc2YLWabOFOyKvbk8+pDDS1oMhw1bVvNptA7
6qdTJUBIc6zWAVEjSXuYg/ZjZdoOi4ucayC0KKwDTYdMHxNBfDpB2cWXi1jMsN+e
vwIquLK6jF5lOAKjOlrtoes6fszQxfw7T/G6fb/U280ZWsqS+vmDUlobnFqJuvxr
ewD6zpbIhPciWo6FIFzEmFspVHyQXNLiCuBb9Kn/6DjrhThDMhspXjHbjBbbJop7
U8t2+4sGbAU37tT9T9r1tFQ3UDtPDVtKvp5NjAn/ZUzQBG05ga70pZ6x0patS9ky
DW6FbwmplGQVvL0VtHj7mCIEMek5L+aLy7IOig1ncVMSgK9LQLgeE5tCh/c8YiHh
eu4OD08ducKQ3lJiSZ6YVwa3ix72Q6SK2IZgMJ2usE5gn6d3BdizGcBP5FnHpCL+
57Wo+6Unn23ZSAG6o6hw8bYWjmnyxaXNDQaNyzwj3e+2aFzAxsKobLMnRwfry3GL
gdA2YZf1t04FoWLvluloESSunTepoSmloMoEJJTlo+8MrQ3spU3WDwkSKK19noMN
qjmLb5LB+NF99iJGpwxMtWVrUXz6lOn+j/8iVoVQ1cWU+5veXc9Ffjz4qZKSm3Hl
UKHmGWbJKa3050hQG/NrXbHJdC6puVK+2dbe5xLBSRC43y19FK+U/i+EaQsO6gki
EdAvPFTll8ei8touECOq4JnyqxGKyCBqivvTmNpGZmR1/+mUEj80un4PssxgCMPC
A4b5jj4OaqCEtiRxWz1jjI5eApqEDg0OLMl/jyDm2kYL+l/OvDWEB/EMjvHAQfPQ
fcbezNvNQmg+pRiT0Yf342FtbKl85gLvFH69550j3slNVmZ2f6zv3GweKN0vhA3a
WqJMb0FwTCf0XBRa9iOv6RjAb2NtS7o7AXu7Ue4PIs6vSBXYEPThcwvvUEWH82gM
dM2hXBGNYpskMAtVv41KT/M5iITiqMg8PYxh7d9UYnOBDTdpH5ll/JfYrxRNM3E7
jW111n+8Z+3E8gO4C5fdrx+jcBOS3nCJnZcay3Hmo2BT5vd/EDvS8C6lbbRbLWAW
1iNZN6H0GNVCSOlUN0KeQCq0MwmzMP7K/4lLrUyuy5i0wlNL0cb28YB03d6c1kkN
raKWo+1PlryviL+Zed8aUoljsK0StYHna0Ngwh+sp0GV8WW4cP/U/xnNnO19xtdQ
/EWHQxV/2hyPclxzgLnUHdLoWUE4wtlmIZTDxGejH9/tFcjST9v3YQJmYIz99Mcq
nTlFNDWFekNx9LGTVX6MrfBvgmBNultPS10f2qWOoznsJJuN0AU8NzfV98l66+eC
S2plqeVDERKYw6NULgZR0Kclf8gAsmBID0xdrLRguWphgE3CfyQnk+ePsNIxGkru
xfjvWq6WkNWuk+N9m9lnpyaBnLbFt2O4LkFK+iH9AlcvZMbiCYsJKc15q9+v8mV1
SkQVUrcCArC5oz0ZtS3E59p/MfkC3vmsjgmUC3WRWHyUrab0kTIK+5r3Rzpt1Dps
L84vpexDGYZPPzAm2/LBYQVec7rxlT82vlvU422AdHpxQTmmnBRWG7YUImUXeVcO
7GetqetkpNmsaDyT0EtTL+UNpxaTY/GI4S0c7NYbT94sLQZYp1deQEXAsmrzcFD7
g3kyViq3yr9fJfI/YtLYCyeEaer7VzRD2K57Cytd4nVgoiZ/01Y3ID25HaFIqGHK
AApnZZdNJSkwkCPKI3bU93bnoArxONrnqc9hxzAv7XE8KLiS48q7SRX1LbMe7IhO
nK1nPH1al0v2qxqCha4OUs2npRotoNkVQ7abqX0OB4mBvQfusPLfRH/bO5HbKVPr
qpZoj07Am5SnUJ4zVWMwXxGtskmApqtBwNvZAFIYFXRyr5p1L1AfgrIAvGxO0QsA
czTAJqb7DDSmzWulnAsylumymY5tTGHtYriKXoGCFVlESDVAKj7Z9MHfsmYskVhL
xziFsanH3JGOZOahJ8Wx4XsVv4DopoRg4+yxLLYk7qmMpNEGEJKAbl3X546Yh3ig
DKxfIZVTXQKZv3CCfhPqBcqyd8SL+E3ekkDxqUFS65J5LHy07P9/0QgATR5ceDf+
UiAJYEkSU2qQZP0CkpLg7N8q6PaOri5Ro3ORg/cxwXFkV2netfVLgdL6R40Om/zP
bBtPK7GNP7Pm7cnqpuaj6J+iQxo2Av7ZA37cTRyP/qrbR069kfcUOICWaj1eP5n/
KZgDkPHO2iuLt/calKgGdVOZ/SxN1lbHCWZZ7N/DgXVPcaiz8Lw2ekYgNDDGEYaI
eW6c4GgWD6gVMcWxenxk40cYgPzKrRhcDjuJB83pHsFK9SefoKKDJ3Y3rkrwRDu2
8UY36T9aoso5yOaCMPpL8ORKfqGDz+LkI+LVxyXA0EdI1DNXCnoh9iA8z4NDqUFg
5szNsazvqZn2mpNc7Kpz3fUz4uuyBmm3KC41ZVL447imQisHeNKytf2Z78+tPN1H
iJmWSRp6z37Oc/TWtl4HsCJDDZ4cBi6AK0t+AeIyHZo44jXQzlOYf/p8pHYaMd8P
XoIbFLk4nbxuHKoLqsjqTmblmmarHd08XH+tfvaHyUzV32iAhVPB0ZMsywN43vXL
V8QTngUUlQBdDq9MDEYRud8K10DdcziTn2aIYT7zldlKtgexCEbmkFV6e1OLizX3
/IbtbcMNsxOMDw9URwIolf2zeO0WaQ6EyKn7Cw8246bxmBJoUenqiK/7CM9d8GN0
gXaDLuHgBQBe4sRDCBE7snsLaTSTmwfdCjGa3WqVi0KZ32UcjFjirL+baTBkZ08E
DQIWEka6n3NihUuH1CGkllFQNc4m7rJ2q59NWrlPv/v/g3g72PbqjBhM7NNBU9gx
NLBnXWtVCWrFT3NJKKanHedi5BFhxgM2T6c5mMtdGqj10Js2IseOf2Dxw7LpPCjq
H3oAfNf4u4mALu0+z8QAd9DfJvnGRflQXz3hX7KfENGToHpBqlshtYcC0P3AHr2E
lLv1D8YKmbzILsouIQYCG+0dTSgS4qxWNjzPvVGXqTsMBeTzFFo+fyl2jifGQcrH
3+N9ZzNx4ArcJzVSqtLNpdUjbFZnh02pIVrWCVpXYY/xvkjhTOzD17y6ymyeQgJr
+a8KQ4ZSazBoektkjDqKnXPXNM3hyHlqyAiA3UwasdMOdoCdsy3QXuXP18PoAspb
t1upIMOTNli9NnBKjUP94xC4+FHQCUFuSoop71Pn+IoZ6uBzVKVyc2Oo0y/raxqP
VDlnxlbg0YvowL2GyVddYnMZ0qKECj/xocXf08RWjTb4NzRUz7cPpKL10MAdCoGW
oSSpiLbKZRe93KTx5ofrv3qdGf5Ijoqfe7YF4aHwgcACVtExT+AjYFOvzTs2Y3V9
x9mGTB6LIQgG6YufqeR5pf18aKkHyKxjAfkyHD27eZ6z/qhme6Yp945S2WgwLCIn
Xqjeesk3bb3fWNXwvozjh6krrm5684df4Edv3GlSFrVTwaSrAYTbQbOj2JNFFqZI
YFrdEaR1k7UqvKw5mhcG92iHs62Qy/3KY8Kt+uOCd2JXK4XP/wHu3LYHLh5At8WD
Wte30LaFvCdqG+WDOgV+MmEOi/edUE3IgGqa60wtzMCfjy88fyBN3vY/VtbCQSRD
3N100BxpeM1dr6tRmjjsLYEfVy455qh+4IS4pAH6RzG09UP/+JvE3f5VRjazAmOQ
vag7+cnHw8sfw4ECChdfeOCMUSVV5c+y/5LjqnV09WcWkwH1AXRW6cZfvfeWrzbk
a2/KhHF3eKymYHP3OmbjTokFPaNuHWLQYde1ht1T3mOb85vuu0Zv/NDWZjIgDGbo
yPAEmUM9WrkzFNB68VO83QFeiHWuyk/0ptH0aZSuC6wqDplzWbUSih17Ypqh32un
2gw2LjqQCN4AeHy2SvHmfsp2ogpw59pSYS3oMMozSr7w1unuSHtGrJSEvioR6cht
/OSvvU0Ene+C7ZZYEEXGFkr6BaAk9yB+0rlRvJ0y5tISHQ4DjKm2AcV7F6vmrnr7
0YfKQpZ3JJl8T8uKO9zuStEDuByzCNZBJjKWWt8DP7KyBbfvS0fmIwX9YuuyB46X
nyRJ0n+AzSUSzptJB6OKvKA3C1hlTaeBQg+mOqXvEAb6mSgjYqDB2P7yEESqEuWN
kAjJ9+Ls0lb5S2U+hgYgDXVbS/9iHJ7VLkW3aw4BL7QH8wIyQ46aRl4LHZzLB/N2
PzVaZZU1GxyZJ8UaDPOcg2S7B8odaKUuYH69PCUBPqUZ/voXl6XAzCrp4NJozKRh
W6UA0lqjPikL3vOhjsypzYEg8vgPcNt7mv+dofktREVW/0EZordlTYCYYCpSJODP
PxVmAckGkEW5jU2ORiu+F87uSXZst/mi6wp/1j61dkZbOs/aqGD2cngwk/s2yfLv
PglZCIoZqqHKnbT0/nw1lNvNaPidsdBt3z2YctHSsZFhuxXWhwlk7JFoI53dL9KT
Zx//fqLTPDOL7iuPq6YG8ivcr4/k8PgnlvUWAJpPL0uAvMprJWLsxyrijUASA4kh
VeFr2wsTxH5c0D+fgEqRk6rh+h44KjntE6XnOld3z21LZni5mA+7Cg6CHVi7WSNR
F5j5XXCuSGEd4EvNndMNfLFv/kjgepqRCYyCSYNkXvWvVJD3FtJ5UDUi1UHAkIwv
ced7la65I8YvKlYT+uQzWlEQTVKvyUnTNFsEniOrgloG7G8J12adMsarPzhPymZy
1lDU1pqPzv8xEIZTJN0fFPik79OSYD/+APQi3clwXDsxjoXYqIstD/AzTy0MoeUT
4gCWttvIWD65+fLHdhVEu+M9W5xvoMxlsqrRscI8jnH3V41ThtbXRfE11QNViBgU
5Q8QQBOa8YxrsrcIrQc+I2oKYKLKCIcMp/0AV9bMCAtcChSJVett0hPA8eZIDVOl
CxlTOqdDt/AxUXlujoyf5ad5B+kwMwKHfzxYnazdQujtJL11eeqjYvQ9Vnd7cqHf
Dc6CFN+mP9Qj2Qik8Xnxy4jTtlmFg6mtgWY4wwOMYJWTHQw8W6BCS4VXqEiuFkAb
OEFdA62zwav5qj+2lKXCYQYufKAHViM9sobPCahjBxTyHlwSg48JWqmX60JmPDuP
GRQ55nQNxO7zuVhCTPvigOv8l8P+OOiztgUDzhBurgN2G62RIYBSZSG/Hp5kzUox
Fj4uIlk0wk66M6Ooh9tdApOZhNOz0M0dUzRunwVannqmuCrEtQOAOppKbtaePqme
BFApjwdx9iS/UHbVVEZ5bt2rzsHXK/mt/XidxDJa0cAIn2mSlhTJabD3WWLiHRQp
TmO3S9/XGnhMgNlBR/WyfwW93vfNSZv28akBljqzuMosLpAe82+1ugzqUO69a3aA
sWl/XyNqPvTZlCa52uMOoEZy45rxasJpPaPRP231QS/4TpuGnJBSwqrs7UPesTM4
gUxvKp0c+SCDb12/+VyFXfV56pI/A7mO+LMGFyM/wUvixhjgUuo6TxckkxPT5xf8
f4x/PrbdH5rUAPORSE/q1NTdhwhv06AL6HUjN2wfo7DNTbv9JkaOuc8VgFzdwEy9
TbzsRYdnQMim94mpF7/80HbLtlGT9omEQxoSBdDFKzEtUxkUnqy9+4I1gZSW302p
qqlq+SnKroG8+gGEhEsPdlkd5I0EAgS5ROCVCkPvh9CcqgNQY+zn2zmgbVlL5pAI
kGwQzHzyohyRHvCvmYdu4T/0fIxCe8RZQsfm5kPERqYt8GB6DAEUIU8SHCG4hUlQ
4UNns/ellerjlYLbcKW4tgpbT6tyziYOwXwcD8DPY8FnD1GQU/C9Mr6P9QBA4fKZ
wM4+Z1+LiqJJhK1S6biXJi+jxrhiviXPG+d0g85iD3PeaMKs9XhD+D9SXTVnDPxn
C26ChZp9i6cSren0lImH20a1WJkOxMprQc6nwJfUrLqO7JMNVuTg6+BJS5Qct4Gv
vz6dEu8N2BXUGQIGZKAJJRCEZWCYYPUwfnFSRAOSBcGvYOjilGbLzMs063+EngBY
cCO9PYYuMPhywKSO8Ks7hwJvtU1DXwB4700Z5LrWKU12IqHZhxy9rUbPpqtxdcsn
evx1bI4vgoaJEqGATtWzXNywHihvwT3dxxPhasI9VRJYKXupxFKWKku+T7FrDOyD
exst0CpYqvVJ3ynjUoNfh1KgSMbGdsZVFvHDKzFJ2jeOif4BOyOEMuf2E3PmlkEi
NY04PYPUarmH5lCj7Cv53C0locTkqaYjQSqNheqx91ERUplpaDEqQCWoSQjZclIS
tJ5sdvfhSVfxWPevDiPB4YO8zU9/apfnDFrbYem53pcM/VXFVkEkub1InZZdBMWr
cdoFWF1KdOJQenY7W0Sl19F3Uzc/mBBtJBqPhrf/RcKcTTgWgeojQu4OV0nolCr4
y0QiNrY2w6XvkL2JzpKq9ByTdgmOWkRM/77kCUbktiAQyMLtqUtmNR3S8exiyy+x
BCKmRIin0p9vWJozD+D3qw70y7BDVlO8C1ngZj+s84tlZitjDQgjQsH2HDQEJxBp
TaMkijBrJI9BWBUCZKRlINLgu/UqLAHi2z2xpb7by+nfnccxSWYMgK19hfAPbm+W
3b9m8YlQf0gvw7EPlebYgc+CKvtmsHJRCm0LIzO+WDn0YiPdOGuG7aCn9Q4EfbmZ
C3ogH7uhhI/0vde4CFwOdFwjEw2D8TQBbU7DJCRk5PQzAVKbeABIbCdJdZwelTVR
8oMJErBjdzbOhqfRLCmFg8jxz3SZ34iYW41RBp+LXFmW8emkeXD/PZsbWOhFIxhM
o4CGZDLwCBdoyvHaeD+vsJk+bLojlDecTTtPDXHPzQrru48lJLW70emihbStrsP+
tGFk5177vTKRLaBpr73RL34aS0Y+jMgSRNx6yixhCD4AN6zOLWmwsCsmJRr+XRAb
kMGpDYKrT72M7kzrbRLS5UxKBiiV184+8Zh1+Tpk8cywg2qpEeQ/FKnq9yhEFFez
RzLg7BUhuErktqHWteUDNDvuza6t+JI5bWT1mNttUNhTdi/VcaKFm+Dc1oM3z3IX
8B9ciyRwVEhYndtbToui5bQbz/4oN8HsGxXc/xBOc5usxl6oN2wdbBgCu5Wc4Krx
b2xAD9fYg4/VZiDIUZXa6+xKrMjamp3TD26LV8LlrwMEBLf1V4w6nJ4B13x321Fa
yLH6OCL7PcHBVGR/XqJZmQemxP2//Qly9H8IJ+28JDSK15VJnk4HRqOOMgEFvI8b
p9DmXQRoAddhZiIRIIfZ3cjFiIxr0J42ru0kQb5xsBU4GFVOGUBpMxuHlCqHgGkg
u2XD3EIPovK+eDbU8KBk3YbJDXwJ92aJyt7+Z/jdxDwnQD63lTCtvA1EY6n1wuA2
oLPmF7g7/Da8/AO4KBj/FZOc2/XBevr7FVQoki5Z1n5vTGmns9BuOBdIEyCeOuMo
HD3U3cBXdFikxXQXGwV4uqJLT/X4muAIaHxXrCDEcKhMpOmBhjCJZmvi8etxB6+H
r/0++ro5LTwSjAQIkEwbHZnARB9H57Cy/U8weICxIp3767ELlL4TOa/krXmOpvlF
nilJlvw3U8yGIy81YunlY6UjAuNU6WhKy1m8OVhWi6KEn2VL7AHJX+LTjNINx5bz
MJgkIqSNOjRXHLUS7xRfDVuXZ2BUVF9XswTjI8sCkCLX9bsddWgPdKIQUWSaQCcb
oxz92ho11qoM3rT7DN7fiqtyU/NJ3Oix9OD+yY4wrq+1YWCkmvg0Pd3+JZFNTNdN
hZj50i0isgbg/ZHujFyd56n6VHDQVJ0lDc+pcNQTGKI/UNldPqRMvs5K/uWeM45S
6S7BsAHLvrG+Gix8hdFxWGyYiNfvxHj0UA6lH7dsHdx2kXzoiO8vIWZV4Oh9+KyQ
PLyNAXytuScarrqc09LJ/SU876gtNtc4bbqvmOqteYwnjWDG5XBc/SNpFOjc41f3
ufVqM5FkX8tnriOd96WJ0A1us3MCtS9O2LwIpfeYUi22gluEsW20ve82exfuIkDt
dnlrGdc6Hi0bCalQdE+Wfn1bLLIM8siUFR/4Q37U9l49u53kw75FgKfPRJX4NMCr
u85xcKEHm20+ed0y6XOlmo2HxnsPI+l7wZksGAkjNsjksk2UX/Od72054As4OaLP
AjsH8PG3A5XMFRX1WgFwunNkuus7aINS7nUbrezVA38bN/9m9EPRdN7MD0qjsbjI
T12wXEqKDmxvKC5Titm7wVtz9JwBuiyArx9KSERIhD5uWIplTa8hHI5jeyKqgS4q
/CeEkYDfhpEiQy95mRb/7Ypu2s1gwN0cIWMrVQXug81aqkKYnWUBFa2GF72ZD20k
DCcGzC5sJUSpjptEJPe74W9AawM9SWWZm/dYxaX/H31v084/Ev6qxJEI7trCJj+N
lpF5BrUeyknRliOJ5wtQmhKnr1QPfMrzrmdX+VDfeRZffQk+2yBsIb50jWFlqc7n
cM9v38EjqFP9kulFe6WaSewhUmaohsb5CArjgFwyUpA9DDPGujixJIwff/v5h/0x
K35ttkXVswVgSj7BGV7K8YLQlrO1C5Z7GFSeoJIGtcKlsTinxOKNEBK2jgj1MIPZ
2UyPTPv/w458UDUJ5LiIOdhKuVCcwM+wCwAma0bDTp0reBcglmKpAkNl/qqTF+hC
4sCisM4Fs+Uwkg5ilaysYCitQwhgZHUbULrYnMlojyD2gkUa08hDL/RueCoGunQe
meToOqs8ToTJp5qAPPLEMsLg8u+IupdWAuNWAiTU7p3z8MRq037d9+uh7uL2nKSq
JeyNEa7HszhyuDl6xJSHnROb3dgr1+cW1B8ftHZSe1EzbTMQ70PjyEWllV+Cqm9F
m23b+DmIAa7Bvk2Qi9GKIbudxglwbJzAFRlyfzEKEIdsPd59NPy/yVArnNgdhZCd
D9D+Yh5LSPyHUhbOG8evCfwJxM7P/To5HyICaJ7HTe7fhdITE3zGonRfWjFEjpjZ
gJ+MhaXi4n35XXt6hwXw49txqqmO+9vrnLJQPQB1F5ySozV47o40eKC10qaqU3Dy
u7vJ7T6A98SGgZNWeiE/n0Yo3OtSYprsZzSX+okCLUW1RmacDSBy+ofPpFv/2JpB
sFAkLo9H8hpTHECdY2g8lV1B9E3Ad4fKeyDlHyNtVxPWKw+v3QDYjNYEgIk4birm
yhnPClhhC1pPwinkkYZ7zcbYgcMVyAL092jpg2hr4yquMdn3WkzI7gW0DvsPNpX2
xjEY+xJlOu5mxRkCUZ8Ib2BMepcg4E0bMbKj2a0mybo=
`pragma protect end_protected
