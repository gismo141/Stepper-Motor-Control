// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
PaiNACs4iJP5KqIkf37La1MkBTHreLwG0AI1pCgMkB13vWddlPlQFc1aQdy4xj6PTNHhyUmiBm9T
MEMRoXhfkQHMvKEvMtUvu88wfu5fo1Vu+YmibiszoY/783quSQew1IiWVtq6df7CX1dexey8jJ/D
b7nRwFGXMzl8IS8S9rFvHwhE+gBvzla+XG0Yey6JF3PPlhkGXZCyS2D3SUJPxqrLTe71xnIqEDiz
l5HE/M6MxXpJluPZ/GwZiFl4Ifhat/6dXlLHdldTh3EIO3uMGjGMceEb4KUePnPFBJSClrLSiKih
Mm6mlE94smbG/0b8xQmVrg+OucuiXwhr5tCpfA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
YkqduLD4oEK+/ZqD3wY2ThU3Z4LwfwMH7Tw+p5ILDeWnum/1XImX6lqueTIIHP2PTqjfxD2MteMe
9ahsPDn2WiA1prNelWMHD8aatj4ywrKlMT1CD23K2x2PZa9I0Wa0b09OdH0z4P1V5dBNpAUEhEy8
Fr7DxTbnv0ZrPE0GjfwIjfAOXACtgfQ/3+DtW7MPs5nrDuokyKTfJa0Ic4BGb/HMBW9LzFAz9A5C
nA+X3neOp1i1o+WwXILs26aavzXX1Qy2k2BeoC+Xgt36yeKqu6ZxVn/lxZMnMNUlDN2pCxuAALQO
43damsKc8ulzOn1GS7Huf7GUXR8pskJMikymdQC/eVObqpfCNjux4q3r6lSR58wPwO8rU7HjHC39
Ne041Nu9cnZDEy5fezBWtad7XY15XTu/XdnoJTqNUsPohjDiPXT/TOix/2yD9qdrWCJOUvugk8Ry
TkEqdYPmhJ2CmwMi5LLdhu3aKzGn1hCkH/eUVM84oHEtABSqsi2BqCFTuuaqZ8Do1DtwdVaYTV3j
r3DTGWz64ygy48AsuCPtdpspY1iaofoxYhK1x6OUU/MzN5wvTm9iphGlTnZRqT5R94Yh2cYI2IiO
Xzj2rRuV6tLLoJ7QV10vUjVFZl5ax6xVGhnFSPPem/E7HMvFdLZtjjuO2TxoF+vDoirreLA4HaPn
z3NcwsOzrQqtwRzHvw95SkjnHrG3bwJCYK5pDVvesAFCSc4d8xJOz+1fWrWveifMveZmESDNqcw5
BIJdDysReoW/Jks052Y6hgy185z8R6yEyz069mWjDgsigBJGpajYl2GnOL1cBCIazMfbnMPz34Pv
d6SeVKSB5FXTItiJvzoGbOQwZh4sYc/jc0FGTnznU8mWySAHnc+/pB+V0pemjzSer0JzEU6k8uGW
Yk+8Ci6Yx+SJQz0SqVeS+1dNd8+eCP3xyRgsfIHQNxzwLbzTpWB+XmyHM3Q+C/M0TEiCNChvx28w
fQzzOV9xR9lD5Dv8nDSy9JjrQhebONpu7oWaI65l+RSBsFPzSLumDw5X3IE4em1SCRJ2iAq5D5xr
8+5A2XCdbC55yZTrzzbVlEqF8Sa0lUEjMJh9QOGS96eWx3saWafZLl19KiYhskNBGPP5iVXg9PMe
1Ir9sUcXXDV9qNWAlgmk8u++321zT04PkwH66tEIysyTy+0wOMeMysqiPGSiXmKlovDL5vakuDTD
suAMka8pWJjLClFc8ou9k1xYJ1Zc1G56+aj4y/JqU9UBD5x2TCQQQ+fD1KKMfAZxke3lwQYeaFSH
0+0Hdi+TOJvr9Bf13qg34TsZ691FBxQXUhwwZVbHFRi7DUFIzCsjBSZfe+Ex2E3eEtnhUbSiwxnf
sv+01A5CpFjLkTJPqxicvPJG0+jNh77d3M1Ws2nKUcs9hgmOfTlKntLZkzkN4RtEYAajdiGJwHl4
sFHwAEDDdMSUqQvq7oVSa4p5nVwfz0e2av3wGZMBUQe1oIYn2svTAunG2qqkFc70Y+PNQ/G1Ptsj
00vYyKLYHfVHo2qgPJAFrCeEZXsSdXkYileV6kxtUrUF8r+EvEw/V62IXYrxx3YT1chmgL0wSHqS
snoJkpyEwtO1zvFHCsnpIHwk7g7QIcqEFqgsj+o6EHlolCaLtVFFiug7OYOh9eizsAPFZQHn2jGl
vz1haNetebjyP6u6eRZbFehxfN9v8sF41J0z51S2ty9HseC8InUC9kHr7IenZuVMf/Fad8ioBU/Q
gZQGg4DG8c0tfBO+/BtUbXTkknGIJ6QiftzxX+DnmFUgbrMzDUS/2GusA5HENuIYlG8Gf9mH9E7g
2ADC+7MC/Qk0XDqyxM5UawnRWZDBAIEq5afeYsoRVyGQlc6XXrRxWacRJXX9v7+uMdX7WdMMRwYg
S23A2IycUfHG8ua+awDwTZDMnN+24GIA7dwlRTg3ZPaRcQjQCVvJPXEqUae2MJjQP9wzBm2B5exb
LhsB3K4TYo/Lva4/pvDnXfRxlB3qoLODNb+euG16uu1a/Yk/ZxpC4bAKgueyKBY0xihnuzDpB4A0
a5SCy66kUoMWA0v02yKGWdl8lX9BrILXAD2tmfP3352GYMX75jol4oM63g3wFh8MQTi+etIsef1J
RUX2jzv+5l76JrwaMv9Dfk8sMnKe8WEpR48qgBeMS3b9vBZPZ07+grGXNjmuP0TSdZTKWwLiV+l8
s0r7WHHwh32DsEmfWMfOcFBRLrLsUawk+pUPMXJvNGe4/6AAMU28RnWeknzYyipB60evSlfyUuMl
sHe7RtXsc7Dy5384DmlhgyD2XIzxZNcB/EzoA2L9U2qq85CchalCTjHjRwxAIVnnHs2SET4qZce3
tyEnE5SIBWGHQoBl/X/mCGsdAiTP8JqO4LtCuKA3oR3kd0iK0y7ynG+14qRNzopXdP6BTthW4ggn
Dhay3WPB+VfR9T9haPHiBfPM1EzRQVnlfdyY5k1iYTSSqV3bD9VHhNYTKbQKHRAZvZIc5RUG4obX
oaTAL/e6u0yBMhtR/amhkd7RFbbqaYgCpxCkLp0Av0ZekxwGY6MfjKPCF2YBiFh7Q2GZKqaetNRi
zOMFRhJJiRK6PjHxVxZLA6AKR9sc3c/wZBH7Nm8lLtNxDVyGJ0wVQTLzxWMnPcahYHTdVmIkqJbC
eNJlrux1x7MdPAFiXLcUvWjLU7HSgKfp6p550c/3Lbd4SLHhZjOnLwQDIGXuGSt5S8vnuZ3lrlHb
KMsoSR8SaugL/X2Vg+eWglAM8YgIkee6Ndo2oGs2FQ0CveIpdZmbtPXMq5bC5z711bzDCleF+SaV
2XazrzNVFZzO5KdBej/PR9Jdal3RoC0T5QEwx2+H4VsI5d1AtEo+KLCmAHO4co1CgbdJkTeUQ0W9
B/N9RWab6V7NNYa3InwXA0IT/pMcDCUzCous4+4QvUlkKZgukqHydaddNiH5WoS5Wi76zBOf4e0b
NzhXjIqEgtJtY+eLgsqPJSzZlZXFsZWopaPlMIGMRUI1IXO/GHy+bGX6KcDeu4MrYMyk7n5htgvO
ZHJyaotlUjS6pUutr8On3Ic7fpGmJbkkYLFaaDsoQoB+LgUiciSwwcj71NqQZAhn0nSstuSgiMR8
Bk2vuPJUX7JsuFJoaTeNhcZs1UUZlAqFiD0OGJ1DX+lZoLutCgAA/SAH/fH2taMm7luPWDEOrpXX
U6bikwAIt4PEqR0I53fDSmDDD3rk7IkR5sx52hgBVp+NFOmjLFKq/jC+4l8a7fsWW29OQG/CwyNb
P4+aXWd6eB6vToTBlRhFSIVt4zlmAWqE/FAtr2+htfO5/lzxk0RKpbevXNXKxeLO9oRQlQsIJ35f
TjAwMVJ6a3MxiuEf7zs2omMKlH0HxSr1hH6dbTgs2nZe7Fr9vRq0t8gBAkdKm+Su3OMJeOKwcqvK
zV4Rztoa/lM7+u53VQqtcltVtAP+GXkG4qgRpuQMMMum9O0BtSbBzt9+u0ro1UAjCkR1PhKKfW7y
ZSMh1znuCPBb0rNOlyi5p2CupSaGVERp5mypapdBgOXOALSYbBVR/0HxW8zXUp0f3Jxlvl53mIbs
VSKVEHYd7PzFUzpk7ajbIHHWeZ6rWr8As1/wcM6rrKT5tQhZyvdGiDRlEyNO1git+k35tRcuAkMo
l+EN/f9DE+9ScaO/meY8QXz9YLEQe2A3Yyq1cQ9P71LaKF+GndHQ5bTz8VLa/sCN/YveicSAyOgb
PEJQ8XGIuyDAFXTKCWOPyyjda8fYk9Uf1GmVSuXaKk3dooFm7nE2sQBvvOmnXFLOI+RkCQrD46SY
E/kG2KwYnZINfTu+izotrCBVUydsJ3kRu6nwPCeqF+exXDFsaflxq0Ckr4yYNa9Bhgypxs/7XI+Z
k7TJA2c9tSyh3AW3cLfHfPveYVvPB9QoBOyIgSWgwfIRbQF+Up92rZRaNxuppuAhRhC3M4c/x5gd
5YQqulD416UdYgMuY7f1T7ckZRSor9XDlGKbEonPJplhRskygX+7yZkTBBhy2UnfhDkrqmvSDoWj
MhyESEjwmDK7yvH7LCSoK39EPAd5pIWFQhHOCV6cwYONZgb1s6qbhTDFmByZnSirv+mJKLV9SjXU
IJ4XGy5JXd+Rblh2qgUDRQiwb8BtyPwILTaGjSJbUK0j25xBjU6k1vCehUDIPasvzjdKaWVHsv84
ez7MQ7pAcPqSSJme6cGWTTUHozG6PHAKIjfHqZe+COFs6bjO3ZWc0XYOn1PGogavQ2f6ONDg7X7t
2ggMAyULa4Nhp7o2Q6nSThYhNoTiZ9WEcMgcrw8jN9qTtcXvrUdy6wCCDaMlLJAC55y641ExqVv5
dGZxhvUZdL718y0bhKzqHGwHEPVJiuMq1QSBNd4iOE02jqnulpien6+gy5GDIp8fFIAsxjTWwZYF
zdnzt33vGJQ/Si6FeSgIA/JGgLFPVSWACiglQ3ygIbvvQ3qH98iYGbdGvwyx/sHmeKtXUVc/iUMi
7a01nJ+g/VjGMLEbuR8OfaWAagXryjP5MTm4am1TsFbFcYlbfejXWuG3olG/n4uYEtBtV9Cfx+99
udTLaRi9XRH8E6W2Df9zpAQfUEMXoDFScNmcD1XbVsGy1SbQWRTPEVI8/RBWx0JcBW1dLjhWgy9u
p/FJ/QwviLAicM35rCdeJmPqx+9P6VWvFDKefvwWD8sUBhoSYGzdvMcmsc2oZVpHI1/FYZe1enLk
z27JuRBBdF15m+ozBlHwWbjkOXX6Kf6gcnj4rQDvwf8INOiDBcs0e1g730+IAW1hxpPI1UUUtu//
7IuobVZqE/xoCC75gAfouV9vOZM0YfNE54sPrKInQcOFHysLqayFS708YMYluXIQjPi01LforB7R
XVaPlUnNFYrTUPAVrDvnQaaGfdhv9wfzDB/MrA2Gh0YAl0haW5dT1PDnHSgBpls/oFmJAfoIdy4q
DHXS6AG9b2vqDXsvLwDSebTejhP3m1GDhYjTyveUmjiG4ngcoCiYiq3JSrO0O6sqQ73o7KTpqVgy
wrJC5fLROidB2YxkrTwnZnCR+Reqt3dU08WBXRquUEKPl9uRMH1xGdgaVXIKuoHIkzFsOap8nx8f
+ZQYiPyVX/JZcK2XxO+HQzjS0YhZZd2S8RSHC2uA7twVWFjDl83hb+NxKRaAX+vVvb0mudLk9+pi
iv5XKILRWXhhwkxNpg0H/LF5fYg9Ojvd4KBORTZCCbM3eXLeQJLgO7eiilET7d24GZsBq9u01LhP
BWQhxI6N2V3RKakCG3ZxV9Kr3mW9jJ28vGjP6jg+FdagS1AYn5+uH8nIo0vtHPUmq7fs57BUGIcz
qoAZR3GRvI6p3MOezRb/L+OWmUX5c1MPrOQYENyE1lozxo1o4RAFRNxrlpjclQG7pkRO8R8p2Zyr
QxXSieHYvTHrblVXRPaN39n0q3xYGWI7NsPzB6zhwj5CI96L/Cqc2LwArnieWwqprN9hAIFz0PAu
3JOTF220pZ9v0PBYPaJe1e9M0j693zKd0VA3/Og1ofRbicRih+WGROPM6ReFnCIltVphEaCGMkxJ
FaUJ11pHyBf6zaMIu+P9UYx5px3pJtlOWo4b6LxU5VVIjY9ixA4yrc5srP/VSd6fFmmEGvMGnY++
RloLJVeL3Hk4/JCB1JH/laXMR2/FYjXXqgqQNKiiVp7a1P4zkSAvrv1E3/LfXbdTam0mCKiDwpNk
chLY/UR3Bt1CIsS3stKIKnG6Kv5VwnTxnfPLH1WaTVk0qxPv0GQuKZgOt7VQgNDJLqiLDBXaBuHQ
zw4uHYV7L7AEdoUPStBko3ieWPMM/HyD28KuvIoedrrdxAhhYNSnt04yGeElo3ZMR5RbEgDxorDT
Zz5NEVIZHs8pn5iNDuFabviQzOaqoxigcKkHGkMdYWcCdeHQGAZblFEeP8jDCo1Ynt/XHwIn2OML
gFA//9CHCIQb0pnIltWiD2yehqixX2N7MFBoq4wB5Jog85lBZDJyRLLQYyHH83gkvVMRm1dkLpQU
JwmK8h7ROmrUZfBhVitQNGhdp4K7sl7TJbFIGeOr9kNIk8stdx8g19PreTr1APXYqZ91qLRz3H60
bnNi7vo06/7zUkFyzYekfMjSpc9PJEE0vSNDjKT282iY2hHwqzkaHWjZ8gyVrsSlo2X90fNt2Myb
ge+2he4OTftLEf3yFTES8KPRpJYt4dGCXKn5v/u0ZhSvQ8a2eb2Chyv8gRhRl2SK/weLtcWA3s+q
arxDT+dsGVpQ0Fff32R2C3HjFsN+gUAl/Y2ynYuNeOiDzM9cbqZ/2bxm8JJx8OLvqv5qffDURw86
fWuTz+t2Wpw/HyjDmhvYHKy3q663O0oO+LLmkJXfbBpl2WHru9uoa++chbnvKRvCwPkgwOVHFw48
eJSTNwGhC6hZENxMTteZRdQDXfpN4M+NadK+L7muOwG2lQyx9+5/vjTm/B696vYG1i00UmpwsE9j
XZlF8Aql0DEISGgcrgV6ws2AECvGK2+1cxdVJ4iPB8w59BcmCuWJuOfze5lSP90iEeWimUbIozC1
2QTdpdWgFL99svcLT6cy53hkKVuNPPPZXsw0x7PQp94wf9RcS4pFgrcG6Cg2OyeezCmrWeYdmhMi
2bgVi0/aUxH7HRea7baNTOK/Tm3CnmzVxgBzYZpD1l+BNJ8F1gpMGXiLRIiDJ1vrgxrJ0pu5lrrY
YEnf0ICw2rNEQkIj7OTsOetUfCmP+pU1iOQ+zUUDJAIplWCYODggemxiAaUrR7JGVFO3oKlm5aeC
B+RanxA7dbUU9TIZgRlm1gWta7k2HrXl8H7W3zRdrEaMxun6zinVdXOCJBo61wt4DKwLX2isDIhO
REGCY0LuFIqyWFNW4wOiTEdfY3IYAsmMeIYktINrQsGR7d3dHp88azVm9qUaT1jzKWkDN03TqKXX
EgnInyT768U/3vVaO+tRbFbIoDYFrBI1qO+HOEbZsZjjENOZ4jboHBcWBoipV4jHLL4flxndqK8I
MLt76ioF1KK2gk7/0zaHfisbjRR1/d0s5Bitz1CPuVr0g9wbk3CzKhvtQpnGH/mdU4A2AW8oeK9u
TfJy7OCcKGwjPIyPgrnENke7T35BJQKURdxWdyF++uV8+ALJHU6V/7Wda23yVhb06FBZqQJwspgK
mLWk2kpUdYhHJ1rxMZ6pwubh/YxU+JqfnJOcDmNzpjsr4Broz6LtB5nCi/LP+VDIZ9yDL9PLDRpI
XYvjviz8rcUyFSdeG6Tr5IX+UejdZtIerqdMD3/9akz128eIF577DgGCvSpfY4deTCC4kwQ7IO3d
m/6aIfei1+mKFYdg/oQvKyn/8tCOn5BA5BKZBhy11o5DJqcUV15NGYhn3sb/UZUCJ2VrkrjEwB3o
9KaPvV+w5f42j+Aivm66bqImaZTrMnfka1UeQEDS/51PxbLh0/A61q71XyGKVebMeShbJRiSfgjw
8EjknSMy5D/oMA1yQ0FieIG33Baflq3deLiCGCwQfUR9azPYPrV2K7x0E5ETzJFZ/aCN5meEUiGi
BwcsTYXySK7akUmCC3MnSdKtNeWIiNz+eBae6lqXHjoW7/+iw/ZOfx2dTuKug4aBUFJKvLf9v83G
Xmcehb+j3od7NklP4/JblcLuSOT6hmABpwQmRnl5HPd+33lltY8WVgfBSAFqCrZknH/U012g1qdC
CHsc4wMnEen+c/gFtnSfesHHcJIrl1/8kXIpf5W6MxyS4dcvMNW/vaGfyckPMa0Mn0xgriBIoLpq
prcEeY2kalG95QGlqGSiNVJa+P2o5pt84CzQviNCNzTXWECAQcE9CHI10xVSeWlf7x6DTP5i9kCN
3cy8pLbYoVutrsp0BQxQ0KUAgukruwe7TQqFXXULqK+D1f4T0cuBEKuXs2CMS+V6nDmM18MileTj
bOaiN3I1xca9JSPuj9+hShHU7nGsYaCNB4IuDN35Zdpg4Haiqzoq/C0jB6ST9u/pBsVGG7SOr3gK
KVm7gvzF7N7QYP90qg/zvgNPimzXRAgGromqb42HGNIbog78xgv6KWygP7yhpqqMOHuWMeomEVL1
LOM3yK6hWEjTziVcVdM9DI01sErq6KOqRT+c21qSCCefeJbCQL6uW1ehvG0q4jtCTLnrL4y2ZECl
OCW9UH/lHNFEr3iZKXKf1ybfxP6XZ25HzhlfbQ7es+Mam+I3iS5Intbp+TB6nmvDJK1sh2dL6XZA
1TqGl8t7cATtZ5JpDq/DxH6amIMCVBDmF33OAu27dxo9/38nWNwLmTSPK80KhYiIglgjw5Bu2XD9
aPMEDGx1cyBq7qK3NpYOYc8IA0FbsjgddczcOcon0pWXhXc4SNzKijebVk1YpyxYbH5nYZODYJZX
twDjSIUK8NhgRLRCFzJnPEX8rzee0l1W1O4y8dcAPm37fxTkottjUL/uAk5Wb9vWt1QdSn8VuDm+
jXxcAsnSq/GGl+FsngD4XKXabUOIRvNnaNlbWRirtZ4cEZsnYyJrz5Gxpc5X093xwIs5zzOVAU1y
6ARp8xvD6OaoBo+ky0wupzanZ1A/mZMltm0tOM5SdlaO2WRVoW3t0gfWL5tLIB6uO/LQSdDg1w2L
yuCDPBSAOMMX01yCWYSex4AJRviRqiY5JUkfnIKaNRt01Us0BhTQKVWTCK2kjd2w/JsqpNAIsyIP
3e0E88SphzGogbfAMJrYjDmsrFT5Somr1jl0VFCyvL60F3rn3E6Ge+YDBcYWu77QbiYgrAmQnz84
9lP2iiwQuxRFv62zVn/NUKMY7hYhP5TAgv3fw1DMJup3gfSX3w7/ynfyb76sjZmCP5cXKZyUigS/
elwJCTQXgpw0vN5eDFG4Ni3nEsxyC8Xv3YuXWDGkuXRQmfsEhC7KN1coSyB5KDITqFjReRfyiR1K
W1aWCqQJbcbX5+/vPZ33pssnBg36ZKrkV1MWsx9G3XICFXIZEH0565I9SO5HUFDUJB653noowSui
C5eMZWQd/mVQFgku9HSGTuS6zU4MHL9wbmbtErEaD56d2l47/+mBLvpnpHZoAE9P+TMJllGx0FtZ
2Md3NPej0vxqBnEy8kQCjaU9zEXKa4zWc15GSDTanCypMAPIHoDgd8rOe0X9Jef2BHCsprsLY/rj
z7HwB2OI9GiK2XvUlEygHFmBnIiyEWdNHTV70Mtvwit18GnLZnykX8Mm5DA/avwnl+QOoAenO5p7
IW7XxcTTGpwyLipzUcI2AJCke6t8S5qXtpcGBShUwiPY7LOLvd2hcTeabtNxUNAz/EM3kbTqNXgQ
fNL/7Dfdx8c+nq18DZX6/FEHkRfCi54cpngdqSULCLRVX3fNHORyR945SUzCQNywFFlgKOGFfym0
QJlUTlKtlopuSFLtaaVGnU0ZAywo6k0usbpUxR6meGMekOj8dDxkgKvGm57wzg4snp05F3bgREVz
v/EtoeP1/7OfiG3/HhNbBRKWSM3DMce11G2lrFEErJDi7VDOHYrODsgMW/2ivVAoSh2VAqxRl/TW
+0Vp6LYsvMKkpoabz/HDFbqvueAoYBYtXvAPZKTONMLiI+88erFgl3R/BSTkyxJOmvFbYKbbK+VZ
IbXKwNemFOH5lYon6ruJlgK4KqWhzX7zVJ5vS67V0FeQWIVfOjRxECg9JmyTJVpNdhfw1zwo+2pE
kgd4Hpbx/xaS/gdfO1QyDl/G+yJlNognfhKd90z5mEIxWLWnzu5c19MHa131YL7+ghDo+n4jd68y
H96y/KbN2w2/TahoBvMEk0Fw86dDfDnE8M/3Ak10hSzKP9lEdYGAstiPTaPuzCkjJCtyC2+ZGpsl
exKAUIoIYsPZwRSs8meI6RPawYIKbEfA98xWR8dtyRg/oB8OkcvTq6MYgWWWcFMiNrO5jKAL4hLo
+L0bz/PGCn11vL1lyC5tDilQByA+/D6gWWHIWS8gSy9XV7X1qV5e07tL/WCpdLNEwATBk49CMf47
Nl52N9j7/FOLkDZtiYwbS5t5HSbzFBGlT3gTeWjqEtyOeDMzNlA6ID37PCAMUYsRPZ9p831DCQWL
7G1Kh3mWlNAh86+m+SXw1S7vlvXulzg3hNqK8PaADJWmAhrSl4Z7BEJi3zDohEJ1tDBPdgMluqJ6
GBvPkCN3REXBfFtcfJP1aq1KFiXnXh/+GHrmwm6kmNCG8/QBQBzdGD15JyMZBiMKI71zf4g2bGsK
cahU/wXWsZCeoV2f/TeryfCJBFt72fqnvUr8ZyeLTYCyhbT3NymZw3XnZ+75jM56YCpoS9O5hYxm
Eei3kNZi2GLP2GTzzZvHB9wGD1xmVO4yu/cEfDgcl9cas5vwwD26dOqy0+G4/oCTFwlqc9HTz+Pn
3LF7hINRjJ2wFF3/jgzC6XIx7m+gq3/f7UWAMAZyfPQgssM7a1HgRy1aJlbkXQhFkgQiEpLKm6k1
D9XDhkSXANAGT9pMhR4fSdhPBMQV8eceqZ6u07Nxu1ZUmlyy/xf0nLw3B7cgNAmQ3Qev5xD0q1Jz
hTFXQDn+DDvZIwvg41imPt0ldN1lCu8sWz2wrnuzWJRy/iTjIkAUMKzOhs0SB3pZPpcTEVW5r+dw
olLgIgtfA+gzBEQTNYQR/ec/bCnUVNAX9tQVal0BqgEJHWBb6KIEBno5p1Oap26Ejaj2vleCe5dN
C6ZMOlywpqZRiHB6s/NJCFy2EO3v2EVogsQZFLkEBI2t9htOF/xPpqHqpcdMy+dZ4C5Q2bNPafog
hwiZqNi9uXCwvSSA71KQYQAQw0mSVKcyJ/kEwXSAztItnwJvM9I49Wvg1pwDqXpvr4SHu1LuBxZO
Z5qDyPzDZvemP4JDZEsMjZcdDfmmu5OBoAsVeL8562C0A5f3iTFK2nSFNOi5OKYD3QaaumIb4Ryn
8fYXttFaT0/sZ33d7X/lU20uVXNbxpOZVUtCdkc+z0+AnHQhfIR0yiarFF+pa8T4Zx/zAFj/Dnxe
IV73IYYLG+4QMpx4EvlcklOZXMXvrCNYj1lVisY9TaW8vQsTKat6RWpCTeiilCLZOtfsJxOlgAid
kAzgu6qb+Vz67llKqYp9Fqsp72mfC2phEEoUwaSr54JKgjz/xqy6UCVLbI5pEWGFxV9IghK4YL5X
/pW0KqeHCmRLodj0zVZDxW5VQumunZr57p5xpDmKTVRsCBHt2L/jKQmY0Y2MWyEKwe8W5mhdGViq
iovagAsDITJ9OooibB/BJzWhDDgrhR/IUseOfGPlAj0afUyfnCzxDiMN/mEIk9ENMnNJnvghNaSz
vgfQlw1rYFxSaV3bptQa6Vif+WIIeV1gxfFhHfUh22jQtKUuHu96LOa99AHFM1DJBsc6tqUaAEPM
eVDD05xTTdaBCGimLnCez4s8X7Pxs5ajPR8bRI3aD/1XQal20Aezqx94SM4ls32pMP6Qy44hg0nM
EfzwN1Q429cY5GMCow5SQJHmazo7T4ac+tNUS4FiBUy08t527QNyv6CDXZzjGS7IFp+4v5onF5Qk
u8ZQ0KfJLd1w+Vvr7gJKonfOW1MqoSy/vK5G0xgisL5EmXR4gv5voQH76elghK9HmD5aCORfI+rz
1BInUtWChPcvR18v3ckisNkuWJFfYPhl+mu9dlR26M9JrnprF0NG2j0LOt8WHyn3lRW8f7jdICQy
xqmg9SIAXqB8U89TravvVzqRgjIW0b4zKLr1fmKn75yfgAv3JqTjhaIBRFVHwlTdadhzSiVUKbzA
v9LTfrUKo2PutGRgYIt88Wqi6u6tyzH9rONNtYox79jqrXrPxhfzZxNwKmqbnrTA1oBywo+m2itZ
cm3oQwvWAAD/pCrsbrkflBkXM394YyAItQ/5BaAYBXsCIn+V8Dy9xh2H71meV4uvBkzc1IRZ13jS
lF3RRPfKUunXCVYaLHGlVbrkeaRogs43f6pl2BgQn9izm48hSYfn+nS+sj5DYOkR8gdNeInR2T9S
MCFO0zAxF3ZO0sQKN3bjf7IytR9LyPTvMIsdOdkyj+m/nQHPF47MC0lGLzasu7PWDftRqgVSPkbe
40hOL9NdqPpqy9RLaTiaPw+LGJ0Fkp+nFcbd2Hyoq2VA4Gkh+/epR9VB0IvTvPur7oZBBo6+zN0Q
R+XVi3XA+Yptpw3UuZM9e92vNPQ0GSDi1MtjQZEsuA82P7G5p4bksnQjJG32a3NIFOEOkVvxBKCt
uLG9gu35xUrFydBUxLPMmIZ3Q+FKdLAWUI2wvmGk1cqx9BMuTSAFVwpWSo7L8kljBmFFK0ogDOIQ
P3a3KdUShXZJ7L4cIIJI2t640Dx5XWe3dLBQMkFvXPLzGM/Hj4xLxIUPNth2G9uazLelZFbxEmyX
4GefDlt0om3DNLfviTXmHDxjQy0XsVN4MeYaUewyb+xfarNp3MuDhMc73N7RdbMI9lyp5748b78Y
CiOmhoJha2nplMSQKjDhGxGTQa0kAhkrfo+4I9a6tL/lxcpEFIsC0OZfwKGfx2u58LTKi29/wMzz
O7FaFCq27+q48LVXw4FCfaWid6fKCSA9KTimw5f95ZMicteQk9vkPIVkS2SN+h1cVFzlCzGSZTNy
0whdTrrJTikzeSgMW1FF6IkAKOnjhlPzE0luJb/UXAUspFbiT6QDlQ81c9f59Jo62gKbb+kDOTNW
5Z/05NtwYM/ShkloEOZ5U/uVLg7cWwyimt5pBJh8xwewHsQOhEYhaMbnEBQaqFPkE0JKq9z/4TtK
5e91dLEJ/oKdO5AWJj05FLoqRSKFWX8/dTSvHzqJ+vMG0JgMdd0AdeW5dUynpSeo2wh8hrRgDeCm
aRMS/mwPovQl/7PqL2DKI1RyTaffIv8k8DyV2K0+nhnDYXPunWP3M9qj6YPAalU5jG+j54pLKSaE
xXPXrCVl7DgXOdih+91MA+GFu51xrgGRQEORZ/15FX01C9fFz91rBQ7cAVhuFdOKyVIOWE9VGeSk
OB9kpEU+IWwm0r+mv29QtaPik1nxmy1Sg6mL7c/xnmg96Ft371iEuthf69ghoXgSqDrqSQENho4U
t9yCaPkvp2NKmSX3yrmVMvR6++4WxP367eb9xNHzpceFl5LHpJe1OHepCIMfcDJVqd5Wkavkhnsp
WRIoT9cQUykcKtoM816fHo65W0xFzORdQ8vxEOZtiBmBHsT1oI5Bok0lIf/KU0vugU3vf2t1xqOr
boJv2RsIOaTO6Xr25uDR6DUJVi2EnwTiVboeGKkCPKVpU5PGkSY81NTO2xsrdKR0oKl74m6y+VPs
yzwYGkG4VZdOip/uh8wRPc4RnLiMPNJIcGYjUG5XCRIKQX2930CJnSE49UJ18uylW8jxypSa1uhe
JneIlRmXk3ByzIL2dmqp16BQ1s9U3GH1yIlSY1rVZhuyGVNmKln0GOp559/un4Z/6qpJFL1qlfIO
0l7rCTDRzbQnoPUuoDqIzdM4NfdSxRluQOj4R+PGj7ayV+1zVVd/5fJwvSMQj37+pjqNTf/YsfnZ
i8uo7mP72Y5481Nnm2+7RxPqfBlE6nuiIZ0NqTrBIEBdePyC2GjD8njJxCVQlmBOweEeGwfyxzMq
8yFEgM+xN4U7bF5+OJcazDgV7shjSGME+0D/TIspwpBh7P7eyylmpMAwRBBGowT8Qng88TL6k2za
eBzmaUP59CSznhASd7wJDOaYn0Kzo/MN4p+XGDA/lS8KTF1cdEH3QOz9gmeYt5U587zBtHeeAS+f
bf7Hbclh2Wna6AFFIXfNEgzblJkIT/PJN50ApVooZTaIS81r+UFXiFvbBR0rk3QSYejr74UaSWzH
Sh03JmzK6aol+9L+c8xFtEoqQoyYXm1Ux5UOGdr5G7NWdAZYDbKTs4UiJXfpEwVxStHmc34U8SFr
uR8zfq8nVbdIIUIQwp4PDpr0LxKygMcyALtUG5+VQCmvoRFdCEQ/E5J7Rkp1l/oRI0vNNSpD7URi
JWmyHRqs0uFqdWbEQPWc/JL5eK8sBRkmPekybhUabnXwtqg/DxgG6qqjR7MZxIDZhLEvIZtUKP2/
KOYobldLQsQ++cK2kXYZPVwYsGbWO8x6P9VyLKeQa3wh3voYR74dfqUDTnGOVK+ppWIhw2NGSwHO
t3LMUxYFyDNVQ8OYKwDiKn99lZTeBc6h4NWQnlbJYT7MohZ+X7zu6XKhC6GkInz2NDy+FC5fiw0o
xZN39ZgclT5uCVxDbZL2r9KUTHZm/LOcGnVCeW+tJBg6KBp+7cQYFbQBNAMwgGFpsEzrssWeK0bi
dQw38xTvRTuafMeGsd8epIf8lCRzdOhr7bIa5EWhvnEvEYq/P+qndsaBKuBAWGhu1pkr9Xdwn9Ww
fBvWEO+G6MuOIaz9hjbrU5ywYA+S3P/Sw+cO5NGWCBpM9xV/1+9jl95hYjusr4svuMXV0BgDBw3s
lAIcV/J//lFKOrvk2v4Ey7IKdihu7aM157AFcth2ysArpj8G5k9v3G3n0Q==
`pragma protect end_protected
