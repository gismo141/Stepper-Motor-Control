// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
Tx58vCdXWmYAQoag3aasc6HccmDr4fO9wJBR42xDMQj40pilkPF1znNDz9cx70SL9NDO/WmXLpUy
+wsc6iL2N6ehokbBiiMSxktEZj0WYWZS01VJEZq5ZGb/NSdcCG/C19aLqa6daKmpBgmgcYpFJpjv
DdDrg7EkVd1wZtiEbC5JU4GQ0ZVXQciBqT2Y7Rd57zrbubiXMcMgc7Vn8jLVMvlH4d5fTf42+GAa
PrGuSnYAn/ZLNr8cOY8ttwKKdpwq+dy2z0vjRr7iormV9oMiYHoRECYu36bVYj95NK3oB+xwl9xR
K4hW0aMJfq6kg88QSWTBZd9XKGVzw1FxrsA0ug==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
WKdjnQs53lNERUrYslGVZ98AF4gJCiC0We1F3vxVClaDgHLFKiqAeu645PeJ0Ac0IIRvceow1jPo
HVTp/Cmwp8pbD38ZGdkIRq7pzQfixBkOExNZI4z27PGwj9uZzSmDuhmsMyMKV0L1wBhYO1KH0LJJ
oVrRP8aumQF/XahunqLG8WHLM62CYAxi/aEf+9MdwtGxwfPT1IYewUYKyZUv9BqZxvxErRsp/d3d
ZkuEMoF1lSJCgkgtDCwnfyZyjCzBqT1HIYJOtK6Cm8X0ejsJ8b1baauxG867TGgn6u6Kf42OGdsc
BjCK59w3636JCWr5RG0SwMog3OSYtYnNyb0SWVoDYjsVIiDepCl3T2poICgOydi8tCwTN6cRaJJv
4wrlOmkuiUeEo3pL1nx/LNxitAyuGerBzSym8zT4XIj//zXhJseFaRWuN3AQvljZs03O9V2sppRR
njnEVFXuvdvCO/uX6QIkc9cBP/kovP64M2hPIf2cF4ijRXyZfN6s+maC67z6E4AQ5uKZE65knWyk
8YFA6hMtc+x9kpE7saktBWYqEqxTu2FALI1ItcdKxs3Kng0sXzPmUJc+usKf33bwyLJZMqeVOUEq
/2AhiL+U5p7NiczT0lA3rrcXQ9us2fxiVSULdqPL46sZcl/I9Bk9m4ehYzutix543UO+hwZTAIYv
pTgMZXj8OL9FPntG3UHEKwoGAJfv3oZkNsD/JLIukkBOkMClgo9uQN+qXyC1ko24szbNkH7HFmA3
KkDwJPXsy5LVv7pq9EytQ1VHLDd3JBmu0T1Q+mN4IRDmic74pJWd79Dsha3kItSuc/4+jEXhLen2
kowTmiLgkSZ+czdufIPuObRfcCdqpZKGchQTI1PsQzGtybcZUEs7mf8E+X3MebQcUs6OST89eFon
11++9DBoBvJebeqESp2EQOhqo6YJSIQQZZCUwocSOxPQv9oKBCNoZlT/0Yl2wOnC7iZYx8UOkyq8
7zP8m7ghqU5gkCuzXXUqWF4UBbv05l0EWKTY2kpig0liop5ADq1Ymz29dNkHq0mmAQXjZ4pqf0Fw
ZVeQZPeVcQ79JDvpXzxnKUKV0GbW4Qn95od8MtUxNkT+xcnt0TE5niD2q+DrS4MCOickcQ4Br/90
M9IBJ7YJd/OoWxs3Q/2/7+pUNb2uT1M1WH3lLIYCop118eiO+m9cYD3/qRx7cmEcokYxNTrOEwA4
S6C+tDMie0AZIhFBkTbyd6Xw5Liz9RfBP2D/MpjQky6WxnvE2NtcNuB1CtG7hEa7ksNWqjm5JBtZ
Y95GOLvPR3PvojFq+ICJSGlOhbk8K1kAUCQJNt/xg3Z1XOHjcy/L4Pl8zJpxRjTLlfOhf4wEK41I
Jjfw5YfaANL73i2Ukk+OEuqtu0kPYbpy4JTWDMB54k6Y5zfNqXY/baJGQB6GvZFD6s7Ep7b9aNDY
DI2EqP9RiUyoaD/MxSBm6GWJ2i6cxaq0ysn6rM1in9WnCexBORB4heLct72zXKMHuAREyDZtycie
IUC1o8pRVkX+dDDeZ/klwbMOyfnoM2gstSHa8vK7G0RoThjmbkLN6jQJWAqprwB6cC7Kd0Emkx+K
J0mZS8otpJ2ahHzybY/AShZTlAuctkJGkLPNX5vawQf4teVT7cfgfBhbLjXpdp5JbgSuPhRNTOeA
/D2X2QKntkgeMXM0tzGLjKsoQCUTZb1E/WElR6H0KrPHYGQqDvDrlqBu6IC46STFUOv5C2MegxXF
epSZ3rSBZFlejWngMAqwGhpuPmwojZqZZRBIgRkpzE/tyaEPQb8joGlkv/tHZL+3pCJAFjTbi5uT
JoMVTXPbfVdFsF+lf6NvCoTqrJpsZVe1ulSHl6AODB8lCGxwkT6l4t3zQwTxhJNxVjj/505pXR6z
HsX2NBjLIhhblMhB+jICpE6vkIxv7hoMLg5iptlGYIbyxPkppVgZR/0BPBIAZNkwdFs4dBb0ndEZ
rul9MaljITwb4onOFmMMukac+lpyKgR4Nd1E4UnlC+L457//J9qKraulGD/8OAIvwim+1qe2a6+z
pUjOCHPeBAIehFNO4eQGCyYL8pF5rFeEd0AE2C1ATUTjQ4bOk27k+81PswyjyjRDt0w6crmxvOIT
2C49OAeiXMUHa7f5RWVOHrbO5+z5rC2OHZyfu+R6ElT7fyNkZXIoOyyHzuwNLFMmPrjh7kO2asS8
6Fp+I5uMu1uHNMWufkr1UN9Gb33+56xEX0N8RbHAwWrxwa4gb3ChVH5gaN7nnwkju04JHhfrSPsz
bNgalm6mQfXKYTFVE2HFrskkoej5MWs9z7P65PQi/0blNNgMKdPdBLmiUUGqdgcn6LsCo9Lr9/xM
tenJ3IQcx6HFEGeIXPymV9Bvjx0lYscB3oLA8jwQHvpXKfCUwJiNLH4qjiKsKe1bahq34oPp+/jw
8HDRjAImdqmISdwIOUCWiqWIcvI5tfOHdLQXzCeqw7BP7ihBWU2zxyUnGo94BhX7mUVfh98hpTjM
fg336bM68WQL+GNcrnBgS4R1Yufg7HjKD5BFdS6SyqkvL77TSSkuiLPm7Gy0kvXIvmNprh6HdVjH
rFQutc597oo1G8HKumXjzKwm9IKJ2B7JBXToTLd9FMgUnR6z+Nsfy3cOZD9QDBq4YKDjujgOwer/
RUvD5H+8U8UKFaczqZ40oJvaUWdP9BDi3jXEF8eFPTJlI/1TQ+sx7jg/u2DA0s3n92UwSiH+43sP
kJgwW1jMvpviarFbKB6VTIAaPvzZAJXrpylTw1FXsuNR/rD+TJrnVrRhmPNKTxQ4//OkG3KPejRD
ceoFaqjPa4hr82VHW6VPsrOF7BDk+CSCw1t4FixXz/Cwr/+qpcpnNdrmmF9ISwRujraS1r5Xo0bV
+ZnTrD3euUQtNhMSwdP3wBaQyIjOIN796zQHMZG9jnH1aKkvjupJH7pD2fcqe+5SXkTGBkADCGQQ
6mwamLQTYol9UWVCv1qatPCapNdksiZyjkIl+7OB3Bufxr18DAM68U/mq+JvoAD8m7ig97nNu9PB
1GhwX+yjGxKZ6CvoOiSyLeylyxLdqjP8VyTw4Ltw1EXbCHXbPrELsSHI7B51o1kPLMi0uswk/DAr
UFbGWjBJSFrR4/oAuJgWxEWh96X1R/QERvS6drK18YGU9Q7nYI2gCXSzYPbstoecsV0obe+6E2j8
7dVM0eD8LakaU/Omb4IfajBH2W0KQOaqRe7JuwvAnCQYIfhziQc4mM+QwPQnFOcCuwIKpDEav36r
HFAgTk2z2akSx61vKiC2vO3hDMI89z6aJDXBxV61sDZXpmlJ0tUV84Rh8etMs6a+yMdJrU2MrgH2
3a9mDM1eXv2zO6o4MBaa4gWMcQqeQ/RtCIDd6lnwJ28JYRBjD6Wt3TnAW7wvGad0U1oJFLV2IZ1i
KqOna1G+/K4EepXk0HsoLFKC7J1GeaoCtL1oXQ5b0+IfhrHEXzZ6feKbgGvSQwsyHD9BYXSn14eB
hcs3svZrSNpcAtUVK0HVJvAZo9G4QPEzdBXCj4g1AYMeF/8+wjBGUCgzian3hABpA0pMmb7oWHEj
0KTqXu8a0upVjmlqpCgaUXFvKCKgVb4iFZdzBfmHZBi5qLQqk0HTvqJG2PVB3p6Om1yu+xfrtSH7
SnODPTizRJqwfJvEBAnba4RuFz6rmBYnXne+5LhN2MqoasjEEtaF5f4mDbC+RUW4r1l6EALGD8Nb
nXFB/qJ1ZbQoJpnwTIIvXQleDB+V0SxToSbvYSM+ts3Z+r/k9KbI3UkyWMHwhNB1gNHRlcigJY7o
/E7BGAfZu1SVy3NfBtGO/bjdGCWs8XtT0EAWWdodhTJ/P3Iju7dlNDdwY8wy5kpQxY/XzbkTxw+c
RGigAUJy2L7LCd0WR53WJpeKPF3z16pywovEmsfcbVGz18qFAocxSnTKiNnfEQM+kxiMlOnkBOAI
gCNqE14CNN1lmYl9V3uReoGgcZNjlyD6mlR49wsI3L5aGGXRvFGx0K3AkPmtO/5ZqRn0R71aPuGO
0Uo3ERZb0UvkwTtQCZLrvZk/ZiO+hTipYMGHAYVpHvemD14zOwjkNNarK5ccFyD6k49sCzP9SyiB
ZdOsB3/1UBej9zgHZOS+o4tuB2iuu61JMG/vqWPpnvKWMczGPkyZNp2Xk5YHSRWPeDN4TOC5WS82
q/HW+ur4lkRjgM071DLkCPIK5NR6xBvBdJMBOLyydL/VZ7/FtZYmYM1Z1RR4DO5MqPziH7XAjn2Q
8tL3cG2RHl3AIFK209fWUsykq334VbwrJMlVzzHhc2sD+AwXj2q/1OrK86y3fVx+2TZAXoouhkX1
xonyB+5fYvk/KceH1KDTpNSgT8i3jDTVx6KTLxFZzLJS+w8Y+I+CKuAXCmY0qZTrGjTcu+yq59x3
GHtcfEo89d65ABce9j7QRTt2JInaHyuYbjGaOqwH24aK0pFxqGuQtZyOy4oLyAdC5hH6KcweukOR
jeKwf/kWgX13Fm4XC5Je7liiMhyrWDnwxKPkn5hPesV6aicVRbMupy5POMvIkpzY2esp1VGinvrk
H1qOAZAEHz5zqd4s48jXza7JhLREHCNjWGFV7oUWyF0x4DehNllt+6Yhs6IU/3W7QUYhKLxrvPSE
VGnDVjSgZJ0dHjOZPZbhUTbZapyFBZQar9eXNCjUzxCP3awx67EKOl8Y5RXo57O+/IY/yq47kWEf
mS0FLUQ/HrACRwSL9g44XoeFtdrgx/pyozJaeDfAIk6gLtntx80o/XMoI/CYVMIgCIvZ/bJH6mCH
GbdCljk3LD7CuyNXIgE7hnQ8DmGpXjp7fQc+Rhr7kDtwTtXBUXzadmubhQjTXWv/+RnWl8v/vhwM
2/Kada5wJncGUkxi600XcAALLWDhLm9pEMXKGgNpeq7oqQmIgjsaHya+pfS/ZMirvFDZ5YUIgGEN
OQBtJ68ajTDfDC36ZCTTq/62GAiOGFjK1C/8Qf1KdY/9HJRvUm613SgTO8AXJIv6yn70TD2j1u2v
Cy/cdf1U74SIJDo0brxo7uLUvLNG8jxIo5fqJ1SX/AxEYQ5bt71B7cFsV/J7U6Hpo+6nIqq8GiGF
6mZSMrTROkZ/7+xnofzvIwzzebdQEWLB0P80A0B3sOQlt0VIAGRMDNPDnJd/Cfu6DuQffLGoKZ6v
wx2IExTYuESzKSQTxmN93rLRLAL9+MktF7DkzLyVIpWsjU5Lx8dT6d98awGBYAHVFs/HrJ/HSvJ5
VCSwVBIPcs8ZEWgrOVa41O1l8nbFV+OAcsDlZUhgWPnAlHJb+Jwo9n/htQKX0wQZZ+rqZTY0j0Jd
+W4ceBea7qzfgZk9ApehefDDMJ6nGGt3IDSnDsXsTmXKqh0VW9/1rKFI1gR2QRItsXc8F0dq/MNT
PfTMmrEYIF0ZFYkZ/MZkCNO6QBHg/4iI98NeNwT5Z0/xvVf1KtEJvx/CV6Fh3BoSWj39RLcc1ELh
MC3Rwf8CwsNF7mz0PfRiQGKI6Q8sDo+F/i0NNYplviZ0NfFCIyhp9Yf2kBBJEWoSdZWcO6SKhw1C
31i4cM/4Pbye1WC5hghY8ZjFadPJXzgFwT557yrMdhu2f03D5zlLNR9qtZxa3jrJ+eB7QZv5qSmE
PXpDt8tEOvfJIqnp9MlCQ916Vx+J0BwJuCKB7bMPnAneofDXRPahZ7+rtzhykfRVgfNOOnmw9t7O
qYCd+1oQSnnJ6plTxePybaAaXCdQ3Z1TrykdVsfnlB1+DUVbDchLPsZFjyKtdvFmOAcop5E1tTIr
HKB2Cw5Cavnv717V6X/4FuSoin1UIA6SUAO6Zf5Zkbkji81WIx53g+i7Nac/miN3UqRH7Uw/k86I
98PyCSKtF5nhsMWMkcimyx0S5G3J9WExS1GALI6/FQz+wS8IxOrWS5hcM/dtJNpHPEAHkPsPnWLw
xpGEsOY+BacQfSvYq3Q7UfNk8WODgC6BDqH5soUCvZhnZ563gcPM4Z/op5L/b27ZAmYtX7SBKyy2
aRhGvFoSBoKCAZLpbg7dJBfcCkEIaOcwulnwm2j0vJ01i9Qeno/fuMKefEiIrClX1YcERUVgspRo
44ACpWeBZoZU7YcZOGtLpfrIWP9qRVeYhAtHzBTUaWbnKu+xMHO/K9n0ZZEe2uTHgL/ahezZh0ga
eZpTeNRQeQ73YkDESA9atDG6FNDyWT7Cb4ZkFjxYPvnyL0LfGGlyloKUUoW8X/oxkxWE1rFFolg2
qAmKjbJkBeFv7DuvvuINqq9FxgPT914tvca8XdRPNgoLg4RH7a2yeJdNR2Pm6ROu+yTrJUrF+fNK
9Yb/+jc0hja4I1rxCU30I0yogy4kA+q2p5cE2qJY2fTHnD9D9PHJygrA6UbJGC+8JVUv3q1ExdQn
WbNYC0nEp0wabMoxUrlJCHg1BZ1FllIV2DExoKuTbn1PxcielUdTd3Dsb+jhJ06NGKauEnr5bOAd
0koxU3il92hbVmUi3EpJyXa39vRzlEVlvqeqkZti1Q5a/deKdomovEB2a2liop2UTbkHrobBBB89
8DZjHY9MTqcj5f8KvIewj+e+InCuJ+s7sp0vqvnwRwSK7iVPZ9pdKHRpHRv2KnFPqqQTS9bPyCMv
Em7g1lTeiJ8bsz2iwBn6B4rl9BYbPzq+qTEKI3hClXyMDqG4JJC+iqrBkAu5ujPa8qRQ0Jc4Rfj7
jmpiPalFJ95lGPXe0DoqniFa9IYMdNjnAQ2jnTWIsOR3gAPAzZW9wrq9nGD/hZMAxEbaqgvWUYC2
MAH4Tod31lIB020qQTXwRn+MxRL+gxqa/9qZMHEog4OqUHH7evFEvvPMmN+vFms6fgki34CgxSIo
ub44M6Gf/qPYcoQ8xfNWqgbkVR7Z74RSTFhOIJ7aPqkfMHkjRVsiNr1qDUJVVc8P5235GfGJuhgf
5VfSmqUNnFUJXo+ecWZ4fhYta1f2/VfcDm/DZxsH2KNGml3NfctDNQzkg6BNWJq1wBVwMOQMb9l5
IOVxgTvVjEHFRziFCoJA1Mp1V6snl+IcgypYZJs3NPtNzk9L5KQ74nyrUaGUGAy8+lja/3gQ83iv
Vg60Z6snv0EMONQxtpohqrheR2VphEtDZbVYqkYzuqE+UKyQv0q0Ip7R0v/MXg6w+V83GyqzLSqA
ngiNFNt4qQnfebRMOH83bGdMjGg9A2U/lk+PC6TCyVT2qr2vEDZfHVoiTgRL2evFOMII/nUGQiTL
3h2sbRl72/PNpqYPHbIXbSc/SJz8agxIc/NME0+Pkdoe19YRWlG8pIMviLcT6MO9nwAVN8j5yJhl
NeIrhFZvYZekWU7g7J+LUA==
`pragma protect end_protected
