// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
fKkOosjY6UW3zyFgzaSzTtJPU0+YzNIr2yHst2dW/Hj0/rtNPHbQEpqkWQB5ExVnk0Hcchhh2X9T
3eaPU9/svLObgRYQ1IayH61K2KX2Aec+ICVgZqFeaGPqv0YKXJTF/1IC0b3PZE2mGwcfUjlmnVvB
pHOLuU1+SM93hhu7MFQaDrNwpUifEkhzfnDiLKJTfMl+RjOaxYI/1YIZz9y8lxcr3CNGP9YGYh4j
8YyTpCT/NU4jqkmoxGHNpMSGgOnE+SB+By5Ivu6XkxnS8JgDeIuW3lKyB7j4+kTPu/6IPV/x+kUI
kwejsqxUF9LHytz4ZnjfhSyZGhCwjYmXquQrBg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
jmdHPrY48lzGl/Ze9h4PsfHH3IfBdhUUeBws/cVroXTitYgJ2A5VKnlEnaj0HV90hhTQWBRFLMXj
tNLdLu4Dxwyy37eGhTT3106NWNxSVLZxnwQXPdFDMjomroH1S0hVa6Y639OyaeJ4l3r4CTmXoQKx
b/3NQqyhmMp0WVyVLA1xXu232yUX+ha+sH81fbFV7jA6Hic9/0BOeA5XvurbmrqBodgdAPWpU6Ta
KRWJTsEWd4MF0KOlQ6WEOk1IshPTUHOFyhp+urL9ICibggn0iN29vW0xF6hRt6N7GMzcz4AvVhJy
LtIvcA+LCLe5fRk3NWDyWKLNHe5/xEiFBQwi+oDbYYxxiptRBJiNlQFe124MTfdDAMWjU6XPl04c
EsW+3w6ysXJjgo0Nmhqpaj+vZrk+DQEhNibPfipgFvsU8gPQ0zOTELhLBH68rnDTVyZMKwV72hSr
LDuWsrakG1kVp/ZRiSqKixjaFsIICwyVX3RT1XZvhzyk8U+DAmaYgCO76RsMnIkzxfb1AjnpjrmL
FLMVwLaYtGL7nImJ8/T6vWZhpzbjBO651jB8rHSaW09PdhyQO3STWVcLTBO6gsKEU9r44SByrgL4
fbJF4d4dUP3YshbhAc/+P7rcx/QZJ5WVuQToT0mxslDFwZ9ONswSBce9Wr8HAaQnBdL/gX+/7FoU
WgqcO2aHerFsDV7asuVxDGO6bzcX1CVgRr/5y5qlmovTm/5eL5p6EJoVFnzCvxBDnqBUuNhZbBhv
xa//tSRQcLr5s1Js4PmwmOolh902DziAzdgIGCNnYsgJwM26sXK/TUKB+Fjrii3tFVBjpDaA4Xv6
r2rBLhZ8Q/W1XclY49YfcuTRqehVCXMWQbLQDHe9BhKNb7CF4coviojf1247vpPfrSHvE4MVuez7
AQ2mTDNaEAxw8ug+veKQ/HObmn1Wab2qZkM4X3kHXtDzQAYGCAVWVhFBOjK6aauFb6JSgHk38qud
0xIHgo1NK3aohszAWYs9zfEJVhirVABZCTVpAG+XI2DOma9ADTZpK5YF/PdrbtcgKmKvRG2fUa0P
MSJPr4RWuPPSvdNOlM3jMeCZXBvANZTQXUCpJl1VT77094JcbC7Ix37mJ+qFk28kiw4u95Ofk1+v
1eXaUX31elbQpe4Ydh2IRDi31ucss0rgtYC68OxFUzEz8Lp88ejRApd9MiXOnsonTMNj0qcsI4V0
Gy5Ifc6PKidgNhFNt9cnNdEDmcVtcK6bLCmsDwzUN0BeN1c7SLYKMuY5KGQbTOJBsUum/eVWqzDI
1TeerGa5p8nAey/7IhLBtdiNVZFH1ofHXhCzhQEfZRexseJD9DfA4i9Uw3bU6AMsf4TnEoAqXNja
c4xcL695tvEM7uEBSg589c5XfMjLXQtWPBIoKsqT+1tCV5i8wUg0pi+eiytHIxRPp/6C3FbKd1xd
AL0TV/HRV6FaB5KHeIjm3H5SWT8wzhRWPbThgtZr2PPeO9CfcBgNMc6Myw6fzdRldLH8UWXrwG9L
m4kaZy3Luszn6orC+7U3RZnjW5h4vt8UZySAzI8qVFWhCuXWuCg5k8Dc9cowKF4V3bUyGqy+VD0+
Y/YEG6+yMZMQJV9B7gSV4qGB88DJvKKvGcDvPQfRconXb4jJDv/ue6XaCw7WgiBDZmsM5i9glAYf
0Uzv1x2EpFiv9AhjjufDjsrW6g+2TVCyTC0DCqQ6O/2By0rJxSpXiHU4aSgxDHV28FwsLwIMlbva
4oZAzCVCc9XbWcIrcPKXn4ptZdgx5kjj3EB542YtataMijsN3WQhnQiVI7TqOAZqt6BrUzDHUZxP
hl7cYNEmMXBpTMcjZOQNSmxBUimtkNHfXJpheOxGyaTYcCNgnd1TLeiN+3CJK73+hC7dHR5EI1wz
YF2fv29F4ax8qJ2LX7G+J7EknYR0efa8OnbcCInggIAWdH86n8KxFwkh412+o2QRvyl9CDWZbqs2
aEpEglDJ+jSiVDut2ehzulCdU3qBcIXpZqRqSl44/+XxMeOliM59sTf6rRk9SSoCvuuKt7NQ7/t0
F5PkfgqCVZE6C8PkSKIDPMBjaMymaqRqHuAp6JrGZwj3Lbx/0eyPrRjMEkrKLXp5zvCn2Jac2f6k
Y0q3ualRIlROyicl0IY/vC8cT5pPli+lmfHFnJmhwBR4/G2j5vFfMTvSIO4qKZcbi0+xy7Uc1T6h
YIM4XOCIxl6/XHn1sFyDOrZYp/fNJEZNNqk5NeoC/kzzixSHdFKsrBy6SnaLAawOasN/QFec8UjH
mlPDOXYf7Fp7w5bhp3CQjukafiBH84PZLeWE1qgdCw7zmGbvuKqSGROsHnO35zP4M7pUe0juUz0m
1Dtg+rvlMZFzQFg6HJqCaiscAdhIi4u/bjuo+oj7PiC0snb8UzSmOzmnOILiwIB1xBuPbDUdsRTD
5EJWKkWhv20nmrW48bOnN8lKq4itybSZaYrJRCi8C+3fhcW4Pr3hCe1OPWX/outsu9vH6tdtd/PW
Oxegtnin8ceixmq+5j1d/AcN/jsxzDTBrJLhedURsqLlhbTS6WInmPWi5BWF1Sa5/oZ/uqQ9T+Ho
+kJmuyfHmXxNHiP/tvvJRECSsl8xeb6G62lL0itqSjDFkjMGWecB9AibmMqVGwcTn19aiquMRwxw
LC1572GZNgLO3JdN/kW4Kma/5UUdJTREpl1jiRcmneicokUQmRWFS0uNhpNTxo3iFqdZLAeHH9rD
FdVqTL36R1R13AhZXlG5CkOqkSr5xwTf6eBATfGSkInGRRvvZwuChVDR76HIwyAzjfttUJ+56DxO
7+itW8a6zO6RdNRqbNJRIHfpaR1iwsO405oGnXCuS4o0jpJOaJQR4qR9EMmdn5Xw4+bFv2w+zWit
9jgJGM4x6NxQLOeGjdoMyXixLVKXCekqJpBB3ZK8WEIiwED5HamTJKmuUNKk9zsdOL4gs7Mbcq+1
LfwDmB+kPU/Qt/7EXyKxIgXayNwELn+6ae2e0d5dTzHCUJQo56wP9XT/cTZS9tX5VKKZtGlinheV
EBaWon/8Tuvdhe0rIL4sBmsl/CcNilz3gSwpttLoDK4coMRr504w8i/dL3Qcn1vVuNF7ZHNm/py3
BiCNeM5QgWBFPsoqG3dY12e4TKlqx3DHu/uZpkbq1k0f3qTMsYsMMSBw8JAtACSJ5t/NNT4TLlT+
9iqOqfoKV2raDaMflE3uuv161l4ALi5StdyT3r6VZ47rm/CDEBtuEEmIJrhx9uGKGGvVTQOqXSE4
nyaYNx2ItxC7x/E6ZXGgeosZ5rXMV1Bt5f7IIsOICbPZU9dyjAXTspoN+eF1xYLZKZXUXxtU06AP
xDN0uOWFFOkqB5vfrDUzFpOF3F8aIWqlxOCWhuDtV5S8j/kxwz3qj6GmSI/vPsasb1tqTO5fZtsx
s1cOomhHhTwBAhGBx6noiL1dQXOPIIpyZphaQYoDgjs0qFS+2Ow9yuJu30PLf9jE5OUHOihd2065
nXsi6nJPDhFXUnuI4737sCCoNUxWNINv4c1W9pDdVKO3+eFmbWeoCaRwWRbvjziUXKmBZv0MZLwB
rUIVxkqCOBl++TUyaeiFM0f1MeieKNXwNzWzLY60GraevZTD9miTQ85RVymGyyj84GVPvM1AFvn/
ecb8VJyAVBkL1MfT0mCIbAanIeu1cZYOtBd0zNgf3BBVvv0m7eHtOz3VHR3shLpUfBR4dnDanA8g
d6V1XdonsKKM19JrMGjDPkTZNz769i60BehT5jzLiHqnJgztsfIOcKHfd1ARxbgf8zAqvM8E0owZ
4AL95u0KpLkaPLnxyjc+jcM6keyjapsDqyH0e+P1KjzmlcolANLpPlcYRydGXAW9qUVfVg/npkAU
Xq6D68hRpeI8YeYnMoqMQbLUxHJq0q4mlGEmdWC0l8v/3mA7O53IIN0iyicOLwsolwCHWF9wHG7l
gUrxiKG6boJgneOh4+Vr7hCXfCwiHljUbQUrh5IaAS1e8Zf2YTkVAVzVcg3oSGJ/Vdk6diPRCh8d
ORHuxRe3blwuFW0sfHmB3HHrJ/e4ayknp0XlWH5Y7qbhYGhl+BSm4I4GxfYAeuCCda6eCMzGm4wc
a/jLvEyZMyUqRCmpm9ICSL5deSz1vKTTbjKL4obHWog1cUkG4H0kgAfnnJSwXxzaCHSzlo7X98mf
APHuehZqIdiWB3fN2EBEPTu/YQA2X+4v9h6RnUACVb2D2z8i20ZAhZS0M2J3D6s4GPAmSnYcujSj
TYG9Ia5h6pqV6Uk9oJCLXUFWdrqntkiQOhadsrDXh+7gjzLbnaWJNRWbLRevHoc8B8OKFVTTr0Ei
gaVx8rFX8JfY3MA/OHIcHNbR+V0QzH+DNYZ31S8StUZwbvKgDn3qh2G61/79bVtdMDYGP9tkhFCm
eHsDfjrm3RluXyNN39H8D6XC/DoB593j4UZTehWEJtOfAEXxKIoLIeFDYVF/wVeuwRjKtFmffZWC
exjsm5YjKUBPTb4RJ8hS5XrP00SVwC/Mk4hpRnLZmcDAquijwHREXOtX3SmMUjqPVNse8WwERX9k
RwZhitAdmR5BevFazObuF2TDf+b6xMw8O/4r0hweHeGzTrLlcebeEfjcY/4QWH2v334bZesMFlsp
fwDuQQ1PqLU+65zPd8ROcHlgc8K5T5MF5D7l0C+uij9ZgFseii3jPJODTSq6mmTHGnrijw6iSQ3c
ygY7HXJu7WODDo6DZGgNHUUcVBZQj98Xe/HCK83JBWeA5oNR0S/iBMKDj+WshPvmV1TnMMb/6irI
P2G0klbjoI6az2cvYQKTg/bXhq+8Zu9V3fmgknZSFmIdtWzaqDP6XVlTEXTxoxRpqVqraysCNALU
AyIMxal4iAYit3KRn5ff+4qYxyEtkHWe8usoIRb7MDC2aBDCCzFjWmiLl0hX9hGfHnWolYTiE2W5
umX9Uj09s3leiLH4h6YPpkYJq3SGeqP8uxTMItJMb9JFQw/xyf66eIhVRTqTO0p/yWN9sv3P8jj/
pCrNy+3ivILFplarW9j3goIEoatJwqYia5jhk7hC/EUYuWQ+dSFVxBXx+yRjPwJM6KWpbPxlIWrI
mXwBHqXeEfVEDcjOf+qqD7viDAiiU2OvNgsP7q6IQGsQVLERlT7hWDmfphnzmSCHpCbV4TR0KqCP
fPG+VKEH/mzYxPQ4MU9BFjn/E+Gzvs1ad+RJez0HY7rlXVzBCV36tmcxoKGogneIopPTS8JBC0+C
QC7Jq0DmRfxfVWIKEdoL6Jhqd38AfL/TWl+/THCAEtI2mTJTNcPExXW/ZPDJogDJDmv7FkZqCNjy
ci/q7Ggs+slZeYM8y3e+4vvgsAZJqTwoO3p04kGuNTF/aEds44O7/bJY4EMkO6lRkGBskq+JDV8t
BlXB/ShLoo4POIXYiRsVMKW0AHB7VPcDc2FvraAueo00AvcoaxmQo4WCkLZqQcNpWl9eB1SGmGrj
hnFx6RX66Q7+cqLmeW+xeaSyZ9unKubVRx2fFFanBrnQK5ykyxIT2U30w8wHcG4C5ze6Nawb0rQ+
cNE5HLVg0ByoyqJsYnaMEqPmHJSv/k1MYygbXBE3dFydHjqKRQVNDCmZ8OHe5qoD7XlNIzWdk0TG
i3biI6Ta9edG5x1gD8B/qQ2n0xMRvSrvQjtV7a58iJp5njpjeWvTZg1jXQgUSVGBf9DMIhYg1+ow
EpCLhGSg/IGkypXDI9uxuy2WvA0a8RA5Gd19TT3brRcTsuMFTdZKTkmTvHnoiXdSkCecGS8Jsf4x
LxO6SlpVgj5RMO8JkO1ACWgcqtkrRQsjs5nwNsNKy5FxWoNXu1DRHQhJEWoAb9AJNd5tqnDog9cW
tK1M1UnYrFe0WicuYWZOyB05uDlXzwVVEZzfm045iCqs5g5njUZ+w7WtHf9jWTHse+nB5JN+p8DF
M5KaYlYbeMMXW//wcDkD+KzPDdkWZdHfuARTrIiYJgyz/YFdoT91UT0uRh0lDIWG8AeMQTbivJLD
PP4Hh1Rdr4iORdgzOa4DduuCIuATlyrkYvaeMPPxnwLxCmYzNvpn99DB9MyxUCTiafrTWDHBiD1u
xmGTZTKCUKjsoKDMBmqq8IU2JsLWU57UAEg9WB8eVD4QvFsFTVu6INe6/9PV2ehPKcQzO+leX9DH
LmXPo3mOyML2eIdQ58OMe43FPo9wejdxuc4zp4YrlD3ICi7nE2c0KwHbWfiafJGIAWPpjhpuojL1
158e9X4ocu6v7rwDq7E/kl88aPr0w6rItA0UvKoQ/xb61c6xFtwQ3dTyU+ERWMOGCrzq9j7gnVUs
PFY6OG5AWslNR3fEtNBTkQLjE3+AyoE7R8f3rUWDWB3Y8JOpJDTWniFES7mNW+3bzJ9MT0la1xmz
1jrU2WwwP2DvdNPftK3m85s7ciym+3XnCIx1OBj361VwNW/BfOJ0aFnLqnIdA4GAfVdLtSFfsJKQ
ydZ/Dwp/jCJTq2vsKXVHMfMCid2mdzI2ih3Ofsysu0BEDTWRRH08U/tA8Gj1qnEw1rXEI2V1EI+r
ewHqtPRxzA4yyTtyvDAgEVm0Qpic2f2mAxpfIMt0YNleE7oV7Tg+b8rI9YMdqLFkEhCG4EhiOcn6
WYZiopeJyUsaw7eSYgbHuLz8P77PLSkw2Ei0iruRSbnvBfjYh4Hb5t6NyY26bE7XEvpv7710ri1K
n79Vax+jZppbVqc1vkzdLOrDpZq3fzEck+Bdkn+7qGQ1+ha5p2sfvEme9SCwMVZOBRai0qtCou1M
z4PfDcspJ0NZQOiGGiIPNuPgkiWTVstXPAizV2fpsaFwEiINjNQcqtm5vhhORYq5p3dvS5FglTte
yFHiqjWSACrvxe/lIUzDKscbYW+xAuXIZSi2ExsCZWhH2La/Su0sB+pDg7c9NQKsfjiaLEVNrbsw
IB9ll+aa+UYW6faI0N8eJa6TDHf6992XG4bZyyGDdoYP5PNtCpEaae+p+rK4BToomvvxbd0Ww98r
t3tBsXgCH5gZ6El7LzAtfGZ07exNOOva9OahK4Q31jl3ngIs4OsaU9GCfPCLIjLI9P+jt6PZlW9f
ntdBu+da1eaZOCVApAfzPteHXkhCqYJAYScA1ShtXtkHfbtVpKppVlo+gktW6/1XNBegHUkDGsid
CDtNcPAERUoPQhTbspbvPM2N9VpJxJjSHLWH1o+120k9Py3ALydUCZC5/59G87lFG+t4nnT322wy
2mL+UGqesFh10iPqYEjgxACEyJnqRxJ+ZzA9AyhB/iSDrRUhAyjnIAFlFBQ7aSUJtc0Q1sBvXr3v
mOkRNSgIlUcw201vCp29iO5HL/jiS0rrbB4jBin0ugmqfD/OZh+WJlIsXiMT4iwep2xQAWY4ODsm
eCbffqh1h2POoKdiWP0hjs+0A4ojY6jgg/KOmKS4Y5apPmtzwdULoPvYgS5RKKo1H2EX4RE6IFpq
K6C33N2cVb+A4JG9EWxCJ866Rjdxp6G4swoNdqgrmhxV+7MJImHynSZgjtuUVwnIpQIuAXpnbSdO
t8VZQh9XWSOWEr2GRLrB5DBfD71B2Fe6JfAL2HdXS9/icgDFQc91B8SaoHcoqvXS8sWuuy40BDwZ
vdCImzv8ZeYYZjxHy6+TXdoul7k0gJZyWjY5rEYF1Gg/FIRGcx/I1wBnDCqfvdqfEYaljStSD02F
dWv1dbJFIiUVcL4drxzdHSr8mQQ7hdHBiX7RaQR/X3BrvYEReoQkTrbhbTQk+NQlYPuepOmPshl/
ovuUFYPKww7+GD6y/cj5q9lZo0NMlbGu1iX0xqALoHbGip0UyozpCpFAzgMnKKzm4BFghUdSFZLP
mtn33twXuWPa9nAzYDle++lAjE/8BWg68o3D7FdkSA4cMfzV7p4QD3QBmCZ3kyw5zMfscvapgCit
+l9GW+skua2cbtgbQqE18/NiOtApeyKSZqlxI/mEyu7wyIvwoj7Si+PCYQfoT8XE+9p0yvXHOefo
VZME+8SPRJ3IzUfMur8/ZUoVoVHdwRS0uOf+s/IGLT2YWZQjUWcN7ItCvWT9AV6Fn9bYkhb7H6Mp
ttBN44yxqCtPxWDzZHGcHQOGZMe6NHZoopfRsCYD7ZqUqWKBqIUEXk2xYt2vEXb3aa6rcCYsHg/u
Nk8yat8/fzJfmvoH7xZM+AlAtm2iyGbyykGGgzeVk/CrJVm49PYJKJJ2p4P4VqB1SOhTGej/b4K5
tKmuj8orrsKIa0T8Tf/sd4pi+eGf8NqigtLpfGitkVckm2tdJam3NTXAH3b5Cow7u3biDba0BuQy
3JzmDbsMTDvicI3jsK/yGy05l9QqUdCfWQXEx8e9mu+GucvhbIpDRJyQyl/+IBA4fjt5YwMHofda
ZB1MSXH5rI4BEsQpApZ7EfYOn22c/RG9HNZW80qBua109LJeppziMVxhi2umjJQHAkrCYk6YlgJq
Ox2UZ9yZ/8SkwGhN8qGnr2kJcOvN+N72/jsC9Ep3aDKeKS/l3/s7BnmKieUVV4TY/D4iEgca1pm+
hnTWeULI+wgPUMT213nfL4hCDDd1coj3psRLbC2Ar1/zCdZbUZDYi5BJIYqwtsMo1t4VOSO+GH14
Nf9uX7FfaknF9YZSGq1FJw26WdpKXfTyKBp08jsdhoTuZE2QhYiu2NyIgDZyYA7XHF+v29j54+Lx
tWX2R92+u4dH67mPqtF5Fclm2ECMwBbt2Z0pq8BFRrcJwd5u51/uRBdnVcUZtcneftu2zzjE2k9g
ONsdrYmWW9Q9+VSQLeQR5h8s8ONuUSCT99UE1whdEvlDiaBABf/6feV0XxLsQdYv0Un3pf/8GaRD
CGkzKbeQiQdeIRreqBX6vQS0hL0nr2IKfatsMSd7WWOlUM9bsQ/JjHFpWS48cUwhiWoei6001XCX
ZjZyXqrMj7u1Q3TRUGhQ8dMZ1nfIN09QWTI5uBajxZWJVWU3ljxRwOAycEYPnPPLrz53meqygUoW
CvYIjmfYJ81IlM2R5NTpMS+DOq11K52rC9Do2N0q7nxGmtPYLltM+m0Ut+1ccoRa610FZl1sV/px
JiILRZhk2Cr4dYrkI41YZxcMIfg8kcefUirid96oSpZxgxMyHQ5ItEZZSMbOmKMj4cIwRBsPyS3i
wU5wUTAL5E4+KFpmDnxrSBqGUxuxD8vTOUk2jcHQ4TCrI38powZGQvDkmjrZnehNkCxrxSfm5BF6
BL6joZ8tCv4Xuxk8laRCtA4mQiTCvZs9zO1SBXpvGwfqFu1I72VbSNAuvXPR0kkec8E/mAHxrUn8
YWYhLUYlt8FwUWkFMIgoDgmENzLFOlUuyVmxP7pQqHX0H10nUL8bPRJLYp69VKeCRXJQwHncFkOc
uRsE2QAMp0ze8ChLhrBPTLuEQhkLCyDMnBG73SCMNSq1Aymala41+yyudGgo5TRi+z9eXihnXhiD
a5Yd2VBRNJSx5Ed9xZnUtGXdU9AF+/MdX0XW3p33NjIJ6gV88IMOX2P6RTeAsYneCklAWRRboMCz
cWE/CfYEo2PQnuFJMbfSTYIQOlBmi+cG/0/E1iRXgnyJOg+17QdjBg2e8yKWDO8a91b1NcPLut30
aQcczk3T0I0P5gLbYYvn/8C9C/QqooL3yN2RjHU0KihOBNva7BLXZAqpm7kVIyqEZSQ4RPP8vKwP
u4m3sCg1fNrzM6fJpfTEuCycD5awG/Xh/DMYVPdzr51/l0Tj903vkaPSYpCfnhTK4o99nmfWe1g4
iOnnRIfrPyC+tZbLwMHFXZ9GkcWFvUAz8UtRwUIOF44hg5CskzlLK5ky7Rnj7S7NCXHIxB4/AeOD
e0dY6wJzdUpQ3VB5deq3789TXS5xi3z6wEwN+0pTe1juZwL5uyEMYvuSG65cWf4N+4cBjKl7np2d
R29BCGHan+FMvpAIUpaUU3tyl39vJqVWX9qqalwWXW2nexBtR2QG+0m5QlZTMv+QfSNl06R01UNH
PiqFh3lLJmEB8WKMLJnMz0/234U34JkPBObWVwG3fYVv5OkvIJBmOPULT39C/s4r5+ccoeo1lE2p
JStPNlHFl/GCR2Otu5TyIBEE45zT1Cc3a/xix88YdBnOuCH6/Fmlq9PtdU9p86XDfjfvXwDMMwYw
Y2QJwYGm46sX91Ns3Ez+mH8co9qAako1HGDWRW7VY4x7jT+J5+fPBkVxfEo0lNvHwuw6fAnPe6Jx
FQCp9H+hX4ejBJhOaByBaAKAAJYGnehUw7y3yCLWWVip5NJdW6sbj54RlybqF5da3JJmFmoRmlZA
eFW+nSp1EnJ4xc1z6w9sqAzzchB0AZrZRraz21yBZaNxo8yfiUJnhF/dnqmn8Wv2QvO8QvjbR+pj
hwakcGHT0iBWE1VKrRhfbU6IGFn9L28R3ECQMHVOWNoglBZ/wZAi075jqWIJFZLyEDdEDkKPL0uw
C+Oge1zTXHIP5355IFuDwhonlWtbayZHNtDcytWhwZ8TmgC1wHyAzRFUbTn4cudjwvvXBNRBncBV
jSkMPsZWju1Jr9da/7LtD9N4QpyJSIT6N4XfplU3dZd/0DqnyOyEg64KSI3CBVO1r0Im0ZHnJLUl
GW2FLwkVUAZkWPCbfj5sZtAzpQGmu+5yxCPOqnZyRvR3dYbg4paY1Hoctfbk5vFd1zeVH4JPnkSB
Gu1gcS7cDCjFkVIuFjIMEvDRJ1OvAg53CSi1ekGVMnDA4pcmI4vCNBMvJbYQY4GVtTDUrlAijEFI
Jh+mK9nEVGlpIbYUGFhPtSot3lzZK6AFMrZJ7QCVg71wTRsyF9BGFuzbsAo+u9G/Ue0Pk4aPNVHd
TlVDUrEP/lXwr7HTvgSZw7NrmRGipmscreRDsDBvDedcKIfI5DMatfztmmPyNAJx1bHxibj2l0rw
kYGDl+1CrkjPyZRedcrZ12vM7NwveTFCdDp/ffusjkI4cV+YYsRhXgf20y3bC9UyqxfuwxWVNY9M
sIlNs0DRtpb12u51kR3JdanhU/5uYiR/GIb/7GWwoNEw/LLcMvRV5E7bdeTjoF2IHWQC4iAXmndW
bJpzECqhPMGVHnaX23bDlDbkUGGb2BtgZ1hqL2u0aJFuSo+xdOVjtpZOUYJ9DqzUSaupC7K06E1e
t8acupNtskRqNoZ0TOjop5A/Jbo/8OMctnF/hYNKbqGg2VrYl7zvwNbpff2HrNxeqCMXMBmkCxb6
9au80OE789xjPz0aEbGeNUh9y1tvkc+EworZG+3KJ5fX+kG0p2vuFWrCtaJ9YZge9fpTMPnxfB4+
nx2EOddWysJqm0iUDN6nAW8OZ7Tfk6L8TimIwXht1Fwb4RvFIpFy+9p8hYhatG6PuDN4FE5mCRvo
oQ/M6sgH5w6fK78C0uhgvIsfVarDwaM/ef6wNxe47FrC6NelASof4uf+AXDh+f1dyFZIFJIQZooL
j32lfUUquVIHn/JkTEDjKLMGifAgJ+9kin2aD8FTdHnbdHT9pdmh2RTqygi7xzQcYf9qcp09o7mz
U+Oy4FxXQ2NtSWsmzqe3lH54cGK4628SveVSlBkr/5e6+7VOh/RJTYpI2sRAnYqiChbBVHuUj30n
o5wFpUTHvmH7PBbzXtLaf14sbQdcgYuv4wOPkjIgTS19KEt7GWWeK5wgLSb5wQbe/FMU1vr+STGf
SQnndfIiRadzBNV0pi5mHAMlDzSjkMxovtSIoygaDMFjybMdwHPDYrYWk2CQGbF9s+qlhVfVuKdO
8sLxtwbLbpnZC0NZSVyBtFRaNDWEsYpDZ6jZwrumCMRR6N/2pfAOYRsFheZqknfcPhjU4MwAmPck
4lnMkCybrSA/vhP6S2YXdCflGElJOS2thFbTw3Ve0ViKxyXhjb3X5kaspNTJRHmwmczD1o5oXnFT
9+r5do9wNn2Um9OErx0TIhlBWRbDJCVH5bmm7qrcAtgXo0WuKwTc2DOW4TjjcEvwc37fyXAJXkNM
1Dz5AcnRiFsyvXIVG39XN4P+ZYm/W/YRXatnqtR9mmrWLl6Q9WX3j+I9EkBUHk5FQqLrKJd/ZvIF
usE+S56EuHk/zeFFY24ZCwW1OkJX0+F0gSwsqzubU8cyMPiu2qGjIuLpZNWtYSVBJlXLSSJrCZZY
QIcCLFxDufJ8CGHw6zSgdmtiUFWAE8sZV/ywSU3Ydnatt/RuLm/lZyprMfhwkPoYjrKtpr9f5Oha
9UgTPlTcSvKlblscSc22JeG2OhVQn/VCSZ6sErXqxo7zimaclS7r/wzdeqQJ/3f18RdAHsx4f3MS
RK/I2nkokbSXgle0aLy5j5kr53aJcxsTKUU6XrM5uoDClM1gOk1mYHXOY/UjFBPTAm4CkZ6LAQJw
dXJbtb6fX95RI/mdAHqV+zufZocMqOEQ8L7IiNdfjQIknfGyIvIsYpmvPwYS66lS/HjbYVMk7SXr
62jW5mumdjWfJf4Kf/lkNhsf2kBihNIk7hJegL6ahA2M9l2/D+449igs6fpenuYvUgCSnOKq0MAa
Rta3LqfIrHn0KgIt++WZey1FiQnSUOfqvzeaNJwYj2TbeUUvf0vX23tbpYUfCyGsqCZySpzEvy/d
6iVmfxZlt5UljPCBV0lt3IkffhdYXNCERKvxet4JYvb83CuoL9ws3f7dj1mMm7nLCVrstN9OsG1e
PrZ5cVCzm6LnvalFnnH7eO0RkzH6JpS6gcKUdljpiM766VtV6SRhQXrnuboDprjXlFCQE0c/aQeg
LfWaEkjezKyNAQ0+bXgzBZlrRR39T1wOdo63Nb7ruGdX3skqjD/0L+wHDHlOQN9KZGGuhR1KDYVe
QVBHDnb2Yz5EVsyHm5Upc9W9E5n/jSS4NV+4mfOXL/nnx6E0Y20GiEWk5msmvIl+1P72yyX6cCal
66XfoJgFGKFjmatwAFMaoaSViEsCtRJVbkYdT3z34EpZOjd4EE69DgykdthXWrehDwY9KHyMR90i
iMCXJpfGMT4IdAtRvWQYg9OQmF1InlSTqaFIwGoxgykFovd90aN19vRKOk5uEiHGcZkRSmV1SEFZ
CLUTrvWX0+9StTtvJOVayXgcx6JtvjOcuxdlqX8epLjNXNi3O6iwOjJ4xVAMDhNbF7Y81ugPH/N0
4/iAo4dMDQZEfW0QJ2grMWCqKuURTHMnLrnSGpI0uutPCHy7JRXWVipqPPa7CvIhIvvsQkEqeHGd
boI+1sPsKeBzqxdWrxXO4wlbm10Z72anC4ZAFUZqeyEVGcf76BrAmzMdcyiax5Ta8klEvllYCv+4
Dejsh/M3meHtpxoBv+hZzVdIpaiLLUxRgfB0d5sTBelJfXNgmaJNMQCKiSDIXskuVkMj6XQI1Hp+
qgiW67Wgi07/cng+njHKQYGDvY4VJFxSonv57P/kxGljMk3ZYsuVPINcnEtSaE+fNSbE8otsNSXK
H3D4shMAdQjsn2sq5IX/d21MY0qbshdGs9Nm7I9Zd5doBRFAvBAdPmF3xS7l3aOtAYnpEQK5mNhD
pvG0+dTYL711o1q2zFVi0OprqtPnWjqkhfdugY52gMHoJDSRAu3MNg19vLzNdv+okAotaCkbcE66
V5zddAJLAijzN/qL/zxu2ovQov36f/zIQuEe2AlOl5NaHwgVWBuC4ES+RhQ1maghYqC3bckuNpXA
mBiO9KBrjODjNJw5QRPldqGmbaD3o+SU+S7HxHrcFTsbIUKC1YSF7JQRl80Q/0PaUoMGAOnyqxOH
gBv95dSDdakJUCh24zZnpH76IVjxZZXzR0sj4V0DTq7RkG6l13Uglyl9eCJMs3Y3sIFoHjdC4Csq
i6BrGn3V5hWaefkM3MXZIpWXJeFn9nSWG4NNybgRE0wvRVCCcdwxZzBdE8siGNLfPGiENjDuLnEz
Vkb4T5M1DQKN0ropwU4Gzpa4CCSUk3QesstERm9rVNI/mFWrbtKYgOqko+I2CB4r60F+LOD7Np/r
KeIF1I6CBG1MtpBbK4OcLw1ckSETwNd2uA8p7P4DZCJMK9a3SA2mq9Ypi/WgSd4Ow7E43eGVOo3s
LefZm7rDyz/6pOKIX1ODXzwSEuE69yOHaQJgOx5OIcjfW9Q0ZIuykUlGZW29Yq1U9dmn2Umk6WLv
T4giBT3XJa2MCKp7yUC5UpW4NKNEDxL8D8OPa+piK3VOp3JVDlcoL5wbPepYk2a1tAa1XbdFBtA3
fa7qVa1gx5zAbjaQKgjgeRQBqFJbguRUS9bJSTjL/zgaV5nKKxt1EnTTl7kOAiAEHLB9dtuvClwc
FBr/ON9dUL0SzVNDPePIZoaJVaaq8s3LUhB9Uhweo/2m7jgvIJaQwoy9nzqz6ubsYRbN0FmUOAay
CZSWx1o4Qv65pT5kk9h2WglrKBjaA+xaVCZ2YvpHkOnAr7P2sRbxrfTmKtcnFSi6YRMS0iRcWDz9
MzYl/11VmOkachswHSzefqAnyN7kLTxjKNJ+dpbVSVj23/Pkjh4MgFmSsRKvJbchhp8eotWn4+om
yA29jnZffM2eduB+3vgYQjdk3Qs3rlf+jhXv3xBjupeQjHhTQPHJvV1R1Uw2eS9ZnQYh/c7l7ZSs
u9ffs33QBy1xxnyyQq0SfJK2taUVlVXte1gspgLgMS6YP2nnmQ1otW/WU7dB8WQlHCU/STw9hzDi
hM5fxCedzE7l5HEUifRhUI3bErZSh+vKnPp+pIcDKf5FEkToA1jMwFPP9+kJeOCm11+aSpKRB7dO
o56QuSnipZ9xhc1oU1cajkNfu26Rx8SPIUplEM6LAMT8B+iH2Jxy+ILqfMFfxSKZQImz1aC3TZoA
C1/bSrZSusN4CrHE3QERshR3MUlJK3z/Fc3vf9KAKABFcyxGY8tkLPU4BRrcSWwfZjjk5pup86tp
aVp2vcna+qL1n22Gsv7YCCkV7PJgroyCLiTpYh2U38EAe5edVGu0B28nTg2GcVf9GIQMqMkoS5/3
YJC8QBykQkEKfUVfqeC9HPZt4L0b0iT4G1c+LZMFc1QVN6XqjvNGFb6/qpSz00kKBKFsr1sxi7S4
vOnCogaDgomfipYx9a9Ljr7w3G7AxYdHQ7gcW57opieMa7OMiHkH2Plik/AEcVuTCON4zWNneP3h
EDzFjLSbmbiZa64SJCp/i6cOgM7L1jNyLdXTsV8EWqP0MZJARU5CmAU0eAt7bmF0mp8UetW6KUBk
e/JTDk/sPfYZEexcoR/SYWCCLmzd4Dl0/k6amDXrOfQPOh2VJ2uKzjnZIOjeJkP7iZDozXCNBioO
VWBljXYugq6AjRGIsQwiKR96ypXKAZtucfjXApW7IW4qBzipYG+WGjO2hRNccdBLemnB83QF6aCC
9MjQIPPhfc700s0gjCUnSQX8XOvfsg3j3A5R44iW2ULaDqmxZGT5n47Aja1d2RpEmE8kGgJAVMIZ
EsBc5/AQpL1inFZOz3RsjG5t+SyK5UScUyvQgKksnVj578VhMdunPhRJjgb/vYWQgL5RZvwr744m
GmVs1X+WwzE/ZXb1G7PDowdAhzbe7gKWVMYMCV7FRZeIrbCcJS0x95TJd7w2KBwFs9YNSQSVDzEN
6RdzQEigZkfcQpwbQtIzRYjO8M2Yoxe831AQ2UGiQcAj0t4qh0nmBbBdu9WcSAo0/ztFprjRETSg
/QQGGbDDiQ4e4Jfl8gShAQPMrBF/OVPmpTrxM7wHrClgUt3yVrxUQeHUJJ8SqtXFu6PxJ47UYZqX
eT8SIKSqDLOJ2b2N0W9fm1MbmL8Ful2PpedB30Izp1k6QVSobKPy6PIrplLuOywQD9zyOTYcjwq0
79GgzAeaqYU2zQk4tvFNr91Wk0JeB2eR0X14jaP36LpyzycY6M+t8MYrhE1r6hX2GR1Qa1I0IS0P
d5bfrB/MApV9ZPxDIiqTKneJjVTrcdfYRj4wm4HS2/bHAQNlE8c/gFOYmn/pdwpRlKuISaltyro7
/rRE/YaT7PRgaNCzhSaXOYIrOCbZyjTJcpVjmrg9szS2OzLVRhRwNZ6VFYpZRckvjBdWXH29OIsA
UYZmhPuK9+98bQSn/6oAgVPn4OjhypZI73bEbRcvjxhiwOAM1yGN5fzbUDl/HAqIxrAfX8nRQzWC
odb72A2P+s/X9lkg4EIg14UHDpR8SHOJuGy1sdGkEWE7zRjMuR3urN8ufC56PqpMfrKpaX/UGpOK
f7qYFiQg+/yXMlaDM47htarDM2BiEiHtFNY09PTgY4WnwSlyZiMSv3QLISyN9eWDFkXslRb9I3Jq
73eXmQJqxF0VvtO1yF2xf2Y2gYsTyj2bTAdZlnFLm2IjmtaZeDPNVHnXRtTr/QSwj3SuTP9Etaa/
Py/NJMKLuZQ25oay/SluKm5qAiH2MXVLSsGvp3tLqNChlpCDVr/bfUC8OIemzcauaz0gn3B7Od7j
gXnohgSYStqAAo8YMXzKpYDNgZDkaF0lnEZhaEPbE/KW5SxQeteoRYZOCBPwyVW2SrpWx2h/L2IZ
FfHpCUQ2yUbOMs6DMJGi/XEmuxRuvAgJ3pSasGccZZEjlOxTupfb8UzAII7rkXJJMf8ThrFSnem/
umCzjtLDQq9xvs1MZO/t2CKi+PJKzuZg1rH5PmucGBmPREr7QdpW987T85GOpAbVKmMH4JcZzbAM
QTEftGJCFW4BNicS46n0Hz6C9poztoWKtaShGXc+VquUWLniD0ojA+eVlbjnEkkQX69a8Yv8edJY
9R03SOuRNN4knzRSlWNGiIU0LjyB7Erec2HmaUTrgazygySd3/3reRWcWNH2vOpMQOGtozcDoT7p
D0to34f5umaRqQOtCxvXy0U8ys9D7wtcCtjUMb+gMBlUvB3TDHUSEPCheOLf1M2pJIT9pCNwlr8E
I0SjlM1K2XJ8fKhJ98BXR943rVn/O3gBAnvF8ams0PIS0dp0V+XQOpKmnDSz8j5I63sV0TX88WQp
ZevwLH4Vx/iLp6JddLJm7k8LyKsE9tY9xu271RqZO6BrXesZlN4gCkqNaGGlfxKRLxa296z0+LJf
G5fj2K+6DGOyjiPhms+yRwqYsXWr6Tq+0psiMixGIU1FM0T6sy2Mxqcg9gIIYJoZVxnDojUpC9Ez
zp8sXLD45GeIsc3ruu3GWzj9NkASJbk5GAAKoCVBt8ByYIpsjodn6vVdtqNCJ0RjDOlQm0i8Ry8l
eNOCLQWazUXE9b+SNdffpECQk+JvTh1Zc1ye2vkwtJCegDYAehgGc41gX+LIKAbgjHA1Sy+aRoxy
ggZGJoDL77KCIGwGgs+tVFjjcjATTS47OPhrBEP/5u31ihcxVlHlOkQKDNqLpY9d5JWDedinPcEy
HV2GeCx2L+g1T/RJxFkb5ATsWrMbYTp8lYKW3VIEKy1Kt9QN4o5J9Ox+o97eK+P31W9sYaMdznzH
nJgimV8PrHKtTARcQIKjJpccAblT0O8YmduiNGd/6zNmkrmlX0A/T0b/9VrUPTA0WotCXCyVRjG8
np+dKQTWC8afukRF4roMHyWskRkTART3W9N8GWaOdoXrU8gLOgUu500ux4EE5X6e+0ROFrlRMIIL
Nb4WFm/ExOeQ9IiyGM+xE0tAy/VOkiCNwVfAouiUAR1SkC5FNiR9x6z8NtBFFYDvc1yCNGPw9oBd
mXP76Sh3LNLv9YzcYp2sb9pGuLqf3kYPXFj55sLk4lFQfJxFZ63pn/sXObMxABmkmsbrkw6RHhn+
ZjFZCU5paFKWZN0+ikfrsZl8189s2sDS8FeuS32mXQvB/2jAE/vepqqv0ibzl5TG1mWHeE+A+8nj
Tn6h/mZG5yFmL4/ktVjp2J7jjyBLeulyQPZvwxHzULovAM5ZCMQ77uLnMVlQYsCp5XOtxbsy+Qj5
xbA8nTYEQQjxmCykNGQialJZENKy71bLwkThvY9ldGEYKrqlG5Ml02StezEtzno3Ig87KrWFvvXE
TYxx4+OvXCEE3BmHVjfkK0fJ66Nv5Dnk2pTwdltnUq4HNa7wIWg0Ova9mVdQ41LUS3JwAAUYIMJi
hQsqs+B4l2cHQe14rS5TYtt0rD5x8HgS753uQOiy7vZ41qcz4Rja055BbD7Kepsz/ajdMPDh0uBF
TCwtHK4f+m49ehqSCqmOQnDndr6jIqsFzf/qVP3/EhYsFCQP9xgP56VhS1RbiOYkw7C2xwYZRZW7
VjD33JZlFhb2WG5iYfFhGzjLxSfrCg1Kk+1r+d4Hi4YWdPCf68bawY8iNGoHJUuXrN15IWETS++R
XjVj8qlHTYR/SE7REe8M+WF8h8gfY/HUhARBHWsOhUL8spGuFfbWJQiSFj1y05rOfj/P/9L6uY5c
nw/+9hP04NDmawrVPRMWcx6jfR3gJX8IDUT1V6IudT0NTy4X6fFqKGqG5kxeQ/PKLrDd/bpW5yIt
xn0XEzwi0tB/sjB6Rw7RlFjMqNSAkf+j7HLb7FxGfLM+tQLvAcbymYNZUm9l7p9h6JNI2Npm7js8
Yhxo6B7ZnQqqbFPLKGUiyy0FFllM4OVfWbZ/iACF4Dvjx+x8OSkeBTk8VW0rbgfMohTVaHP9jNv1
u+BueeDjDywRONCiXr6vv0KwPv5HFr4emFuTpxpqpoHZFdEV1g2Sr5hxWq7b7jWdWxkj8EgRDyWo
VcGKpA+pcdsP7ksPFSDBipI1lr4/R4a2aPvh5qCezWKpo+TrqpBlnCw1KdR2QSZWjjUxDR1/oSTq
09JImM/6cdDNPXlnXTqvMiMybflChj7MgP8mejvt7QKK5C1Ci8qgh+7xCtisni/+yD6Gp8e0gvZ2
h3u6OhNMehplUVyGQRqhCLJijthxs6VKrOEPCmwwG5A+2ZDA2YKoYMi0wXxHxIYMd1ivV2I33IBm
nF6YB5CMn0/9i3O+UUxNtwEX00639MqU+VE1imotGuzoKJMzTlbx/tnmcqKzlfpMyZS00hd4lpOp
H3/St0EEmRetEOz/mcm4ChBr2huUepP3+kx4NlJ5vN6otaacfMQyVLmYJm03mzhV4OgZQaPCF67T
wMlkmUX/T4PkQkuw656EL8p7EMnYUda/5BAaVNfpdpeHbtt0hHrZw9BdYpfLSP4pHRKsjA04+QFh
V9kzsyxk/jXsgXtlEdUfWAF5g4d/GAl7AFgrEA2zkbA2aeSueh0owgz8tXfS4w0ynrlz4rleBTKZ
c3Mw6yegeW+b5CjpEZ0FSi0LprdmAcqE/34F8cpQ+fuB5FRcCVngpvSJICgLXnAr+4GmF8W7sTaS
xZRrZnAsSEgSFF7P7K293LFmdBdW/ghDEc7IVzYfoYW2ppx1WQVVng14uZw+BYg/FA+cL5naOzQV
28N3fjDf96uvhutByVHOlQt1OvJN8XK2F/Z8Cb4UmGgvmODdUYki7d16WQdDmT70bo0Hdwsg+eGD
KK+xrX22JIEiGiFQghwojwPmWLahCqJct2BrPrKXBaAwZnjD9IflnMoxtEwlrAkFP1h6lBTnjUlk
x3cHRnaNAHunwqsaINaLM12mekOojkQob/ImWmE9CecYnvzi4tt2R+f67SgQgauKoSmisthqKQPZ
Ci67IJj1GCLXT0BMZFC4CIg3zmUnPzri1jLFEyhtLdm9uykYQhlLGqjtDa6NNXlYt+k3g8lcKlA5
VoB/LQf+lY8bi3ompk1ZV4pYBxLJJj2xqtnJYmuYHGD5fl2lczkta2oCzIJEY85N3hl/M2HAtJJ2
gSXjuKMrStO1N6RvenlMSKPqEjGqa0HG76caeBKv+Pjz5hFkj18IiZdQRSIC4iAmphNihiZUniFo
aCCtberxjZtypCmatZummElAUvSEyOpMg8IavlCpA9X138fK8o4U8h8hVZTTq0o0ja9kF+DPMYLl
cVdPs70am8amHLWrS8PoVH/epGf1m8/XlKAGtjuvoqTCdT0ozJctOwiNJ1iKsNgCEfHKZfpxe264
vgf23qqmWCXyesT/aXIVnri/c4SlAAQSasuZ+XUac9BhxJzdt+Uuwa0co3jU/uxbvu/7LHqFE6nn
KaZ2sLAyCJmnMN2EDiVpZmwT1HmUkdGHGjUrU5AfJY4/VpKhkBOx1SrPkSCyTDGsWkWSszkqPum8
aDUMbquJB8VaBKVN+5aqrp0WBLC68U/4Lw/qPUGRQJyKPFyof6xCtzHVOKvxfjBn4/Kkm6jOnuh7
NDOesLOcvXZDW3wfjYmOhXpy5TlwU2ZLE3mIR0Mpc4uTm+Z55bfagERq6V+JV0UEZQgolbIu8y16
6WiEOMQtPwAm605+MpDM8DUpm6BVZ0PM28ShdL10Gx3jRY3WT6+Bm4M2r6sghmSFqpFt6D1TJKs7
Nw9MmS1LNsqxujnjBAWACg7yszolNdBh+bOt70WWZB0bXge+pJ4pxXgcBTJy/Qa/ClHd/wcT2qxo
zjgRdszoodR4ONUmL+h4MBgrPGx2h3XsB81XrtL/xwXK+n2RG5nu3i7/vSOKggrA0aztJJwM0myt
Bqbwjbk6lTdSCY1MBCpbM3438uExY7fcikJ/APYvJGFcpEpb7dfO73b4o1IVSeH0nGy4ASZtFj1W
a16HBzFuNwV4lsxXgLLHA2xsbufTI8ZDrXIXGXntFFK5DkLRXV+VS25eFmtmo/p/oSTPqs5ro+tx
l1mFVuKHo93jqevy5pRGa5rcYMHBI66RxYnuzhJWQsr28UoDfqKYGoUjrcFtSx7063PdfpubX2ha
X3rAcZA3FTZXSHl11odXGSe06bARK3sQHW2I09CKkStB2GGBohhyImMd6vBHXkzYDzjGwA1bCrxf
wCnyXocenOpZCMd4d3SEKmpBtMIqRHZuxlaSaxTgryz84hwymsuKzap6WwBWcxtp44GyAiAmvFkY
ZdUXWiQbEq9d3d57+XMnjPP0Kw30pKTGlAlL2LRGFtx/xUWr01F2FtE7LUQzKSP70BnTBImCrqBG
Ieo2CmnuOOmcae7MoiXJYt1PTswaHEcV2kShkTNxp5vIUtYnd7owFsO3td4/VBVy2dabmEn6SYBs
ho/dOVduDITcnVuKms++o3Zh9ex8XjQBND0eXwAO/LePLGSU7W28vTKjSHA+wojTDFaTy0IbYWyf
o6lWqXMeiSTIpk4xsiBFKXD58xdSV89yCQ8H8otJp6IpBIDgUCsHglXnBLS05nqGzWMfDO5xzmhP
zCg1evrStsN7WjzBZjSU76K3LGzqJ2eDvv+It+F+1bhWiyNevILiBpOiy3VcXUeOQLZfw2C/T2+J
Ead0qS2vih0Hpnwx01P4YEKA3u2McnNzIZUU4k77MDWyS5pWA7gKEtHgZxf89nG40226G5RNGoPr
OLuPY9ZcV/a8sl1CZefhpEkpXDAMnp7oSkaOrjdxBAHxmEarvZf0Iw5jfdySmmCVbBsc9HSrlBz4
Ge9iPmw0+DLIhtES1dft2v+eUJB5hJDHBH59uKw3LyzhV+d3U9WgPrg7SiOmj4k2U80Ayx/hRE/n
0Cj7VLgQPN3wEGBLxEYiWxbqwOqJ3niYfOP08JdNvnP9BDbSEJcL0gwdJzJ0LFgm/jVH7po3I01c
EJPa2/GJ43P22jWikTI4SN1te7wrkqJH+fDkARw8Jjxm5CZxKNXNxJzElDSqgPfQQWEa9ogmeUKh
pLVjp78Hmp/vSoXyUQSdzaNkdhkhbJZgiAmeyihQiwW2bPNJewNeSzqrpvGnTJlbs21v9gHhUHW9
/87CNWdILLBfGslgqMBFrsGUuza7GhBk3ttzgtORc3CYBivtprQeCBqn59DBs+Ux0EGc4JBiBpJ9
52T5b0kYNEidgBmrQ2ykJLI4oZxiLbbGVDJ+yj1p+bziws1e4AOHRGeNPaQ08M0RZQlQ7zlGAEMn
RpHwt9z+mAV2q87TxR7U7AX8IOpRpb+CTsN3E86zkHtHBsQWcVPZNAtifoFpew9X6Tule/IWAEZ4
D4R8Ts1kU90zCLoULA7MTJcZqlZQWOlGfvMKzYjrabsFK5JX/DYMPdBVlwcXs92C7Wr0U6S66XIO
py179lddEVNW/UB+I4EIDHcAiY8KHKJrQPUMdeIXdcy4N0+36eIfGRWdWZTNl0QiuokydpRIjkko
6IvLv0pCub85ueFXo7Yjt72HWqz5trb2VL4BtyDDFpio89CHG4gnQyVVj7IlB0XgnTPlWrTlKFBY
++3Tp7flI71/BaVCVkgx7gCNn9kmA9rIoYNX60T7MI+qOGxO6LPA3XRJ1vdxjbbmTQt7UQpEtxCG
UjidKJEzmqNns+Jzxf06k1J/KENQkGF0Yc/px91/gqCENorxDndKkriq04CydC7KItIJUSx/eLnz
r5o+HUntZ+5if+hAJJkzrsyp07vfIWlG7C1v3ytKC5T5/ZIy0uEow2KUaFK6VvkYrN3em2vF64O6
QHS6MeKJupD23ZV/+mkZoo9lVi8Mcu533X1PSzMonNCgKAzE0199NFaxrNoEr7+MQPCN1lydeTVt
ip0IETUrPZowBc00ZscCET8wZYE9f+0LOiZl0ZjUngyGF1FjedsvPgISEdUamtFvmNp71Pam/0cy
NJs8AFj7S8M/LBsNP8Kw9fKdYkYjEUXDLGyzvVvQoAy/wE71wAAQMgznqX2FLV87jwJwQv+QRdwx
xcqC/CfJguSlNmZS6ehEyYc+BDMHA3xhTS033JNdvv+sLtr19TiqQOzgWpErZC2lbEvmwsbXRlQF
ytxQd+t87zGWYfIb6lIeOojf49GU1414s5g9Q1bp3XX0lNHq9Pyt/l4XE+uGpDBbiLOBS9yC3PIp
AkByuHNaT2wBamg0MjS4yfxAGdIVb5hNpB7zuHfEKUOUIsDp5OBF8ZwzDPrGRLwGe3QglgBmjcvl
lpNgxMVQcZwkhdgglUhttktRAEYaJmgBMCKWVJuFo2lvIK+Q/gATrbcobtm1ntYqbN0k1bYoOO4e
lkq4eaDB+R7WYIGXljHXi9Eu2wzgjtjAuqGGwFGvQruYkjNjAZ8CLegtZjZLbXFhlf3SKMUaqa5q
9OEJpU7gzwPPDNtUoRJ8YBQR46pZAOAoDnFMHncn7F+egqpufPVokaqiehQb2FAucK8X5rEkTrXE
se5wkZCxqHKH10BODHG3YQ8wm4BF2lM8qZ4B4gEjDmOd0MzYuRe4pLmsHYBhtthG9tMeUKZmAGrk
xbMienS+mUdrnEYoAhtyj3WbM9sbKW1x4AzPlH5GaOuyv55N9MzNN4Sypcjdbg9dMhYdhizXcvrI
nNzocWVOXrTRve4WtL0Jg+XRm9sydmRTcq5yQeZhMtlp3s8R2rrWt4zmTwcl1f+GfOdYYP3X850E
zMvNBi7M3LqewDgbK+ZP+kyJASvdTlb+H1ELfN3nkVsdUPPNHpmuwmCLT1e8Vl1hgy3y/XrnTa5f
jqN52ukzntcqCedh8/fw7VMdiyxhXI9y0X4RHnt6nG8bZl1vVOu9aLPOL+SdzixP8K6VHLaOVl5b
T+hseWEAX8xW0S2X46kVMlqGr6enLhFuuFn1X1PvTIVsTiN3m7GOeDqqoRy+UWBkT5FF/VOgOwSU
1dE430KkVFacrOUOI5WbykiRcMAfY/vSDFp487mTjj608WYSdiI2W+5zpM0rUPgEGVhyq/+vjshR
FRiD1OUq0p+d4lGwEc4hJ4vEOhy6b6j+18yaaxglyEba/OURMVxT8VEa9OHchYMIBl0FvRA2NO2s
b67bAZIzPXp89Ycnx1CJS39Ytst1HYESUqhpguPEaUPRjI8G+nD11cyOZGoGcCkGgHqwV7NjBkz4
v0vKU3V6Es1tsSVPIcTJ3dy8pZYZ06ACs7ui+ajos9KTmRBHTsxW/y1vNHmPmAPQ5aBijytBDOT/
XS09i77yTCTNXsAOryNdUDc+ZUDSxQchcRRaJgTOI8eWJGqkePYppEb6whMBXplGctix+3GqNI4R
x79EkgRYCPIneaVkF3Evcg5cEx6eE9aQBIFijAouLy5dTNjJ5/rZQpsufyxs5j1NasDfxrwXuBKY
4+JidpbQvVbYYveFUFxGq18wNuqao4VU+0mAC1npXP1ObuHpktePVpJWxOFiCw51PsW4BEqTE3Xd
ZNtib3jKOIGpVQHznTEe4x805uQBYkJ/rHg/9fRHpK5aalM70Bxyduclp84jdVo8suHBEwrkP9WL
Kn38gpmUGp57e23Co3aHCImKaazujA7gwR+at2sH0EoaP6rcTajRoOel25KYYbuJeIIXZNprMKCV
E2E66mbeC+c+stS0wbukxhD44Tv7RmF3aDmR+xicu94IFYhXXIIrvfVpngBiKjgMQDPZ0CoE/URr
3ie9HhdrLBRv8xK745eQm2WqaoLTU/hc2L2ixo0zsQqUKRqvihKq4UmPGjZ53WOVahPo3mh4ehiK
mbqJ9ZIPsQot76y06bPRz9NxWJ9Y2bZsye3eUYy36yTM+iDfbRPQh0TiNPT0gSP6Y8enEx/cW0FM
EWVvrvhMU8bhbKb9quo3/RNH9h+HaHh2opKqVVuPqDMVz9G5SiV7rWnrdV/ShjOZcxSsmzcSypl7
lMDo45xdRdUwlIomUhIPjKAyWuZBBRwwR+bxUFIg8r34PiNXMooO9+yh0HvGPu+0TnWWKhEXVi/L
IRvNhKVxeJETuy6dr8o8N6aAXxxujoGrWfTjPvoQUPDpNnr6CA8lHFTWCCRVKi/IKqbWB6s1lGtP
qv4+Y0afywKZY5xhGuVBd3Wn+nqlZVl91WnlVHIETTBAXUbiT/39itMReSDBCTS0OipUblFMqUGC
mnp4VGW6BdoELvhgTCLAtOCb6n+UfGEB/M28UjZZcN5yVAJmlDH/5Y1a0ku5SmkdFgd/FVd8HLjE
nVd82i0ysHsP7XXTyvN6QjFHkVVmmEIGDJyTBQ5Jglem1+Vd73ActN3ISYhzDyCIhQfpZVmRGiBC
dhMXhJMtkdNNZ7uENDeQHFg5XWWFssnbht7dM1ZsLX19PuO1EuQeVstCvZ/m0KeobU94HQRAIslf
tnrnM95BFta7yLk4+a4tXNmA88yEDa0iHPc/ZUZHj+Q77sAGp4HsXwgk2QSW+YnutoFzmhZXAIno
KAhnGwsVDQNDpMxcnfK4QXAysAcJeqwUGr0p8JxGoH4sAO/VAZbhuhRUla7El8AHj34MyM5qBqut
C3AYU8N1ule0uErccx8TyPUPdrweZZadk4639gxF9TYxT11+syhQP6qXtf8SrpKP6qcey5GqPsEp
jr2LY0E47czxvtZxHy/dEhR0rDynkmefNFJ6XARyYPoVu1JIdLJbbK2Vi6QlVYt5sx1YHD//d7ei
35ScPWvqBV6ZrAhml3hal084P7mvET8eeROEEKbPkThaSWCIE8KJ9Es0wE7bpAEZsVaT+xVVVd2x
fEAlAoJaP40SZzLhafJVBHzRdBjiIl16N8+kDLLJFBMnCMi+UhYKaNNUbGCzOGHhTh/YvRBApA8q
kNfdn1c9+cZdo1vwNfE2SmK329j3yicCT9sfd4/J1XnGiaVoPpMEJzCFC9DgvdEoYqcsU22sYrzk
ggcJV+Nu6D6OfDFbNMuR7QAAtTuHyBqq0cIUNdDb3bYGKeQCE0omQtN2Nq/UXt7zZn1n6sra4sWZ
Fi3pbKqNv545ECdIKTZYBEnonbQd5gJ5asICoxmgfDzXz/7HHHW6tYOha4nAZWvAr/rFTMn0nWTf
QAeZ4EJVDspXqDuquaLm33lcz8xfxdHO0odcFpYO91Ovh/Lgx6kvETuCSNNYD9vFtSWjI/RNT4S3
6Hyb0xadWLmRN+G4B0wdoDdNX76rk2YOq1Uw6lQUaVlrDgMKkljVVXCkO7D/WwD3lq04qD7m9Tbi
4qU0UYSG0ku4qqdfHFtryaKzbM9a00cJAK+b+icTRh+NI9/MY3y34YMMQgunbMKmKVVempjGjTx9
sFrm7zgvjVu67B/UHx4PA4RrFIghLPPYvYrQgfC7HMEet/op0T7yv1CWWPPJFC6GLhuXEjsUpeg3
WoNXjLYOFWeOJfWvRhC18/CofZKh5gZpJvi8iHz6trw9B3B7T7gxlu9+Bi6+1Tnfz3DWbH4Zb1i9
wz4tWbOoUt/v0yQcmPdP64VYPcekJB4rBXgTqhA5nAtPuGLdBD0TJ6jEz/sHvr3rYc3mZwhQefHX
5+nv2DgGWD8q6eB+8ucd41qjc+O4TAXIsRFAPFOOuUsVLR2zfq1Dgo/s3p6QMi0FgSM879IFTGEA
pILIJFnq1tTmrmC2k79gAVK++fGzu6+OR4FvE1Y7rWh0i1Arfs51RIQtn8N9/URPSj2VrcaDa+u1
g1MjLSSndWnBnqHtZQ2c4klLwS/CuHCOxgTf6u6hn0sb0B2UsDx9pwsvEAUflTinCMYv/YuedC4m
Cvp8o0TYXtFiHkdGrc1lMVNsR7hv2O5Ojn7nhIeS++L6v6feE/COcXVaCFkVdO04VEYD0TGFDQR7
4BCmf//vogQIKHvdhroOY53eHn9DFQF7NMW7qzk4NkjfzYLT7OuOO1omga1+JRqXmUNvz8qURb38
3kRGMk/gHO+6RrvPIzbTChF8tNT/1ia3AdU6TpTVb2OucUcKSAUgX6wYRvGPRPATJNVzX4cRZ9cs
+UR6HWcalysf2yMc2iC0c/EfWgcOBSP3gOOR/Fw29iYwzQDbVMVv7FDlZDNzyr/VU7SXgwWGYeey
sG5RF0AG7LYDRU+0lMGBPp8w5fApHHvZEko/8VP8Zi8ttC6SoTZciAX0/J2tL7N9eU/dL5zdmbyT
UhiupCjXkoR/gWtmmpjQpjlsDIh9uxasJGlULxkFsSGIqHxPyhJoWm+yuwnlLTUZcwUao4JNF+v+
pgLx0a6ooB4CYVXZMthqF3dfPA4/KiWfF5iAkvUrFYLbz9f420NY6eoY+16E3OTEV19Bsg24Dls+
hrlpsA7GNzV8wVfYOT0pTNHwhdme9PqOI8TfUIAto7Dvh/JjNnzsPwbthkDac2co0YzKNMaHVyXj
KO1cliEkgJoSe6muC+xdKiLH6f6u27izKh2spTXS3m6+XoGUULF8v1czitC2Thm1CFw6qUJWAUrN
9ILHR5b28runsPOAc+7tn5ZzI1mImmFhvYIVuVJC+s6UimMdkKOND0XTo0ArZ8NFRs5FOXrQ5x9G
bhGBCpvXnd1uhYlauEfD1dabaH54XjvwLj+Ar3OwA1a5jjkEa2pfpLUE3rOqYnNikXMQ4lre8eLc
3NvuhyHoBM3NQPXr0otksXEv9ooqikNa6TIpPDqFB2eP3OY92lYnZfgyE1jNmlmIRGDGgKFFkfwh
yqmc9g+JjWuYaxoCiflL1ik+8VOIkAXs6OlSXNd6+UXulKqJMHY6zDzl2KCYNaZA1YIIOe+nSOyy
227jnaY9hd+TGYnNKTGM7aeP4WuKmUMFc94KjSu++VD//tRIhLeAu8uvX1nd3bQQXwELyzqS7QRA
RIwRqupIBJR0k9bXjyuMclTnP0tsmeq603kduquNzJzNZFc/OTx9h3e4IUrS3zBS9RKvpcygeXJd
Hj0HrEJoWTb82htaq4blOAf4lfGOLxWMtD8ET7ACqJfvfaUCfvX6bfgo+Dr5X7ffIF4qiFmpKTOd
Lwnu+f066wsa56IttpDq3xS5akfcuh1f4vH0sK+zzD13QVGERIe37r6p9ELkPbQ3dAmrb4SAuPzU
9EakNwy048NIVn76nbZV6+gamPRqqWvmFuGv21VNQbImTwIMNHJ1bu44CcH3VAgTGtynF1Rc8USj
8yIsL6I9tO/V8ttrUqLHIXj34QKGxIazttMNJh+MNYScha0HxsP8pLtpffguhIvYptUZb6dfN5Xn
Uvqlm+WVO3UVo2J4t1a7bfkKN0zkDjXJdB8lt44LDFffUzKkMeuJURiAIDBL8OmR30lAY1BAjAYj
W5xpodgTPqSfLjW4R64KskSWOzlUyveB1ndz3haHWCEdPLSs6YtM4AJKrijoKS8hteqdM2re3Kmo
QvuM20VyaSiVzxuFD2VHm9itHILa/nBhIpT2QqNh6Fu9nTyRqOpKKw2t9MhZ7CI2kyu3gZpKLMBr
4QeuJSReWU+CVqlEOOLlkjNQWM4ouuunpcVifUVEjLjen5LqC6A6daiqThkegv+pMeMemNM9obVz
t4UaapXZ1nPac1uR83BGhKNkekw2ZAhHT3Jew/yo62nMm1RHEFyzfgXM6lAmek9XJRkf4MkbiFY0
ukYwBxbbB6Yx/N6Pr0EvUGKfyUuoePZE8KOnHkbKkT2eqHq58v60+Qr6W8Kl/fEIR4ndxHkCtrIs
wmcBDbCvosYH3Nh11SKGvzH0hRRmNgMucZ0ja5M4MJiSA2lzF2rG1otaqMag5XwUvmKTRV5GVhsS
Cf/3DWXdQuhN5bIPLVSmYY13hDqrqVWBLV3eQpCD/RBit8DMEX2NhDlviKSL6Cww7af9uzm/BoJh
eVfqRHQTWHYDyEvACS4kD+2+RGxIexYtes1yq/m4w+4OP0Xt0FT2hP99NVBA41YUjH9CJtv3iNxJ
Q8rvbsYO3pxPWkxr95fvTgvt28SFJ7NA4eajn19wlo4R1wJvRGQpUmV2cJINQoaU1Vyqe4xW8kvT
y7xzgxylm/vtMdfIfjcdd1LLvPG7PuqRgkhgpHjVsyMIHH71guR6XhPNbzQHy5JaWgI7UBPUexKW
RdlyK/xuNIcEO6ET8sdPjqRJMLKHrtq8VcLI6XnxvmGldM1ggX+lCf9J+FJmovehJcnowOjbpQwR
4OxKbGZlAvZmqA/DvoWyYBQ0MvjwyN2cOTXYuNaZuDzvPHHSuP9Xn8dgTuv7kHk3/L0asaSihQzL
VuXWxPDgH8AC29Q1dHEkS6S4dLO5C0d0gYJ7Q0xnV1Ttu+EHSJcCLJy62kHZ04FbyCbwBBbW8zuV
Hhyc4HccVsRBpYFpJmPHB53mZ2E4egaKLlFR4Wv49rAfY+yLnjkXhMA+JrYV8fmSu/4Hz7AyyRAj
uwR0RSJwwYWXcLqFfxaWfAaEaIo6xfYqZMOsrkzuP4eM6ac5zdDP84HL3K3u//dkI4EFoXc6CiLI
eruFQCZmUdvsOkTxu0IjXnyAX6PB873AQjM6qW0rNuXfIAQGKLNCTXW4rZGZ7Nj+dPqqdOUX0dZx
bi0cN8Vh3zGOdq1X4NHxRmSPmKACQVpN7p4nr/NerVHn9EUTw3J70iDw4Ohh3XaMkiGR3vR0pv3z
Dt0iCW0WVlOYLlzTXoNSC2rHLt80nT3/fkRPKlODavP/PgjdK4ugwrvvarJuSxT6zcLhFQfZ8w31
QXzEANxE3FchZtiwvOi+PJOqzzuOHGfaFxaGnuCqlMNfkWtO+sYFnLl42DDVdnKvj+1hRlgbuJyT
Lrn+UqKSYhcmHAv2b5tRkqLBW6dGhNWSxKxacZGcI2INRWE2RJ90zZfZF2tUaiUsQVEkoHMw6VX7
pcfQjc6sPqqnfcTLgHoyCqLcGQDbhPPaG5xyQ8pjpbTzLDTo9g0HPHixG+N3SUiJWIcW4XiwjMsn
8xNevRCu3DvLTMtPAV/BDFQCwI/qkTQTBfOGDyqS1A+qXOzYqMjBa0/I2uzrkeDaZGLYCaafKu1F
wSllI1cgaykRNFKg9pGhrzojGSR/Y2AUoCrdf/yLZmuqO5KnELDgEivd1OlMgjV0tC6OdHYoarvF
R76CBzOTkn+pWzCjd9XTPvm0O1fogUakP2kItRu6bg3WF5XHA9BTtsDuCCQAcbxxnFIK17pl3F5Q
ja8aPmEA2T6wEWdXIgJqJ08Lh/w0Lo/hKTJKJ9r+TRFV6lAVuiw8Qsi4WvQ+tXYaVHwzUAp8E7Kc
nZJVUkxhSNkFWGufpd6958ljH5UckCIZQvGs7FsWuiyxp6w2hMOv2zKEG5Furx4wuL8BXy+2hig/
gwRZSKOsGlX/wPi6qzGkSjuLGKPSkPQxBLYRtVE6FU27lRQ+x/h6y1SoYQfAh68oVvbXtolW5Eg5
DTTTKfzQDOwHmsSWcDW/h/FT7v95q7SZC3u7BaaK6YMvKxSf7cj9UpT/eSe5XT9+4ibawpKT731f
kfvQfjXRz2GK7TS5349dbyz9USmqGNl8xoxNRGplesYnh44RGDbkkndweyMeWqSyZimAJpjjtQ4I
1IVWXyNQmXBQM4Jlg48BHEA7O9ULpTv2f/j+3p/4kr044gPaCTNyogFw1q0CZ+NJkedZCVShMhto
WVO+ZMKjbUNQw/GnoiBhDaJO3f/HM096rWJJGAxXCPYmltwZe+LM2HvdWY2E0dloR184LyJOAjLU
jw3cWk+j5xmzWp/IpcF7ZqjgSAhZ4WECJMu9vO+BgwSJghCH930EqvK1EgoOquvz2q5NG0NxKeQS
D6jeU3k5FUCkj2QvT77p3vAvBmehmMlHjl/O8w9164bJEqY/0PP/KnOAW1kmZDeOYYBwmJo5EQeC
tV5Cu6A6ok4qbk6X9ib7SrRAzpEuXKZ9qVciXO8xIZ1PaqixjGh+FtjCZHn5eNVhvwxeSEnATuEs
VRH+ydGLqtUAhIY6ph4STNbeJgYrbajeNmWsH79VlnVKmMp4wl45+nGfgjDHGaT8uwgGV+eNC23Q
ZQYrN+9sBS4lOT5Mo3mmJdLli9jEY7+3uU+WwE3a6ySF7eOOFvE5o7YDNVi8ywtjkL34jr4ABPjc
T9Q9zxdyhqgiKqVkTzrsdoxHr9m5QbmJrVMMZb3Y5+cPdWzBNLbtkj5OdWoIv0R9XhyPhcNtkwok
fzBiM0+bD7wpI68az4EzWKIPoeAOPZP9n7vuDKa+VeFxvfWmBKjOMiQR9oNHDGMBUjZ+nLHPxeV1
jd4ie4xW2WQ1vK86yAJart+xh/6Z5o2F+OKsPivDDYsfd3jp7Hug9U9Q/nskWPVMyeErMuo+s/xa
fpGt6+oJ/u77XESiVnnba/eJNf3M+tLtBBM+yh3byT9iPqEDEGeuKb6zX8GFhjAsA2DijpwiCAW4
4jrZm0b10YHzYuuXOPTInSh0y726jxykNzsBNh/PkJW39vVlPTJU3tlLbEkxyjSREhNHU2muFcCX
sO+F9FzhbqgxLd8dj4yQENMppQUJkVWZFbi42j99/7Y6ER0c8U26KQMNpTfHJXL9tqCtUGSuFUI2
s4UIEs24Bp7YEGzTw+aYlI1LCfBEegvjkI+gVFNgAlOwj960/HCpGY8Fxf0o7a8j272jox4RE3HI
bpkB9b20as0mpzFbG/samJ0BVRG4pSx7RwBK6/9Hu2nhQZoexSZrhj8bjmcfpP6rYkNhlfRbP4nU
hSTkLW4bK/ZD9gtzGfe6/qCXgBPnRGmz9/OeCu/evk05j8EzcomdXaKiRnl2GuMuGcSO47budaX9
fV3Gugv+zvyx8bRIKr6vkjDqrODMj2m86VujARdXc6HQ/E7JZjG5E7KHDqlsZE9ge6umzjVkROYD
my0LMacJtOnZ0ccgQJEsKoRZIthqijYQuiPp/PCLNYbsIrS6Qj4SHcXU8lguhAC9RZweztFltkoL
AhJWA+JpAUMycnh6/tvw4j97PoBSNtgM3MbiAxQ+znuf0OkrlsB4bgkBlrst9ytueQocwtxgDcp1
lIXkidbMaZ2lgRZpIapaL59aeFd4TG2tWEbi+yvs6xrT0Ido6ibAApgeRp45AzGu5VEHdvjn2eCl
TzH1yyjk6zViAGn1x8Dpgta/u4as/9dxDfzEy+v1HjIfol2fxmIIniF8ZnVbgst4LGRi951aMBD8
sYpAM1IwGyFWpx+fhIOOxlTQb+jz8uUNNqBjwTnStAFxGno4RxK44olkn+mLzzKMBU3d9k5F773/
eh3kynGPNKjU0DfK3vOT8igZFuBz54x/NPJ73P6oDtAVowku0hKvQFlAFL5jQCpIWtesISnfeZq+
vDa/qvBsjtNdlrPLrSANW0kTsCIq98kKeDxdeNggZyOx25ZiPUeFIYZhlUuQiBi1YA8na4wC1VQI
q4jWQ/VCyPXl85AbZq1SCJv+N0Iqc1xKv+ioDGybciWPBjjuHihuD2HsLDjyJhHp6+LZYpmypoZD
3NV24z9hKoS2iqI7cvuuqH0K0ovvk9pr5FscoEdWtoZqz9Q4YvUHMGD7PiY1npQdjGGBNFogehjy
I0fW70jdX3TX1NHJI0ie7tX2Vv0VJgBEQ74CTBgM2L428Yg2+Zfm6zCsKHz9voMDog4uzhOHrKyH
5Ds21OL6cHEyOx0ZCuCTZaCPKXIrV/W3ZKtNN7Sj8hn/CMrLY9aqIzRequz8YEqGD9YLc/yL3xzx
YPvw+IuZXl0Q8ADo9kvzyl56nokNVWUU4La+E/q2EKJ9na9jWoMgQ99e2OS6m+rexFo1uBJEWWxE
lnGF2G/lsbJG53+x1WJrj/5ecVPb+tc3JBRRZt4nCDb/X6wJzq2r0yPMEBh+7CQRXzQe3MMJEO4p
syQ3XJzKGpuXG4H3VTzBtpteAmSCb9JIXz2Dfs5MySFeXUJ8BJsRPB43719HNpKfvmctyLiN7105
JG7RP1eP3NoUxYOkN+S/XwMxGAjF7ZuUQ3dHDNVTLD+Gxec5SwMwYzrsK4Z+5a/s2/v764Tj2xTu
qjUIveKUzjCCZxsoVzNCjsseR6rzKYsbgqMmLBiwsHoRqHijIlnbTWXEM9nNX/hrsbh+/mV9ly6r
47WOj4exXJGv7FeLqWAUuE4Ecd1N4rshAPDSmyErdPUIdsELPKOwtuB6ULg7EffSdm8j2i77s6bH
uJRPk2SW/rzQ4iY9AykqEw4lx4vsi3GSXk4LebFAofM2Cfqz9jCRDS+YHP8m0YR4rw2TXThgLTWR
7zcCMJ4yYNqljq8XHLvff3gJBcDXaDDMwr2NM6t/DI127pMuoKaRlDHdnNoWo021ECijacPNqa1Y
w9UN+FNvztFYB5UiIoyvqG2FvQ0VUez7bPQ21n6NEeQ3gEWQZUzfmHKiM3dXKfgyWsKfVA357YRK
sqExI8N8rODhw7tD7IQrG8y0wazQYfNerzWOeks4EdYCNH+R1T+b1vfGrjOoIKCcXoJuzSVOga3G
t7NRFFGYG2wDFzq8yzYPsUA7Zdkqe+FuFGJZH9S76h+yQi6OYd/1FV+7j+tceSvlgnqiXeHNyKb8
gHhgmb6EvqlOExevOkloPVv72dc+6zFYvhtS9limJceEGG/ZH4mRraZg+xtBp71NMxOIm6sGsvOd
eXYxcaciwpzjlUTObaV7m9LgQpTZeAe1Mt/I3g7xkY+IZ+dVW/4N0DD9x7L+akOV8BoEwjCvfZwC
8fLtYhgKvJQq3U53lKZLkWII2qmBWEpgb1DpFo8TQaFHBnmw2GUtLczoeoRAKflzO8n6IzV0yNdh
Cwv6qeDb5YEZO9l17nqTEcTZXqvwnUAkxdUZKeDLrE8U6ClBBJxXaS802Qc55ZvnBW+PndvOO/mQ
km45No1BnBA1LPpFi8W+lza+a18HDx3i9uDo6ZM8x018j3Gw4Wh69Bfc4r+FACl8pHfoJ8Yaxe2N
qo/1ds5DmsFpG5W5DFJpUwqu3MZTier9k21FeTpGMEZeoD0mkyYH3vs4k1MHoFebfEijMCfo3/rr
ux1Q/HGiIAG1TRNHCnJ1SwOEKGiKtwdwxPIHGbltRL6Qmj2qejHzGarRbmuFFVOe5HurBo8zHrqb
/6zDAyzAebKI+7AGCxjr4bUbBONkuysC7h+H92mKaM4+KjNWWOoksoAX3sG/btBodc/ZAu/S+1Jr
CJnTNS0kfUxToym4ziqmyyb6PQht0bbCTczlO4pIG2zzFDOUUMGC1h8B3JEpXezSAMbQ9jiPwRjY
bFaj0i57HrgYqfoDiUyoVWzHzY/L3bdNrw5YCBpMMIqxoDxwGxyVkOGrWgul3iL0eJNMpKO4fkdh
pIBo9q+xPeIUohRT9jV95a4rSUfeZcg6fkhu7awVBqn9fXag0Wwck2UXu1oPB1Yy2TUsmr4n3YbE
yFtUiobHn0NUC46PuMU8VDWBcqEHp59noln1h/gc/t9PffXzirZjyGjGtNWGJ1IH6DOUvxjZhvPt
vpuORPWAxkg5+nhetxK1qUa9pjs737XlV6N74RGjynO0asJwY0iTEhOVcSzwHpkVio5diwBGFnj9
VBqX0A3zfpPyrV6C1+/2jgfdKobeD0ZXueEPo0Ex/ugXv0VPnIHDeXuIwyebSciFSpVGbrwUCz63
em/RHp15PtlpM2C9rweiWtA+QeJMa/qx4qLtq53gIJH3HAg/P55dY959+K1fSOEc0ILog9HbS9Wb
xUjMgROU+N4rYoegnwc6J9XlewpC0oTfBVlUylKuZOlKlf1vftsQHtdE6ywj2tq5c8wf8pZtO0Vh
DU4MtQQDysAyS6EOQwmBf7SyrD0U27xS2Nttv0amBECNdypZf57E1vfxHEAAiZ0U7Uv2zmV3Oehg
tfgje4lWUA9QYt/IKO6tvBJH+TkPabXAU9WDnVT8qhTO80iGHPGYo8fZtr7/reZoebTyW8BJHt8e
OhKXMpex30gIStrpyIZlV6TLogzpxF3lPxYDLbY5OnjpgOAO/6SkBtOkwXmCv5+wA6TDCvAjLWCe
9YNMgP837AEk0/+9Epr6r1aBNkvXmDZsVipGz654oIrGzMk3cm803XA6oV4W3U3RBGp/iXguZCo0
tJGdp2kF07To19GTAOQh6Im92m5kzUlQT6Qk6Ee/QHBvs7q7FBPWBQUpQnwaVFfuJlay4nsBI8I+
BX2/pHIGznRq7v13IzZJKxaodvL/Ici5443+iamMm0OO1oIZky28L4SzgSLqJ0kQsabkgKwfaZ1K
vNEafA6A6z3QZCDnsGl46Whhd4BGxxT40n6k7oCEH+lolsKVcvV6YoaotS22E6QXiq+wKYrGFzn3
R3c8E3OnLLs6mF9TBKZrazgnAWJkTWs6jSq3RuT2WMlUseYAI6qI7/11XXKrFV7VFamO2zwzDlax
t6i68DsYbV0d1XKmqtE/uGOjymj+J5vYG6HakfN1quCXWMs24qPz5FlAnDQuMAUyqGed/CW6d5C3
37Jy/HORriAp33fzueaXivN7jW+uqltNi6vgOnwznMDbieprj1exWisF+w0dnIHjaMrkySPPtdWH
bMhNX73eU92XTGkVLJEPAMKIfnmD2n07zkeNsbauzkK+RSrWTg82L+7R7/r3eRtNnjc2fMBtgXkt
9I8+vcNWHPvqokQkdBL1q80xyqTMX3si2kl1dTC2RgpgpdFU3pG8TBUlZQ9JOYJ5d+v7HrfBuy6E
gBQeHhWyCX457A1tlpm283BxAGCDSlREIxDoBazVy5oaPQeE2LqntT1Qbd3ZgF+nwbo6SH3I/dYS
pguX+qyylLTClkLjmokthfpIsyDwLUKWQ6FL0sO1WukuyV6rt9inH/7wlF8nGvCKQuITIS167DFH
1Eh9nlk2CsHQhHfyQq8pCw219tOtqfx60qKP5zejcy8Zkak588Z1NqSdDJNk/P4hIz8LDnKXOII+
ASSJU9cpcC5KDBopcNGUFZ1PV8EZHkNNL0Lb5ocxqXk3ETY0IaE/SCxD+940rIhWBH8GNJxS8dSN
O3+r6whh8mlWdaeQSe71E5XKmYGppQc1E9MSV5yTBo4uz1mxzHQpxs6EZ+72imNYqyqV5T2w1kbZ
Z6CwnCFCM0NFrBxcx7eP52v+jgychJpnWCwwlsTrC82mu2MRwub59V3mQlm7S+1meLe6an6oY7rQ
lFrsqUKp2lXQWaBdkNA0Eum6m1guWEVASXGrELf+fzyFT/9T5l15ZDFze+OH2Rt5hxJ8Oc5qJEFn
pIKbtzmWkt1jUs2jJDTMUXRzxvQobIXb8RruEOkAyZIwWJSz++OdlQlKJh/KNc6xCkhwKb/zIzSg
TlA+Afyej1XxrWTR0EP225ReB/fkIcsc5uDlT7uyVW08M1kTnEtWQI4giwIBEryPnb/C3UmzBalz
JaBgi+I+ry9gvQ6OQvwhfGzU+NufR0goCA3SKU2mcS17Eada4lhoBTxnP4UN+86vNl0JJh1VuOWT
s+XlSYdZhRzHigtrc+njHp1+wn4UXsbfRVWlNpQS9pt5RCkOAqxolhZcISPAi4yY0+Q9cma+s3pd
uVZIxtfM6Na2wPnPToqb1pi7ugSZ6yYdf2zbvkKAqwDdaWYafOnVPVBwo+aE9Fw291DsBZ6SBvpO
Avcmcq1ezMy9+pzYcNMQfNj9J/KHF1BVbOD2GRsbDIobI6sSwS3g8qcMd9ewtzfbpy+jNzK7uo3O
9ATnWeOnxAPA24+p9r/gcBeZcBMU5aemKEtCDBiIDR2MVHcZFRFAttfGHQPPrvd85dPM7tzXZdeU
WXPkO+NEyUrQb5aihjHkMR2o5c01zqgEGzTGnEKDDDv6XsW0Dtqrnp0wCwzLUEsxNt3qytWGcVy4
78XRoX/DDC8UmLsY5uCRjBu64hZ2OxxGU7Id7a3i0XRFR8Yk6dDDeTB+yv5eOQseq98cDMSEAHlA
xIBgZB2bOmY4Lt2BnXM9KI8xC/Hp+DXfQ2/FL+1jw/cgdYfb4EDkrjuS9MPgfMU95ExgTYccxFdQ
m4BQz01QffKQOJsEyMpv9Hgq9B9mPT072oJMUdHU/Ag71FMJ2TJ0NodivN+pciq0XOJ2iuMv9AIy
00YWh1KuhVwiBUq16POjp9cgZ5+TDF2Nx96L/Atqs375nCy8fbnyBm5ZeQ14xozXv4TI9PvOfiZj
+rsTTTNyovoR1D7fwKNB2d20Ov6tMb61PRYePkNoN41yfGz4bu7pm6v165rRxMK1X97AePiuE5eB
lgrr7D0FhHQg1ZI94KEFIImGdFmjIFilTNJqS4CgDQLl+BOX3fZqrcjS7ajdPmood9r1txF9huAk
rAjkeL8PJvfUDllesAnd1HTZAiCp4co9wvwP9MFvR9t8TST5TcQwPvOUgMGbf9XxuNvne+Swm44X
L64HRcMZYlB+Lx15E7CL1ZyURwsFUclB9iZsciladiR0F2GWieMTt8DpEXlZJNpiiY9x3kMZ/07S
rPiBC8s9m+kY9OYt1ynBYUFCKJfDgTB2duIERnDTiCoUHFwbhSUTjUATvo3caJsCjfiV+gKbYjO6
7AFIuDgTfUTJLq1ufxP2JVnWd5NRmsVExc0TnpKtuk6RLEPJo4TgLjFl3MEhTEdguCq5ZErLGhqR
IcyzXU0Ueu3gm4P1TeKTKQXQcyPmEsYpB2aVichHXA+kx4Fwh/EJ00F/3brIwE1J9j8wOwohkgDG
tqys9dndcNjbIDUhj82SRivFaQnlf9PfX3HaqfZYFWsxHNRXMnFWwHFPNdGMk94SHPVu5rW+qLy9
0Q6SlQPG6CtgT/dD+NvYDU6Rs7DNdr+OCcvT1oduhE9EpmIPk9xtENAxJLamdja52zxsD8ip4pCM
qv4yr3Y+MztmOt0wAPwaqQV96JXVB3E0PwjtUuZWVoFFf5882nR34mdz2/FO6F597B7cI6KqIUGr
l3EGIsONeVj0Lg8RtA9KXTihbKZWyzkgb1+ZIsO3a09gBkwRkCrOfjq9Q2r2Rd2VMcMSGSaOV9Nb
jVL5q1szd10iZc+Sr5ZiaY9CZhY7ec/XDW8Qk0cpNVyR5LDqBw5Ejf8Jt0RgyAJKhSWTuKxVUjQf
2+4X0h3yn3wPsN+76c7PDgAMAcqS+p1xF1VYLnm/ualPA0B6Pl/f2vHNbDzSG8TzSJrr1BzRU9lV
mtP5xHJiuztZxry/kMUueu7EMSFRQqodsZ2EK6UEt5urzCJl2s94OvtwrqHnu5UIFCVxwUIiMuwB
9yTWHK2Bj5NVlC18Esbgtjxcpa4Eni8Ad1Ks37QVJRn6i8P458lRPpIPIaEsYY3TnXouywRZ62CR
XEg/PXUSivPtnXRe4JA/poNMrOtjuBCRLr/ZGCu+s+Y9Z2CPkfIqt8C6cOjesGxt9pSUYWoLlF3E
geGymbPcx20Uy2+X0krPYais75Fg1KbzAGH04RMS9OnujjwiC6PDUaEIN+5ezGEJVext7/Bg07Ha
y/4fF81oImGANLyC127H5oKDrrOSOq81rYRnHF80sC9NWE8C5j6rK3Jh8e4dUyDZZS0B6PAgSI3S
+VYmtrk4iyzC15nz4gIACBhim9i+v8E7+0ghu98B0gNigFkbu+KnJ8QkOYhKdUw4Lb1sSQuSMpDH
AlXzsivh5+CbKROrOO6j56S31QzN46RnwyIq7Xevj+leTX24sczY73XInINEjEzjkjM+PVe703+7
P1OYMoJRKH38WwZ9NYipYSXtkHiIq7vbWq+TyJrnmWwaSsG8hld9ZkeV1xeSZ4O/q9tq14vpu4RH
YYv9Iuce7HdUSzMpU4cOaxUA/6ooPpX1ypxiQd0vITTxncDLf8CYAcZo+tXiSs9WB4Kjncqe5enh
HZLmnlx32xfToIQMgivkF2GmX/1AbgfJk0IZkkv8sSBAqN9/aKv6TjBTZ4mkP3zJ+M5ue4quZwZl
7X+YmZqQ3a1YA4NxPu/VRUZJlQKyyJ+E5qmYBdBD0pC2PEXohTD27yQ3YzwVIQhS/2dqLz9xxMm1
37KExyToekNXl+WrEBzTmOLl1/vPI1vwgjXEX9RGt8xrOmvOpnTHvvZNtZhEFHPmz+19WsrP0/Ow
M3bYuSKru097LX9MsTGdcTKCc4D+8+/hKpgMRFDfcdS4GWWfL97sUBH5bNaMdDnTRd/Px3y0F99O
qKIJtakMQb3tocfCqnBK4XuYUux2eWzxnw8umpie9PYWh0GmxA1n04sIR/ukRZASdO1VHHCZ9u+m
StaMRfCO32emHlgJWtkesgSWN/xSuykh8iDZH/poxR8i1wP9JLNbCCckc8ngNUIJtRUt/oji2hZn
L25W28igKvUu0TMbtMBjygBpnPQCuOLqIqVR9yi32NqdYfkd86WCi+gm3kQdJhnjQyv6EHLSnTSE
bGPu/koJEdz8+MpilZZAZALzpuYPnyh530Hx+zpN+x7cBzGPKG19547CXf48/rTq2mogsCGf7vgw
87+/XDqAW1PflscwbT60IZODJeej3P0ZHqe1aC09Nwn+Sj+5bguKEw9u6ttJ7910mTrDl4cBp4ZU
cdvBFPfJbNCDBqnmAJ30OCky1TCWo6XHBRUKa/U/nP0c4fk+pt9QW9WkiXmThUsWq4QzS3QuUn9l
0VF2DOvnCdY9eq696uyuFQaJkC2g9qZRMgmzmKDB0knjOIrmn/tA4bP1t5a0rksJgTGlrGgQXWme
9T6XrxAQj6+YPNoiW7Lai0B7j9ePV+p7zxqvoFT9eqJVSYonsTtECObKK/TXCK2/52q4kLnxTJoS
GDkemEYaOUyT1u0fR7OMcIMPUgQtX5JAXY3ZijUrZczHQVL3Yrfb6Yju3bxNiU9GN45q4pUTjgY6
+S80aZUByt31yL1RmlBL7eq6O0C3eMXiJ+CUzOAWd1vtWAcrqYxYJSSfAJkf+0ou8K2S/o4RrVFc
EJUutNuGw4eA4HKss5DT1IuVUObHJbpqEIA0uLNB6C1d7Ms3ryz2ozs6L+NW4C/9GaTMgzftXk2l
CxiIRvdqZyRcr/LmL5yjLbSkTp0Q/RfLzeU9G+cNJBr3JT3p7HtRfgYLWmojRr4Xf9NcsubrRiZD
k0ESzr1G1hPOURmlJha+IS3o0GpwQoUwov9rx0N8ecrpyTPeLkLNjK/1EDuH426RXm9xMwxYC+TE
Tn05Sn6uv8Ewr8fl9+64KytZZfdFGKWQzTrLozBBjJ3qOqJJXKEvN3q+sHXe2bwAARXHPvqCFWKh
p4rFiH+DTOKYFmtnVyZxsk9Yt8Xnjvi3DLD2asJFQT+Mk9NyaZBugjq+rYUZoZEaEUqgwjr63abD
WKFdOkeOPkVL5GKPIr9RwmEIFg2NR+KQwb5Ia4sg5KeXqacCOhqS8NmUjdsR9IzFcrx7MhI5LePd
Kz1O87Sf7gBqVTmMsPuBKoyttQ/X2KWammrCyyhqaY6O8IOr04Ik8pcZsu09GETCEsNlauMmt5zz
bsUMzN+CGHp/XaQMxBfMRgV3235sfw1llhc/hjS2DrVUMuBbrbVymOmSS25LxSJh7+BaIKLCbwER
beFemcdMkncvI7f73ZuPN9El5wP0ftWP/eAAtnHa9tOvjUhkkVtyGCNly97+cm+iyp2igvEAiZQ/
Uj+Tdbm1NWDgdeZZUhT+cRSNoVfUeiTeR+m/9esguohCvbk5+34mb9s55bgzJs1Jv0gJ4VB7gFf7
9yMHG+KYWHJbdttrxW2YOEb5hQ+FhG3d6R6qFGTG8a9tHoSUR/LPMYj7zPthbIDpoHdmfLYrJogb
Ueg9891DoJOvxwM33aPXxfxQ0tHzbAdAaXc6h3qiwrF+xvyUdc/bbVPeGIlz8ARkyvddok4+UfFM
1jxK2+4RenYvj52Eq8YI3Ds6knQnlrRUn3ueDOwzrJ7ErvL1dLOlTBmxhqPfuAhy9YC+YzNeZgBx
9atSM0oOA+EpraiW4gVNwuxGdXoNTyMk5NQzLEVARHLKWZ8gA0v7iUb74qX5YTECPYt2YkWGrO3g
Olkg/rbcK4QQG+h3L2QYZMRbCNU3ORfLauSGWE8EIeBUZFz21IEcJELu6aTaNWoN3hAtXrEMCDVv
Dv3O+IpxWtLWvaDy3lxxqVRaogg9bJlqVaP7R9sn3A8CrykkpG//fvUTDPuvJeeHfaUiteSNChnB
7FbOyngAMqRmuq1P2rfUuDhXuonwFSmWbZ+BuviPErV1TEYLsww8itBNmvX7yCoNMi4Rm+Vw/uPD
LQ558MS5IdtM6EDZHc9ztQ8M2T2h1bMdSY+ya/Oz2CmTu3FN7T4Ldmt2+ypPgMiGNMo4WvreMND1
iNkt4ZLRSi0c4fRPOpVTejPA4SVjjhqb62VvlUeXXmEPwbm8vSxjEat8TKvXj0pvH39hD/XQzELl
Wagx8iKFCKZkjzJw+RrUkSWEI5OLw845xMdvxCfiD0Jz6eGnn8capAPzy4x5n9FyRgWhVE40YkA8
84dAjWXZpgY0M7U4gm524ny4BMVFdpuASw9Oyyxm1A34gRQ9NSni3zloG0Wps9XQDRvJHNRHqX7K
/vZ7Ws/hSTXRESQ+a/EEjX0jw2YNOC5EG8KEXBt9YLxgnym9uapkdaMHZuAg8CEi9llmsf7j0kyF
1V0PzPU5QiDbyOmjPTSYWXZ5euMbWV/CjcX6nZ46AI+WgabwybjTldo0YiHGNe9CF3TK2SKLIMYN
5ncRcvk48HGpkzend0cB+a1cIzxbVVYWw2oI7n68LjWwV4PC5KnuxuEfiPYM7/j9NR4HAI50yDnB
UvS0Xc4B+Ghl047/i/dlH17FSCth1EbjcPrMO2VHJNqpfC0TvO/VkltvmdhdM8Wr7L3UsybU73p9
Rs0zVh/VOvIEF+IPHADYxv/afUQZf32a37IMRkA7kxSDv0ko4wUwk8cdDNZcdktjqrWeD44LL0uP
oeByswADUopCtc84ebAEpxj2c1EK7Yn7O0P6A7g+/U28j96X9XqXL4/DehvNohyF/mAn+G1qpInc
wLP9G2juy6vEOyvg1D4Y/GNEw8Xz7u6L0C9U+kSHxXtZ93NbE7oawIroY7WY8DOM9qO05uLM2OTr
ZC43kNC9vWMtRhZl8bZONkkRNK7wpWxWYSIYuzeOnnHoSfHgcl8ptGc1W/tcFPRFzbzPIPzMq7hD
xAK3xGBK3OFOY7K83/nr3S9bNfpVOjspjZ+N8F+FSTyVrHNItApMeJXFj0qjT6zkn/Z/CJDtsKKT
jl1JEg6H2jvXHJfvGXqlB31BjYfxLDRKVX6vygyCfn8GSwyAR7Fh3qYCvMathn3RHxonv8FFVm4h
UoSCPUSGh6kVtEZaAajc2SRTbqZNYnHl3uwG1NLeV5Ft9UzJHnyiuhmEaoVIZNW5qS8TFUA66yGL
ojkEKuT45w4jocYypto6ktmsfpOHcXIK/I0feFIw9twNjowCw41MQ2w9lV17qUJ6iISj4uYISbY6
ePCeKHCHsWM60f315NkBALtFR4XbUZpvGYdai93vzvr/g9jgOEwU0NoZWZ4XYNWDfu96SGauWrxH
eqp7CCzNE0CbghpVKMX1iqQ7wsirjKuT9TmcdzDPogUKeaCejOm8P8gyJCHy/HxiHKOlST42eAzF
MqpTIfbRWHeE1BxsFyVywtInygvdsrj2k6eEFwmdyRERVxN3jZyn5kXXwbLRBPSooG6uI/ZIHi05
7AXWmqMWEqatH+wBa7LltdjduUjQrLYbLOf1vJyPZkyKCLJnznwRSgl6X1gnNHrXbn66sPxlb54z
nBKAKAJhchJDrBg050fdQ19Kano0QXyy/4pUnug/Uf+GpWuHvEzF+dxsCt+j4csGKGXBbeVPY2BM
Ge3oofhul36NTUBlZRltgP3QoVThKAHSB9Q4vkiU4LpHkKxqJkLX6vCfOwnC+20iH/ZlVGzHLlwF
UHqvRx525ztnt7NOV6sM93qc+3ZDO64LtVScEa+vqI+Jr5G4xxps2h+cnCCyOW510WW0O0dFth0s
//xNZmYuq8qu9XdqYxjwXb8n6CIw3qy2oQh4NdgCo33VTFzh+Tf7I3RtKZcNIjcTndpa9PurN0iU
Ck/EgweHnfNVevrp7ajFa71zTJyPKPHj+GT4akkvYW3NZiS2rKypiOKO6VK0PEeyluuSLOpkuO1l
tFm+SAD0pPUFdSZnqgQAoxNOuXAwLxa2p4KaPWQdnVjtqlidsQEvtw1bGh5ZdSkKYb00uR6zwmc1
XNgQwlKPj5tewvoABY+HRp9DuZ/pQrHlma4FGlURvKY9eOsyHQrrWW3iqZPaDnvbRkpMh0JcVc5/
BUfrv6mLvwacDC/yr4a6ciekrbmq4og7U0XF4ZbaRJobPPcyTTDu+nue012nJtH+L8ZApLcimmRk
+oPNHFC+Fpxi8OmXOmd4C1ajYMLIIXMb8iOwTjBenuDLH6vl/wZd1mT9GuzLROExl9BJnHfU5ja5
epXAzvQeAt1Gg9HScRkD0B/Mp25Ttze1kMBZAdJn/hXIY9o0OVdYcuu6C2cnGD5ilSYLzOE5ybKP
APytVoZrxAFvk8p7TKYhwKj+h7WlAx0zEIsnpthNHSPBEnD8hEOmhjJ63q1C9ZzwWFTuO2OPklDc
xZDcDnyyjAgX5/dmmbex4qo92efUmRit1WHcp/09ZUj3KIQmych5FLcDITiM0RgOK7b/zNUk2URn
SJiReccNrTmWxDqL/jqeKnuZwopwfcHsZvOa5lvtOX1fO+U95kwx9G063djOTbApZK7mU0oh9ol8
gGrgy4eKgC3955tJNDkicu5A6NFPQWyMywyL6pp21+06w3EG7xarxqbAuPdUwr2IxnEMVEdi30cm
FIF4FWcosCH0ni/foz3r4u16B2PwTEfgu7UY5KVbW65EsFy347AgdufoL7TKeQHznT7Pn9l6s/RJ
x38p9gjh/TSEsffVbC53UBm/WnHZfqTrmh63K5HFCWME7NXy2eChfN5IYDfhtyUxuf3h8fpCS7OO
4eT7rGMeRH3jguKRCrVAvjBcv5D+SSL3VYlbIK82+xi+QZxh/ewMAWRHQYaT1AFJnRM1tt9FZkjR
KtFK0WNCz5SgAskT8Lc78zzjY+3WW5rZcuGnp02h1ujEijwIMFekzxfFgXeYRG4Be9gEHOhyvmER
kFildSg1grpe7IYlar/MnG8ovvtOuBMi5OsqK8Ftb51/IJIOwPAh/+pPeR78wnwQUNlcxYrntUws
5wKDVorVTGSGZS8+iBeJ5P8AgkpvlDHNpfFBHEC/v0+JIv2rMZCnBUdRSwAdlOsQXbpfn4xbfv7o
4gIb1fzUWj5lNOpnJzfiTaVESu3mPy+CVul6GWaoBxe6jNklQdTPu7qdpdH/ecF/ICaqDv1igj4A
Husplq9Bcg9TOFV0KKwTE3oVcWAGJCy/8Yt7ZDvMcPb8WsMy3lmuCVVhb13AENVGSyQ5RWvqsDo2
8shoRQL0XN0vYaMbnEJNIvbVUQIyY7pUMdXQ7I7eWpDNDyaxIh+wskz6qdV21lsmu4Gz9yZXcAwb
1ZogahVEq7ci5vcPErqYItAjrZcK/xZUmZ2KiFPwzTF1VEiiRs304Kgf2CBXu/CFuYngHpIRJ9Da
noR5BBaqcUEV2lUM4AUAXDLenikq8r/wNT//gMrQVWhIdCrp2digPn6ttcuXucRhB5ybQTAxyQqM
6gO0BVDRDsghM4/lf8JSix0UMaHv/SD3nrcBxtuRZWkdfvODDRfAiY7pXTDesNeuremU3gcIF1fd
AbPr0Yy2FqPq/Ikwyk/j001kAQ78sh+0sN1jhx+3UQwuV3OUAKYV26TXb2joG/6onFrM+adADLzr
lI4M3g8NyqmYFCE89l9lS1RihHlfj/MnJiE+V1RrrueGXynDyHkoOiNz2D+3CIhwHkMSuPlhOOTG
8yXbCmIgc46OZD58MZ5qhtOtdeltWKBicERoAiUc07l89RSmmqPpIgWI7aoSmf8563/22KTT44KK
p65qeGcPGGSymOY6lI8EcKRdpOXDQx19JVS6Nezuk+rAe3EBrCnvvFWlEn90KxK8Y2Bufw/2ouUF
FevUHmHzNjtpPQlG6JX7aZxvGc6Rbc1l3hMmqcIz5ctFnma6HcsL1NGSrUNGLlrtJFjCLEt4wp6/
J7iuZZE6Cedl56czm5K5ktNl9ZTgwL52l+Q6trTFsaNG3aRDAE8QUzKh29GmuDe6tVGUqwfpOM1C
+PZ8G96B29KLNQ+50no8u9WpWKwmrl1FPvYsrDuqERsxLOyGJavO/FVFlVSQM9+z5D1VUz5qRDng
d6iYBFvxe3GeN1PuDX/zdq4fnGClZzN/wtly39fVCmN8pt2YoN+4zvET7W20+kaMKWSa4xJpyXr+
yVwQ9hS+Ofq5IlqQZM/XFDVHv/N+54hGtrZbewGPC8VQP1dqrI5jDlfA++heFn5Rr1LnQJoVMo8I
8z04CEwXmv4x54NgkNL5NN4tYZmw0+Qt7hT/mgJHDvwcZ8ExX3u5HBwUFRMqcmjvDWAUZMDQb2rz
vfIcZqK6ebkX6YTsRhYTK+lGyJfz1RDOLyL0CqvcKy6I/mZjuFFTlLWmWcHa4WRfR+1rIRYShw6E
wevu/67xtyv/nF07frzCO/LomjiGo8nmiaX0LHdFqh9VJH0urs5yG7D/Z/LFsL4nIXAt4b5OFnRG
jEC8nofPsYlLK71l2+G1klKiX5HMsJH+GexF7rEXrrCsVARVgclsWK2hR3IvBc4wZDcd0UZDT/cC
/8saTuLNDRHx3gKpP76bX9NRydfAeSUwsSXIOu9T9GY5kBZK+t/9aCxGOVmUPe5iO+/Da4XmmH8B
5SAoKgoQXc/p7ct6GPEkojyv2cCqTNDm8IFXFz/bDhjV4z+9V3Aigw64Db1PJUOGwlNv3Ae5QYpO
rIEvyMaUflqaF4pPLMm3RvQIvyIpkCEHFXjI6gq+uyGipiH3WGGn7tIZK0W5apS1Ar65qku/Luug
EXXftXZ1T54w8WwGCB3z5+ZzVKlFb/jpde11zULlH8eL9i1A1XPuKzH17RvC/2fA7dggomDNbXJ3
IWo4M5B9huaQ/qX1BwshsUtOfzyud75ir779so7GrJ7QSu2//t+kXlHH5KJHxpmWHcCsSBzUnzpi
NcDBWLMJNMp5CuhzRbaoOkBUcDKL6xXOiNNoiv+Hex808JXEBXFd01qnYpzE4u3UcBS4sPa/NgRn
VbA9FQ3PKq8HsSsH25A/Bkh/7wZZrPtqR3c9/RldxdfFNqR83AXEeihrLS096xUpCDQS33cQ2Omg
BWgfb82HjmhE8vgK3yjR8qgptQ8wTQaCQaCmU0/6HsLkmsTuogpP1QBLx/c8Q8ySIRrLipGDrQTA
fGyujZwMMGWFdiMtresqJO+iCAQlc2ugrq3UCkdKKsxDDli5FbDvD5qVwWortbmy2562HsUpX7/V
4FlnASV7doi8NXvrBkN/fkh60cE2ugu517bt52gVpCByZaYU+xRX1ZxzIPhXBe5hOzPDvCbLfHGf
UeCjVRlxR+nra9MbTSRgdQMF7c7byr/m2GVQgZOCDUxFNvxHiRqdYeKEmjQUhHuVuL2W++Ia2/7B
kdd3ZuQK6pLXwrfX7QKYU4R1lNvc6dSjBzjbu16fEMBIMH2N9nfGG165oqf1tigen6bvyjrhvwXE
2zVK/5fzNdT0V751pBP5qMdEv1/sm92MPcJUJwXOnAx7ov9yjvht0zyjF26iAvXREXuKmCBDDIXK
DOqfkW3wjoPF2JgN7LTzKNGaLHpljyOfTQEc5jeFiZtdKiUydc5z+RAajYgjcXQR3PsIQRDwsG6U
d2Mul66pYC9VPMdeMSCYwqeXDrc4y+HvwdFIBOJ9Xna53eMArJgD/VKbs9HY9YfVNTz/a82jtYcC
lG3Lf2YI/EJPQRh+neZPoY2Y5hdhvZlqnqQVWDk7wqx9HfBccitoKTvNKhIU4ftgSPSYWMPqFG7s
cVGqD4sYiDpWFnzP7YNJKzKjll4h5+9husVhlqryN4+fgI2S2PxQS9Y+md93obuHH2ZVST4xknBX
WuamlL0t/3tznLsaJn0kzYE14YEYnGjiZxohMXdXTAxPzSKZREJXxAs6HH4KcqG+NonWnOk1okfP
C0Ap4D6nmvZUQWYbgnxoUDBnQJGPMAT2Tiegwjb420gCgmo9Nbhm7g7TRMKpElnRpCjzTm2KLe5x
TomP0ohFSZAEsY37Sg1bCy9wTGgT6/IKtRQ5FwWzfHHbHwn58UbiVFRIbUqV1VGjjDPe9/vxbuZ9
7m1I2aMqxdsWLbWFWYFO2glVNmHYUXQgbwTe6xbhKhnkPlPwqxGYFXLlp/XshL1v47Tw33qGOPnH
zK0bHF3xyLFsnQdKWKshJzeOfYa+zPFHIVmDURHkMlfhiPP/dvlVk6cl2xJNOxPe9tLypVEDx0qr
gBEqV4fXZuH4YVAw/MCm0Ysz93gybtRnn2Tp13GQQs/fpipdulf8XTQHKtJSr7sIi7Tuq0zkyLyN
0lJsoX5J29IX2I5cBmsyNN0d/FLLT8vC0BRynWXYou2oqk6vR4cBoWpE+2x1XTrSsUojnJ2la7dw
jtRSCONMK5JjHti5e7jo8U4XTv1k1wSyJ8Z7imuHqOFlskK6KvGLK/lvHlBG1Vka65kmD4RXNY7o
pgFg3ooJ9UjnctxBiBbJyb7rxVWbwQwRX5wu7X2+HJnuKBF5NAifaLQJHneqcobQReSKHNsnzPkR
zpZ70HWhjl2ZEKjRkEVtYFcRKjqHAcx1b6C9g4rp5SyY7eFE0lqarhCQ4JI91UbbodpV1ubQPCye
lxMRCN9/BJGf5ag8fWV8wIlgaedG9sRpx2+2WUbXhNbeYil5nmI0bZgAj+UhpZ8ptjBvb4QhCVFe
/tPWcxNAoWEu6qjIuDH9OFbwXVrglzoT8EbP0Ik+Oi26bTDzo0S4QQTlWBwT3ScaPsaakLL8OXKd
6oo34pkmutE/EStxuDZ6Wm2Q6r+KsIp0/Hdoo4HecH5BM30T0Oo318mJtt1Zd4g7DgEnz5IuQHXp
UXM6G7RHV7ukslPO8jTGHjVrwiNbA3FL5H8SkXh5smgZSU4gwXRyeexS62aNrTb1HFxgeYEGDQQ7
o35WkwZ52hdb9e+dfXEtDeSIhllNSTrD9d7gljy8Iyxe2SnmNQL/NA8TPrfVqpVHNkOZi7OITiR3
9HUY+8dFMeAGAdnW9uMbFSJScPhZVipDAPGh0mH6hLxYUf0wa5MfM8wc0ZV1F2pTDZs2d/0bHlij
J6GAkansw92LdjO061EXlsZAYUpohJj/WhuigSHpiRO0zuAHOSlgJe9L698iNFON4Hh47rPqE7ar
mSF6CUJOOdxPpmhASkT5IkHn2Y1Qa54Fp3FjPe1MeQ/fKAClpLoOe0bP8oVeE9f1DGYBOAW+DGEJ
IPZ4sflj7nLYAQTvTDBcsZcSYI4/tab8WT6UJgbtBg4NuC4r8Zc3gFgzPfbj4R2WYn6yMzB64QBm
Rfxfco3+P8N0U5HV0W6M/tENG2Ug5RCz//cqPQU0lxx5FVoR6Cx2BJ7gP00T/55sAbHRK9+rGRtP
UOU0tEyzyUoY1+3PDrVeXMDNV1sh3wQMUF/DsT12qGqAAfcO/48XEayC5n6WhFEKdtJbu3Z6jRem
yGIGzRyGdtofwYqsWMBIA9n9tgYFG6f4kbmMM2hvTF/kgfwLzYnJ9uHp1CBbT1tOhirH6ahN3cEi
mPNqs9jt2TYA7bWoiveJJ1kS5XgjyUfipB0IOtFoSCw3zaDpfajMy8c6RlwO3jjkdH+UeoECoRz6
oEeIKVvknVP6kpghqjiKHH2rdjbsqquLCSdVUSFrRK2XZJF8ynOm9RivFGhbKyPjmZ3jv6TbDMj2
1WZcweq0k+QMC4VTp3+uAghn9Xl4CC9sfaHoYrgeTftYd2iScgQDgvXpeS3xOM0vjl/HJHg3gB1q
QmWYtxK60a4GZlPd7GiN0FRPnmzmslup5BFJLX+EmpJRFjqBe4TOrrLhidX1yzJwS9XoaTsqhmcm
APW/UHC4hdEI1vRsZMjO0AlaSQwaH8aQrEfOq/ZfUcz1/YHFnU9FsqnevrAzGnb/byIxFxPUIUIp
E6XLMyMbItqz9kv4XRkZoDhrLF37LCYj1JJcCpyND/0xKSKgo1DWTzhsnqllfeV/XupkC9y2SVok
qq6bpDaRIgz5pm/7/RIeNiWW2M6XftjgxCtTsfPJYaCvqPlnXy/lJs75AneKftfw0xZQjMqAu+J4
Imbo05QC2/YiHxr5HEs4ltme9iJMeyzSuZqyKcOZUrnwp3cfwnGr+pG/KLBtvDAH7iaTGnVsNGMC
JcL1oAGnER/pDEsOvtBlfQSEvnvzluTSlAIpztcXFNr/fXJ59a1tqUUSXPYufqr/gPtm7EqEs4Rk
dmMrk7uSWu4gubG8e+m9ml9nx1Z/7AUxfH2rXqqufju6COU0XxT7bveCX2zWOVV0kmNAbZtMs843
nLDYN8PNrnrxgZVpWk1wKQs913h7yS9v8rZRfKLPQwVNjw40al6WVZKgU3R3ljqM3CyFUzc4bB0D
Sbz0mWzyuNfQ9ekegYX+GqA2IPKjBn/CWZz97BK+H4HtaScycqrFXIebgkVxBEs19dW5B80sTkeP
Z8WQAfEornivQkI7b9Px6BaYQyDjpZPYSR7Ev80ktB5jMI//srulSudWDc3OtwdU9tZ+N2YcHuY0
rdGUJj1Pzdx3GBfTYxfCyVlnswXc9a5sESH1R2WRBzRTW93W420WtCBTlYwXbVawHB0x66i8UQIM
O9llGM0Wf4ql4fULoaa6GiLw7z3CyiXjIeKKSzD/+fU8KBaokFU85U7wyR/bQ0/ie08Mfm6dPJ3U
BmU3PnS4MkxlrPy/rwPHDTZWtsUKuDBA8ZQssIMmWg8a++pMDxbmwEhf4Tpw7UmaPJaub7qbs10S
NEDt2xiVS27oA7eqk2974NBRPSVSW9nbH0XPLzDl22zUKArQjN+4oiC7rvaDR+V904EhnoIg2UJy
e/jcO3zfCWhLSmq9tIpYUcZN0jQUjnZ6Pe6QnPgCzFdlmlu6SDE4J1sXqN2vYQMju8cYvwe94gQZ
yMrF2WLX6ypKWAdiqNR3hNCqfd50sE36jVO26/4tCn+yOafng84+7TDBLzR2cgBooKxliOwEjt6G
6MBmTwYUzzhP6pEgukc+CCqsKq/yglHYtf3cIRAerQ2aotopwd6pKjZ1Z8i5iDiV+ZfiOkb8YXLM
gbwWCctotkrmSu24xTk4+gSW7BFwgRK+d1vy3znWCbTfyRVccq2X27oT42mNZSewWvWCwfdVLWXC
Ci3EYJJnNKCbX3M/6b4xQ+Lmr2dUxlSdrVuuuoWKpFp5dLXlLwef/CZXG9HXYaicx+cydGBj472X
p3FdyDxX8QKtOhJ7svndUQiEPzHNprRP5liiOE15UHGso1gwwuzVretFeaopqvqcZ1chgsPvaEWJ
FQm2MgZAD73HGgNTPrx8Fc2lat/zrni8q0avJ3t4JKyja7K28T82rB/SrQYJzPlLx/45xLZX2Zid
yyq6JqzGSjbUT1ew0MiRJXt+GRpDJYODC6NTWEevmgRogJMYorXbO7Stb0v/8Jsc6Ejv6mqprni/
nPBtEwiyeUoIycbkU3+by17GIKz7ABn6jNbzaJJ/34Pj51vJvVho341HCK1MUPHRwsXthplnNqcF
foatJBmIo8ixA+kPQNJnWbiV+TgnT0HY0leQ9I7zjepA2+UlOQQwPuHdocic6t6KaJH2iJ7KZTTz
uOBgHde6vIfKFzSAWNkzbemt0B70U3sVQFbIMLKBl3ik171j9rG7NyqWR4+UEPAanjvfOUgdb5hu
LfkV84/q2GJWu0ncBXU6pBT5HtT0DPlb1RrYVcTiPafBi1szfWb/af2NxOaVLwx3NeMck0AtXf6G
UvNNyv5Vwpb8UwJKuso+uPxOxau/K4v+fCyBeIJLSrok9DqZ1nHFQI+SnBiCrd5q5/U+qaBRuhls
WhXxS+LPwsw+uFuKuQR6fGTeXl68TfS8/94ZHna3fOFoyAPwJme74WyfFHIC8o0qX5LFoKr1p6fq
crqvuiTiB/ObnzUZSWEhWiDVaqus7v6JdAuRCMtjQpMjtTT6F+VcT0dgVbi0Yy/q65GnM4nStlyT
DfOJb2V5SvDfj63dGWRobJcTAvYdcv28MNYB4+tB5khGqPAytzRwn98px/7mcdRJhmxbMS8Cc51z
dRLTeIsOsrXlS4P9qMtvfQoMaOeAeBXK9/K5ZdTIcafQKimXsXtxU48S6T+SDRwukhhriighE52i
ekhDXFonsj0FbNDy23TGVBT+bYjB8KqpiTOgmzGM987BjpN0inxRihQDzsVc2D/IkRqkNosRbgRE
pBPhBenqF0JgwRrKwu0sgYUkn+o+CbiDMMx37S2zXcsbDD6lurU1oZ0z1JYX3YzXK6Ppyz+VGTW+
yAVOG4+tN5jcChcVMm7ua861HnDgOSfwhxg8qJBup1yKf7/eAM0LzttBgPFW70ezLyBbxJj/7I0B
nQ5yv7soFi6xItoM56+Isog/xvAr4Sri6f2y3QYxy55+7RKuKDzSPLke/+iQARG9mgOSVRc7zlUj
V4shl28lQduHW2XH47wb+0EhBl831KuOt1y7l08H/WV4GG3cZTHNChLFermrmR682QheNMr4+6z7
AlspioN80tnmhVSX8YY9J6MH5JZucyGFTe913te17+SYlb3LpQAB2h9lopNSEJsx2OuD4GI2DvGV
KmmyLf3iPCGJxIC8uGhgN+vI10yC4HfJ9qFpmERBG5S9BNByhsaXtZ0M58nQWnW8zfjPFGuAKxBN
UQdf1Sv5Rlq+YMiKS7ijgVQQluKgrSIbeC6zPHUcPgO6++qWytuG2F3QV4eZStygUwFxNI4kZwq7
t2zc14p5Spk26ZXqEunx/mo/OMh8LWPux432MNvpxFXKQtx6RNF6UhrlOS5Nf8LLPtHKV6xdBvde
ih/7hz45d+3xMKft30TkRFcaphFD4FgkBgfnE4EMSoE+jmhq0c4njzFY0j7TmO/2vbzxQIxjlLt0
dE0I8YO181amIrHfzo0DyCNjB2byCcxGkX+Id+iRvnlaD0gzWXusovTc53SIFJqpYzKyq7OgJNLG
gKQXWDmTUUXzCBkTjmHoqs4QEtS5dFBBwHStVvLeV9e0LTgWWr1FJ1d1QA/8QjNxfCyAMGKXGZGZ
Tif/y6nmC9n7J6DNIg6JDTPA4Zvq3bjaq8rmnL2+jjTXGIpQtor4Cvug+auxLDKdCX+66rMTK2hQ
fN0TZoiQfHYsNEyda7GU7rMT2uGlzhvXQl55IpMb1HZzHHHh3T3KSDoCXF/4LQJo3TP5Nt7ox2IU
9lcREtwo28e0eZJbHc8yloJqKCfZpD8e/DY0DzzMptwu
`pragma protect end_protected
