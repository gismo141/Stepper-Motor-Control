// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:50 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
IbbgARgA7A1iA2eGzbkmfWUeweIoC0NB8Zpd42INiO5RInmPKjgR3Fd7Oawxpqag
TTqNznaBzUYl9fmU9UY25kZaWtwV5JLTMfpXMCkobbb/GVGIaCrlwvlhLYrm4/Ty
MQpJ3vLV7Dl2ZBuTHToOBi7CQn/YJF3AILy1+iUHRxQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38960)
ILidEPUGtxEl7098Q1hwbyLf0Gg3jfupi452CIT+rHabHKpR+rcLdnzwg+jb+/Fh
Kxy9pGma6/tXdkA2lpUgd42HSoU5dhMLfXD7I/l8Dwz8EcCBtmcppsIV+AGH1USx
XbATy4NC9Z5q3a1eS5IuETog7s/btfT2YlONvuSMynnFojz/APyN43XiG4QaEbqu
pCMfZMKfwy1zx1CRiFS0pGlm/qkifsCZPqk/wpLWdhj8oP9VNWrzBp2jUztCrtwK
cB+qp0kuZmSWm89iyFinNbHzwVMNckwu9CM1sFbfzg9NmKnASQEou5BrWudbsI5A
HJ06CTGf6N+o25vXeFJuYIXoncYBfQ1N3HgW3TUOfDfM8EYWKNo71tzhnqbtvmFM
KioA0YXGk4V1XhvFRrUJmLnk57GhBvmQEigPgnWK/4O8DMLYTZP9qupSzqh/NwWQ
E3OutgCulSmhEH4K4m+P3+EG7zlpuF+SYBiolfC/F4Lb0gBTDjq2ayQKlaoKZiD1
7nzNguurLxIfWVztATe0ju66God8Wpxvw86Yquj3eXnSFg/uxx2K4WgAV2J4lOM7
ePVOWCVHXIZZ3TXzKLgKFjLdtcGneevtSzXLzRwBjbyc2DYI45IlRQ9cNj682PUg
k+NbwOechZ2vS8lTnvdCLXEE9kZwffoGy4T1ZJa9Ac3WWQQXWSNvEwr6cQS4sV8l
6QNo1Qkf+nO/U1j6AFWkfMvQIqLecUMnVspYkDrtnxnYlsvgrOz7LrnIShyypGHE
mCOvx+5BDQWKrFAE+vSDiwJgm39u/ncb8bh+HpUXseL9xbUCiukI9zSZzg6ICWdU
r0nRHVX6UBJg0NOm91DkMB+ITm4Yl1MIXa5KCaHIfPA2XDArng4gsymHZ9SV4xV8
7vwuOSEOj3NZ8/Gui0JyAu7bQeOIXSXjlSY4nj5pvtCRyxPXs4LWFNo3EV8QgNks
c9Ay2F8Rquc0tliWXcw+WrWlMeHkLVmkp+B5D03ut17gstc7gQ9dQXqcP3ROy0wg
f52Iuu+IGaBYVUU/qaqAg0+oVa46nPSHQGi+Zz0TY/0nKff1kX2s9IPGuDSo3gTF
dRYeSmZhV9T/F4WT/N21uDVrtxftx0nTjkUXVu4EwAu2J+82s9L/+aSIaTLCarkw
eeDB5WYr63YQOh2+WlA7o8mj18fMhu78pczNjCjegrTQfiNt9kpYIOReo80P1AJy
jc3ugvKQxdTJ/H3tiwihZ6anS5hLupERgGN1oKE0ddmsW+9rddeA7fyHGH0QpZ+E
3k9bTd0TCa0Oa3SzwzMyaEY2OhwFzqUDJWJSaBgClwGaCqlGAQWosTmL0Ssug363
pkMRC90YZ7Hs4CFt5I52bgiBhEbjV7SOLnuq7O0mH6UzanYcIe/0DfOVUhgxs/MD
ybWqjXqjaVNLwI3q/YYkc+80esv5vIgv0VvqFfj7E3oRLZ9NSPU36rWtmmjtcnnR
KVqwPSFgRik3D/e4WJYY7V0IyBpM8XpBqSxtSJeFWbXBWiTkGJGD3nS8p2mR9kXE
8GG4hP8dmyLlIvTlbuMmPAC6SZVoWccUJik2khGbawoH/ZpddZWH1czrTcWse3Lo
UHk4SgtWkOA6tHafrxJYovM28DWvG3QLcO858Wb/0GqRfh+zu5FChGvo3WPmtj8s
IX90fWoCbH1Vb16vk0QbzCfxcumVQiEEYz1RIfGwxZ6pxEUFd++B1jqNbOuw0G97
LRSAS5KeRkpFaOHV5SjAg0FExQzDw7ZmnIFv38aoC6dRlvJUBhZp2CqeHMPeAGwb
YR8kixv/GfCFTabjx0yWj+7ApqlbCsdMH0qRGvfk45MlQIOC8VaZHeneeQkIn1Fn
eDFnkM5w9NOjHgukWN/fpzIVwwbqJ5E15Oz2R83YzbTvW6HUjVkWhuFxXGEdrf7x
OVrTp6Dy9LY2uTDxN8kws059aGH/m6KZ9neqRywXIYtOo/mvXtmuF1NmoNzMHVg7
hvncaT/5MyF69v8+5p5dZ1skz7DxXj2tNAQZOs6ZVr4o5LYwa8zM9WqQDc12eaEk
gy1ayLsG8HL7a0kBT4LlwFbOz5c8qrb+NNQKZS4RIw3SFNLbryVl+GsnvCVTqcDX
SkyiRnuvfWtmIH3OhfhnLcpd8MBRd9PRByr2aShu3JCE7gbMm+4h6Rw+xqfxDPbR
+CEbSGTpGCzoeO9VcjIAOupNsPrNI6TpVvpPeZOb6zNTIj9C+4NbFjjXAkbs9596
NvzewGgAmCKpEgrt7AZHdJ6dsN0YhA524jiQGSL3yxUi4ZDZ6wnt4VXOPNHySLIt
LBD6BU7kc9ZXDr5kRBQcMkffLatycn3GVqht1sbAW2HRooQ5cgA+Uzneeujowkr3
0Bq9kx/z+vG+9PGE40fnAXcL0Pp/diYsAfjWEpnsEn2S2D7MjeeVfoC151z3NWOe
zx+RO4+Wzx33x29jWK1j7i7Z6qQKMEg1EGJZlvaY+L9mLpD6PngJWKxM31+7RLLF
nDdhnFqcSV+Dfnx1EW13Fh+wPZI7HZ3SR/P2HOLiQzNTKJnnZjTY7UON3nOiqjTm
KgCtV/U5TYL11XWJvvEyS6lu1dZMPk1k1JuHXsIbjedEoghY6Ks2bnX/cHEK0aur
qQWS/aGxH6HgO6vz8xv84hYUV80PZhQb0kdkoXukIXtDB6SIf/rWo//PuayhmOwj
EwSOUCaDHJW01ML5HBO08xLqBKbScqgXmvHnH+F7JZdWT5TCyPRhl9gjadil+R3K
c1DxRkeixeAZcoA9AVhiSyoMdqyRvqJVVRxTKn1o56heWiLk//wXnEy1LwbeTGP2
zneH3oExgpC2AFTnejUU2qUgZExWiH7Q40zw1FKoQaugMGUt7RdOd81Bjs3WWiz8
PGWu4zXqfQ3fyDHj8dZ2qbsg9JEL+Rstfw7J+lFIU9D2iok90329P9QsgFK+pu2G
mU6HPXXrqr7j+fUZs5a7QKNOBOAUZ9YnSGrjT7Yuy6S/cWLKhDnPQux8AmqbOIeR
XPKaYqNWgTDVNKRuM/DG9d/wEhpcdMWK6gqoqyPGpPSEY4Sk18SPz3dQ04wCLJdB
ORKlLzigdgTfC5aNACotd04vMFsKwwBbrnk3kKZheT2AyznPef9optiCgExVOcWt
/iZm7st4n31hOnqdOiFY/E9UhBzllzvgUyr+MYJ2GUbojf1IEkrA24M+N7pX0TeC
VBj/3YRlO+mz8mYavI03E7i9nQBYnnM+Y13UAEIOT+66L41AT2/qPrS0FmhEt1cF
mWd/dg6hzpGFBcfk+5oEQirKBc3+vyAY0AX4ks3d/qXcojnvncffcV1shnbYLeOz
nTQEd5hE7JImcH6OJbQ/fmJhXA3zDjPdbA1ihJe2RqfPolEo74uTqTSVaTSq9nDP
XJOtkBkQ57LNro7AgW0pW58AkSy4K6Hf4op8J6TGp0yQnC5QDRp5iR0Ies9sLXEM
7PBDzHnTQWd5JWTdhS3fEoXZ+BSBrLLBGmvziMCmkSTQTWy9xE1rwya7UXPZNugL
TTvepKmKsbruz5pVAO7UVoUOoVBSnDk8dlup/8bWyKHlzQsZwq8Y0mZeueouILMD
85h0Q8LWPyyN145JPBH0DNb4H4sltBxbnnHBnS/x0Oi82f3VRQbYiHX6oskiUaa1
lGC7nU83Acw8y41R1I/tEkeYJhGw1UJCyK2BR5jLcO9QFTGWfLiFkQnUT/Cw2uSK
s0mTzY/Rrf31LADZ10nWIHM210ikS2Zp7SBU43x1jYk2Vzkheo+YsVzWtqpHC9Ng
h0mCDPriSTIdZpZGD3FqtTYpzPakUXWx3a3QaltEbk/dk+XVBxh88QYNQkASktfw
HK+V0R3ySUPoQSLXLi2o547V6QjW1GBKVTRQlSTO5yTa5GxvZz+1KkDQRhhXssXc
TI/UWT4CsMOOJMySOu7zdoOv/0Mmg0oCUJQKruHq617TteHRZKH2bNbfG2KlgeDs
AU1qRIVRX9J/xS9fsy1LUpUiLKQ9IVwBkfd3GBQSGEnaJf+xiCQJ5bO0TPUXImOe
lO4n9WWOAKcISVzq+Rp2OtE5Y80TNxk67RVAbpk6jqSvtshMlu4KmrixXbVEcTrw
DR4FnLQEuPPkDdp18+zirXXKGeOPHvhnoFRY9aqWlBffX/03MWJunmg0gApOm+n5
4XdNUJpOoL9bmKG0vIbZBYN2NEnt4km5Syv9ngOlg1UwbkD597TWpieh9lxFERY1
9wnHgm/FwIrnddsaGEO8qUADiFzwwYyK9R0kxS4j58azy5BfBRCvFSRJZ+uz4zn9
Q7NkXzw+RvyfV4iBDgX+2AVC3pI6CCQi6JT/r3gfbZfYrofRriAU9SumD0mEbADY
l9pq784TfDQMylr5Nsl9YtiaG7haWew7Q7X1wral+wGI+6vf1T0L/etWQTtfvPXx
oZO9zrP71YZZvCTihn5LvwttH29iMfD58XegBHPlcKuSQDP7QdCDMdD8ckjG15sw
dtbEnaZ2SJSAQBSW75WwmRMvFm89tLE0u7FkXOk9z/R6/0k7JXtUXW0kbdQqhEfL
Nlr3Zh2z0s7Ezr646rBZ/lIQcglWQ5J/JiHoy5LsAVZJhUzP2SeM8MvVexwkXhks
A0k2Uo+NUeYqIgdKlUQDl9SRHWYQm7v4hSBvQxf6QaoNkPWxZb61nedxjBlmzEiG
IIYaNbIAHXTHZ1V3hYuEjPegtWre5hzFqqB+jFG0DUpa7E+PEsVsKOqe9O7g+12X
dD+6rBhP8rpDJtKES000UmGQWOAA43UNgyPlK/53zxRS7ZRWbah4niKJeIAnb719
BVV7RZuOVvLWASlKiERX5MbmAmVeySXFXC12ou1HZjOtWeKm9gBvwRsRYpLNSGHr
Eud3DgFAYtb2UDj84c7YUCLXnFtxpsBU1WfzMZESutm7CthQsQ+1kyBI1rw12V4P
Gj9ARVPt1vt+2LFk3/JNiUmwPXWm6CydSk5LPcXrJOSYsiwB5MgPrSQbXWWIyF+U
56QVIeDLGJlQlisUku+6JnwGtTszClIgUI3dRQOvuHD/NjNFnzMkjLp5iQN22gzF
SbfADNBopG158dZJIlBXS08jlu/+gLLONsQcD+Ze0sjrp2yUOHziUJN2JhOivXai
4VHjJrDKq93Gtw3ZCnIXgmTMGsRc8JhZJY6n3Q082+vG0ujGSwucS2Ldmv4PxGuZ
/sIhgxwajrLWEeKehBBii77tePIL42aDWRCXaXiX4YCLY66aTPouzNf5hJwxuqh0
EgR84eTDCKuilj/kMEZPkXweLI5w8A4ycYW5KcH+rmzSgBV6rjVFxwAxySYitboz
warCkPbae8KyIRNsJrClFPe8iw9DauYxUlB6kAMiJq7iI2+9S6T+OYVzxFOnmdS0
Ez1s8wceiEC9aUJurrSkEEBP7sZoxEwDqupX2qncCtxpbAtcR4TX0mOKTMbEfTOr
SVTIvKSF9Uy/zOAB+yjaBxIEmn+QPk04SbUwHi2oFUjZdFWUPcCIM8YXYV0Xqe1W
mOQRnI9rvzAUl304XeqiyuQAimaCeUDSDIAya8dYsJKEmmyLuE1BGRdroDRvbFFz
GwicDAk8Vh8aq2LbmWuDHBYZdEomvz3NLrcnFvzMknWe6NBID2yflL1oF1EvHo6T
RVr876FShlgwqpggy9yu5gMMQ1lxp9moAXOVF1hfuu5T6oAobpxtouJj8q9n7GOZ
2yaS4oKC4xiiKPK6SmnTFODo7nK32OB9ZIqpnMb7CY3+yUxFAH7xHzCbTEaQ2g7f
CkWOka5eohpL0DuZ0bD1JXbL+U6hNLOp1LTusEzZ6X1sIhIZLQAhGcpuFHm4Le5K
9kRlD3i1bnJiAMdvn1rzKSxqzktZO26mnEwVv27K7uD4bV5NdAQFPemKSuLlgDRT
jMNsuRGblgGGrOi4Lk01TCkxj6NPkDYR0Y749y6sWJziQF7n9rl6CeJx25wIsrxZ
ZtjSLeumNBDGYN00vxo5AO5/JVMH9miQKoAYduvDvoC6QFyHKKPBreHidaUe6xrP
AaeHrCISbQXBGgGgH5CxHm2grnFSSvdTPGUf2BYOqdQO1T3xjzI39spN4+OcZ6vL
F97k1MuptgQBFmgyZC824Ix+cKmTz83aNC5igVaUrYmNertPzxU20EhSA4VSgp6S
w3JTKnUTme8wln8dOVIiWIWux/wc7boHlkSpiL/Ruu5ngvbAerk7K17/kp1a0SKn
K/UHZtSFhsSw/wMNUp1KjvWYS4XxmTuda8bmiXJOeuNEpMMUqMa3sM7FXm5pmtvi
0k34aFRsLuB4lJbusndfTA2KlMmF/2guuYlzsHrtWnX3OGNn+/WmrWYxYE0nxrCC
6llTRwcDLFKpPRDVlaKvaDvzQdAuLcsZOHreuGq5cAs8wfFNXWNKKONGA/wz9cwg
RwuVT/lE60QvbrqCbzBsPvChlAwytYIklxBOeqz59XqZGSl+mC+OMI+hWZlVonc+
dfVZPqT4DQWBavRNmcADT9KWIHB2f/ntaU1iLHjjxpfgxHGtGFtYD5eRr/+xFD78
BWEvnGh3GwZ5f14NXWMoGyMgPsiBYiX+yDC1pmNMEEQn7RZP+wt0dx+Lho3Ip1ba
iqQHbomCwyeZA5u5WqnG/23AgHKBPwJGimf2zDYoUN2KCeXxek04H2RbQJ2Yso/M
cc4vd6b6J2LL3YmbGqxAOXc60ubZNngjPJpPZTQdkvtCoiNdGAl6DqsDzaUtXYrd
1tl7IpYLYiYrRFcv9tyonoKA0zVvYyovDyvc+ih+keiwwggH9VPa4zmD9/H70sim
KLeWLb+7SGO3CHVgu1NTqMAdufC7BmNeh6A6MLytkrAadzlvJnUPXuO4d8keY1N7
XjlfkL1677SdxvJKoLhatmV6xjdMQO2Ur0lXjhdPHUD/OsApxykpyH8g9tm/sbqY
DesD27mxjcjJZv6pTNSNK+jYYwm6jtRlr3f5tYLA/j4qBWqKzQXWcwwNnPtyg/vh
jy5CTpiN/AkYZdiXHz8PfmFsa8j/NSv76gk2g2kBCW7QRsFtzf+UzTfCrtZz3Bnp
WDadpKhUpain5NI7z/OD/RF2tQPfyjJhSPD2kbgBz+Rr5kggaBIk86ftqzxGkwSj
NGRdTJNgStyYm2qQHixKlIhdx/mQiREaC+0bcuAhFQ3JFakfKNTnsdGe9gQ9unWp
og3pWPztVajVo7o5CMlqZj13A8yIh49VMUIhJ0yJE8/m6oKDWJJBOuKQgiSw71Pe
O4KME/1FE0iCn+KN1KZe+E7TZ/GXGH5lH4ws6Terxgv5s7juW+4CQl63M6L+UDxh
xOYR0jwPEVFTTAtFJge3P4qu9Dyn31qDJ4rjYvk97cQpTM3WS3MHEs1l+gLjwljC
Nh80hoStbSya+r/mho3Bnc91Kh+WNACxmHkg6mIj7mwx3bomAmyxnx5lYnsLfve5
vmmAN51uojqKkGJolP7KO7PdL9hiZ4F3HaxNzjczGtATVaLnnvYfIOIZ929pGg3m
IuKo+o3HLF5V0spVPq4zBk2kwT7ZGtoz0btM/IP6VRrl0sAb7PEVvceHlD/zFg61
0n6fi4wcvoRC0t44CvJ3z0YNzz1+Q+bWzSlU0VMgzsubc5UDCzc4TsHuH7SjDk3P
9y/BF0wSd9GfPelk8ZVJUSQPEi/LAYhgNBBIxOtPrzdcRCcOvDxFsQKtXXT4U63S
Ypnjqus50/OHIpTVhCSu3FxzXVJHW0tyxuhhzl+a1qqyh9UMtwVzpDr3auvU9dU5
UluAmasRnIOu0Tex8W67cm5908ESFYfW8XISC3D3HDsPwOVRAVzbZsDs2PK7ToNW
3+Y9nhx6KyWNtaopOnBqrnZluwUU+4MiDPVLLYHX1fJhH+rRYai7VbQe/YIKgA2g
UZ4n+IDapazf3Ci4AmyPOpVZQr6XqG5t+RW54alA3v4MMS8XLksu+Nm4qLgXJxEQ
+rvCrmaOhYolh7qVzvQqR0JqvWTrFNbz3+5CDyCmgPhs6aqyzW2ZadTuFbf3hojE
reyZD2ajMZC+Mn+jD8pNOxFEljyMcLEh4BthAzS6537qxeHAjZ62RXpHxxJ8ZqzM
Aw1Yic1hZpm4cxj0Eey58H7VvEkjP5zGlMnmtAau3u6Hf5szD3WzR/x3UHbLmD7z
PruhPT4Hf3GQvvpzEoRXv1UBdAmr5TwQ7LRdCSk8o1NoNoRSY1Vgjl5aMW1dOmCE
JiRubgfShE7X/C+qNfwDk16SN1m1cWBi/S0CpFt7iqyiuehdyIBuLVQcwknuYqil
kF+tMfO9CNTd5KeZAxNkwwA0bB1/lJJkEANUuy4FSrZLtu1wrM20DMMluBq3QhYH
y8oTYpGTuB9XKyojcO2a29b89o3Po5wWTHriILL/mLXUIeB4DJx5hUzOqFXNnqra
9ncioJ3GmFt/FrdsGRlHbHcgpQt7qNg0aNhCGf2b0dHAoN853Od4MROQfpZeSfjL
QmD8tfzyGtxR+cKSPbmecGAx6XBE9otTicZK8u9IaB7KJlYIIUTAUQ+bJk5E8oN2
mkwWdlAa/kRdOFEB7CwsSkcp0o5NpJ3GGkCYxtWdrB7NQ57NUXnGKOZe+gVFjIIh
uB4qh7XQQ1H6mPScNXzFi97lu0+W/NWu0vfdhqxEBwNnn/j5EVgSGlueJ+prNO88
0EXxf7Tb1YBDHPhLzZvVqLzTrz8iSJ623XJdt5dxby48eXIYx/rAuOAQnAcpNoyO
scx93OofFfxamhl7c8IguuYlEdiJ0SfXyVwC2eqXGjN36uFJdwUslqQ01Glnqst9
xlR8jUr3zSp43EzyZw94q+SnDiRVelMwsupNFWkW2ayixvGFzjT8TVaInMbFEzDT
AbQSiwj87+m0l3piuUI8/qT27YupF4sjJwIkIUYqQKBlMTbC7rnBvcyS9snAaHxI
LO7zOnidsMIvOZVKvGnIulz7z03V5Bcdcl78CnmteTI7Ay5oFtV9X+HTodpSGcdH
Xq+X4AXso27vbiDVgd7GD0Vy0+T9Dpg4Th4rTUIc3yRIIUDhJeb+0hzmkPAML1u/
Lsd4mKnNXYtDnDgpzQkIIZwuMmYN2Cjd20RDYf8thOLD8lWZDo4VyVrvgjqbimwy
Ge8yQuGgBmCuiI+wY3gCKP8XTkP3eB2Lfy4B2UtuA9CS7q0uKuBWO+bHXgxfEuSs
U3AQhKnX8XmS3RTJea5MtiDN8v2RHp2OKfiqaWNewYA8ugWQknbayDHy3GqY2xCT
pRZq2ArXX4umSswGwpsL+9yi9wKfzUGbExSVHMIbVIGbizhNEmQAqdhS69KqHoP6
B3nu31vjLPmjvGc8Wo9PyTW/wOe3KAcvLuR6liI4taB297wDTfOnqQmsYl/miw0N
NK13S9ACpV4kt1zcwpi4SuGkSFL026spU2nxFPENurygdAO9NmnIgElbYutbZRii
AHckP2K5GTOAUs3mlvVw0zlpbxUXZuRGqmfLNHqXFjmOj3vlgC5U2wdH9OooUC0D
K7cr8UH63nFcf9bK0LF4RsXJA1hCuNc81761X1muH8CAlxJqmmi+M3h7bM24/7hI
Yheh1P/xu6kNy89Vn5mfp9TiyBchIZsGDFoDyrBsW8lOUlBSUNPl7NpZ/koku78c
1RcTpZYXC77PA0lk0NmaykbCtYkQ9fjm/ckBh7arCy61/uIldNb+nvnokXQfmLk2
Lwf6JTuy8jjW3yGAOop4mytbq3coYedfa9FuZgLnreIrE6/MeDFyHQDXmiQ/rlDy
UNINt1ShqPgtZ+ngS33XnqEDCdmhiBKpRMFLHENFnir67Vd08nGEDaRZyyMc6I0k
SfhKPvl1YIc2gLt5U687xGNPWw118vJhz8yFTGEoXptRZ2rwVFvpOD8OV5TTXtOt
sKw6sBAMfZJAVUKEbUtJh1b6mvGtebYj0blkc7I/z7N6HQSiw0M0aRfOI7CturK2
vLadOTLXqvWN6pd4ekJw5R8GbWQWB7+wv/F2fBJo56qAXRoeElqnVoHRRgChWnRT
YMPKGzPgQYvfbzeLpUTTtvj4Wby54nVV/8WVAnLs2gB+RKRyTZSVL5c8QloznxTL
KDYAscwZyBKy0LkaC1lBbi2BT1OX4PCTt7YJSkHj5lydhbAF/Qdljh4aS4URHDZ+
maSbxhS+EIGuTA8xGo0Uprx3UpLYQIAkYquzoaJzSO3bAQY4m2iXlMUld9L9jny8
+c5iVtli2HSt3ThSAfTTu+MS9no4P1ylLw+myMy409+EXHNEljVAOnRQIdyURX6j
Rfu5p4ifIKPWYOq/YYTwaCk26i6R25O/RUgOUWdvsseY7MH5go109Vp6PGoKYyow
3aB4g4J09jBwlpwpcYJ7lk/rbpevth01t1dZ6p2BZmTxz7NV7YMurkAZtxLXNQe7
AT4TCRzz1D65aFj8Y9dSeOdfEfnw62NxSPtaT6F9BJJILK4uf2NWQ+JU2QdLBbmK
Tnq+g0fq10qliRjlUjAnTctC+ClfPTeWBIH/AN+QbSC+ybNBFdR2HFA2xVflbyjz
X2oNKLOJKUeEElfFzAzHqYVAXYbVXy/6nhmrDAwq/7PG2fFHZe3OUGdH30jbCJ4A
or+Si1jNvXYnn+y9V+uRKFhzs3AkaZ+EgIBqfFpVVoqNYhcL/MrUuZiaCNC+aSBu
2cTtWxjw6tOVVo+/ajRI7pkcjU4rWsg7QhFY7FAhq8yNGTin+oMACq3z8wxVK/WH
AfAptJjkCPHVA2A1he4nK8qsB4orwfqWK8hG4Hr79Hb6xKOqe7i4WVuUYFmFukq9
bysAgxpcoePpny0yXlqu0A2bK1sPcSubekSyJH2mPloS8HlpiyVUxxphtvshoXCd
2KNv/Zq8UZx6aKw04PRkCLnSHAbWj42SYUYyHL5F3oBpaY8wvGII53K/HwdFqP8T
qtlSJmE8IqBCspDDA7Grpa46yZ4jifVwRfdV48sCbq+I3+SWhRX/TECCrKkmxUkL
z08s9j3CJhtFywNA4S8zaMH53NWeMmII2HNvdC2NoKg/HFSO4/ARSTL3+q0tOKKp
ElumUcfT7Zu4IK/HNitSE05skOLUC9ntxZRn7rXLQBqmim2oVFP17qrfau+XGkWg
LEO5+PEv4zBm1JZNzlgaMPnKiTWUT4hjd1L3N50GP6iWf7kVMR8zSl/Xm8wD/Q0D
SxoIb7+HbN2Xrx0IviI4sRN+EU0Sg5yR1UAnrhyGpkhRqzEOXFCBJdoTboSTjOtO
AyzN0Vjh/NAYV/LQk/Y9jrTbkIzKTdTUToUpTfka2DNwGFPHc7WUDVIB30Ikk0H4
rB1rP6cOLyz72HCusb1+8coTDgxUlEsIUFkzBHJ4kC4b4TEYdr7sVmY54SAF5CPV
YqUez+aDtkEdYNfBkdSvbO74hOYnYLUfvU75v89139iRD6DJUykCrsWUSqg344qn
SUGUYG0nozu+IurJi7WjR3JpIp92H/QerTgknfRdENxmILEl4vt+o6oh/lJFLWwi
/7JwPrzRNRdS5tPQFscVVtmQHdDnwP4X3b58+PqoJxNakSGLzOsR93T7PWZtjiqz
/bJVI5oewv+GLkcHxP9a4+0zevRa1/vOObpi23S6uCuIaIIiXiw0KqBWywn4/r1S
Hi/o9vT0QsjbSLim/vb7Yh3q548FiDebd63bIuYyHyGg7QaLXFcq9IfwcSX7HfAT
zrAj4GG//9yaEdr5dCQLxvBKZ2Z5KLZbo8t98I9QChpMAAEryGxa0qAMXjNpqY6Y
M2yxlSODGIYodJnMzF8es4yzEU0waMLg5jDUpjhuHJrbTDdCofpEWdoMQ8Qj7M1K
cidDRZzwQuYh4sQiZfggETlowlFvMN7eFkWSmQ39knAu1ruNPMnOIy+3IQyX5zc5
MXK2CkwVcVzzH0G66lIDwebN9ciSyPWUWjURWpAs3ru38NXsmpBLbH7bWDqybyMb
0s7STf+dtLdlxcNRM8iNJdu3PKc48OwHEeo4P1Xp9tr1sOSJIYlMwBwCtUUKIT7F
+RXVxP2Ja2Ym5tNLY1laWC8MuAp/1zSDKIbMWGOkEFp+lvbsK4FSd8xk90EzhyVG
AVUL+ys4Ps9xHHyiGdjzh1zh9bW+mCxHiHMQN2mCxJTtWlgeGlwrzcpqb7jtVcAI
w2JSXphCs/XXfF9kWsNtfTL05x0ScJV+ICfTRzvbRLQKow4ZZAC/uU+ME9YRSrRF
hgEebAzmpgwvQks4G3p9n8VhcoAfG90JXThvALO8k+FrLxosw2jZB6TlaFANhgMm
wXowVJYDCykLswCC2stHT9lRZY4tata2sJ2tXOy5T21gV5qtaWNCYG7Gr/f0AQoq
/wTmJEZ++3HjyR/o5C/uzKuLKX+XJ17s36EnvPhIORPUISE0Xg/LZKSqxNoc7ZOi
2j3DaADZYUTV7ZXjgSr8Q/IHmg00/2Q9e1Ib/5RgUyPrzTxs4MVFKMNDLwguYF2L
Y0/+9WyThwZ3Q6MFlHUlXZuaq1E5m1Pc8Baw2vbgtQeXMlFWALrJdKjcvxC3dBtw
dC1dlI+DZ6lWgW94zw5dx2H+cKNiE8DukOQzU1Eqve8a5JX6hQxwljY0hM/qCeOo
bLpNUYR2M4rQem2L9r22nVeXzwCOgbi5VeN0Ik+Ffm4bBFPgAuRhGsEcflmNwjVp
mRTmV+Yh8sFgeHQLjKvGLStyNvgytuHZ2rSXqrzHwNunZ00bzO4CLpfSyYTtZt6l
YiE5baPQh0d8ypuu++gzaZcxLG/d92P7eLfeNuadgx8m844URwWa0B5Oari5WyAr
wHN2Y4TOt97eRKaEvvlpjj8QmylL1PzdWJcwSc6+N58MoNH+52CRyddrgVxO5H/I
43U/nRfWF870/eU/tvheYbdAaS1WcjOXqm4lJfqV25VtObprituYQhkUryrvaChA
TU+GuSpZkFET6XYD9URbFaKhOBMnJkG3l+D2QBu2zKdTX9JCqT4nFuIp/V08ERru
B8RxXD4a4RO4r+h2+IpCBFll+UAnEKTZ7L29XhS62qYCnYW9+Z0AaAr+YIA3We1s
00/XPsBUmu93nHqpv9IoaVYEzOtFs9MZgfEakgXutx2j8ktdGCnuWBY7MZAYqalY
iFVAL6ZTCgs9brJftEQGVt5cjd4pDLKleKcuEpeCTK18TgPqfdvcUoyJuvyw2gDg
9GakbYtIhlj4/5gBvQltoSABPX8RrcDjaUIYydgMspnWRf/CY5wSDceswOjnrVJu
xvg6NnTiWrLFvue9iy+luGOnQayY7B/r5+wyBcCpOU/CxNjjK77bs53EDEF3/e8M
abbhZQX4tE5q5tJ88TWL+i4mbfglb517yiCgLHlJWkUtEf9GSJdy/MNQf3GAOgVh
oWUMxkYXdect0hmpEmwtaOtWlv0tVrggLAmk062HUbxHe1gmMvsRSlmgfHC3DRyM
DLKlzVnRDyP6+QUQ+0IgJ3pi7RnG5NCtIXqqdG5BUsn7P4crIRaFw2nKytmMZJTN
I2UtDe7i7vnNyAgBzkZqj55ZhYfOlVcAzjDHYU9G0qYMu42IqKq9kHjOwEvD5ivs
gRUfA7n3Daz4HYx05Wxen1ZvR2R+WVYSasdEmGsGmVEft6ZPu3pvPU/sKIXi0gbg
/GK+e3gXaypIv9Dk1OeoRxWWZ1rcVjXiAHINT0kUrE2e9fUUO18dUJA85XsLNVCb
vNy9/IiceO+lUpdVRlzvXnHuNSTm+1U4t/4ayQiePVSa17HzPaqNsvBqLAjcvP5G
u92z2HUq0hQROijTderr+urZh38/INid79TUi/y/G2w7WJONBixHni2hxLVRRnox
OkEhIdUxtP5SpISqPZNJaYvESR9Mh40fzDJUt+7BHQi1zn43M411PltlPJuE2wpw
EyPMuyq5OIASyoPRVfZ+QynyyklUqcIbB/V700hNP1kM9UBK2cXdE8kWijPAoSgf
fHuKds1h9MKOyOAAIzCOD1f79BA7DjGzoKwrzOxUMBS+ehA20wnCT/Vb2nIFPj+w
aQaWKGZXjZHzS4KAMSXrmLxLct+zoGzx/iDHNKYWzZZaSZj10o+ZIzq57Y8gWWQ+
HflHIkZTLi1ku5+nh9DkWM5SCf3KSjFw9phFKeEHj48pTZLeRuAP4WkKVccZ1gRV
NCsDK9NWcQq25S7Cyw7ByJYr64QEhkuJruqkvCOTdiqB/1yp6arGhBKkzscm6TSj
T9hVl7ErLWxfSDJRnpr/JZdBzvJUsD1+Y4ynrKfWMWIXLXklGX0HZ5P3nC4uRDf2
hVci0eNS4DemIzbbDKewITeuwwxg52MwRdfYO1Luqzzk09Rm/Apil0gQ6Wfc7dt7
98L03uTvK+F+2FuS9WBTWN2PFjswDoo+iT0Hw90ImPb9FxGRUJOdxNFUTiwDOvvV
MMWSWmS52IRkXrZGB1DLk8AfMrv3IibQ0w0T6P4uSf4FI8HozLQH4sdp+VRmtNoy
PDLU4z3+pjxqsklYDaEuybWR42jF9fIBWzz9SuhFBRspW5wu0EpiRj8cQv5/eLgr
7mQ2i8tkrsNWuMOlmXkn9/2YMPHTknAyyZlFINKnCMVfDicMkJgbeFNt1Nh7kVUX
dSpSXpWu2po5ck2IkCUlgaGjJfz6GVpCUyXFFMwzjE6xUUpphSnvbzlEBUB4UMd7
Iu7+tta1zzJWmiSaO/hROmJQ5e+XNpWib/1JPTlf9QTRx55ngCCmuOK3Gb1qxkhx
VreKvG2AQYySVnWSRKGpRYsn8NeDtOAPFRGQia4CYhSWCqPoL4b2zEkVBKqJfM3T
fWeJF+8kqy8QMrkskIp41+2w1tp2IonbEfBxA8iRbSe4dc8gUcgjNfmnGxrC1qLi
kjjIWVcILwzO6y6z4/LnvO/4s/wgJd7Ur284DD86RXFHet1zcv2+wWYhkY3B6lxx
ybSZumotivLqs/hYZo3ep8Ak1T62HI0gs/kczJM3V77J12Q1z+9HaT+fUyVi37T1
GnOhmDm2bYqljiV2gSBjkpcYiag+OtYR8n+CMBAvYn3Oip9F5kWkbBHyLH4rODA1
dedDNitczlZnbC9npdK6JwDYxSB+mdkxUZ/BE21LCEk5oGqGDB7T2E666ZnPLfdp
FjDIYIiqYAKbKIAh4/xUNEY+wUQVTVW8K5P8UBhvtiN8h6XzRIRaLTGA6/N0PDed
QSstzKSjF6u3EVRx2aNVvWHmTyLhWMqtir29BfMGyKH2ctWEwQYmlQhkbryf5fFz
DtHqPR/JMOC4qm1D3d57gtUaymRcnTf4WxmT9fN2tz/6Ec55VPD3wC7jQtgWBdcG
cs5C+ZcDIxbz/vEP3OO9XMpNosKBDGi/pfAhAvkmys4bmmsyaSmpOa1USuzg9zn/
j1GSWsN9sMYVjfqbUi4IYgigqIDU5HVnKnEStL66niWYF1NOsW53oVP1uRdxxMSF
zHB13qlVDJ2uiPlhpm6bOx7rkY4KGvT0KT/XTYrMueQuEh/iFtijHCt3KN2QE8rH
x4O21Jhv0fV4F5EZNockwfGORjAiJd4cg4m/F9gTuk30S/jiF0+mHEfWZnbcOpEb
6rDhZd2yAsflmXzIbuLocoORsLHnzzoTVSfcTLKvGyhkdZMSYI+IhEE5Kdq+3fAw
0Q6uy+TV0XKPM6Vo+U3GsDcV3aDQ4g8ymLenWjOgdQ6edB92O1y8c0KmTopi76Oj
0N4QmLw2hTAQSNy0NJv7/xO9OB8bTn/qyE/3dul2XWxYT+ACqfzGrjh7P1IARA6p
mmDBMYRkaxRrAK9cb8STV4wKGUVQAJYfp8DFD8O7LvLfTmBVRZtVqjqvJwYwA4cd
SO5t2lozncK+uhSp0gIwdSZdsb0Scup9dfA2nuyRIfsKLS59JFBPtghYtH59ZNGy
vDEiWn1aGrzPOOArge7x/rBr7Bu+LYSqoJavhgaTytWi63arLd16gJ7FKHpe64nt
bwrhvAXXk/fiCFkBbTBjtm03z73xB+LE72cZXvbKtWf6AhSmmBZBusHRbRGDotaG
aTKcyQDmkf6RZObNOgU5SC6yf96554IdzNG60am14nsM7Rgt4I5c9HVm3Mceanag
UWim+4XYy8L9zcps8ep0amSxW03pE3cAiJhXLhX8+Eo9+a08EhUQssfF7NFlQDmt
119gedmUVdKht0AkzzIrExvliI2v4kumpRBcvS16cnwftk2+80cpGVgi0HJt8dWN
ToUzMAPlkIgMrm+IR2eVCdkJP64S/EMVttvgRZTzzY7TpglPsXQXMDqAscMZsqmT
NgiMgQlNLvEiHe9rePnrTc8SAdfvMO4KrXQSsm/m3Ts1GQWCzpgh7P/h8bvp3Fzh
5evNAbWu4uPx/5yhF7DdpLfQNBu6OGESp0RV/JEzxyPkdXszNs2AgBIa8DxrixC4
i0LI6OkpNarblcTWYqKH6bxqiuYqX7h51WNu1vr+Q4uq1eDv7Wj2bjW/Ui9rAcWg
sHDv2bf6Dons+BY8gs9p3C1uXCLOp3sbDOW/AM/nhbepiQ/L6WJC0UfauAju3m3w
9VLZXhikGQYxhlCrhLSnYjWOT6u/syaAJvf3SPxmsf6//5PP8cGrpec9afk3vTZu
nn4xEhcQ5OzVxR9YDAaG2zvgSu7HrBGtk0sx5eWd3rVXBK4zfHwOHC74tSpGqo9j
+6OE3lO1DDqnOejO4cLofE7iJPMCNgTWSeRnu3ngB1YbKYyOzm3qW9pOnadvax0s
32D3O/5X2CY18wdExB88cbZVBzrnWDzkZHErANWdkk6MzpB0YieshJKISXvv5rO4
boNooZ/N73Qa7rsswmh69aId8+OH1VP5gWSGD9ZmwXtXZ3h47nC3wRDLhsLiNw3m
L/j5h6mHEPA27meK0EMD2VKCWoEtSbtrQylcI+6KQXaOO3KADVEsJm4lXmwFKQi1
BHpobpkY/wCREwKreB129PYXqJLNQKl+rRuRFiupYh4o2ClTRyEiUS884lqFF3+u
wIvl1tsfnn9P2GVbBIB9I3AYupGMMJrvjtARADNQJeivEfd8R2KM5anKoKg/nmcm
n6laNpoHJAjuO1e34a4ukcW8omzrSDDt8J/OTfnJHkWGuuJMvZjrFFWH4ZgJhnOM
4qCZfVI26VbDr0uyro9kE8lxN4CzUBY7I58osiim6rDxWBrVvICaYZx1Ba7YhRLe
aVTChFlBQcIsV2p/j8K6wPRamu6plncXs6Mv6rLyCY6XwovAZDPqZuI3XP496bTW
qNCPL4WH7ojwYfC/MjAwNwByEfLI1ndB9EQpwoAVe0CCjlHrILlnm/ujbZMaCmcF
LVRbFvfZajBrxOUOhwsaYoX0ObdLvlzeeucYpfLf2MGy9gNkhkn6wIGfB1yVTHcr
4KWABwyYel5RppLzU+DUYdXJ88weVyQLm82Pis/+kgB8+S3Rmf2v0Ug+0GiaEUxv
IHoWASZeeV/oOUUWwCX7TscOXlDTQ+K7+Q3sM3W3jOp92vBLBTdaTW/E1SG4ojOA
+XYz6A8OHIVuzpux6oI6tcHzMNYztCZX1sqlXeiHL+AejhmnLnYxggNDsX/a4Hwa
/c/z681JeaLA5K1hDon/L5vzJa69xEtegRU4jki6vjntF9JYDfrjy3N/1FyMpMsp
HjLrpI8dsPIdYub88q6tCtEd6mXvby3K3Mf61q809yeCHL4ib42s26kkDzkaza2s
Cg9lcquxq/QXR/Do5Y74OCJ3TKcvFUFFBoMQf3eKOu+SucTy37Nnv9mkVA+bGFRb
aw+rPobDCIY2DZ/Pr4n5Fww3ffgMGHBD0fnI9efFg7D2B34VfS6/E2+/o0mw7Shv
L3ieHkbuBXsdm8PrervVY7H8NWCnS6NUkJo+hYizihrQs08FYTEKN/J27Z7R2xma
iCta212a3dtzpK2MPqPKXAo3ghifnLN/OWiwVlMSfqiGkiO2YRmOKLSu7INGYiJO
n8yBhcuOi1/dWlfnPRVvXPpZSo/mVn7XHrnthGBwH/almzfhJEE3boGr/5/GomRZ
5w8Qxs1YE5Db7ImPE/ObuOValX2UWqhFbIDtDP2PRhPeLD0BlJY+ULeAFXmqPNCO
d4Yj1ryGPCUxa0BsenarB4ShTMUsftv23gL/EcjQHNff5Z9VAsnnHnWpTaTYIEoi
kHxAS1zAWgnHIH8jS9EvjgXBaMm7blOBHxy+s+kaG3eqmwwwQRtriBGyyqtr9OaV
UO7DzZSyH2opinzIG2lv4aaB931Z6c7Qb8aqVeKswOLcs3f9nxkgnOQ+HXJkkLBB
EYeDqqZizgtBupwWem0M6A5RhYqrvC39fu/BehKRdCnhknyRjF9voxzAt/VT4MtC
yRF/J6/GyuImg5cBAFNKn8kIrxcCtbf6fk17aNci+EpKpfngDvGLweax+e6yUUes
H9/BSU0v/pv86osGOgL3hFE2DSas+hj2HhW4PB+ukrJVX6wU3PFPU+157qhGRjSY
xfVkVRDxIY1RAvQRo+KP73xWMgLZH2AbkX0iylKGwfdLRBtzORGgnxZrlOdEuM3j
4vMwUIZMtupO09FRnE4HNiO6h5qV8Zx/bXZHf6eP17QiJwPpa8pYe275fwkOO0+Z
n0mVt9gMr5aNRIGcSuYv+8zHDILUc5xeFPb0ZnCJvikh2VNB5aee1PSkjfbvn9cm
11CKCSttsMmnt6L3dAe66e3IPLkgbOS4T5x03CC2aWt/F1iGKmlJdFmDSKHWuArk
ugJuRUVAwlXuizgD1OmCPMUgb15QntKifbz9yDL+yJZSPO7bnl2PDuxqFoBqFwm9
+RibM0i9vA3Ht9xfCEiS7dC4Aid/0bSdYz593DqE+thv20BMgt2QAREB5uYNNELi
8ilfbCydqlt9PeptmS5+XzLY/3YRB2XLhMqCqHyOUJdMCBpy7IcZEaV6xPyI7VS7
44q4HrW+b2G038L6YC5phpS9BR/tsGJfqmRYvuZB0ETMkqRLx9MCCiherF6fWeft
6KaCnaHt2d4hCYXhFIpYIh+mJ0hBj5sHaP8WXaOtqeee8A91bUnLIJLkzCnrSRy5
mmpggskHNXeQ02Vgr9KWBvGdf2QscsBSjeOscWm/hjdPAH1RwE8aCUW6nN0S5vHU
+ikywXrhv4muT1jyD6f4fFBAQwR/hN5INc9zb3speCxCUx9nd3CC6nBNScqz1gx0
7WMz2FArB5oBJ91yghdYoppW0S4xIHwLCtTxcyXgAlmgl+6HvHXtoxeoQEIIgFtY
m0LJaZ/Hl4gdkvJ/H0SAej+AwhckOJWekrkoI3OtkJD7FqEWFqgZEn80x1oHiyjC
Qav6NOncgZY4oDUuoLLOe/yn7nmvtjASSm0jxiuc8axBlWXaHZ186fG91lJSBrGk
0IU0FSJXDqC7mU+oPHR/Undmq4fnU5TpEalqdjZYTE+rqVHY0NXmgulcLN9+7E+g
mQ2i+3cH13TXUEjgBkASP0YNSVtnCqoyW8L2aapBMf00AZYP6WPQGrwDZSUmD46A
B7rLckWUbkKCF13tOH+feXp3D/7hkuLM/zFOyDxKh0yBmepgCF3EMC8icKphS0yu
PjeqUEIsaSWlHc17g4vTIQqhcm/8sS1LtGB/+XguB6OOUc9lrfOYY0Q4POG3pn/Q
L/jnlh1u7E6Eyzj50TKESRdqgxdnZyVhETk7Y9tZdUPA6TfB2AXBzKTROS1HdgcM
shx6Vu5xxFB/iDDJdmcROkjh5EbHWFU0FSJJW1a37VbEsYiTo5KIMBi5TBm5fayE
Yf+YEpZB1r1u4sCK8OGDwHfdUElQEzy5WFxlaS70M3kByXmyHDlBIvO4y9rDr+rC
rAqxwz43CHcVLjynYj+7Lkh+CbqwbuR8Jmmk5m2rNhwgU2E1eT2QjyJvoCv0bP25
MptenME7Vrld83qD2YBQoz7iVUuhkpLmUNj9tdu0FOH8XDZK5hpCI62iYPHTCxuy
WT0P2ZkTXS4IQVFeNL5IZonux8411MX1G7p+suOZ5rIveE1uwkh5zryUdqUO7KlF
FYJ8BlIghSJyowXOrjM3ambOyJIHDkR5tToKZPUQxYDkGNkUDw17IxH5n038Q9cA
2T9k/23u2XLzH+RGK4GNDTu9djvLtHPHqP3up47Mweb8zw4Q8BYs1zpUiuF6FcNN
62KMKOp0pmB7XjJzXQfbYdBxTjAthmMEygDcUjUl0ZfGj4tXB/j1KQ9F1YalNC9w
oN2pBwAUyyrRVtdW3sW4gXJKTPPTpWfxAHyDwt4zTvTDppuRafH3gsMv5hkw8qvz
n46J245mfpLcstP//zVLmyE+QO/JUtOzCH5WNRZgg3j1ALYT9WryBMLHkonWf0hv
77udLzj9/0yigcjW7lhNqwZSbGKXIUSPigDq2AvyuBeBp1JOQOKvTg0RKx3kZN4v
efrWEUwiTVydkBSm1OfSC4KTOPdMTCsjlNKmJ+dvyGGmz9Elqe4QKGQxaSx0qtoi
Nr0xjiOoIyHAo+LGEW9ooZ400gQIazh+1erprrO9Iw8HWENf+SGN8Lz7hWteietN
ztbjSgklgu8YeIHozqQ73ZWzD+kTp1jfpas0nIUtnd89gcu1twTbUgdsVOnfqv/l
p8YUOyH35WnRPPzsZhBZ6QGlf965g7fWzexoAzQOOAreY6N0FFgWwLXi/TYUnfwf
uDSqcWflcJUYFPCJGMbrfHpA7rJDS+oylMpNDhzku5XVX1I3CnPmaswJ2YWB/KCi
F0lrwo4JyT6AfDMdwKZDHaywJb4Gtp8sOdSk35qfEhw8qhLSbHT6F96aZZMBXAn8
2egCg4V8ZzIPifLhTKpXpYcUfYcAqIrLiBRXlqPQWrY62Zl3njN95+Duat7jtG05
LMEd9JNMGAF1uZYCqGnHu3ei78golijEVCjCHUi/9NCTH6mbjJW15Js28HOOyIe4
rNcK10v6NTrb2oA/ySDbAk4MmvevRNrS8L3Avos4BX9yPUgD24Lx22S6Kp4w+dIC
3dhRIkYhu8O3+TblrT9BfGq3T0CAdvDjX9lXlnAGNzS1aUXTXGiFML4sgzCnl6p+
iGF5VGmj8NR4ddWAaevkMNR4KlBSS0KgsKheDjtUNm+bhrY9J+nOIelUIi6E6kp7
yEKURrInlTdSsHAVAGzi+ecQCf2URfCXUMThyUHi3IYsJ4ou12+XsvCbwtkq1kTq
xkA/Je0EjfG8pAizcesXmbw779/Urimuu3kODIeUc2fufFA3nXWLmNVr2lIVZUKi
hnaFi9ls5JNTjupxYyTWsbOpO/OQTDVfCPIeXHH5h1y6QFOOSKf+X+aojMGS0ojk
a4lIyEoWL9q/QU3i97NkT+S3zt3C7vsBILL3ra/E+2f9J1VDtJ5mM08OAiBhSEPs
2nSY4zLaq/N1yzBOdsCdec2g8cAENkndBbPhK109JhFSAp+VfSObWxz0Sx7BxwMS
wGjBhxAagIb4qNGsVyA5w9m+4U35MiKYA8040/MW8KabxQFqw31vRp8r7wjO05hs
XLHzYNFB+fT81Opb/jb8XpvfxFWdSFKjYV6g4sPUA19RjhlzbU8g6W8DoPl80srz
cyrJVG/t/bDu8mjbhIGd+j2LuWS/M8pe5sN9T9xhwVzwRzGTQJFTmjyHhBTTetPW
eUNulC2/Av2pNPW8J7Dug3Y7MGeJbzMa0NRtEfCh2K6FeAJi0t7wxT+BSq85dOuv
EkgsvnRUVpGHZXdSEN43G3psJZaqxPvHKyFrvZIjNeQn+SMrn7Q8Tekv/MAWlORC
9W7Ut0WU+S3GqOAfCKE1RCOBMTGEclS8mGnOkCEr1w3TS7gMO3y3I4zIqJoU5M2q
ffqU2Hq4zz52q2EXrIXAO/k0p1Q5kZXYKvM2VQs77cuO9BkNJsSKUKbbHq1E8Cfz
dj1slb3EIXTZreDISDKQojbVtQmibQGNvmWIhgZ3TYsE4f4JT+fpkqm7qC2D6hkM
spOYzuwXU8CgrFmxPvaxzCPdugZmzkLxgYLJZcs8eKEvTjDUZ/Czj9nkjxfKKqI3
CLCXv8Kf18PDw3PAEn3POHLIiGVDAiXFEEF5cEWqrRoCdasKofSYie5d1akbXlkg
O3k78FVYoN4zdpEVBd331pZqGToS3CvK8nLZwF1u1LQy+Hmp/oO0Nfl03Urbkhyu
4k+zE9QZAhJLrDnBrbPVxihEm7qTGyA5H3NmaR0WA3gPWdI3vOpsOQLCCk26kY2k
AI85RmToJ09dKbjJJQq4BDzP3MF2mNZ5QFmiHl5BWIPw3ZGHcnDqwqXQeXwfNP66
DjJNpNrTJrjQxAXWpR0LANBMdydwm6b4EzccqLbh3e+1GYMXNaiCoZvfmdTivFNj
LLpzgzR5xbnjRv+jHY1xFzOH2k8JoF77Qjp9jpZDu/rmgGXZY+umgPqZNVgS0sNt
v0JozdL6L087ABlqBnUXqv7YROOYQzQzUa4dwFlul1uTUxyB7l3hxgKw7rNqkrYR
2CBLyd4RSrn90bOdPNrt2GknwLeLWmI9KaHPRKP9ocDhPgD33WT9wXpcIHVXSdMM
DlTHfHypoEGh0WAHA3AhxZoJ2jiwFymhTf36WxOU6uKWLN2kLKR51ejBQxHLSu+T
K3INsnlrRsiljf8x106VSG1oE5jQsItakTYAjH2MiXr8gukluTcfTr3loCZwSByX
pRhavxWJXcZ+EbuEi4eXp901qldjhqxl0c6CWbEwcZn9Xzd+Tnt50wNT7rro+EWV
2rpn6NPYh6BQloloIdSyTQT6ZR0EZm4FlhNGISF2wZEcUIEBUTFlINe3KY7mNWTP
jC977MkxS7YcVqUsv2Bd3WiQjWIvV/CqBqXq+kB3wpRHo2EuS6jfwX6qSw+V01dv
2wproPNuOQgrDbdy4zpCHI6tUVHYT2KOVQAT+BipxSchfwXYloi4eoRNngP+T1RA
QlxIms5uoa2Khqtze/ftd4TD/7FIegHyNC/OvlOJNrgyADMxhWDg+V8q+oxAvkt6
UINgu/mVsIAqky1eXl8X90YQZOmymHv1LpwRoI587EcIF02bTMXSypI+VY89f5Ct
aUi7y/uOhtLsXCjYro8hH6oe2BEJRfLUUdw+WKu6elSh9yvNviUWPMaXoLMbyUYv
sNEaq+qzjSF6tazAMXuKiH09idgzi774VkVBjYJrKaeJCFNZ1szBCFnwrvN+PmER
VeRcu8j+EdM+uoguTvIAmgzJijXefoEXiXo0W59p4YryOgL5B9pEEn/DXiHVqsfg
iQQ3n7gcVxmuLHaPmWFB+6WFva1opmCEaMFMNxzBD8FCKHiBTqtzzlV9XZN+57ni
WASBnnahM9qK9CNFbDROpIZz559xhq6BIrCa2JvK9odgMRhcAhDEE1jiFJpQPbX2
SloM9zOpmjo0RJ6NZlzPS6iU4bhDhFY90pMSpJ7UC18+kgG35cKMLk1Lw8+fpxrq
svesXfQ+0y49xQsfv/mO52lAXHOJ4lBt7ksYkp3WZz6ikWhws87Tj6c/pxv50Wik
9JP0hyGqhmhWBEfKxChRzBXNuaCbXjZ1f0fNmxmAeRli9KnVIgsREPkyMbatN5q7
bSNdSZkrSipk7xbABD2pU14QwARc4T9xNwN/vhLinq4yUYHzTXiSVdbpkVHgNzYC
8fng7EtwAku2jyyIM9/lVRx/Kvwvflwclk/lOhx9W2iGxvLlK4h85vzAFJYtA7J6
mW4iluNKgXkQM2ZVHOp3qQnN3sbpK7KSz4mkibrFhtENgfV2uRErA6SFAcbkUaJR
rJ3fbTCPAYaRdle2srlgCMTdUPtQhuh93bprbMmzV8vgU8hyTjJF9o1vOah0ut9b
IyHl/XRRXBUIlaocjmd72l9wKxb5G/BKXnoDXq9Vcl+DAgaOOpgrt3G+JkBMIdcc
Egnivc+U6zLYgPC1WUfCgeHMGp1KrjOZnhWscFCkezWGhpuqNf3mlpaRVXf1yuXP
IFiIAo8+LUUHfbjrhRQ6cinVNMezSE/YGyLMVZ52MTL3nXFIKwxJDMyi0FL9VpRG
U/bXSjSD9H4nOCNOI79BLnbJliMZGxinIqhZkBCeDivrgHGiW/29iIGcOz8Y4VMF
Me9gy3ihWiLA7A/ofFvNju9TgueBuJWqMC3pbAa7GkjI7wSpwKLO87gwDjGy4Fgk
rzono4FK2ZztkCcJW+ynTPf37hx2hIi15gWl2sjS2t5krvu4tVODMmGb9QZOKWLK
Nc6kf1Xg9DmroQr59LGUT6Ci8z0LuEMtiexF1xV+gjTbRXwKxf4yVissfh7zCJxd
zZXpKXYwyww6E5M5Drv+L65MhL/yVnz0zEPWb7iHjHA6YlV2daViNpE50qEZTjz+
jHACavJPsCbyBXWPmEltKKy1DYblcFQmlFiq643CGTL8nyp8jtUFPL4afe0swune
PTmmdEitKe8kqoPaLzYkma0SHOCM1h17ypTU1hRW1YVs3xXoX4GS9I0q++agx+6D
xvcTYw9BaQ78oG98Q7BVWw4MmirrnGVp0hNaKcNEaFw6XyJ2eyx4f8QV+YYJexzO
syGWyX0At9hXjKsGpga9IcLVSUWJ85fJKWjy01MhQyACIK4CQPwsnr4D05Ni0PWX
NVfkUZx0jpxdBtiFRnplt86y6yFjctoy95Ht8F7NNC8789cB6UY3ymKV+DrvUXai
b3aksqw3nQl+Gu7ucU47eMwDnyW1dHqM8cqObzmZFW/PNmTdlPTlbZ2A2+gObqZU
FSMyh5/5g1h8gjcSjoSzNSZH1U80+7gNhxGt29NVciHwc4SdumMkNBFW5ftN8kHj
fUDwOYWrFqn01JY6oLwmo5alA11G32F++R0oVIVxgPggMBeRYbVaV7y3DOsD0LZM
PvE3I3wtM1B6sfVHILx7HrEKhnzu5qRckKBigiENzV8KvEVOgiy3pxVaX72AMv2H
SeXgz4sab3QjJeiKwiU3W4FDx+gZXgCz8BQe4bmscsLQhxc+UG1RRMsjxmLJRGzC
hePv5ZZ4sm7Qm/tQodaYNbjnV/a9PTpQeOlxk/joGR8NeyyUk5+zTkhLD+NxBkTI
nifOobA92zUOkfLB5A/z4MBNiblPjYh976H8dcSwhIipt1hLs/bzCaysvizUcIHW
haxE+26R8+NApzB5DK/CpwGaFZY4gqbDp77js1taoZnK1pbBZzE6AfULtl7A0xat
R7OeY+lUpgb6JZivljIyI1YzSuf+mbLRDv0fIkTaIVXuvTMsXM4wCdyJRYbakOAo
pJ6aotPtJpxRn5DcZ1G0G03AlzXJjhajC7MUI/PLoeaEYJWMXN/XPuMzPPaVmu0T
EWTD6NBZj9tKUtIOucXdZIPKYfGjy945Fg7s5FNJouezigQZ21CPq23d41P67LQ5
zYXu90Uy3mnE1N8BewIkZWgWi0XnoApdy5GC4O0i+bQ19yefC4nyrv7LGdFijhoX
bZLsSVEqXPNXYTh44hZssSLEL0w78PPyPMPeSnAGrLnkHL6uv8MHzNvz/yp3pexQ
+yYPfINP9gDkJiYYP2TOxJ6g/Dc/pis0Rr/kSh8t+/Jcv+JlPauZnPQuw5VjysJT
T0fRVslV2eD7Rie8ir0MO69RMT905Xa3Qtcdm/qGy70wMvViJ08XAEiZWCQ1PTKf
LO8kvq4QjJIwzgG7FnfZvlWKhdPXnYMgbAH+6QJmA3PDB1wb0gt21otosUn27UzG
hrZJMCNPKYJUrHdKshHQJhIaF3poRVINWg5hh+cSlWiPtyFp69lVGz1PNMh7E7FB
JVd6En5Hk+fl7OPI7Dldha/6ynS5974bI0FD8A1WQY5zhed6pEWcRNDjZsZUCUCz
HZhAMz7jdi3mqUmCkLa87R0i4rxhGoYLTQlCzMBrL5yLU2JqGqAWvzzUhAEhGwHk
WVDJigp0Br0f4s2j1WXhE+xaHhuIfL00llqZexxNVztBk5w0zFCWTAsDC5jSsA5F
Sp9iWvN4ZDdUsy+KvKycjEWdPcX0ws8AQg1KAKXhmdPK7bPswei6VGU3rYeB5AVL
6geKqVjrdjN3TGxz4hCa+I7jfKdC7P/J0+Qs9QVCCZ8s0njznsouIumsRST3VVbx
QLIfaWYhbXb7O9jwrIovqu4yiDpK8Qbq0PVAuuIaXw0Ec0+5ee9e1pwD80vJp9aO
DXGNNNMEaS48Tc+rIO85cs3rYjYUYp7pH0CgW5ZY2stxmmgL1f0S8jYG6rtVla+Q
j6/ftWd88cNjFr15vwI6XENvCd3LhTSsrNj8tf4TwWx78Xr/3VpKoZ6+yjUkWgiZ
F4LZArcrk03VRC0vVBJ1CNc+8qSl/trnMS5QLjf5sjAbK5RkQTplxMBkSF/Ll5Sm
pmRAHJo7oM7Q4D2Fy/1XzZj/Qzlii21wsfcaeem9gFRsLw1XJ9KGxSVvHTWE9IuI
tcPuqihEkNdalmXzWQLTBxlzrVexc32RsFXkRD81zNDz5RALuft2rOtomQicOQad
xguoqaQpcAssjVeWKUT/RkycoBD2HUVLeNynGe+Tx6MsnD9gXA7RkGS3OA68Nom3
Tk9yE4oRkeSKvVEKiAIi6/LNW0Dr8vr+ewSFOxb4tIu7HlckakLxLire09BtjYhT
qqj8lHKb8ehWe0YOKtCL0LqPWv6OYnR5lyCjod8Cyii6ay+RMjorIYsBN/SuVITN
IuNZbhUNGwVXyhpQl8aCYYgn54RZhFm2qeqFLlXJl5XhNo3DC67TE01MLMeJwQx9
0wXVEQCkzxt1ODwBmyDlzLjavX55g5djkjUE7HFn8efGWir84xFmtJFQFARg3Doo
fLcbqfg4CWTwm05ZktauXoGM+xbKS3WUvr7GSzN+YidQXk4DnvS03iIzC7ulz2nD
kxIiJRpAQuSmvlBhfTSzW833eqnQtVPhFOnKdysxy/tGrEndDBgR4LP8l2u+QaAR
gY2W9CotQiwBMp2ZZluToX6oU+9is8AWlm1B6/RVXB11vvd6vy7Lmu2LMtMRAsoD
x1HmSdQn90MtEge2Yi9ycl8bCeQ1E9ZgNd/T2aIOI0Cx5Ue5FE2LF3s25SpJQDt8
EEAwoDcQXa3vGLaRORx5RyrwvgUGwcjwXgP8Z5fus7DX4dawSYa0/MaGOaJWlCQy
sBduLJTT+/NZmnsZQrh9ewlvqimI34SnmQzCHWa7zcqgFiwHQ5iRnOuv98/fM6c0
qvOnxEjCH6rt8zxN5VEhn5po2Dm+lQ0con4GtGn1/xcRMWJJQkr/d1S3dj4//y6B
UYczBOR5EFgP6eTCxZ4wOw02Q0AzHPC2g2Xs2zFj/BAN9Du70aCI9xPXDnxhGsvr
A35xBly1UdfljgZzrNDOof8kYTiW2B6ECbSGV/yXdPoKpgtqajY9K+2kZwt2PL11
q0kkZ3/zKku60+jv7UtlgLQHZqJbHgw0KBc1hk3kVeEAz4A1NLbLMRH1mLsL/OFL
/8Dwp6xDF+CslcKvT/+yez9iLiDCV/q/5EUljV/LTux7OTOflAfbXRpj6gcZ9TRZ
mNacnlQ/a66839YJYq6zhWxbo1Pkt0k+5uWGCUDtJbgpOxDZMi7sQD2agiIGveh1
VCo51TiZgm+hKIea7gXMcC4mgSZzkYjmo+UFq2dst7IntbyfXG3pfvxdO4PeLVVq
Kg3QrbWkugNdEE4/uLDe0X5350iFi715pfCc4dSVmDODj61pguOqV2AkwRrFGd/y
ISOCarKwHmTJh/yIenzGvt77bmyYvEAnfQVoM2yHrExHGVk8objXOCHUpXdbW5hl
dQ0hWZpoGqqgq/oLArYoYEABoju/7cShIWFRn8ZO9/qNzkyTe6nKjtJZNeNYsqk1
uvBITdQpBQc3x+bIz1gDEYc8AgAdqH3zvlj5X7GNUQpVdBOBZp2o9lrntv07yDof
w/+7wIGvKooDP6T4SJDSAbKrSxsstMkg4kwOKijj5bcc3ztiqN3IdN8yITJij+Eb
1tKd1xV6EcfFpE5kLXNpu1rglRKUEvj0/fmdbor2Sv19nnCe+DaBk1bsCAAXQmMC
gB4RoPk/RnwMkvOEJSU5HG1XZc20NVLOTVZjJX+m1Ui/ZSIjaJH7Fha9h9uOptNF
qqRtHm70axvPPFxhYIsiKgwSHssA7SDgoHsi/xk9zGkBoeoWPcmShUn7ekUmNUop
mfxML8iNHHNO9aahS81V+uLypRUBgdrLs7fgy7f5S/52FjcW49IsAL4HcTxCBn52
2z2cLX2pbku8ruu4hE9p4q32PKdlTPctNxXI1vRRJwXISlvvPVkdgpn7/HJ7E8PY
1gh4HB3cfUVEp9pevjyJ1W9+NpbTIe9/vixHWqsHUowVSGN38Ag37B+j/M/dv3TZ
H6gr3PhY4xKfUGsoQT7wkmx0DEIEnHmFl/CMpjeVadN+6nVELp/ha5AHwGE/6gxs
YnPoiWtN3sCQUzpjEgguaAeHOSC52KrRELWi9QZL6ixxCuELv9No27AnhhsvUvSG
JCQcqRPO1oxeSZtsebieIj+LQRHnFEra7LF9X9ArLyQuUaEHYTHodsItSaAKCa/I
+gXaav4870UDV7suF5C1+SCaROHSJgrz87arFddB1ol0tva8bLAwfaIeHIbMi9GV
S2PhcACLBvechpdbbPh/bbbU+7cjzkenfjNPmIyeok5oP3SXnEFQGlBCrL+tX2iu
tDSflZXLkjo9shErPBvp/3052OOmPnE1bbg+tCtY+UzrRQC1N79QcBrZSJeuIk7K
jCG7EKgpf7B+AX7E8bnANhfUyfxTu32A3uoRLVgRFQiax8AlksNmHwC3V6LnbfHB
Rd6bB7nzCZAzVYwWFg4BXws0u0RYac4bNmLV4A85ujXidDL6Nd9wPk+uwfYIYMRb
I05mX8wRlvUK31GmzqmEXtDgAwaaLpL7pH24bTnp+efjXS2cuGR+TDga6RhRomi6
54ZQiqMyQrgbeGMwqJt36U+F5rkUKxgpX42rRXIoL59iS/46IvpczO8U6BeqSiIx
qdpaeZVY+g8QvfItt7U/H9oiiKnoPotpjCt+ql6Nb398zhr4yTkw2Yb8BhtjI4b0
DeJh/Ey2yMJ2muL4GXL1yzVj2WeA9rlFW4h1PrfGrfwFVrysWzDvwbmx22Dq3cWS
B0klASKMcurRnN0unafd2kJ/X+xEfb7QX6IanfqXxlvkWkXXVL132/B9WF3vR39R
P+A9dlS4cE43u7u5qrmRq37itsf6ZArglrESmKkmyy8KM1k5EH9cCnRmspk3++Ru
elKW3z831WQWLCAptrqivd3AZWvQSV/tter2wUcnsXXJFBmaCwqivZGsPMxQ9G2k
P3MZ26q/ifXcn3V8kMBOQYfhV1fzg4Mb4/xCAdWlSU6ynR7U6RLV8onkZ3w37lJk
xWpq0MiCn0b/h197MiFXeLcPA/t2aOm62JS+DqgO7n4KMWr90K3H83T/Vc0lShji
DV7R4wDy9LJh9wv/zyPauMZuyTi1AJJpDNnp/gAxwWYTdyhnukY2Uwi0JI0i3iap
GQlaUbTSRW8tsTuCU4AKPeR1RY/P6V2/gHAh3CZ2I4KUtijVBnOKKI74R81fABxt
+doy4Jv8aRdbDMcClnvt0K+Ezo3upmTsNCN5iEjBVTEUWkT7A5zRsW3IyPtCph0z
XBwgPggLiQ/M2y99kc50cZqDfzrCCf+9zFGTAol3vyO2dSzMVhisjWsdc/nAARnl
TDkkEshmSuVMDbTNs3I77ywmn/cp8ag+8afulCo9z1T8gwOJ5JwuLKIGXJTW4T6l
CYrPNYBA7TO7uz4+bdvGFaAyV9TaR8+OuW8D0Q8n48ysCAH6T+vBFwF/w77x2w6n
L+hDfY/yrRBSCZT5IY31Cqh9kNUwj2Ncw7y2rIE8eMsma/QS2+DqgIRsWGUysN0d
UqH1Y7nUIX6ePGouCqaFeyRoOPYpcNmYkCl3gE5lNh9MF4SlS484xUv+clglYiLq
6Lujy0JiHDjlKxUNF21R8YTydclcOHSeZI4s+mp4FD3tph7jO51tPrPptxH3OwUr
GCYjOlfKZNFnkAlJd0uxeh7baqyGTfPnZWGtCHLq7FjEJOWaKcaN5oHrpHwpx8h6
f2TEeJvSItxTaFK57aokJEVWzD6iZ52skOxZPlcSrU9EVUjJxhjl1HmJpRQrEOGf
oTveyi9zvEA/0VzyZnDKxgjSUswehKBGOMg8VVQE/A7yLbMplRtCyDCim2ivc1vu
s+/nEgQYOdOWjJ+OnhY01oJE6j3J8F57vqiPagMVe0W5fLLlJnCYOsKn2HMdOWys
UrIP/cbjBjUs1XiyEA+14Z7G8eLT/UHqpg9Fjzjdo5g1EV71U4uO+6Tzv6wCuRR4
sZvg01WebViM/57N+0oD4VAg2SwCcahSF9zFM1ulCw+rC2x1iFbCloDlEu+0WtLA
5S1JjlwITYgGTobz6Xb5tqmLCSPx3u9tdT1ZdZZJFIEhbE+RTWrUmZf5YO6Jm4Zt
dcf6+xvZdKNFOEMqr7TwEIIpXvg8wSLq0CasPZInbdcjK/zy0jjzTTVcQGq6ucFo
sx1+csTUfJmwtDgabPTswHkHZ2pveXoiMRlIWnX91z5rVp88q9l3RGqiWWpcyV3Q
I91MSk1f4heWXZ2wjjzj7gUh37hEjiiBIgtXt7J9UzOVLvEnymmM1V6lzConPJWC
bJCo3FdtSZEyFkHCH5diAf18nhq3x+9FjfguzMD2HNKkDUNYuKtRB7tvTfgfo5kj
lFo3DlBST59/ePUe7jVTFNJ4KeCCkubri7SIbM5YMIDVauF14bv+Z/znWrrate+j
kBmCLf24K7nbUnKMF6Gw4s6iysUnLtIUBDfYtkkT3KDyTYryktEGvcXxYceUUTH8
at1mTw+hv3GqlWqBJmWpKlKIAJed4Y+IzGXmxusRBiu2l5YfzQmhvbRvV3iu9cDy
hMqXxhwh2DF3+tVZxyeKRkG+0BSclirSB+amzSlMwRJThp45WcLAY8OaxT3L0iYz
xvnggp2cm0p0mHeuukczEFWhva4Rjp0eDEY0BTVd5SIbgurzScaTbnfcAkElYuLo
nL22V2pJTct9rDFEbl5+ciZlnox1nSsZu7AqkdftIfj2p2QRNZ4S6vQ+UzHdd92p
Xty1lxsNEY7oIcMGX9BjUgMiQFzqjURwPak6RAnrox9SadqGj5WnshqdF1op4CIr
jDtNMfgqTnkkD4YxBry0pFkTkrm5y1wR0QXSc/V4Qgi1eMXkhwa5OY6A2/G0tSuw
XGm/s1L1kDZKyOTvGTqSMLRcMtgrTCblr9z0L6IyYSugyl8bdhxGWo6Dvwnj47AS
tXv0ZgqrofEDiqRuMBDBRt77cBFVuXVKEu1K/fBIRJq8Ii1um7KtE70m/iCSgL4S
hcX3D338rX5qqhbLU11brU4wXWxGdSJDonIgpEuEKk/ZysUPXonF38lnlFXwyn/I
M9CA0r/VEurkncn8l3ySfg30SnbL1IkmzyJIqWBxWyZ0BaEvoczQLsprVQulaasZ
uRD/7Kh8GsXjyaBTs5cJEldnOf6Kbu6VVSI1+dK5YFP1akB7RZ2hr1miyYlFBMKj
53Y6XgpcA5jJ63on6IgXyZvypQ5TJLl4RPC3xm0YQNRHTJc0ID2tCsJ6gltmIspY
jg37Nyw5Xp5vC92PcNfXUb6gZlCGl1Iz6fdeIpMFfDBHI/mtRDPVZkFnzz7wW6RG
r8pI4udgCRBFeGtoLD7aUj2BdrCG1eduOEXqx/bbLrr1oxCHzh+YkqAfHzXwyU+b
ilXaVrx6HnDCCqzOFDhLUEA3IlUoYahlW0KFqJAkYakZdxHZyecL0FlcMGVi1J3y
X6MmDyfDs3p1CGJApnYXPJQejCnR6v12P4xNntdG1oiETH7HZ84C7eOf0nlcZouv
mis6FxbezcI+P+EfYpokuLxZz3sjCc1l8dMDwHzUiES1N1+b1U/MHlJZZipMULrf
1mNhv/YTuMYAPGhuHqkESzI6mHoCf2It1o9OpbrmtUSaFfRU/FzxgnowxOdj3/Rr
FhqcHHcnuVCc0+Dul5/IM8BhsQoZnofOG/XFOjqDNyhM1AhluIGOXmJloTXJyt0x
x6KfCe8qczZ9s+opi4Z26xgt/hm/rU9AAjJW/42Ach/OKUVEiDqFsQobVL0BBa2L
zALcaiFhYU+RWDPMOMFDbIsljnyRa+BT4ORK8ZsLo7yDr8xgAdABSam1CvkLkMoo
PpHCym10D3PGLcp1s6VBluiq4W9xvIjh1XOK+3t2OXNmVYylaj0arnOpfY4nps2m
Vt2vvZHwRajgLgfcgteIJyDOqt1JM7eGKnxa8ALPq3F/5yCOznxxMCNmMT5xnDLF
1wZv/9tv572ysVFGUf0kDbMOCw8VzJMZzxjLpQKRCsS4brd7BnT5wkBdXynzfR+G
VmPiSSTK7pLqhb480ajie1ertClTikMPSSH4b2bqWiWBEM+SwjIbBoxY+remKddH
TSkCxjOPd2AZXtOYGKYz7I+GRhDmliiKBEDnD+F8XMHfOyigf7ks1M30ULYzCc4k
H+fWy//kexhcmhonvYxKs6euvDQcLzlpeYMAFF0MjaZKoV1C1i7aK/b8elTSUnaK
MndMEK7agoWklyg1/TOM/qp0d2mLvgzNwsap6f3hUvDTHgMrPvFEdS9ee1sC2zin
8AtGNrTJ/A2rEkLIFo04vhL0YkrjCWwPMMj3meQJ5Ykp9HYCtxfA0A9WVmHjsft8
mj+aRMGG2SE3HmsIPZA28VE7f/DD4JqIK3l0KiymtcEoLkWm7MMjvBs++u3X21UP
a0JTiT0qXbz8swdyHlBKCG/djkx8kSEbI2vuL3wcNsjmwp4m24inaITieI/uZRpJ
95PnGLQk9MYv5WZcdXvFaa2JlfM4WIFvQ9Vhd3/oy8cIKMCw/gj9Zuhzg4CmNBiW
OYq3UH/bGCYYMMMr5OTlf4J52qXEug1SylsPt9oM/1IS32aCu4TRQRXzGQGuPV2B
O3zZ5/E+SmXcA/PotgjGq91yo81r0Xymh8hkVsmOw0+Pb2nWzg50pGua/t2thfVL
STXVmS/ue8Wf5XU3eVUOqHS1BnmEHbEIhsUMSQAnHsrK0P9ZDzNBQV0UQtObuTK1
F7LpYNwfb5D3Bjuxqf+fNE6dPiEsfGoCxo1cHKcdEgNQK9EruF/42Z4Hdynx7qax
XvO/FIoU0C8uKs21YmsktyZP9auVLgy8T+zg9LDan5xiWBJ2Lv3He9hs8wOzPd9R
EjdJdiBEHo4604of3A0zM66otZsct/+0/rcPQF1G4mfHxXs6jvkdscOQPUArtR6q
98HV6SguUejAX58Quyz3yIRSpg+ObJBNQ3BH3ZE1y6fb2jC1Kd5DX04g4ofmu5XA
9erlDsTjqTn6mKq6Hm0cTPC6bGbOMq0R++HdSYiAQ+6o/KgDp1H7lnnN5g7hb6Uu
/iPGTWhB4buMk0HdE+JRh2ZCzuy1UE3zoLYpf75RJDu63A8BSKiojWjPqHHJIY0Q
oVnISD9ITfa9Oz/Gxo3I1x+g7tOTdOAElF9nPi+7dFGMyFZi6THZHjgsQxJRgawg
FABDtU1oK2RL9SVVPt5PeKMoXpuk/Vref6FDPlAtGeVdDnfa/rTXo7CQO1dx/b78
A3HzQBUDYlf6SxARxPcFAC8ikKokjJAHQovAvtqgLQ0env0PQXeOCMLPPxRK8cgw
TcKsXiq3j4KNLCAopgpMskX5V5G6iXU6rzA81bm2q4mrcKvnNWg6a4yKnC3sF23l
J4lLQiZ/om513FmQK58JK68DFT/NECnfOU/AV2XquQduimPxE9HzPdu7vOcQdwz/
07++8y4A7gSgMWM0W3kd/dTKjXlk1NopAHsyLMRuQBfoLUnmgPrYTBQBGXezrdRo
mMmPqPgfJlxhj3jWb/m9TWjSG+U7CPyvt4jvjd29od8vLcVIqlE9RHr6lBFxlAOv
yRaSwVodLL9vU1hFS/JHTynxPFfWrzK+NZteVS6RqRY9blwz+4IJ51cbYOe91lPR
BqFMINzvj6gFBWROFhAHmpAYWmx0u+f9b18ZzkiUuXbUVPLc3xaB5kYSZ3sFejIw
nPCCRfvr3i0TQBvuaBxbGUGQ22TPBlIQhkFs94Y0AO/7/2yZxvSDSOZIaBqLXdvX
DQ+Cn6TOZNurM5BjVBcin4lXmQLWwYlVjy7SILupnKZ+SjdHLvY//8ZrAyzbsLrY
R3dwJa4Dgi5jbFgxPHjxnY8i3tdHuE6UR8WDmrU6MY4sD8hkBhaKfgTLlFny3WFu
ktONZ00n5Li3yWNJjwjQWSGz+/phllhqsuS43ZNydNbN8jCLBMyf3KwvXAhgJmoI
aOaCB/ru/n+MR9tXssxUcGARj4Zv/BIGX7puPMm5vnvgkspe8zMdlCYLoB6rwjUP
c5z0Jk2X11uNkuH0+BXodj3ibu2eEjgi0yefguPJfjQEyMN2QNm+7d+l3EX/uy+3
2wCLOSclebpLbdfekPsJbCrlU6kHdRoecfBXAt2P2FKj43//6Xs4Lin1nUxonmH2
rR3+zKRfGdwK1ifBxVn8/uuBgX5w1XCiUEMCbpGy52VlSj1kEqkTWoniSrnrPyLo
1IIr4oxi4Hr8WvyFecZIUBoQdp3jnzO79wmhjixT66WziWv5EwS0G0tMwgpuEHBq
c9/uzzCPy4sd/7oYRb/+E3dMncJXVulr5PRqY5pnZ/nyIGZ1GZ5DvIslPTmsp6uJ
u0gblxhOIHVxd+n8E0Xku+Y136Ws0x3JFYb1P4DQlnBOPmGflvxCp0SHF1fYZC4F
ir9Z/NZZ49IpINR/tvar8xdMsDE0GQryHpOF0ApHLZt0vTdTGsSqxjYJQ9NPW3/7
qOQ/qhX5H3qe/6ViRV/9N1LCPrjklPryaWuuWOUpx8gGeszM9LsZNqqVJx3KqHuC
ZsNQQsokFpZachCmJ9C9HDc4Kc74dhuwWDkL2J+H4x44Sbor27GLRZ//Lu9MqSlL
xkciW44tMPVz6cpeD82KywGcHo1KWzVvlwWGAJKqZ34YULvsdfgDYu/zaHsXP1Ij
24E27PzXTmRLrw0IYCyrzjYpj4lnuDu8sFJxxiwl9wC4Aa3Hl+qOT4aRhF/8C6bL
9tN+KwurqtF12lU+ujz0+VPdn7kfgkr2ie0LIlo8tQC2IeFrBbpvZiECc0llEg0j
pOvGCzR+Ls2o1m5puPAGPOpd//Sc342UwVqI2xic5GqEkqRBo7tQEIa2WIBm0JuS
U3TuRmhp9WCIf2hhBQxs6boF3TATps3KyKGIC3PzQ0tLOqb0QInj90NNBO3jdJ3C
43PdKDDhd2np6nqeeGA7fqnHngO1AENqdvLDGdre8SLWHEdTZhD6t6lGwfyhHsWz
a+fC8+rNn6R1e3ceBo6UWj63fYnIXi3r8efgf/z6bnLAIuC6UZsOycvSpziGZ4ip
8Bj0ySFfR45M1DNYh6R8Q519JCtCDBRM2xdIrQdiTPNlEsXUkKGMB0mE+7INbP0Y
HnIOoPxrz8tUQtsPakDcqYD1aZODX3r7A1UkvGDDSNLDUsmGQaOG/z/zGWXp8h5M
pXBAbBeMPHS52E3/U3yHFRmldHe7BBDEZQsXiLsUt4DKlkLAk9ZjwqawOUBHHdW+
m197FX6+tLTbQRTe8VLUHfqNu32QLPgVsocFegcD+EqlTq9bxaYNexn6KvVg7Qyc
NkX2Y3RQkY7RRdVD5Ry1d45caxeDJN5gTyy0ttEnRe+gvmOHgpTrcG52ToO/TmTK
f41I6nbyWv8dPT6Jubu6/cRpLJGCAqoG6C4gIT2Ld+3VlAF/yAWMnbPuNHezZSZV
h7B7LbriSvfQ3cbtKnTblttaYymUdvH0YdxSjDkPVymYIexlqV7Ceh9ezOLLTND2
Fa8EqQ5KD+uAGjsMB0WIC5/Fpe6LPpwn1swag0IO/L9pGyOXsQeSWfB+vvHBR5Po
3+csDyChJnTvamu4GZ0orFn/RUt+rggGlIQ8jAbcvfVWUh80na1oJm0Pm0nAXIaO
NZpvMERGGcyTtMRmuepMD6ylHUI8JAIYyN2r8DrBiODx38VysA7zllgDWoQZMBp7
s1rwNTkF64izZjDzmzo+gdmrHp/54YPvpuhFoAywDWmXtaq7io1rtyzG3g2uEknM
PB2AqEPEFnEa9mgAqqkNAuK0v5QL0DYaGaFDqux32pgnHp+r6KELxNV2Bu6MvOK6
FvE8An0wYJt69v/dPjUyUJTiC0xhJ5+5yR0KJYAMs2B30j+cJ2c3xJmQRinl9M3z
ti/Bbb8VcePXp9yUczxkZRqqgXrC0o6/SaZAxOgz1GQeHSBZons9/Rhnm/kQUk97
m5S1yQBmQ4m16kL22flnZJ97FBxIgZleuBzNyp0pqrdPF1rlkawB+EQphd66MRHC
OdWRmibHlvn5XM0h/23TJk+B+DtVKtGkSmWd5/FDrfm4eUr/L5rLP4e2qBsvlctl
lx7LYpgUTFnHqFAGOeXXydvb7G+DhgfL2N2MvfFOkDC9KKBITM7rqG/9JBo+2+3+
/3td6w7AWzJ0WYaKxZrDmwxRy7jWVYPF+/BwZ8rxwEHqgUjcp15g7+1q48mbB74y
ZJ9tVqEofUZrWIMZXvqLfyasl0aNyBCat9nFGbsKkpvH17e67oBPF8wUJJazf26T
b3MLRBepSd38JQb1rga5uWnuaE+myglPNM8Jezte/akQ/McHyDR5v3xVpVVgCV5L
7SMX83cc1Py1VLshNTtQCpMSrtpu/zyGoNd9eD8xgscPTd40eQMvWDYoDdrFe17i
JI0oPgVTO5ffJhOnTESZ/FAy5W6xQPN9dtRMJ+jud5BmtmbjHC6/OAevX+hlfWVg
Cns1/w+L9gxSH7m5Nsb9gAfHesBwYh2WmB5cf+n2uG37dhy4lIT4vEEKUI0PlN2G
YCdaENnEGOx36u3DvBhD4oVglKJ1jEzg32az8EApmM8OJBm0YJ1dCk8UdRNBKD8g
Jrb9wRsbRC/MtN1MCSOzTdkgh02i2kRiP/jnHEiHkzU3/DjIhbiiU3UtYWWHKLDz
fxV9xiaq/pPb8r9uW4ExfRSD8KP2upPdRA6n4OwCTztrr6T2XNXHySbCPDTFm2Xo
CCm7ZJmnqrHQNrMdWEoKwGI8FKyGcNruBZxH9Ad8w63jDmyhPnT0hzRUBNGC1Nyw
Q9aiN+GGeSua8WkKtLQhOZp3PsC6ilutalQvDSInLER/hQQmhQ4HWuwXtW5wFfOo
pkrR7Tj4H9/KWN9iGNk38KjqWjj9iGTcvQ/9ZiStAoMdnlaHPD5t0Md9ip4oBjPw
F05AogBl+qwFfaIFydlpczDiZMWhoYKnKaUwJuhw1AWblbU7qpxd2rQ6UdltCdUz
5i5QmcnNhVAJ91FZTJ8zK7zKyI5Oxn6JlvWE2TgymPIeoj8RlyEb05VGUhESgqxq
VJWPcun6q0x1jL5EbskYBOcbkbiewFhF9AWuweaF78cK+/XPq0Q+2ws6IqOqPH0P
MEVtfp4B2uiCTvez3T31dwKpdxnOWwb76tyPOJWtU3wyxujHB7hfZSwDZn4T2VyF
YnQD0WCKVvEa+pvkm21tZ/ZlwDUOoVn+ueEMwMfoy4qust90LURHYxRX1PF0inCN
JWSHl7G9DfiptGN/DeJNdM+eBG+4CXAPTZEpaxwTK4ECck31OjE+q2gJ6hsvlrMz
O6gKm8Owvj+dC83u8wY8krWJ/afhRiXwEslyBsuw8jC/FSJpKdEA6x4yXqxcDO/v
7eO83ULHTUs1seZHK5iYfjNcfCAYYOMU2o/+q4Yck3hKhAvaS7tVYPQjJzZGrGq7
ebWfH5SH5hqmv1RUXZuUHW73eM4aUvWndCCJhu7jNc+S6gassr9HUgdJFO0Z35oJ
m9NAD8u+TAVWSOJ3BznA1EOCyXmx2aEaK8ZnP62Si2sityjD+i3DsFzLZc+5vvoa
4p/JUyRVTIoQ6TclNdyx7FguHWuxGs9cBTh2UqOK1PSZRv9ctLqlpRL0BKVGp30W
5O9G4wFU7t0OfQZ9eGoO9rvm9l/UzQDVt0DhN7pFekgyAzbGcAa/zFgpiDUu6I1z
H4yJAGJjsJrJ9ZTar/tMggPqpleClzXWhgEDTecexlhhaZp5t9MeAEDste2vILCE
KJizp1EUIitw6wucMi+WVs1gIlqmnEbR+h9qA9RxeRePMPfQCqhYAhavpAwmztfr
bsJwzKucaFhYYUdBTMa/QRlDc8z8ZIplsCqRgmHDbLX1TTI4x2kQ4ow88BlVNcEy
l2ZV1uHxuu4y52KQuN1tD62FV1/eBe7ksZJY/6fiHky5InMgwnMebG54K9giPa+a
2toxgYtkCBgEOegLnbtBBgg7cLso3Vbq29dAHfX3GUQN7LLiq/ost6yryx+AAH02
IuefaZ2jlCWNKhh/dGQmvErYop2TB2DgdUc0w1Iyk8aj5tkRm6OYNVw6sk387wp1
KztPQtmnTzUeobOqY27DgaZ4hpfp2U2BnAONUWYB5z+q1L5tIbLyAKPAFIQfjt/y
uyDUvKs2xobael11XS+LT9PUERtIJuZKNvv4VklqS8bLlr9H3yjfPrqXnVdiOSo0
k/sYdr/fPJNIv4YUfKV5RboV4WjURJUTaJkbYZMmdCy7inxGV/38WtZB9Wv/N55/
9k+n5Oqj9ZDcS0Ln2zGB2EsnpRvOOs27jN6h5m55shLdVszHPp9FjD3nc21dAFlN
t0ivW/D64j2sunnlrT8j6z920pNae0Dns0iGxfUjyunWsNaj/XHo7EcMXA9z8Kf8
rr2K3feRdYd2CTYxDAq0ACkqLefCfzuNHN9aF+UtAxzGfC8bZEk7e2lPaBAg9yi4
2HuA42TLXGqFF+cJC6fjlDxwBQZQjHUtAdrvezRPgHWrPA+JjD0FTTSJZkMYRVh/
pGHCjGDAmNazsQgIP3ZbWwy9qP+JBFaZGWNGDX3HY0Dxs+eTBzjoGmsX8pOQ9F8j
NQZ5Bj+2F790CEHRtVDMjcl+eNUshSLYdfZmtqi/JPQl8lEklwbixIxNzR2Eafyn
1VWbAEopwWf5umZ+5rLnoifrAKkSnlyAm2cQzaxXOGmcFBL1bYhgd/sw789ZbhH/
2HPC2pK5PLvezNGx6RgEk8H4sXr4eSkjoMsob5JkL9tyLkKs/T9WiSladLaKzu8d
aGmS/3sb0suBdan7SYyjhkAWnTZpMihQpPel0zLKHG3gbqRD5Y8VOmHVKTfG5BbZ
QJcjPYMZaW1hCnnR7gNt8hCEnVfW3fQaIHVnMZbnpgTpPWKKbb/FlS0vH8CBHbsz
E3qBMHqCw0qH+zAtcV4Tu+QAjzASx+NjhGOuB6cxwrcde4vAywISto/Q4oeLPF1o
UBH9LS+xbFzDZcv2L9afCEHjcEml9xEBfHrXRlrMzLNMJNbOOAvLiFTIEPCcN0LQ
s9xHfVwnRjCLme0W7UBNoDOxJ9+xos4+0uEAHoJrCh4ZSy8q1uhjxfQTMKMC+8Kh
eDdA7x3KJ8bVpPoty7C7DVBu913Jfjvwtm+dflRWdMk4+GvE/QmCFeexSkUOuBum
HK2o/NBf7Xn03S0ecH6V1tZtZnn0Bsjsn6rx9QCeDyAR3g80/3kjTB7SYlJ26QFX
fSKPCxU3uCCzR09MAPCatlG7LQ2RZm/d+B9XcGbqn+Mjmux+ATueMKbfauxmrsc5
WeMputxbSxyk0/QxKaMH6682FoXj0/CaWO3IPp+lTrubS14LVfc4jnIAPNVC2IN3
DOwuiME2f/7XmUdox4n8vS/5Q9dZREBLOEsD2H4Tk4tyd70GtSKzeiN7A6C4fW5G
I8lng0QiQLQed0u5TZSI+a0h4eAsC6XtkOvm2inyWM3jujUJGRFsHHiKWGZ6Ivv2
Eqbk7jy6uOXdw4W+VleoDjjWQs3FNWZ7OT3nCZK7ct+LK5LdLeQMY/VYdU+v40xw
efln0VjyV1rVNk5sZvny8ZfuRGhCF7y+0GmRCwohzkDWJ8xEr8zgeqi3vmPW/x+D
v5Axoio7M+Qo1N2hIkUJtuoQ589dI52tnwF8rILv3rFatN/2R2c5K8Rcjtpaq5F9
zPV0y3UUUKgsTlwHAB1JYu0Lkkkge/gOXCiryQygb9u78vQeQSjthmH2dnOP2sa8
wUJX2SKwBbLwZ1B+VHbWUv2MxS0Z3TKRpUVSFdaiY+ypnnMiAa0CmRKsCVhGt0kX
6xPDJMDo8ZclxqA0sru49R+8FN33x/k1agxPJ9iL32iJci8if5H4AD13XAnpk2Es
s9BM82N8WQ4gu6DwsVdOp5gaa0Q1bgoLT71MFi1jCJIYgwYTA5D7sNSnf0xcqq1D
6gn2afnIzlVLq1vx2UpPpojSk0o2/q3fXhWpU/OdgpN46ZQpLQVOz6O9MDIwpOCe
zNi/mqXmBZwVw/yKjRw7u57QuGK8bADUGrBnVyDrReNWRMDdReVz3oJE/5oVAqgV
utCV/my8WTf1mi67kkFkyttgmVWLCP2aPVKguyU9wQXBs8DiGy2dAMTa/M9LhaCn
Iwapjafgl5BIl+0r4o9lnmhKqHWcNPqSln5tJfTdTkVh8xRjbCY4XyYmY+ofaR5K
zyFbXODXWOipcuQI/REtXPRIgZEYLBZ5dyRFH9t/FoGlfgn63ghPJYSCJcYdA3dc
mv7ygLfC345+p67H6JYJX2/9CuxGU3dHCP7iqL14+PJql79y/qFf6p3jxOcCw09V
K9NzbWx7pYqMqG9LJ/TvyLBgPThisQUp0FzfXyDSzDHPr1hclbl3uPSstc0wPhSs
fz9XMrxj5jVU47cY75S5b5q4TLAzosvIIfiGl64x10s3usnh2NPVbuoi+sNpjIoa
LfbETBcCRaYaJmHI2fdetSgVl7r25t1q3bwEufihbCGrV6d29QmLFn9LirPtQCgc
BdyeylAjndTSvZ1nmZ+8JkKaI1tWFfJqT6skiQG+x3EV5J9RUV83Pg6ucFQGpF0C
Hl75Wf5BcZtMVtrgRNph+CYJ2hCaVKBUIFJkg6hYvCDFgKdyzqt+uWKcJrk9MIhk
7Jule7xnSwYSKjMqbj06w5fcnGqhmgMtoVFigqV/G3GGg5sJ1A8rTW3Qv56Tto6R
FNkd/EFRZEeg2pjWYTSCkJxdfCODsnBI8/A2r5iBrZ84xGqIsIgP+AGpJVxLxlWB
/Z5e2UyZcYqKTfJYbX74f0zBVeek1lmHpwhGZGJZFeHdT142TfrwtokLYW1/KvVq
XwG55u/0ZK0cSLQ7aCTxEUSidAZTSDQLd+6dBsKo8xkY/DqRjNhR2AeuZhjv9Qm9
zR5pcPhEK5nDqxjmaUv49gLGL+UUTXunpDzslY8by0skkLejtYkXVomGwA5TgnB5
HXRRBAOWGg4qZTwDHy0EpB6a4JwLLszf9IE6lk8azCABQFXRcP6wul3BAPvRb/fd
6Xoh18ySe65vuLXAWOHen11/X/rF0XaXQHv34OI9ZZ96JMN0yHSChH42hnnNgLHi
uXYGKNlN4g0M0YWve3Ik+gRvkCw6lFgjEARndVec4wVdY8HRRcVE6OcKS5rN8cAu
XWbUfEOX1j/F71AlR0Gj8iKIgCXwxpniIJAe3K/tLCsTYdPmvYqMasL00kO68B6G
sZsmrhQ/IBiMaQd5kY7uR1r+8adY892OUuekxFeX/daZd7Tp9TE/zefL9suMdVcc
FXvuEcLO6Rqj1JVzyvD3C+COHhlMIqCLElQ8CQuKV0r+/4py2PIiyEcahr3ls5b1
Ez2dLdzaHP9wKTdgBxe2zQK93BxUau7FmbpYrQIb/OmuBUcxHrzd+e4hIu2T+uCm
sTfhO7mFANNUPQGz9MnOgPgjWj9iuyajGRFAjnf/15YmZQ7VAV2tfvFp2p/5kqdT
lzKhBljbRagfEqUwPrZ0wqe5syg6gU+1M9s9co/7ffhqaR5fWC1ryHQY26e5dzbG
wMpTMNzlavgKPGO3blfwx7wBVZSX7ulC5TDfzYJFoSqUXYKXx0ZAQhhksbr5Bb8b
Tbr2S+L+vnwMYIw6BIikigDA20nimKMpOQvqwxA/UN/cF6MV7heFUJH1sIC0UxZI
7+5x0OrFvG055WVarsRxpuNt/1g1wnT/1U4oQSbRZxO5xUWrW9ApCTx5cFUkYR+2
3xEalhpuGStQsS5S0lKMcXyS4ymQCw+y96LTASPAPBVxC6qPo6Wsu1/QDm5pBijS
+HiWxaUbNvWevtYtBKI2nEETuZHoc1W9RDgNCJAmgiY92O4KHPUtqUeZ3rET2SMM
DKmAmf7WElCtHcaVH8TS/5yGrUAaGLw3H3Lufog+vGTHdNOabeJF5TlOIglEGrMf
WlPaA7Rh4iosGKhpMjyRww5z/pOtFual3C089Hj8Zpr9nywMkRbLYoFXS0N9NPXB
vztnloh4x9pWjMqmnmkCQxBzgC9VA9T9NBjDmVfKetjLepR94Gh8U+3hntZ7N01n
wcwhqe0+oEHC+6ZlrS0VozfY46wByUspcxJ9hbTRyW6XpF7LaAi9FaqY2GrD6Muz
+Z28iB4AXZ0PyoWzrHRsCLOzTjW9QTtCQS+OYROnH2HJJZgoucO1chSgPzMx35XD
D9an0EDkyw64VFLU4YzZ2tDB2sWxxfHGLOrJaLSGbJfxFL7N/KDae8HL7dOrNafB
KTZCg5NtaX5q76rMRPbq+Rc+A9tJHL1h1F58fUoBIE3plrspWBXI0cxNZ0zODJFX
4biVR2zUQBKfwtSyh0WWdxkBmzGRufN01POAceZ83fr+ORlmPT1utnJZgD6kXbZR
KYdKXTWFCEpSMytcLXlotNZIT45SMJwlwW9Wmy7s8+X9lPspJvds1w++O1lMiygI
m/19INFs3fIeyNxh9UlX4KBP6pL5dSUrkuOTC6imi64LbZ+NpiMhqx1i9twuwJC1
7Z+xOpVGpDdI37Hr/9c3wCQ4CqpNCNyvZxhhe94StJsAsKcUSGez3ilMCxDdwYAb
NAkjqsZdsYV7a+eN3hQjWvwEtwz9D6dqLeOPB2scBflbdfOnQ5WbDUuzWUFWQfJz
9TicbFsIN6F3tIkW6rPi0Ftrp1ogxBgiUVfidolyfopqS1grSSmO5uh0BIHy1AWs
hY1zeCS+RNbX9ffaScTfgv+vAmKWh9RW248udBSVkf0Bq0Mo3rIwCtGiFGUc/dHv
xMDkzu1fZ34n3Mm/z0sczVDYNNkaFIVzQqQVZ+lQ0M7OHlNFoRMgmTvp7iC9lWeN
oRhInZ7nud41CVo34LsOfpHB90T6Fq3lRK2DwLVOjwU1f52vLNHK/JBoz+w3DFRW
0PjrV+QG64j6Bqysq2pywBnHiDWEU61V9lwG2gOR0wcnGqRiOC0fOEPNj7iV35YK
UT83oyPPeKklgCWefbMIsWIGe/AHFFuyj7iXhI5LwrKQKr0rLdWzgXkgkzif9Jj6
4JhhUW8xTvhaXmJrofS5kcW70IkFnRNbQQFB8tGKLcdcjqUfCaf//D9c7wVp4je9
2T+qJX9U4K5ktTk6LdEdlcQv8zz7AyA9MjoKlWWpXpbg0B+mxI6IVx2ODPeLqjBM
7GY8EkyObiPCMh37vsgKiog+J7+SbXcH7AGw0vd1Eh6QJd5gWcs8oXpQB3l8b6yz
XG+uH5jeHAMQn32x/OfVn5rhDAV2tw9ubH2C7nN9qP08yMhV6SztzEHUGolOW/UM
Xe9KTXvjOiT6xTyMJG3KHIBuBw5jdUskwDmDkVGVNGTCW4wsXjKOYs/4ANuTRP1s
U7JtLTKWeJE0jrXOSOrl/QN/bKqqcDGfAos+KG825D1s3sRegAXHHhKVSdsjs9j4
AvJGnbuUVQoHphF9iMeeamrAiGE0lHbdktrXuFfDSnK+7Eem/DwEfrxmBDeAf+DS
IEDw41HwnAr0P2L0MZu6JVGTH3Zi4lcQI7dbWwwcEP9wcTJQF9yPL7Ut6a4NN7DC
tjhoiBcMNl9CrrJGD6TsgR58vHfcsn+dOmdqnVCDhXtpLfeY8Jdh+zTKOuRP9KZJ
PSyZBMP1M2jzN4vr/lHbOfp8eAeXwByLH2Ests4q5yHUNu8JSdEvRFKf6avknHhR
FsHknz5A2hTc5TKcqpMSwYyQSf1R8TxTAr1eHeTWLv6lTHQr1UoZiqrXfUJvrdub
Ep4LPgQZSGmOHRWDE68qjKGmbxKR3UclB2mJUxrF/dm5noeSU9fveJ1KMT1cy3hm
JQftrOSTyzImBawtbjxCieFpSA4dntOxgl3qAJwkRmxDObcqsvE21QJ7ERqyn3bo
4jIi3zUsl2BuZNPwVywiTxEdirNxs/sfMV07B71UgK74Dv4g9cclQDHHXO+toLRj
r20xqWNbXzuoJo40nhhNSairIT316NFmGtMhW0go9dnSj42Qt+IrEG6QHrcPBqWf
YApwzGKT4AViEKPl90VO8l4UCdmxNxY0AH9Rda6tgBPlwLZ/DFBuXa48mQW0Ut/Y
FHHEkInTl85IIc3WQyZHOUzdQCBCuIcJR10joq4JmfsrYvOE4dkUbwpkGYNPVtQV
CI1xADHHeqoAw8Mc7J1TstZN2NZPPws/uiESU5NzvUKqZF4+Dz7/HyygA55JLj2c
+2+mY13ifNAiTomrfL4QrgXSbikRjrP6N/LCJm/BG00kc3W81SL+IV0tqDxGco4a
Kp9LAgE7bWuDO5e68OASp4BuG7Qi2SCvc0Wpy+jAGz2p/Q6mXkVNqoY1kWDCMkIj
UM4yyn33roWLaZxsS+koKcTx13Ck3g/pJL+FsDFe/uelxUqmcy8pgV2+yd69R4MO
MFjuQ3XTQkoATSJe0WelK2tDiLngf2DGAFt9E1JlehUtpY54xUfGTBDxMcWDeIv0
6JK0HtycbKulycNfcB2gEeERwPcCHtb6rpXe8t9W8mbx8kL01bW2nktyj/WZaR6Q
W89XrSKGeoZFK/xmo5DEUtZwOJfZ6RARXICW+kVcvhQmkoQYVsbRj+axJFD0KObr
J5v0ev/XjBgO2vjKWa+dBXvMj/r0YZccmvD1N/Ht3SzHrrtLddfecqkTvJV9kKeq
Ty5iudsK7h+0ypFC68v6QG5WroRc5TrjHe4oXE/Qw7ihAEUNyZgIZR60253rXYzC
LtBd6SExcRj+RHfwzU0FsyrMMPQkvQGfrsrgqp/qYiklMHFJ53XEKxVT0vojsOZ4
1KBTrL190ZPsIa2Zr1ayMW2jyfZWqkiPgkVof2+ycpOmTwzGvRaXjPVWuWi+o++M
Cx7MICOvBIG+ZhPFXG1loI+lnWrig0NcAGr3QzHlSyUPaRa/tvN1oA6WrvhVi+dv
UYzct+SplM8Ro1oLuMOEk8V3qsbXFvI9OHhhGGak9aS823bZwlgV51PQS+DuGIo7
kd8+9WYV+Ouqds0rbuLCoK5plsXU0vxLa4P7XAM4Y+Mm+p6d9wVR0g11C3WdHKmr
Fd8vnz6xhF95AhZQN7pgjpIQBF2HUA/dCW36/kgYTL93Ij9dJLqZI2qA1vUPJasF
1yaeLz0JO+KqDpA2KUD4OOIXpXU4w3h6xu5fOrwOmJwx2Q8q1euDrpFXGLZpjhfW
J100MpQOEUNc5YZlYhcZYslYiBudeHR9peFEBBzYJJlyvXLQnkdFT5jeMQWOnmo/
iZOjk2XonYgGa9FC/32objeGyWs6qNxdw0gwgLLOvvrriXYOp3ZzLdq2rZNQRQmf
xBJpOsC+zTErZANpnA4ySW7iImHA2KXb4i47AaF5RH19BgQnRzmX66I1OT3C71Bt
MDYv0DLOWEk7nLKma70xOt9tq7xAugfSLdvrmGI9Co3I54kbqLIj0woDNyEWSmC3
hf8DM5s4cBPQXz1E3iYWvBgR+uzQVONVpEl4g7syv8xpoqllzn1ArKX534+hUGF+
TBSP9yihZmxJhEsRCjUsJuQB8NDgR9Vv2boMyqCIdRwm6nZrwDGuREw33P9b3Tcy
lZKxhMHnOHIy6YLULlTbS4f6PVXVTR8CQlHQhHp1xu3j1PeCx4gF4TXgkcbzDg22
ByjiTd0TPxKiZNSpcWfP9ljirxU1FYvV9Ohmy32RvrElXcGxV5Zv49MbWguSxb1j
nVMylEAA2rRXE6oavvf1jUZbp5v2okAF19E1RXOncFSq8vxocics8rtU6MTNeJfC
TlgiDeunkozxqoV2Pie4zXWB26TrW0GS52KAjUSHPs/AG5ok8/oKLM9VcojpDREH
yv2hzpx52Dgi0Dbimca+rcs56DlNfz/INbH56a3LmeYRc0BpqgQUqUuk5LTH1XIO
HbsXGNic5jJFxFqw8GbbYf6p58YU0gWq1ctBqMPHgUQ45xAHvonH7ltu99IAZMLa
k1/k+aQ7YEuwLta+queiOgORBNPOujIjz/ChKtbUiLM9H1UzOUepr0ojlSz3/EYs
XLvEEYjIawGewPPcwRdILtsrigrU78AjRadLVHn3kahahdNJCsGXZ7RGh3SGyz5V
CmNrjld2f0EqMWZYs2EixZqFSjAlIsVNoPmun2YT89Zh657143XQqFNkLFEKfSJh
v+WX7K2EJetw39grt3klcfXGC+9sI6CoxmZfPT8/kpoo131Mpnl7bnJXh8wZlwen
FSv8QdfcpF5OylCgm5dcAUNjYb9UfYsWn4XxArsvOZDTMzaV53TM0mxSpCBy4ZnA
J8c092CeRvqAir7EDRYMki6UK35LQAQun1qRjU7EnZknIR+3IzqYRnCr3Aem1u4i
274DFNxnAb/gLRNOMAo64mv1o9ID+ZBFTyW5LzlD+Su8mkX/d5pWnKOPUNCRP6Lv
pjvHa0z/K7gPBnJGQmu2vevrZYqTexYEjkejwe4YllzHrKt6eTsY4CKpYefKN0Tf
q5K+Mj4PXlUftV8rYUGo+2HmrQFTJpl/lBJSbdyJ6lqP+xZIbuPs9z4Vxkf14bHS
WFT5ZpUgCu1bcvLOgza35SNH2kCCUX0HeuNGBUa/o0f1C7/hnbVxl476mDdulcXL
t6Hn81kGx6YzfJ50zbl8KUjE5Sbr16xz0hLDWxkNTIybHfLP3MMAvtbKOyo0/Yij
ZNOBGvyIkU36P3w+VJEYfdJc0PgXhCKHJmgeCklqokcK+jTTykaEM0WusFfICpHq
qLppW1q8FA1jNpvGeUxbaVVJ5Gc5/lhbPPOPTSwLmogtcr651Eqg256w54NHd8nc
QLj4/GywcDbIk3Ag69AsEZ51Pn16Hms4UN5Rbr3XIOVEwRUCOvr6m9IFnLYA2UV9
UrrHyaCpcQEaKdXGfDs1r/mzHJoaImPt5SrKvBySBp1SoazE4ktuk7tC77zCK6ra
8V0SJfVpYJUtD8JflSdLsDCxt5u5lvPdriGPzAmt6RoFAwVBuUrHzvcUS9huATwS
U7UvmzWx+Fk+EFOBDw5wHmIi5p+ibBzG9N/IpKPbdA031SN7NydznNyABe/gfQ4n
oMmnnvJd+dThjVpY2u8z0GF8h8SyJv8zvljzN0UmNQmCjRs6GaYRuTzWgyySrCHz
h4BRKqf5Q1/C2rrYAZtJeycHtHOBk+iLHzTR6UpzRVVmv3U0vIzE63OXY5k6MTKk
jFvt50SI8CQKL3yy51GWAfvI6EG/JzAPfb0/ErWJ1C60Wm7YmvIZDhyw4CLfdWxz
fAiC07B3PFHXCPy3SrP8PMda4bTYJKabOJtC35RIZdooEpcX275M8oZ6JOG1Rg4I
ZPWbURIyRPcgbif7RQj0q6hnyzKqayUWuXQikS4hPNoG+XkOoSubPGrEp9GrTS/a
mnTQz+PWDeEGI6+h1COdILVagZgkSId9cC62EfKkb7xF/9MiO8tuzk9f3iqIkTuB
EprWHvJoIzwGOJHWIDSCFyo/Tq0Nt3Jkk7+LIj/ER/oI5rSQCsjb64+ncJHuVWQ3
FsEtapjjppk2jfpuY+nDCnPIK2f3F2lcbGA68op/u20HcqmsENj0NUenimIDEYg6
bunPkRkzmrHj9ypdpIu2qT8zBZhtfyLCDvm0HKVuuV/0SSNnVI+fxcYrqyoEnqp2
pWTUcwnghXOJAdDwHNvp7fif21zOnc+dFEd7GjxiL/zRPf+duWwPdz0QSzV1vL17
JyiO772eKxgklM54BWYFLNBazCnCEtjMw624egAyJh8Ryho9eoxpk294/Z790GSl
3TeaUw8jM2CRYKMEymJ2ZakSwJvfC2VamytYlJaQm0DaIa47oNxVef7bk8HRXWXX
G95OeyQAegsRgGFN3Q4s4Sl67ygc3Wi+6YPGVkCAb1co59Q0ELvjG4tyFvLLsmWZ
Fan2g+hSZilU8f8r1JuSQ5vx+IywEcHx/CY/8FI1Do+riluOiehd/YEtDBPCyMIF
2Rl+8Tkd9hOlYz3v7tD9dIn28VZtfZy3+smYAutsS06+1fUmxOC69ftQcrbi4N+w
1QtBEjSCjpr2vBHdHanIFEUQLl+KS1S0hvJR9nZUmkk3fGoGujQ5nOUKzllm2lSX
3PDRiu3Xq8Rb1f5TX9gvAPaGiAIY3CCTGI8+TYpsY1GRKjmCzmvy8x0FVA/Vm6O3
T8bKHee8MuTq3t99Zs/fU08BBgHJAU/MgqTwzZWJ0ehNzsjeoDXQtBaY76rVzVQ6
JKIydmZGXGFIhl39SEsK7BBL2FGKJ3CIFwhb/1pj5N3guUhCdWOChtZgqmuW41kc
iTgTiKitWvD3qEEqrXE3YaQhncqjp10CQvzecFukHZboiIF1/oHxWio6L9I359WN
OLxeAhM9EiaXHVoMaGKV+iBCxQevTZYhbgHh3hHSujqo/4Ve/FoNXtPdP7vRjc4U
5F37PBo5rK80s/8pJlaOxdMW42OoY0IoUv5jhjH8w2qTuda+SUG64fZEr46BF3ux
S2chUM8qnGLMJt2acwXAgmtiIhhMsLQYa8rT1tTIt0MlSHn57tb40vTp4jHhHI6Y
O7RltUxddiPMatrWZCGhCuS0cQLnpnsm6jngmMROGw02mycIF//kCyRzo2sbFWD+
+E5Xp3KzkbNOwToxBKNXYbhkLWl4c1G94qsgAGlubtYj1VnQUOgFEd9hW4N2j+vG
LjmA5MZWYrHrL1u5WGlZz+lI//CX/D2KOsAsFxOHIbuesv9z5I7cuuCCv4qmLcl6
x1DmC038VdA8LbQkma58oWtTNWA4ozVvEWEza/AAdIkAZiq/QfbV9DT8HAwo3eJy
NurAO2HlDZ1M1SyKiNoLLWsACPUu98IHxswS0GvEw5U0JvJEyAHGN0lgwFS7bmin
a/oFjvJCp/HvE3yMSpTSFuzYpYC0jr4WZO9gEQor5qfo0Gtn+3/SwOg/al2fxT6E
IohnzoCVEXKuERDI//Lm5cm8985+SJd9EvauxBpKCa0YDo6m/pBVi/9F48V6tn4j
WwMYBfzgSQMpmusIyiST6hpE3Xhd/mRCPaWb0l/O4pFeAzgJZJU09rMgg08060HV
/pIuySpQmMkI8ObFClQ0fAbm2nynsuSG1UT5Jky2+bo/zAwZH9vLHQadFjful91p
7HmfVseqrMTMcvfnofZeGmlZifKnZ8potONULp+QYIo7bYciv+70Z1Z/HMXOf/rM
k14HEUu63li5ZQt2C+LcSEAfC/oySEajWrEfWQtaLneMyVdC3DfWz8F7SHLm55Wm
Xb11vJ33dOqkH4431fmvzymlZvKFpFttlkFZjIRcMqIWWLEWNK8MlXybAjInKk6N
mKhkDORl+sLTKgGakTVFgb9sAOkIhskyMtIw4yrj+I8XlNI0COyCffsNmxD7mpHn
ucVvX3hMhy9SSvV8QL/rAjp+GYQM/iI/jyOa70r3Q9+N6cEB+GvZbIx0yp/mB0nr
U+puW/tBD5dXU8GJh3VD6mSh+QbtqYcT3KZ7e9MQMoHAFQJ2hHBlsJ2I3UFUuCnp
JhVGJZD55jN5FYumXrYV+jIV0aFZYFOxg0sFbQUFArzxOz0wY0hRFVsKxVIyu2xm
Mbkg64d4vW9Qvp8XwvyrshzC3DA4OzWqyJCNylc+SAZZVTO/DgJcRqcvQ17oz99F
lTDmonwCW+NDXxvuq8yihWM/LdAxaq25dcqMGzULk1wVG0sVvZ1dUGda12f+r5yP
r4eBNIO4kMwhcUKWGYhsFFLQzKLbLyhXbe1GKSaXm9u/9nUxStdv+sSOV5ghGIA7
R8zq0tipnDE+XeHgyzAmXiBKFjASDGahbBjB2aT6NrNFlMCH+fLxf3t2Zshh4189
Wnrek/8LdHah6cq5YQTrqCKLddLoo08fHG3t2DgWYVaFxSb/IwQfvKlaC0boj/0a
Xb8VP0mIgzpYBThywfE2v5kv9Xk06TAGA7NqUe+FA3api/Fmizd5WsIGVXGVgn6t
3YGgTxuLzaRL0oBNa2KIYmI9+khJ+Zo3RPa84zKkhbq/ZLDS90Mm3AmMgmDv6ReP
JtKtkQbeLd8ziljxdY9idYv7zVnUiV0rjr4KJWgZTxeIPIkLm4XGOzfTabM+FGzl
A1fHqeZxq9LuTyz3J1FYu+sFyMKsc4uvBDRt/L21nAYpCPD5h+mMdYavZo6KJr+h
9dDfF5Y8blbOq4b1PFSFc+7wwD1/LxaMCfG+ltMADDpY/rOArMlxLGQAZNWmS+6d
Q6DYu6Sy8ZDfkKNYYVpmQmwM7/KIDpgNwn2DmrBH/z2LBh6TpiYT6m109GkSbzb5
Kj+qHDHcRy3qnxc0rUMoYCiHJ7aV7sx9tEIXajjEr8YVdlJwJ/a6eWipeO2zywZc
Hw/HdNAE/uCdhzA1L0DoxFrd2zQzLPv8nAKtAdnRzbdxFTEoKO2l6zf2ys0zoenn
Fa0UR2/x9gcd0ZOH2FilIYZKFMzCgJbJtcQYNzyOp16QuFzkwd/Wy5aNJ0yDzke+
4ZrU1s82aMY6MU30Q0ihZ7Glcg9CZEw5VRN6oGw8xwaBKUzZEtYz1jhsNuXN9aXv
fD8Fox92gcQZuFLVt1TJsjSdfu1obFU1ylQtwKpGjm2AdEm7ZGOBAl51Bqdmm7/v
iqKAXL9uYIvOzgacBZ84WZjeGf0jDhxA+P8kTGowtqApvpN/2Nio7ojy+x98tqyC
05xdMbOr+mk+0OjFYiciiUQL7J/SvbpByu/JBKoBk2ejrFFM+ZaVSL3eQNqSllwO
xAeGImx0dL/K3sph8J1ASXixYr6oOTSUnS45S7AesG08H1gHD1hBwc8EpAomkQvq
W9OVQ2lBZZq+NyuvZNTUdl2LNZTDcHE3f9a+hMhKIbJioSWmbIHO8/3AK4vXeSsI
+ek3OaPLef77TT4k0+K8neXY+bKJGgUzKgOx9hkUErCswaJcfhLtSIwvBd/ZNCeh
r1f/ZgdJT7P1aiwIhObh/r8R7OQUNlZMuXJbb/Wrol+ITYH5P15d8P5wnXd69uwc
n5hMX6l3ecB23TEcM5O1//ol2JGksaQlarir7dwIh3d51Z4R1XFEw41PVzv++WOw
JPuqLidAO7wgkjEAnPONJLm4YfdHIazz6cLjxOFe6RzPfRFjsrd8St7xjqKblsYS
W/NhqsziY0eTu95/Q/qxJPyd+WX45hM69USe/5qfV3tUVleWXT67Q7MIC9rsRLGJ
urcdROOkzEQe64oK9q3R+eE+WW4ijR4UlkkE7iTuT7LkDndOodSGrq4+8T1vTD1q
/KImvFFWqVbnwAMV9sif6D8DoQqXH1R7uwA2dGGHWj1ZjtsnBZgBxFH1s2DcADKa
Kf4zklrxwkK7hY/e6DyMg/uZfoEb8MmxtLkwisMdOImPOopxiS8Gt1PkDpFNZE5i
/C/umYQSt9sjjEFOdAKFGQOKrOcs63A5phukdVoAEAfSSPiBlVMXQruXCaUICrX0
Y6ayaX60fkacPBIipar02g3CwsGGd+QehFalV+g8lYrD26H6e5f+1DqO7yH12TrJ
r5h0jE251IyHbSsjDjRUB4Pv0FTFg3UmxZ4nHDgJ6TwN1spTcWO4VTHwR5LGzciU
htbTMq5EDEABuD/kG8CHKwXTBGGDjb6GbSeCHdSLizkzkvmsHwSVQhdSiCEQWzAM
wTgXIZ/vCIjsdLlZCKRYyAfUSfMSbxcIr9EF91/nW2CCXmSNu2M13ehJwTj/I9Zn
jQp2vLkYpxbpug0wUXRFIabNYrrWvMeM0WciVfKEKqEI9lJqz3RADl8Okzem8kcK
5fjgwyk5QVwPEdiBzVntCkmZ9iZ1PDPYFZyc9Q0jwcN4nxnq4vsKB653FzaebCeW
IZtUeWDzbouzRQTT3RUHvsR2FaiGQ80FSI6ArXj8G9FQwC4rrTUSwpf4WfHK6KmA
fk0mf05PiF53AOyL5kf7+9HJW/oxxZIn1NCIpBagYhg=
`pragma protect end_protected
