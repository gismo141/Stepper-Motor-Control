// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HsdbwPUhEVjFkbTbRRm7yQ7c8smfiOCXon7C8sEhvTk4mrU7cQPZImRw00qFwgvw
GPgAx1w7Bk911kZABZkhs+FtBQhghyOrnRQWzIeiPmPHy8PymMnLqVZk6PBMW3aF
OhGI58cUNU9jz+/hSYLpdxeJCgFBrFpvSYyWiIYimQA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 29360)
eYR1CA8kEvb7r4Q2ob4CIVelFdemB/yyuh3jL0vCEB89iEUyBoWEWutkLdqWfi9r
K/X1/Mi3HA6PIbMGhftp3E2H4YHnNu5fZWgTVL/Gy8zLNcjdcrWaKwlSOWgwZxkF
SrKUnHCykL/tP7HC5G+YkfpPZi70rfFvPe4K/+zeJAa/XsqxukThr+WGzU6YTOvM
zVnIVGCup61Cf8gLmDSnoUwjfmH403ZS0lEQrhe0a2hFAifcT7wSHnr2HtAZbOqP
QjoGCgHaGfhXdMpHuq4Ta0HVmAn4ZLyw0f+aKMcGxNUJ4otLA2nqto8TIOOqklxl
GDl7Klg3MFlIULpdwrhA+iJhf6i0qprsyVgokKCpr8MvpJkpxWJP6QzCnaxCTSb5
gDim//NwNy8GBheWNhT9eEtIrCD4Jtpghy+hdXmDOKVL6z4ChyKwf++ZJMQ1QjXg
RVHhOlkw2usspPjiu1owufv6K0aIRPJiKh2HuOB9Yzu0yVh8fbIFK/i7Ebs22l6N
hytE0OLeFm+1J0wZJTMR9XgLcev0BRvF3SX7iZ0FiFHDhj1PhS7jx0eAt/6ZUhCJ
YPJUa5gIS6rGVcIXPM8RcNysttXwGOODzVtcFuyVCpJ7YIthYoIAHNW5IEzJMqRK
e5WfQvi8X/GbxEIRtoTAiw7CtPZXSi/MB2aBl74US3/fWlpw7bfG1pbef7M3UX/l
SqAEkgEI0dKf55Fbttcxgyul0ZX93vAwDG4l9OXIO+oGKKfMljWEmlNMK1tHSNPz
nucAX2tqmzCglZUPfPIlpbW+Uymu4UijT6sYGQlONtS9mS2E0L1tC4H745FQPNBR
7lvxmJ3Xuz3nyWZRXgu8jMI5VKhRyejXNN5/Y4WgIFpVSkIJYL4fl5fUDaqcIQiX
pfVhEDgQWuj9FMvJdpqRL87vfyqdoQzoVV7n5N+KnDhiSuZGtjN1PYmOcJU5f5F3
tUNyd+NRHs9z9yT8E3X+wpAB9b++tyEZK1fmY65TqsRcRi8KE3cTiC4DQKCRWwNm
WD7oR8wCLqBAz2BSgTEqzr3qX2MvigJie1JSNbhpHm9ngODN2P1QuR74iDLYEwsg
ARAPpu2dSwE3Y/F7AdoL5JCf/2XFN2PzALzzMsx91LpvK0V0mwfFzaaTvXmpsnPp
5ja6x/19Kmy128vR79pf+QhFQpIB4WfiY4dQ2LhULTH3r1G7v/Z5NKIHs7yajOAs
aLEBdS936qw8xdxBpDHAYen8k5wvWbEuYISTP48ciKA7oN2JDMVZaBnQTYwOBGLu
crUU1MSjJW0mx1MgWz6XrVmkKuW0PUYnjgapVwWykzPc/SQhVcyR5/dk7151i9zu
q/w03T7x8ejqtzShdNVR1oFnlmvFu1Vdr7Gl3e1XA4FHn/AhntWyHu8yVs1Kui3f
wfZwZ5QQwyX83AMdmMTCjSnH2bMg0KcNUe3LFMNdeTsWpD/bxeAbGJ3M69yKyJsP
//7I/rUZ/VGtuPbC81nzxytl+hMBrtRXVD5t0QpUI/MqlMkWilxY0gWXql9CGw+2
bfqz1pFzPhtR9l3glE1kdiBMW3q7kRn2i+sv25DjVr/ueGOJhbdebmyRPtNkLp2M
TmD0g9vvQjg/N/knTJW+X8k5wiOqQCee5Ie0rkhQSAhIVV/R4XmYM0jgSy6+71xV
C11hl8X73YQfgDv1HbNU30uupKGFV7Qe8IPQ9c0cLs2d10PJZxsb7Pyn5kPd/kPO
PSqF1dpSElyQByauEl2QiVnjUr3mJlJpBK07MhjRmAGgtg2fq3apRlJNshpiyXzQ
91q8XqkhzP1RFRVxPRKoWLUvspAKXdnhweKru2FTVk4ffTGhRJPmPkdm60TmdlZn
G5Mn3thLWkwapF6nOjJ4ooCCt1viYsn1iubZ64foXYO5mqdv+dvEifo8PKKAt9kz
PqHRgWObZwmRhJ4/tX6TWuN76eApChGmbpp/fqcBdulMhIbwafYn/IBQXQlVVJz2
GUF/aqUTKsNpuoU2sRGiAcFru7f+6tpQpp/mMhw9YPtqcvTgDKfibhpMPmBUJDAy
AZToZeyJUtpCGk/eCbLBYbngUpFyHtvK9ISgzE3AenQZDv51INJCnqtPj0bm9ijH
Y835RaxfU8YtvDKCdldFv0oN6pOdKO5HYuj1aEAok1Ap3dl3ZMg1AUbay2dSBiaK
kRkU+AYAzGqADIArAOQRsPekFSUxOM1v0B30dKUFZ38R2xOHvKfKc0VD1qDNIIp3
+DBeudxGZUNj1rsVuBPWoINu+OIsl41YVPV8RT9PAKdXZMRxS5VqulUn+SvDZeY2
TzAq/ytxwP3c3PApvPfsuuijmfWoRGvJaTORpvvJeA16kIqTeMU6Zipidwq4954z
7DfMOb9NkSFTGEXLIHMEukX02uDwAlAep9ZImRzvzBnO/fu9IUP9yyPBOKs36gRn
xYvQZOwIkTYYKbpnN2uy1WKVKHobYkkNn/l8L2JyBLTIeeu3ATuIMKiMs5S60xVo
bT1KZUbxU+mSoSJ4QeMh0aVATnxT//KbrjX8XA+fpyg/SzL+q263XySl+eo34siJ
0aBpvpVvx+LTImSKBOxdBiyFcjS4a4KF5qosFmNdnVZbG5qhkzN5HPHpsi0j0jJx
i/yjwsMk+d2me+hF3sVKnhEJ996g47mtXcz9aU9UV+REdAs3Pb1wdrEizFx0CGME
CN4BnUgqSl9j8L7kMV1gmDR+uYqvUtKgx4MhMv0+uSr7jcXDBineZ76ALlkc3J0Z
Ok9bXpQqQbPInk+4FrKHiC6/n0GYrzV4wsbbUW868bmEf/K+m50WUWogpBQrxalq
IS6kQcJUAGdtxs7YDjFqsg6v6jGaK75X5aTJlCL1KFCdPCmaCnk/nPsWxthi3yx6
166wTa3rwOI6PHPewdx+9XV91xrY6dSXLyqywLwN91gDUs/p8yoKaQ+UInlgXw2m
PbeM6r2xk1De702ExsfR1WNcjYNtmz5ASeFPvbGoZXBM4ho9Pp6DI4/+7Ku4HC/e
DRJ2Ao2e4rTO5lGSDwmNf8rbT5cGFQzwnLjA3iCkNz1Q2lxIbtkgGcIOdAFQZurv
dzxxip9D3MvxhIid7y5FvJOlkOX/feHAq+IGZza11HJLQmCCC4B295jE/ZBQqC1K
VRaed6GjPe1kwOWoLEP9hOYoADvLnv7thZirkTt4d06a0U8D0KY9nsWdUMocAo3D
cOxvGKH34FDLh2yOC27AwR3PYFFHAJFbWZKPrGln0pOGzYcJDdyNXSfTkQy0uJZ9
G2NN6Kn58M+Wo1fQze0kEATlT8VHXp0Qoo/oi/cbnx9izZPbH7iHadCQOK8ywCDH
T50ttXBI8PsUHcu721csz/4CLps205Uwn96xpVpCVC86TAQelx3bMkN4g3cuokBM
xP3VkCEkr9kpNAvV00ILiFS/1uPpVo8NO32MIMWWfi/ByrwBQKnGcxUSJlTIg+nU
SOfwdO+dF0DYuVmhw35nhALLC5+77nBeKjtWggaouuJ3K7AR6qltSuOtEAwV+33U
yxD9lEoXOk76qrDW7in9GrCit7PXI1953aAAwaY2kgmmkpFRXZR8MHByXhVIpHgU
vhLkcdbCiLAQrkLkH0y5W0OMcXADwsbcyooJUOoJEWdcC2hBFHEK5q15W+Fv/ykS
YD9sFnuUCXXDgXFfRuy879BPtmwisPhmLThaO78pSvbbMQJsoisC3Qoxx6wPrhDO
zJcA4xXgiAIkMSPuaFA4j2BatSNqxylnBsgZKLHE9uysTxw6OeEgq5/N78ACI/FU
xhDGWeIjdqY+C7zI9NPG1Em8sykVniAaa0jdWpnljM1Q7ewtKesNW+mG+BbpHjOB
JlFZdGJkVTQ1E6J/Q4Slx+hSV+U0HzcJ12NaZ9prxrZkyNmO/RXlKrTEum/O8sfE
eWmXoiF7Be+WXP9F6eRxgZk6Q6Gd2Pv3U/BPpx8PAPElWZQD01kt0JbF6jjRqFKp
28S6qPoNZu4oTwcLzO3Q7nPph11DXgpEhXerc57CoZrs/n9B/qKo06wzMOMYCUEK
FJC2UaLYmikOt7LQ4dq6Wipoq603oPQKzVHJQWuTaC2eTKAsOUei5xXjCQMBcQs7
Vt5Kauy/VOvAgXBu+ICgj94b7O6zImdPwlPSklAVeMdCVE/1A356h6CmKOhf2lwt
DVkNIopGTVTOQ8AHnsNstZAFrFS/HbLLONzTiKen5rRKfsnwD0Lcdr80OX2AwUof
p8feiNJciJQn7FENVbkbMIaMpAfjbRilzFZSRW+TcFsi6ZaeNcELjXY28xZLGOI0
da3yf1+uLMp3GzVyg8cqJy5kZv+BYcxy2p7Butnt424/3wKF+tnyeVxQM6kwVfhc
LXc37Wcwwcw9UYnICLMUkmmxqnIuNqRKVE0N8o/SCFCkdu+yG9M+c5+ErLPwzTZN
oJWNajL0Rt/IUx6/E8m3vGO0+c+g+wMmYgmx9Q1si6mvs1WPI8j++T7rmllyaLOn
asRirjYsN75UN8QyezzFExcJDYxRLLCwwKi/E6Mg7hu+KOpo4pnSUpOJf6ujzWco
tFbC9NG5zyhkRLSb1Vl3J1Xo36On0y+gmbDYYYUDyC0hb+jZch6LxhmN7SmiWlFk
UHBRh3A/yhrM4z7P6UN6zI6bwgYHZWPo37TMwcdpcxgbeKPenQtcF9aqeCqgDsCM
LznnJPnJgNKVnCUFp1jftbFSy1u92kAim+HxalinmdBE/Ustcxiv8GQUhnbysT/D
u3rf+UioHS3C+pE2Xq6foxF04vZ1zNO+JirkuSDTzWIDHygpB6EenMv5hijsKarB
Ie4Y+WmmerVVPQHrWAPuBFGo459mMLC4tjInHjFhk3UqjAf7CikPUhqwC2HP9QD4
2b+T02Hkyeq4SvFlLV8j3RbF1gsad+H7J25WS7Kdp/mCaYKTKejOXqvUoGcfwEhO
zDp90aWzDxuC7n4iCjBAAxBqdSo5lMk7OInguB8h/jz9FuW2WV9HZKnn+JNlmxaL
JnVsd1hn4dA3gSfpwTlhbE8Pf3QAFneeLufMX3kldS1CaISgKQ7I2EG9l2N9DiPm
HYssl9st59/y6EYAmxExczGCxcfXJI4pltzvbVeAWZCODZlmaFOLiXgW/JgSv4Tc
YB63EDq+dRIxbU364wCvKcgRFgUaCOJdJf+iwD7kgo+Dcct461fKkQgNghiF+TaP
i5vVzz0IUD2VdRh8WUT9T/9rI4lQUUPFzC7nrBojTCfqIb/4uFikpR3ICpqmPw2W
K31zBcKYbJHjT34LFAjrdig1tI6MCQTdQa3+bVJWxcJb+l+zvHd1KekqcUTBgl0F
gbxmOlan95Eh1IoPoy+FjgJeUaiB3/8vozuMVhZ9ZpVk9ZHMrHoN72FDlZbxxllz
csu58HR1y3wouExWNfqjCeTmWViJjeNVWFRkUeFiNTr5TPbdhv60TQZigSUGWgRO
Ah7XoywJYOIgr3FVUwYxV4+4KejwQNrjTjVYTiwItLgsP81GYUJEagP4eW2u1a0q
0T3Z5+8Jt1JCWCWqjeVdNA+L/nkkkTWbBkMZLmEosVRKpvHs4SxLxjc6Sd/nO7SE
IrHHGYK17TjoMzMN7WZxhFAuc+FaWDdjZiLGz/0i5whAgctHqdCwpQRxbx+PqR25
GEuj4lsYFgrzSeuGDOV7wEoGOm9OS+WyymQ/cKIOTcE69sq/xcGxedCxX6IRPZkj
9LogjovjDxWQPMMRPXTtke7F2nrhuYS5TAgAn7jyhpgMPbgDr8lSn2sdWf6K2eS7
j76URMoiCJ/GULjirEZsMxAHmhNG7+w/Iza1H+VzlF6327VVoubh+jH6trvOjzjQ
snzmbkb86e4FWrJKqGt0L3wBgs8leOrIVWQRvPJaa3r7uBgFxzUMdz5psTGS/NWy
KaxYFXokGOUcS96cJSxLQkYhSIJx4Ru6BiHI9/Xzff/Hs4zPEIjHqvyVY3Y6MFbx
4YEx5PiwiVt5B6DEHK5f7eS2z+V56hmvRPCmJwrSyupKKQE+jJHSyzVce+zxUNmS
3Jrdgj9OJInnVy2Eu+thz9ikAW2nv7WL+B++Sge4BcV13aHqs8b5uEiiQbRcYJdD
aKhmBiawsTpV1y1ku2P0yX4rB6rmuMMdVo8IhnMo4BPejxdIblywi3Yu0/aIOlrx
SiAZSqR2aMWa/iJq0NyDYxiOWjVo1tVjThSHOVA/11qqyEIE/l4dccVQUJr0PlcW
fh8vN6TDfcVWgMPN+HufsvAPytskmo2k9YUDvt7C0MjIXw9IAUwCaWkMGYIfaVZh
Kl3AJQe5pqjftjzmf2ahuhWLuKMnswtzqgAcOgXifKxlweCPXSnEDPN5AWNP66y8
l6kdJx16yDIg0HVLTvERxbAcy0w8K0oiY5YaHrt1N1mPWyo1cxDpHjU6ImYFLL+I
Vw7gT2JBwJlN/b44mQH7zXsogLJ9nYxR7zlsgWX59F1CjSBmsmZIi1uoLUNR4mfI
OP9muPefvUuIGQ0xUhlWf1UZAuEb9tyK42L+BGXgzz6HyRrPa1P4t6Yx0EvH98hX
zUy8eg0fOC0kIJ2uTqJQuE0sYDZ+HBMX8Zq7vUHZfhC5oQ/rDt1KUTnBitwjpAVw
TGlCPZZfDdOINRSVyYuiZdGb5oSqYWzivQtdNZai2b7XOpqR3HCfCuVEKOZW92Ol
PVsmwsFconnTbM4BEXqU8jpAhE5mxvY+Y+OMrZVLx4TSClR/goAuQiyB5ixPGzyt
V0fmoVnZfJxbRqlVpfG0Nz2twpcJLzwEkaANQK290eGhYFc0SO4eoML7v/Tib3oP
vIABRwbKrFFCw0OaBqnZDjuAghFitWOtGP8GFxlRrB69WXR5uVxfj5vblYFEwXwG
jkxaIgOm17o/imQ82qPoBkFdH+whzGvllHvtNIiOaNnO7wkoa1LuX68gU2rygVKG
9TpppRGhToECVG8HUdfJKwG5MWCUJRMXAOK8FMcF/HPkvG8PZR7oiC5lcSP/gllH
fcAXI+d9NbaU6eJ3lMg7W/YmYbwMw8s9l71xAghdeBv+vxzRqlJwx59sFdWYsbot
GmjDZf3V9Ml4MQGB+10Bj1yex5bo+U/9tYrTW01iMDWHO/8Sd64Q4JfLYuY4IBWb
o8epK0lJPKj8VRHq/2sZm/iA3/uRubn+KaFkBlRCzYtFU1t6U5xn1HPGoqhXEzXb
e3UhJnxaLELIUwb6LSsiI6uUnNXjFvB7M+vke1Vu64ROXsYU24Xsap9occyo68oZ
ET6Awk1ONaykL4x5P4YrsN/cQMJXr0+FwN9shR4XKUmyKfl2eJfKQvpDNY7k7XIz
+LmBw2a7ImmUj2PtJJx09WAZh0R6rhU1jmtUjDJyLFHeKRnNFpPg9jms97H6z7Ur
6/cxJ5NmqMAcqOC1qwtOzfQ7ZiWzhGI7R0Y1r0GtSeZXM+/E8bnaRX4Brq7lHMiv
Mk/HOOIpiQFeIjTahYxI39p/Je41Q8w4nQtGPyAQVus7uz1ZpQkigoeqThMkFUkI
SHkUnQYOiqeBkW1LlcrzAfNBLKbXCIO8gneENekGyWA0hQ7BFL/7nh2dbsa3wMnK
EXfQ/P6zWlINadviuqw49VWdQkeUVKu/5V9Kgn5wgxO/TcwWiTZnKcui8UDnM5/F
o+JVDy/UAUBIEoO3GBEvV8t3g04xBDm6y+eyGVnbnx1q2Hp5IBsKzvd4BT0kkzW+
T343pdYWH+56L6PB0W2CyNGstkG1MPM8ABz8IbZOSUBOFm7oBtnWWlKjdc/cYCRI
V9Lqx4jfHq7UGMxNepk/gGGv7t/Ql6s2lzNLpSaxzX8eX0D80Bpxy/EBMZDr3Vnk
0JEazUCaiMSlE93SXPEQY0+dipaxDMaCWOIlDay38iUhEqpfUBhxqfDJm3iyfAPK
cPQTTaSm8zVqgj565/8L8nXKWX3EXUF92mEfBPYPW+IdC9CxPHSP3tiVDw9o4a+w
KTmNfWzbH2u0Ilz2i6KkiAglAxl/WEQonVhHDVAhsuvZ6S8+NAKYj3qVIUi5n0Eu
BQtlo18axZe55DNjBPkzdhsr8jrgXtVhogB0FpBxj5YuXi85oHBLXc0lBRTTG88P
wPbSmI2EuNLd2jlKKxzXaRGmi9ebtNrt9qXHpjegoruXH3aeYj9h+wi2t8IVhCOi
dqYK/fHyf5F3ueqvxp32jDDLVyctNW+0P9bt9tmGPzwcJ1s9Ky/e6+T0tDGd/pjI
iE52CY1CEnKuHLVR/ZF0RXQIzTVXM8lnwG9nu/afCdShOKPaUOUbNbnshLIi78Bk
y+xUKcKSa3eW3rcrR7W20+C1fwFn2fpau5Z5FJmdVdU3TkdvwKNOaaJ6Nw7s0QkQ
UjMNQo/cZpLMc7e15EiWG/48UaB9DZBmH/GyA+9wIXBUGJciOcbK+lSu8VqchMsJ
pM4Qpp7xxZsULESMHC7aq+mkT0HcCMFWhlej4v6RcMcsINNzqggmC+iYE312+Njm
1ToWlD5RO39sm/nx4IZ9LVIwhQXjme73araJ+smJYV2g7BZt692u6+A24yP1IyFv
e0kbM1ebYiwGiGHZwhC0ImDbkCN/+g3a4pwSLBmu4VI5y4o6XgM0B6iB+EfHGrpw
kGWxqR5qHTD/Wd1l2YSPrjuqPfepaFfFXqY2OFHLRXFhxHlJY640wvRoQDpQv7wS
LWjKX2tYKh4JkVW0C08r0iGyMz9frZTMJLnN/wsFj4h+hwWWMMHOCjqSt/7fRBbi
GnK+QWnQAKw3RUipEwZP+geE/5a6reAs34aNC/ue1ecSijAbcJqjTFfQ6VXqIIhQ
EhRCgR3lhGc+f9cYcE6fu7HiiZejeBloR1XFfJvJCBrIRpvC1tqP/8qPRBis2usd
kbns2B/TO3AjllOtc8VJ/0jZf6Rufyy2usUxInbKjygOwZUsxnU8FGK0VPHdxPKN
6zOn6VAl+DTSFxymXH52xpyU6aMqkA5s5rHwsMe2RF9cIT0C/LT5S4BAFdmtjCXI
NzxUuHmIdUfnFAT+IADDjyp2nAsNcd5Gb0MEYfb8QI4naqxSeimx1YjG0MUEmhgC
K4NZ2eTgylv5hpeqjKpDacIqzfOixnK4kzwYasiJcFPzPE0knpJCNOxnWsoqKz29
R7Z47/Hq2L9gQ3pOq/EgC1z9Mkq6kIs2EHvov+n2p8EGIa8MhoKVT6xbxv815tgW
odG7xRGwWeZdsvhi7bQNq6Q0iUe2AtwAT0KBdKrjx/qCOic6j1A3dC3ikYjVh2zQ
nBdlFkFyoZ7hk7eU3xxL6+IJgmYlBLzRJFjPz3AEm3oq7EGxiluXn0yqYQ5VRri4
0ZADCtF1Y8VzCmufrinQjwZO7wi/r43g0ppOvSNSHbiebwJRAgQXNstR68VfXzR7
3/UeISdY5iexfVrD8t1dXSA2clkuFwppBw4k0nltX51HMn/jtPMzes2QDD33HjKA
4wD9D8LFQRuHzP2LYj562pv51XMp0WASGCVsTVq+/2gULKRTSrCjxlJ2axA/c9d3
+HCIJXGUeBZ9UVbZVJ9LOmkFP6RdxyKFV0YTlupzNFpN5l2ocHAAGsJZ8tud6Tr+
KtKRF0ZgkVv9rltT/jwSMJdayOPtr5qK4hDF3Lmbbg31H9W9Pekrne/7k22dwOpp
IKP0H+sdsLtzc28v1h9vCyrfsDub6nlvIaEnuJKAphBYeQfNjEbr9ux4tQScY2KP
BDwB0v0QSiVhuInrRqiJfxECTQbSO8Ts4DelPjU/LdMXuc7co7Gdkc4oDuCqFQrA
uy5/pfZ7fTV2MQj8Su7pzk6DLVCRYWTLqbrqsmV+BI8t1FAhz2ivCyxr+UE3lQPk
yAQ9ARMYlYb7fZCgmQXY38yUd19W7NgBahU1cdI/DKgCbX2ngRj5tl1wjzix5MwJ
oXfhTYF5w+e4x5mLs8EmfozyzucCUKJLVuwXZoZiAU8SyGtdRM5rpFmrvn8ZMd9F
9NqCaMAK/p9mFjiP0xdKdpm6Ol6V+2tXhZl8inGZknMBtyvXfzfM4PfQINUctbUY
yI45hrz0IiAjJVJEAwFAmYZOICtqLrt4cYssf0Di2kmxBmhakcso6dc1/KpJNLaS
svxvMctKsYeAz5PN+P4d9wii+tbvLfp5F3gin/WBuotpeErDEi4BRmAZXwcXJMgp
X3f6tMdfzCU7WuoGzlRLOr5XdCXE/htHCg+dvb3IWhnc19/deg95PhCwRyCJV+1L
t6ojPcr/JQ5kv5Y+dmerdP4EVrLpVqRZU/CoMemyiMsbk/a39hdaNRUR6s//WZEn
VeQHP//+YrPyq54jK0SOMM+vB2VuDBRiZzgoRXkHN9AJ6BFaftZFaWEzzmk2K770
OL9LSR9cO0y4zPbfouwqCJ180lQRnKWCtUiwmHF/n/81HTc1i/MEaV1giW6nUcvI
0PLbajMhZFa3ybIvVTOxPmSn56ZDOK9g01ilQrszwgD5MCZLiK6hfGlljmD76mJ6
oRvtQR1/uMPLJcK1KB2QxttJLs4uQgVaW9Yz6b1xdqCP88vGu+hz3UefSKr8jsFr
RkoxaBzN4PYB9Ei0QEnG3Vp3JVq2J+fvYRliw0GcnU1QRwIWhfKSLUh0tuodfeKD
tkEAfC3U0eC2dBH39fqXuoPBnECUjZa0IjfNqSgauoyVUl+kNmDIFZv7LP3ittaN
bRzehp8nVN26bM8vm3350G2GfZ7LoAMvDJf4EOl2HOTQuomwqpqbR5CprK2WqoYJ
YO83eIoOsz+raq9igROGYZ2tbwj78sJVmrsD2WLk6qsUBfSSB7uc8oDm5ETclcXB
58EaOEUFJf0QToFhCXkM4c0lcofgiNBDNS8BKJo4RWPwTlc8gHmGZkTvGf3RkuHn
XD5Q4qvnOcw79JrM2N+cMzVJ8cQj/UltsWTDDIXRfSaiafNaM2y5grRzutqJ9Pg0
//koNzSauP28Qe3DswvTbLvT/hTzLBIHSPJfhLCtHn0M4BhFRNHHLZfiZJlog+IM
0bWtT6grdqKqaNzmoNkQeVO0Sk2hYXiHgft339sXIRlCkCOyB95HC7mPP3Ejc1f7
BwOOgPXbYJpT6ygYSmkFbPQY8zSvlfAkmIo3626qwk+c5tkDxzVxoP9vXfyBzg0a
QkRfYjIhGbqOOpUpILnTtwTZiGvTgtM4WPgAqpywu90vws72OoINhw1AA2EPvqor
SC7wrdt5Q8vfeaBr469H85IEis2M+kKI4cwOl+XPy81B8InFdrG6BurrIxhHZZtQ
mwWlWQ6D9/c9VTA2YrM7icbGP334lK8va0xjpnn7sQ3oTbx+QzxSj/RDhVd44Kue
bqm1fNPBz/gIZUCG9+K59HacoOaYFFLRABnT50nvZUg9Xes++S1DR18i2Bywbg7W
InZfelDJQMX5JFd3MjLoRhINFh4qPhqmpxBtxDG+eLFha2OVnqlBm00MNpyGVr9R
zuqLRGeo+ERKnr1WJAQs+KsOqy5nNbV7oHikxN8KbsU2j+ZpTh1eVU2Ns+TjMMQz
TqfTKcP2j4fdPEpJn6LRYqPeZ0t/NgNirz/XWdHahHEZvDsaWBohXBBaXQIstEfR
V9NJWSqZiIRer5J4/R47f95kiCzX2StP66+gPDFE2mYENM8KUAVyyB3AHJEImgna
42mF4x6Z0rQuc8SQqelse96XG5BdCEXMsFVnlXd3sdnz8QWLN57xnbU35XZmevQd
lPlnvKwhf0G8ukuIb/0YE5UwNo9VmkiULtRU+IMA49Dj+UtCE1ArOBl6AV9boLdl
cL2xN67/AXIbNsmai7JbDIfQ12+oDnteeTX3QSWpdTqdjF+VlZfWGrJeGSbaXXFH
Anns3pOWiCjmJExYReBJMhj7Poz3jc0OS7XPtCuFZY43vgLngjEMB6a7cpSVF70f
D9ao1X8AekXUajg9QrkDa3Ps2faLjTrnzV+0gC1bOXmsDr1uXbq63wfs/h9AYleS
yzD4AzEU5YxKgxfgqHi7BtrEtXUiaD4z/WN6DhWy9RzqpktKjDzrruMQWAVvUoiZ
KqPbL5y2GvO35P1AxI1lOG2gS4F33w1hifEgHpqKiyd0R+N2RDbhHd0LOR3GS/fn
BfMV9b9RfFR8Jb+oyNUcI1HcpR9xYeW321pUO8YkOFJ7mTiqsTcXEZ1lCSmxt0h5
k54XHuMtxHOdBZqxbqEPvQUQZVO9rv8eQwxr9mHDMx+dkIDqJ1fGRT1noDnFbm7W
YYf/h9+xZFwf1/3I62b56W/7HHCsUpAswJvBLNndrs0ScXChgUH9EitBfvYAdxaW
X0yfl5EUwtR2+XHskPQq0RxnpELyMniX7R1PRr+SyZL2/L4O3atSxcQ6zCwEtMes
xE+Ji04hX+iVRfYXf9UV4US1dshwbvXUspNZuUnZbxyTAIHvUDPOyXIykkM2/O39
28amgALCY+LkwKVuLZoO52YGLX8SjCH0U2U745htHVeL1qbBPJesI2QnSwnEcOje
pol1lY+AiaG/QgHQMmrjK/+3t3ESTB3x8vKMKDkLzw6fUWW/0sbp0JcJEoXU65z6
NYZAeZnp/fEqWxmKRLXvX+AFIEIRlNwHlEMv0oAVN+mTQQpvoLY6WYVM5ZO6gDvl
7DJUQiM02/trHH+uZ3noMY7i9DiyVznQrbx5P3BKzjoSuR6EKcUCMX4uP9gFDwe+
FavqrzLD5l4XmlR+Xzkuofzh/6/2Ia2K9s2ICqdUwOM5DABBdFslwcHAMLBZoE79
8NuqaLvnfQ2Hev0o7P+LKKNMtCvOS8mI5Bq0xhLjIr8zx9nw2hSvtfswQJNCEaBR
qFPeXIeTMnwKq+mHPHBLwuVAxbRPgKiGP5hy/pOwrQ3hIuQ36HMaoj4sLXMwDq0r
IeIxG3mSN90hGXm74bcnCr0PPdowleUtzAa19jtqwLnxLMJnVNGQiesMhi9g8u3U
CvUQDyFGXPXvGlkTIoiFKiWiDTHNcmAwq6kmGdzdWGTFT/a6KysrdpYjmH6yktS6
yfRL1RpKDbOmMamCfGZrh9arqMYCkcYNMzl5tHOlrWFmOQuGc1dZspe1MAHEd7/8
Er5/Cbr4H5+1+9+ALLm8W0WimDBFuLEtEfSvgoCDw52hlhq0VN9awlTO17Inrfj/
FI9dAIGAfe7Hsr2Dspn3wY5Chf4vow3cF2GqmApwM5rd2uUAFDJ/T6ofFg0I901t
sfUYHFkNu3hvu4eSqdUX+f+C6xB4o/yPcZb0R4VEn1FPLuEToqqwORW31yFa0vGV
VonvatUJT9ndXSD8waAM6IRLkQs1j4IuLe98lUH8DCw6bMk6NQqFM88dc+sm2suf
zpRs3B9oNAO75f8MSnqoRT4DGQAiVoqZKveFb0jXV91gLx5rKdlc01ulRIg4ZlrC
y9qD3zM2xR61GMdAX5u15Zlep9jlKmp/LIVvD50IL8Ar1Ev7fqj4BxHswxyifL3l
g1u6D+4YlLFuk62vjvw7WEHLlBC9ZKzfVf9V0E94iep4SvC3xepw+eSpGNTdWZ8t
gH0+NczdPIPS4V4wL4OQcyMjb3BKQlW9vckraAgCOwnsu688U1Q83fTLsdtbmGZ2
FKayvKWSYnTBOe+OdHcjU+N0VIJr+j5pqVOBBSZCXLtPtBK/WH/Jje51zitmH2u1
fP0wOWkm5JvWya28Tb35SDuwWUQZBq8AmaEgc47uG+t0Ls/1mVYQ1ezrgxOGQ0iU
Jykxr6WldpwpTHWrUEEQ9I+CzQbb8IrtJtCFc/Da4Af2VjcSM18YhzrtW5YEv1g+
d4dHHIbl+lXoMXMugtwMznSa6dIzM1yxFSuN/UIAjZDK1k240hFb7E053yzXpsZ6
KnZANgZeg/e5uW8KKh8mYPt4vGDfOS77GkLiRDshO9w4Se1qiQ2mIm934VtuAcdv
lBdfj5Fk2AoNd1dVT0H9N5a5bWMcDbcrkLgZNfQgBVWtblNDB98kUbKo8M0UIjUU
6Thph3HChynxXczmVEEPiEfXV8VysT60WHddJasVTQ780Vof/FiQ1Vpd+gtCQ+B7
sjWXD+YOIY1YfgF+oWex0gvUtI/Boj7BINrMNhpNIQ0/JSvcG69kE1Fdf3+n3/fo
c0PvcMNWh5F2t3g9O5sy850CQv1vod9ClTvQPQ9hgGJaVIcolW7Nm/6AMPG8VEdB
7wuZKeQ1jR8dhDYsZhgR/f8jGJ3NqyeCCeYLyNfpTTvH4lzHl0LI1BuA+LFo726/
JGR3pEnitqPr0TVFxxkUI/wsbv3RtutbGvm0UsuDbQTaFPo98Cc3iYns39b9vcLf
tiCF/hSWj6665sQTfs2ZZAtFPO1GnlBK+r5yBYiIyH0QPHQdX0x1pQ3CV5HNy+j1
/NzJJgZNVTJqM4vmvkCxQxuof6QukEWmXCPW6EuAwNAtFOb1gOBWyxdWtv6N+Aw8
yo8sYI+FGe/skE+fQFW5/ZE8RrFhhZei/EBWzN3M5LFwVYZNZlf0SugzJuMiXjBK
XvG/+TaXjJwbPXApDv3pO/fFWLrY4iLTekuu3x+mV/WZLwz1+A166fdoqhBx4gtz
QtQ/GlX+su8F+nkHXKLHK08heYYMQHY5UN3ev/U/ST/U2EzSUWfBmDlkny7gmUuc
ZQ5mXaXxhV6zAekOaR603NUz6/EJzgvUv+/kMq40fv68i6xFc9L4blug87ZznQiH
zm4WZoAC/Wh1TZj/1dGhu1Z8KLsAkwlmm+MTw4BOm0bb9XvlrdZ71lpLFMpf/hBr
YviYQ0IW3XOr5EO2DMS9owgNm2U13pnc7JkmVrjToloH894yD2xAIfKQCbr5xNjA
yxIHaQ618lGSmzOn89uZRlOuyRUuBpK6fdBymB5y8fvNV6IINhj0rf+4KX5rPfXi
yPguHCv3mYdvzXYqYyPGblJkMBZ6h/n6LijsyGUL0on58872G92WsEY2RkCN28+V
anBvl8pk4dFBqoQVuMbnagC/HgtYL2zML9PZ/Z20ggZWtv+aVWuBPFT5gkigWo+h
sgXWClscw6h+r4Ir611DV4Q1MiJZ0rODrb65Pak2bqNWovS8hmEaWpsMHzki4ZWh
iwtkWpEKQEGd8gyWqnGA2s9sSii2Q7+BvTCfAZ7A5jcr+XjdAUsZWaSwbuXR5iUW
i6Fea2/kjWerT2KWo9/W9iO7VXXJRa9VplrgcWr2Qw+flUD4ow9fluXiB3KOvvGC
pRbzy0Oj1SQrauYmxDdpBGibg8dNCRTu0ahm7N66cRdg1XDX2lWlzOfhVUke3Tub
68OxD1eX0n9AApD83SmygPBA+jMvCQEoCJoAZ+EzYFrab1hFxwyX5M6eY83hTvTE
7IUF9kkHgZCe7uYFEYjBVpoiZgEDn4R7R8eZz1CyowWcyViNrL0daeO+GPlLIBxA
zIKggrcYXhmmu5nDCXIwNnprK6w+ZrZGjmM6k8lKZP3t9v4Ck/V8WizXIuJBXurw
yWulDbNuKEDGzisH2gDeHkd67SNvxWoQDotJJUMl2Q4WsPqzW4KlEnQXF5WNbv/4
EA2810byj9ctK5WI13i4amZxcfdVZSLIz/3Xy+2W9dN856ivsxNM1+VWHbQUwXGe
3vqkExpExHU/A1Iy1pCaehdluBf3hbrwgVIm772tq9QK4qevAXFeEIZuMSZF8/n2
/p8V0FbwCN2CjPrksQaeaWW4HbKQRqd0lBISUUhWcPkHurtSe2VLRyE4qCLhZALl
MUKhjwp9bWmca+LmgcgDi1WWjI/VQMA6gUWNhB6WqTOg/fhHUhsGlnx9zbS/t0NQ
1qrOjiT8JnZoyB8/6q62wcLVpe2o714vPJcGzkVOh/2F77ZRQayzz4hZFAiYX3Wl
g0BguVEJRMA/qiMFbTiTO6VTfPKIws0FnOKDRdAPACHLKVF2Za58p8Lr+Pbg1Ibk
hO6XHcI2doIjIvmabtNevvtJUty5q6TXPBuGVBZRnS3HUMgjfIXNroXbzF6QSwxp
vwXXg9c1v/A9Pil7mWLJ3mN68WAyMEUxMQ0QzS+QNDEcqSXi4jVreIg0KaTZSVrD
zrSTWfMlD8Hu4SMxdC0JINPN47/D2boBKjveIvdFJ2M0ewdtr3OZBfZUWgxXITRX
r/OdzroBnbXnmDynyuHZMo2SXxb3r3TJ5VM4cD72y2hCrYu7OCLmx2md+5VNnWPq
gb7f/yg+bH8/sioIcWU1q12NFBHwHT+0IEejkElqYcivaCMMXIUrjiySEo1aesjo
KYafh2YzwHtl21A93wKkbRw2XFrANgW7iZTDgRXqQ4GEfeoP6D2xk8tC3TKs7QMd
YQABXKVaA1v1XEvCPdli0xuBwJP4tOELuTK35STvWCi5gcnxwjoc2BSitYl+TMN1
Ztt5r1xS5He5HaUh67FuTwx7vcgIjz4B7V+OKQUMSWLdXnAfjebJ0mviayTbcb1j
ei5uSHaAKLfAo2bTisKHB2Fm0wYT9vQQJnT4FoVks4XU7Bhz0JZyRfOPYx8/s2fp
XUm3oN3difkOLi28TKZcleDlzIaN0K3LRm043N3AR8Lhh/bSPyJRcxBHPiM+tuF4
9C/LeAFqSEAJQS0sUSWC16IPMlNZg9K3x9EDTtKD8sEZC2f61woBH4C/T2ZjvOIC
8/NQ5Il7O9YJRHsVS96FpQbJLx5w3RuffkI4M48KRMHMJr5KvREIwjyO4/9RQwvz
3uBS+Idf+zIkq9Z3m4blo+uodfE65b+6DiYf+jhUYLw481/cLlYeNyfTsGZhNeaE
ySnE484x/61v7rCsihXwsrBB/GDy64WK8rNoXUWWDveLR+vpjNJAu9Z9E+ikrh/N
c7a9qQcANLEVLqRim3rXQgQLbYHGNxY4ttvBOoT6lquQLyfT9K+VvBCqEQQ9rP6O
2Bm/iBNwknbbZGs6BbT6XeEWq0+gSTUP2y+ktTTuAhhCDzYpFz7KLtYyHUGJpoH9
IT0YEJ98yf9PY7IYNiLY0/iY1PMZ37YTS8EdCWqI2+Bc52JuWl9pRymyjrchIIQ4
jvoDVY89i1n1j9TIiNMJEmxfo1R5xGluaInoq/hBWkVYozb9A4lbAh79JGjGcnjt
Cqe/fCW3929iYOsOhkC1bBgzlKfhfEKW2N30pdiKKGsk5urb5xTG2v63aoC93gFc
YKH26hsFUuYscHu0OmgqGojQ+PUD5R+U5NjbRgj9yiO6/8pqjYzhDaGR3UyEhCxA
sF16BbFl3U+psfFpWJFYAzg8mPUYIYkt7oYbE3D+YrC5JkGJ88QPmHSDq5MRLipS
zGCxK2B9Ja2Z2iQTniwIa9WLKoBF7PF023HHF8rKPemuhIsg/Rc69UVlNWjhax43
tz/RtXuZK4v5cCHKdogmbQNDggW9E3hC1dIOFSDppfITfO1hZGivRSo8WeFaMcO7
BVrk9cdAVa9UPoFJvhvIQ0SH57io6rawsZOSviyjvdKgkOPS2VkHm5ym37n82ZVu
5OQP6OQFJrxf775jbp8o0Pr0bmsqhXU8P2JpWYIC2oaCvuobm9UeoQlHAEjth8Ws
CMa7EBrDfok+6gmpzEerAzCJh+vvja50GL2mf+JpKcWqopsbq8uim5FU0VpQwb50
ZXrTSVzwQdWIRDpQkVP+oq194Ete3e53ajdVW5wHpyhACihoXzWP0UOA59D1DcXA
Rxf3r5dKVLVmGyHqvtaJ6aYm9O8HUUAGf13+tJR+rbs9BW2b5o2C6NAYGUuOPpOf
0oo2FU/LhIUxZGvSd1/365NpFKzyKpnrTARmwz052QqnGbH/8/SbT9zvmfRPilLm
UM6P7sxMB08MmGFfy0YE/5RXDevnc81kRFUAeiYU/R0WVRBQw1rjR/r7BY2TE3hs
i1aXiElBE38i/dEt1CJXeZELjAgQG/VnyYTqRaIABmqT/qyzJRoiFJ942nsWj1UQ
Zgc/58dJxqY9MiH18dtqKcZ0Fvt+fXazsaoBlgAz5ttk4nS/w6wyM9k+hDt9DJxv
Rwfr+K2lmMa06gi65lBAQQUBH5ixnS91zaBcUNFiHXe84sSniSYs9fa9Q73C8U9t
WqMG8Zh4q93B/ewRMstrf08x8lXH74LqMk9DIax4IHhRMbb/su1/nBqQsNxeVyxD
IeXzIFvb4NBnVmBa24RfZ3Nq2XxQOkmUC10Rn2U3aZdHnA9cRiKSAMbHrpCMUhV9
s27uWhE8oANWz/AmmxeGUdA5a3jNFz0Gx0GABusIdbKa6+g6oQRlq/WbeNn9FF8N
Dn6vPHBFr2ryz5pv2/2Hl9fVWOKyBpVMeVgYOMi5AReVmUCE/46aoD1z4s5d0ZQ1
e+BLzSkLDYZSwro/wBS5cAhQ2VCyGyrBT/rpLGBjctXbcXCGTbC/Z3DSFTR6OZud
MIxVp3C2Tm0BUdD/DBhysde0jSnP2By1Vnwpq3Sz7+dKmDKhjDMRSr/RpnFhWeav
IMOcAGemldWJTlJezuWb08SQEuIOvqPXSMPkbPOY4t4KhM+3riBMGjz2n2CzjN4v
877LJZju73KEURQHZXC46pBcY67btJjYRP2HkU2iNOmXM7btC+5SOGEaPgyClQEu
626uA8gawCRtoWN3v05JKK3kaGE/SoPywAzZfH4s80QuYl8l/1uRDMaLqU0uK6sw
+sYwbuTrPU+xOEmiZ5kjng8Kue/JaMSJ6x8edoVbBi86qxRiHSLU76vrdRy+cZFb
LmSk9o2N84qZhldSTHhOnCtubyMNsqLW84Wle6LvXePdOxt5otbQSwjqoj3hvKxq
MXaPt7iczsjHspmhnPsZm08zQ7+iTFGz3xFHbejv7eG1BZJkKW5rxTrLkDZkELsb
mpIfeEjR+wHmHAMOAGv9+2dCGT5XlDSoj/CGfhvgLj+Vt1mP6Hhf8T3qKRY33swf
I8OfqDRPREVmDRoFU5WaeaTKo1imbhw0ft31Ca01f/skU+pxvPYEYo9oP22fzuWi
283jW2dRdrm4KpCurXskcp/ESup41/EIWqReRa8T3PYl88BIIMKhtL1PmKL7YTlG
5EsK09n5u1kRWGnNQCMkhzDjN1hYgPPDTPqK7nao+LrH135bCr9jlAkjaSUzgAsV
rX96h5sZT7JduRcqaBnUO/TySUHX82nokA6ZQZcqlZGHbLYVicl1YR5MWcU9yweo
UJdXxucmcsk59LXYAb2rCa2by9kKr1iBBimcAA/Q8WYxiuHDpF4ON48TQCVUKG39
a8llT68xQFQh+ku7ogdqgHAaXsmIQYXqbAh5IdtQeyIrSelwWrLDj3RE7SoXjTZ2
R2JdGpMeFZXSWmPocRMun2TRmW/1y5bK7vFUxrqAFhnoKhNtMrF/940gsZXGyyDw
rg5RXuNdjZGCrgNnf5TOnuldvtXtsTYCxDsVOIbCKTBn3MOuFm6yzlIJmffM/tZn
OcPFRa4zlTimCxlM35SdiFhrO/2POcVpEG79nR9SdhHY4mG2zv5kxX6HfcTcPJLq
nvu8uYTuAa+7j/ufP6kBccpZ7K/7I0DIeJsBwkovuOW7QYMp/+eDoHkBgQV9BsGx
in6C7lQQeWWdpkgQ4G26b825TqrcR482nyLTAzvnvX0xPxKD8wSvrcSeX6euM37t
zlR5PqT9FV2Too6aRplZiLFexTv3s7CrhKnzJ0k+tdKjdVNlJjiUH62r0ryHHaHU
Qb2INHchgxnNyRDFqvznB43TFdIiOCLQosP9wj/ej9oZBjjqvCdwLjYF1sNh+JPk
oggyGpORWtqBTVBT8rXO/hTKNtr9CGUrsGBnKDvMoEaSDEB7Hnr1/bqmFp6iBdVe
68rSa2sZSKTWM2gbJYpxmr7fS66p7cxVR5/ylvv5AFPii6YqD3n9rOn+eCsoTO5I
JhfCwV5+OMehncccLBhw2mXCgo3FUoFN5Ker6ZrbSeWeZCRrOy63/wwJSVN9BBw5
WUOdhJbXmLji6fN4HstzdrOFGh8AquobW5zRYxHGsKb8yNuZDDXNXoiRLagmTtrW
j2y6+k5tWH4V2zkjiZppHnzMa3rDS/VVMViodGGSbJxRJ6rtpqBjMcglIyyzW4Wx
C7UBMHf7ND8ozScu2FgMnavnsjyODfrRjVjx0aOpwYiz2qyCOV5vd4jHBViGAR06
beGiestT0MyB8A5HYUELJP761MQYw2D7NLnrZsRaHb2MGWtCeacv3JH+SFjhvvNC
HV/LKPuufz/WAbaE4CHgoCz5MOIBBXr0sWSK8h7QTxR/IP/LGb7UX/3nn3kBV/T2
vkqNmWrJPtGM+X2swiyxZdN6GR4hG8pLv+pxGkS++7kiXBYpcFAOz1YZ9lMk9a9s
7zcqalkb0uWeMPwJE/whPOfeGIn0Yb7FjnPUKz4nUxLSo9QDVjNvuiUgH/x7uLL1
a6VrdyTYW/2o0PMgA5tLgw91TB23XaWjvv0I0ZL3BIsQSPMTg4NAARb2lr4ZkeHN
AT5Bsl8U4Nh+aiRvKtVYnM94AFHJSA2LRI55m9ySuvDs39mn3yKaXR+Um8BCogdo
08RacgLi9kk+RCgBOrKS3siLyNjw5R8/VQjxHiOnkvLrzC81ILeUFLhFXRxDQGcz
zV6gwMQI8YvnG9V6vpjpnB6PVWpLCY8EmuV3AVrqHCVeye5IUHeyGePnvCpw1KHS
EOB6HMqHg5x2F/5L5n4+FtIN7ekoOV5O9EX3BJvpu9zKX50YnAdndMuSV3+50K2o
FW2s8twHl80TYimrnAcSOGW3BIKaGDoEhX9N6pKmbEEJpUhTQX+wMX8L8BmGjWSn
GefCbc+UrZu9VUHWDzVka2xzUDSdicO1GS8Br4UFmp1hNsZIN+3PjYt5p2wFW4YM
V25ZLZOLPx/+fWgJOjE5gCCUXAlnQECTPQv5909wnxP5/FVhdyp6rEFvLv4X0zxh
IECIMlUCSXpwURbAQmKdsDVVN5BhUkR8fKCqpZS/wftxg/Fp7GE+yEo5qq4DfkLt
18k3l163ofzNFINm6uC3hE8G7Cu2jraJ9zWCiYuo9NhJ/GIuQZAeHyoqgWxA7chj
LpRixt/R2GvWp+BzqH+b8hva3b3B0rruhQ+nxUlqTDIjOn1Mx0nQ7QWmCeywVyAC
we3IcLRxDi3gvNX9uRAMxDPUXmwkt4hmKBmJeQgD4HAoZoDdeMFmaE6PAaMeo9pD
CZ/uoiRsosr5J1qxbzvEUSA9fDp434A60+7vBVP6kRvYMtSZJbsIjV2FiV7EOo80
1mnRmf4HpXubXTXGxspCWV/BLj4iZO55XFLbMBWrt/vxrxzCyLuc1R67y/zVoUPE
NAIIWcxPC8OIsP1ifLevy/ex2qkhmwD8KdYQGOihXUFw2jKxL7Y97SRlYDCzGFVj
728hvltZPJCoF600GcItXrJgbFS48nh/8Dr5D6ZEYFwF32UzO61I2NGcIX7GWGkP
9Gb6qEUoJRwU5xNokabqDHMeVDUQRyY+G+UO4fhSb9coe9IolOMVjRCh1035poR+
DJIlC8BGPL3p5R+1S2IoU30DIwe/rPzp3veMeDrz0O1u6LQiNp7rO7WUcSgyjB3n
y2jxiW4WKf5B0H8efTiuMwxkBOiEsYtGNIqzD0TWtlPepHwjun11WbEXnVHaN85P
vARYUUUrhF4yqJKu8sTVko1we4m8vNORQNIiWdPBlpPqluhb2GhthisgFVZjAPgJ
Afg9h0cGpSwSyPCmeWQAXoHMMSTfDuBWPdmp6nF16tIWux8s4AXfUiD9MY0jXJnY
J4ZESWZHLm0yI5pOdy12v2lN6tdZixhQn+ST7YDsbVaEm/50ojCEUSM/FsgBbGlv
Qdt8/qqzKhc2sbzdhXCl98J9KXxWvdTBAUDWBYQT5j2XpRG1YZwPKyCIHNlT5iGF
tzsfej2xLh0F3/yhqwX7jvEYvly+G751bjMlUhkyMUnHm0E9gkd7HjApDtzPGaP8
mGNSa34sojlkcVYP/x1zVtcqn7TCGRAMD14VkYNbA5QxSh9S018RJnMDAs60KX74
KVJykouKJY/4dIxF1fDnAmXGezbId535fOYjQROmJdbPSicBHLxbhQQ3aUiE8HAY
vq5n7gB1Bd7tVVDso4NsGb6bKjhVu+VWBn+BiA0MGIYmDt/eyDODRZUh+Ks+4z0t
NhcHUJerjYjhfwFWDIt50LjyPjmBaXFHP8YE43u3IKo94HEabHOoG5oScySVhj+E
qBVx4uWmt3jz7k/AXmrUEbLpYSaOKa1z1uMWzGi8mAnqfEGgSAa0fy6JP4iM03DZ
5FGP+CQpid9+YX/Z0/5TyihY6H/PQOsgDNVrdTh+IcsSPHBgHN4t3Byk0md5/cq0
8CEnPLSScb5Iuzcoy3Hrtctt0O47utoX0RTBRaEvyG3ZQd+zFw9x1ZV2jTiI3IGz
kgssNO4Ftjh4R6nsaYf4F0/I9sjdgOAbMSjNMzMOfBEBQFkscrBHfxcFO5GYi/HG
tqDTaifJJ0+NW3aFX40UHh/kbo56L/ahwBvVEz8ZOkLO2oOk9hQRB8EBXIZ7ckPo
Jigr/sK1ohyEkxcWrnhv8ekE3cx1wHThmD2qiG8LOGb34+GSgaZ7qJquTnAju9Bn
ZS4t9YSNeRbFOX5hTL0zw3PqIdWVRAXwLU8YbCAEvVQ3seyim+D4L8EA0OH7Yvfs
MqoUDO5QG8DVa+52BZVGEqeawHaRrGTQukmIHTwkas95A0/GGZ8lnfDrZRNKkeg4
R9Iar8NlrcxIAC6CZrkAi0xcEXFDhTDIbC6zs9lE5BYJAi3P7BDqnNIAxSX3IXvP
bMuWF+Uz5kkmhbOi3hQ6MmPMOlIe66mU6octoMSgWfdToOdLoSW0AODe6Fh/ogGl
O+etpW46M/0v5DhJyF7iDt4+ighcnrzcLrqiCVlkRjw9DNguT1ihbwKsWZxy3g2e
/8/KPms9VWW2j7dK/jlpAPA3PQDmHNzEPG6sov63VPjlL3aYo28iTNZXMGfVqmhF
WTmNBU3JDRlQ8x8Q4zxqVrJgDyajKpncR2PVJ+J3FWsiE/5OoU+y3yWH+iZm50kG
QIOJhPTdccsFxpJ4wRurwvnG2X16nUPrlqonQGV6Riq1VKMjVlkfyGcHv9rL4CYR
V9RfGcqbFnqWb5NdsWwPGhI05JBl1g/ZxLkb6izZJ1tMHouLY9UDWxHJI0nGsfdf
POoaIHXsDm3Oy9EMKykdDY3qNjdOHnTnp5ZFtTuAXFnDQXQAfd1iHFM71i0jssOw
xeru4X+nkXptGJVwD9ScRukxcHP4fsWlWOgvndblv/mGkND5PMMMeIlvDWfVO4L/
RXeiw7oo7cx+oN5QBZun4uIYRkVHFN1+iUkHyXaljw24vFy6kkuG9w473kYMUn0G
v/BgfcxsVf2ewUXpiqY6qziQCtjLMemYV3EeX03PnR5/xQNmGYdsWbzHBNZgewvP
rJBQYbx75JKZ0HuLeHFfCLWUzI7s1EiS5KddG6zNXaespCDNYJ/00n13lZyKoJIz
AA40JnGaWMpYGtPlOl5DvguQEN2ZxKuaKZOMLAY4Ae5mdNBTZGL7pW+WT4jsgwJk
6z1WK/iFMaZocBLjMD2GOm3RqKI7WT2YmKtHPvNEVZr9D3yPf1H5I8Br07I9zWIB
ufZhv0AyBguifsytjyRkXSy8m8SYdYGLm5xXfpKhUwHS9RTxfYD/AN90T7zad7dV
dmL+JUFdLT+GortE9hZ6MrZeLmh3cZRoyhrWkoa4uzIFejDOJfgCH9Nj/9bLVgTw
BuM6mcDZrlv5/qXgIO020kmaietSE8BWKNIIwlqy8ghz8HD3G1IW9f5/a44CJLjB
JRRmfSEmHLogCgtEzEXYR2wci/jY5wsDoWE4nTtlHt3otLxfqwfE2W7WQ4BAMO2f
80U6ea1z5pYAcnjveYIcVq6ztKkA9Upokby70Zb+wrYa/jAB47fdE1m60WX8iFUe
cJzW7qOjlDWLOugIHvMoCnDoOmJl3VQCmx9cjbaWZbqXGKpcK5KIl9kNv/hm3RCe
azRpHiuE8Rf8Gmg+Tg8T9cYl2DejS7BzoxPIbh70uc7MNeewd80sm1d9swk67RYI
FXUES/1K+2JwlLGsLJmrXAtm4ZGBbeDdcmaEbEntVQOfGQTcawWo5LNShyWcdaes
7zSmbM8khyFTOLk11Fao0qQo9+cRY/x0jlJoUMSF7kJgOpIDjolyKbNA+rS9V+R5
M654QYeU0FH+E1FoUE1ZWvyFdKL3jIkjKSYfKAHaJeNaw2ys4zKxO7gEYJ/Hkj2Q
frVmIPlted6po8T2Hz/KsC2g2e4hMQdaW7lPv50ML84d6Rl+wPb3VuIA/PDwyLvm
A8hSeEuiBvqhVe8XQry+hbAB8qGrsIJMdF+4wkdtdw6lznkpQhwObilp1MuP+Mpx
MIL9fjlTPYvjPU3gF/3zjU0+If5LKrT2loteECHA0wqjwBD2h4EyAvmuiHfBeXjg
Fm4HKrRskUuG3ggQbhNKK/8F4HjzxX8Av1TSf8iqPRFeLjeSbTOke5ffNYqtezFD
1kEyW3vm98ffMLvUCy9CjVe5Gnck8khi/hC9Rn5YO9SeAU9zOao3aOW9gk1AmqRG
lFfI+bxfL0sAWTL67nC8hNpskSk22w43ochAwt/D/aZLpgUwuX/g82rJsp081G9E
kmnuRBYMWZr+Qnetnn9zZ7HqRU484J/HyK0//1EIs8jphJ68840yc+B18VOIQPSl
kjz1Y68WrS8Cp6oIS0pn5azQw+0zLQB5uJyvuJ24zHN/i8UWYlX6PyE9/w8JqGxI
my5Enj835zmtpHCxQGTely5slJyNNRIVp7+V1cIHlbxmaW/eBzi1ZkBGsrvDvAsr
m8itleA/vtQlrq2Pp4OyDzSFdeDwLlXg6rQ9kV2bRC49g9D/8WR8zIvolR1utQYG
tB3zGyX9eBlfTriMnxTZxWIkwVh2dhPiR+1JiAj3rrXZhyIeJcGrSNGXtsMvc+QB
Uv9AEk1iMO1QK48RdS/IsJeeMTF/n6y8f1KPT5dBP19Bwbc5W+tyvEyeY13Mr+1w
feiSkr521sT+itBKaT7euSQf4iRccQxabXtBBDBhtbyHFkTZk/RXDj9NLcxvYcmJ
t97mHDxocNbnr7MViqk+x2OoYJyZG9595tNyXvhYWhd4juXyZ/o+61x93QN4pGz1
/EBSynk1Tts4x/6mk/YZO0GUdjpNAOKM2NNZ6WBXEJVp+tLkxXicpysniWrUg03o
dtVtZ+NXU809aOon+Cc/f14i6aX/zCyrHvlEJ4GQ8pnfCDNJq9HocgyErftXh0nT
W8qK4igZTpobRsXkueBpP7iF+ONd3UW6GoIXn/zO5zG4WpjMfZZDtafZEXIfeCdA
mr7KJREHhes6OtQBm1jdTHu2VuwGXIauE/Y3ic1lepv9dulJCjAcHIdJbPUjo+bP
gOtaH2/kryf8lasj+QlHLkrJrGLkErC4AXAumprIeVOBvaADsCW+hwiczGlJCxLG
AXRuIkK4IoL+XZCmt1nznCGY3QjeLRCCOxPcBAtRBGEoIY95+FjQnVAYNRKC3HOC
a9gdcHJhFYJLqaHg+DJe3lOO/ZAJPsr8dYJgtgZbLUSMaYa6qCQEcvGClkqMjKCP
0mqyP7EyRAkIrqcDLZd/QM7YtQTgxHr/3kSmsRb3QUlrCNjujgTklCq+jG+UE8Jp
E1VP+2eUh5pV/h9HYNGSC6doYY3Rqk9LRbdNGD1IjliIdaOpyOmtJyX8TuG9KhjT
E3f7xY9T8MsJf9ztVogSLJOJ9NH2nXL2gOKqPVsS9VgXavEegrgZ/b7WSUg9DqbN
qTwaYls8XKm6oHORpQAcMVMffkeAPYYweG/7FW+/4Z3c/XbvMtspOeH72/eBez8z
lTGOrtn/Ax4bBvo0c1zn0q2gqruasbn7hh5Q+Mk4MF42WIFzCy3a3qhxuSFJHMYF
WB40JyftC05Bhgouts91QEZvRLXt4oTCOB0iPbDAUsh6s5vgmucMtnERvhykgaDf
anz7I+VQrVC0L+NSocwD1hGTPtiHcxVC6XFGokMOeS//xkNfRzSbE9AcnmsV8SNl
dH4vXWljYQ5zT38J0Zz19oUnP5vgNS0xMolBpcB8pm0ZSZhYgWPrANWYfOlepvSI
Ib9vijoJRnpEXnuMO3ndR80iayov8RvXFHXIoimCa6piNw9FMO652EKMyb+sT4SS
Efut6UwpS6WLAxCxlojd4gDKF4zKpdfWw76VUQo37TfktBaUjpeKXxsswLcndiQm
0J25T5fUEu/fc+uTpCpbNofO9du3QDwSHWgOyYVeFPSDx8jrVgNf8ONMHZ3Pujpj
+FNkkUjyurpCThbTQ0xJDbqjvASe3f/7EGAIliqxikRub/cwwgDs4Fmus5JEOtcQ
Tk2D6GdNNSEDYKWQu2etTZ+Ivmv7UKAwVfPB/9wjVTdIHFrMhH38Y1dY6zVN/jiE
MBZ/yHciSpTXvxCz4j3iODhGbiSWPlGjrp0LQh6PnSgsE00c5GInbvhvOxo+e28O
YsxQEKurpbTAWQcs0ult+NzMH08tarLTgpLgXYk+PjQtVFhEZeqdV3h5ksBOsx6F
Q3Z4J2l1ThSi0Sz0V4PivX3Vrl6ZSCLo9abbAAX85A5nigZY1f4ejWtOlh+R4zIr
4c8qE35UHIQyRwgZLqcKMORK30LUVV1VgEtEHnC5nrLamVp5qcZEHTntMkSdbw0n
2AdLXRYqYDY98rm4EdthRU3BODSCmG/ya2uplNpsHaPnSpBqWGl4ymneHaRiVC7Q
N0jZRB/kYabOz+WOOJX/0zjJITuQZhRdi6d3zlth9ieBgYca3gWtcXLf82t08ZOd
zPiPr28pEtrCh3xIWIJRP1987ClXOr6hNSYg8PKO4UGooFgstYxkLe6vMXQxknVL
KCxzBRdUk4pq4ZxhJNReNtQyfJ4rB5x3avl47o9PCfR0Rt6eqT1iVF1p35cStYBm
CmSD3vHhP3Z4As/NMv3VqiwgEpgRuAd0zkQDW+AF2EuevwfRqFbjQdim2xBN9YV3
g/2SzFx994SgxaPgUinuQI0LE+6J5mngGFup++xGoTWWvsY4hpoOqmGvRirt9eBc
g6UwbA43eqv6N7crJKEEmoRVee31KLggFS3fgTYhq+X9QVemAw7ZhfZU0XoP3rP7
YFda+KDh/k/415szurIuMZ1z3TuP0FalRYds23uCZhZBySTCk0V9Ujsxmvwn56F4
1szpMhS9NibKdsQ6Plhr3aia5pMrwUFPuSgSzUm/iM1g8g9EosjDL7c1JIiAzwJQ
WSH2Rx745pnN/rkdc+lFmllkGcGiZtBnDCo0UwLp0P8ZscD4YkPvmvkUD4ZiUA3k
I0XcZOD2jjQqma32cqV1cbfMDx/PvPSw+DaK5/mI+cUKpriHiEq9r4052yvnLfzo
Iuw2hz6pf0SttVApNuiERZPcPh9W759Gkc2ly4wfAy/DDDW8VHbujAuX02E/r506
IB8StPEym9sraXuwV7JRtQ8e4P+tLfp1cK45HPmnEZIhuQNTO7S1n/eVMPXaKTgL
oCZhnMR3MqqaU/u72xovGgCd2lqjZ0xMBvlWmnx7xwssuWAEcUcl+JGF2d0Ayok6
ouMp5BpEdSPhxuZsViVLn6N1INTGIPD41+6ETit35dK5uHPd8/JXLUJL2YIlkEn+
qEs04+IG2MXoDXkpaDdJzbx4pmg5vth9lbrTLZBE7ACU0e7tbpESdkCx1heeGg9c
dqzDvpGnq0Yk7/Cb9rKahj9hi/ukx5rXlt1POrS71j0iQXGBtjlU1A0fWWnUu1gv
hIKS7Y/RQkcqv50WRyo+Hgsa2f2XHFPrbvchtzj6cRuFHz1CxS3Dp7MmaPgZ68Xn
YZ5/Ad2/x90yqBvJC5iJjvTiYUIjH67/qE7r+JP+KrP3YJ8wvQ8mQ44fdNWyVYb5
c27XjvOlsGZc2PRwHkyw9nBfxNGVXXEwlUp+EZy1XrShFomiwIvT3a1PDX3JW+bB
gyZ0gLlXEoUcNj+yI7L0spRMlrgKFutNB1cUbFbRM+fNJheAW9i7cE1epHrSY7bK
dB5JOLlah8sguBCGNy8xEglNqnM2TWPyCoOYxS4RKOssIFJlp3J5yV9CZcr5uxZP
xVxMCMtV8NO+4mL/tcFTHJ9ilT2944Ytil6hOk4b2R1q8V/weAwUmkXgEGW5p7ij
A+VCPdTQQ5F8kPYXfFdRrdA3Zpvhh5p433Rf9Q3/aNLxZe1lQvq5B3VxLHSz2Ew6
qeqMNWIgoPhQ8z87CzVm5J89NxkjncYUppaLo8hXghdjJDHBfhsjjQZZweyzK+QC
MBma+Smqrz1s4BN4f4R7pQTpbFREMYvBE0bOR0/Ky0qUSCoZw/oiyXX+fwkxT31G
54lFbPnIeM1ehXRJDbUHWr5VkGo4mbFmc0dGqWh9mEPyjnxdJHmEiyE18xRefVJ6
ekPEWBZAdftrh+Q0T3qP4EMS4OTDaoZiThUfWx7LlfhxNhWbIqYv0+gvSJNmB36j
iPKm+kA4fvsIaM5RKtHBcuDWMvP95gYtfArC1GazLTkDmi+fu+f/pMgDH5ZcplkJ
sIjGGG1ZdzDPyxJ2mfB1Ip1dnFlw8gje/RMJz5yZquUSoGKsIIfNB0eBwY+B//5X
2uql2K7cNbWE3u2vyzoDVBrnBWTG/Sg8rKb3RCIwKIgHoNharEnCXbnAX3SLUXxT
Nu0l5VwVKhoGNfHmIaABjy4o5lJzr+UZuABV1DL/LEcJT+XTs0XYHNxgCLDLG5/4
XdHVQ3fCj5MGd/jRMkt+e+DgNOgJHCbgnylyDS13IPrGn/naqFwiXUbE9XUr5yIS
fP72jJZy+HZGgJDge/Zj5Dl9LXedxK844yzvqE0xbhrD04cRn9YIPRZ23TNjbXe2
69Eb3N0xDIlWJUBvf+aUc1amHV+bUQzdxBcyzKicNAenv2r2dnQUzHxZl1ywqDNM
idUQ5dRUQIZHzxYPOme6mD+Kxc5Fk2uyqOtPoy6Oj5zVz2X3SZodaa1lJu1wHDAP
U8Ie4RQnWXMRmg9gaaAakQpPGEyc8DeEDwVom6rshdM8kMawGnZUS/HwQ/pQBbHL
KsHPa7GRxwbELbz6bTgz/UPg+WsFSCzcmF6wold3B7nY1mcQgw0GkPZjTEd6GGPh
qdKzq22Bu8vs0xi+9UG+Qb7Fto1E6ouIU4JdrojMPIHFXQuQ1wtzCj1Pu34/Gwxf
vmq4qQTKO4sFzIl9ZsrPSGISZBIvlpxEAlFFt2vbkw/UA4ANfWYyBL5qIk3vTkLt
671nz/cYJdgePtG8b0BB+j6k09ha/PYPWGyu/RU7JpBMmB04EgUAAk6Klg4fVuS5
jbVTzQ1HN07zaG8E/5Vn0Iygw49dwny5IrfPTQ0IOfosEhy9Nfv/k1MYtgIW6d2K
cTYvHtCnGKvlKcpxF0NzC/ecjIa52Ot1Lvw0dEFcfZrXa7xQ/7/MfGSUFFVcsKO8
yUjAgtpRzIhRysUgxurAkQXJR7uqQM65B/Na9tpQhWIQQPjqGHrmBuGhDF1GHf6L
g8wzf0645U1lEug9EWq0BWfFVXXneVVQYRa6NUec3qt+UQ61EOGpEmGWj3r5cSA/
7hKEPzRyY6+aRyISB7cDiKqSkxmveM7vl8N2XE3rzZOgB3rF3LOIROFXFKQLVqw0
GEoKsrjfvMW/F8Ti1lizx43PP0NuU1+1vBx1B8KU1/U6eADrrfA/575NMydUlVkJ
LLq14j9s61vTrwYN6Uj+mL1h8yb1NVQLLKZ7AuUDCpqAq5rGxmSkGEExZ1XZf3Bh
IODmf1G1U1gvj8r7Pk+B5Lh7Nc9r/GpQ9Ien/eLaCr3TjOr4mCe2uj/kHWswDNhy
AQa+GPKHgkhb4V1vXZjrGffMbFiYh6aRVigXFJPPwcCA3y0xVItv+LQXk7BPjAkJ
w7I/U95zMIUnTk+XQPoYkepIgmuMRP+1Gbn7NEfZgFoqG4s3FNVLIQrQR3UH4yv0
xD4XheD4ZXRDlBbgBA8p1pU41vhFRCol8joYm4EmE8OS4AE9NXcGSJaeXUCePg2g
pyHG2Rz8u5MI9RYKZ5DHHay9rOFk/P2/83X9ORG9lrHx6vH1DRvHox2Sp9V6Q7q8
/22e/dFm4SnIF/vchYtnScGQj3S6qebtBWM0FhxrPYruYDWz9ye6fBBZV2aubWmJ
UVEmhsBHZ2GlntlBPxzRS1kJWCEqUBxqPkoTEFFEs0R1D1M34ywuEhvEOUwpsCmg
hMKAK/k+EwYZMBtCdhulnuZdmgaAqdBroMam9Ld3mdbf/wlIA+ktYIa1z3C7/NWF
tz5DWseDG34yAy13XCBNBET/oECjeDE/i8YptNaEBAE8GHlg3WNNqihJZCO55P/A
pSZePmUVxOsjt8mwvVswg7+NEGQ68yoY+AXCoo99JdP0iW29uEFFc7r9CwdZoJh3
uVdf0GLEVLN9Cm/8eJvR7teeSsmImJs/L+gnZ5IdOwG5fGxhK5uWkf3l9ea4Jkkk
z3tEVLNnzEsHdQ2w+txgjs7ENmCCtHBqZae1yQKTCNgRB8BI4mbzQf7UJ2BZN11V
483WLphwVmJ7J7+lhyNC0Ggirgrmf+cscddY4Hd65la0sVCQc7/nDXYbgzB1e6eP
q38leoIor/5lMyu5pC7GKkxiC49YBj1R1/shXOl8ZD8/JSqdAsq+3v8J1Lubu0yx
4P3n+KKqX6H5V5EgO6Q6ByjL+6XbgxRzAEMPQSUox+dW3rhgZYw4nq+d2Ff/JTw3
HC4M5VasJWnl9E7kwkVcilsTAQyZHECAR3fKzI8pAEZLXTYd1Aup161ayBb9bfEr
Nm4Z/r1HTGQsLj7fpldrq+jIF0RRVOORrubdbKk6HWYyqyWitA+kTsSbPNERTYHU
Suk7IP8xJYNgXn+5o+BdCeFE73tL1TkzE790yLUF9MuoTePwAWF+xnecAAZElOuU
JnBXV7zma3Ej5f0YXyq7aQuqvPd60POEybCYYG5nGEeAnXSlFxgc8MtC0yW93lgQ
uJNKVpbJfrKivk6gtITrR/K6eVEqaaDrVTMgdVA3+wLgLT4eG90qAwGNCTvNPU3K
8I13dK6AlBtkg3RAJipaqtJuUgLVlkJv4Zhr07dBBngjGGjKS0uyAZtq6HSVusR5
322y4d1BUh7Pufjp90JQoiMyfd4bMy/KyWoxGHncoMfDsxsTmpwRfiLXXDu/XBdk
GOzfrR4Hz0pGedDlv8wZ6Z83RO+GT8ZScisTPJrRpI8swaot2HeSNCjUzSlLYPbF
Gx+fweMaMLBAhrOn2yQcp5Fm/C9B1KbYlElVmYwKa+qSFs68DWpNK45zmhdq7Shg
nw1VMEenUDpk65WZ44jrJ5h+MtoA2uZ45MpwJCm1IhdP2sUZEqOzQrSnTE0FX0LU
1D8Pr+C9Kuw26y0gHlrMIkoz2rYXj2k59qCR8LDRftbjCe5sOgwQfFdKHrtIxLo8
UviXVW9YAFTIrA8UP/fw7m9x+shQKE5gt9nbUVmhpTVMsTN8828Xw4YAx53gW8QO
+CIbYv8iIgwHkSE/bmuR1S7kRAAukZlQqEMVk+H6l79oT9OTscpDoG4i7ryPPS+O
r9H97y/Sk9EHvHd+awBZFQ6IW5FS7RxcBlo4o4cTHU5+a8csmNFNoIAgmtWBSTbx
/OXsaYojuPNIMOtGRUFo7OQ7wmkE4EJaGk3Uu8FGUoAc6jOZKjBUueUIH/XH2RaR
RiD9NHDS7j6WU5GLa/WOcecGz3HjijUyBjYXPARIi0r+RFTyph5KRvfJAA0QsCvQ
bwF0KxqwjCBqLe3TS6cWHPfSNU+RDcCMY84Cr23nfIWK8PEbdpcTBBtHybgtbUSZ
3llKlh+CPxEs1whLvjnGidk3+XT52k/OYc/VJAvMZVuOym7Cb70PaQjJdjj9xUAy
EU2/t49zUeCIv0LxQykOAgqD1DraLYbjztG49/IhYVonDoqCzg72ixpo6HfRgf0E
yD/Yy0VVknjVQO3x3fR7v4ugX9EcAkK9O2fYibKWgRGRS9dehLRvymMDtUjJ/fGX
aDOEMgzrVHFOfS86ZInV9O9teFhN2HJgg3y9lKUZ/U7va9SydkrdhGzvJyJR/mnb
Gj4kUJECZUxQnGK4A6pt4TdtFRt34S44iNvvMHsY6Zd5qhubLRmsr5gAGGCoO09Q
9fS8miIRK6mKvAl1ltXLAsxMtWnCCiYjGCfzGc31ATq2Eeo7X1NB1Diq2KuSkDT8
Ia0/Ny5vycBYB0VLNzxhQiffjLqT4D3K5AQn1DID9JOmPuqk4hgIPxOt4sezICB1
GbvLNvKxB8T+NPWDaaJqRfAP1+BPixu2yMOvRjk2pd2eGYS6sdTJinLQigWUI56H
L+//ncuRnx0vr2eyJcSZwQIXoPa6u8OZm+OJIIhFRi1icSMTLIcj+0MAUXL4e3LN
m1IHlMvQJ4Y3jpYYSTbx3aQVmQ3cwhWK9oMEwFZPqGvcGYus8+98KWWz/vbhzphM
Abg2p/yDwYhTibOJMmlnUv3XgQJLKNCF5WrLevD/BH4M0Tl5nTsBkEmh0kUT0NQ0
oQg0WulZ7i9IaFWuNlZVq5cm6Mw9ar+5T5EfkHBiShMkbUK8eyJ2+adbH2n0qC1+
RKcpBbE/gwrHm/XRKLxhGUF6ft3ZZkc+zdP5fWZpheGr0aAan0sP1Tmy3Wmbbgn/
YhNl42YKfcI/U39AlPmekgUbpIwxYzfjoJtsbro3TI7WRmi9nvBs4gCZ2J538JLg
8U9qIA9IAEF4HiRzwwG21Q8jHIoigec2gjy6anFamHAyNUIl8MdhORoeUKYz4NAV
jG+fNJIUYNW2dE+7ZkQUA0LgxaSamToDBaawXa7WZNpvZGPLNByF2908cAXoy8cD
dtklzvLSnY6s+o32uAc89QyHRw7KJ683vP9Gf6mW3mtBqq4zI23a/CkznQcE0Bl9
3I7AQXNbVYWyuSB3PnVqFNi97rHTX8oEa3hqMdZGhQexxpfRt6LyvrgkRr/ZTMC6
NZanfLLJitDCiCb6OIFkckKkEr3TXiiN0ofPQXlK+0lSlwzUNNJ8juonoHCOJ9Fc
Cn2sdTwXbXhZSAktqDBYXBY0PbOP0dg3ZrgwiYe6vtcdyZv7OGLoIVrwos1HSE4q
pmqQ9Ho51ntu+NTaUg3MDrcudmjlWQxXKlUBs8Smh43JAEuVBVwQWq47/Dgt9Fq+
elYCC4tHFFOvI4L0/FwVBd62frMxsXyADhLgpxascbNGfuAKYHZ983weySKns6Iu
oDJqPUV5zXOF+h886ZkoDlD+Fm4b4wvaC4Jr5uYnFxw6GlytXD4s1G/dNE3XPtRI
UTPVV+swzxQ5Ruw0aZBX63Tn9C397n5FNr0fC+2JkqViwidQXMq53K2Q13ghFMT/
35/i12HaZEHYXsMX/Er+WuW7PRHytCYARE0XRGkFidSoRWaMButGW+y9cg8x3Hxs
A85Bb+AkeGBelHF5BHbSDGaD3mfhVRH/mvSXZ2zxeg2kVckMU8BVTIMx4curZrai
rA/T4s6J+aV6RUPUruYRkwPJlmdms6ubO6jrAVZGhl+g3I0gds2hchqC/cLk29Gi
7NjEavg1Xju//ofuawpJm6bTY1ny78uzAq+2d+tPygrVx0yA5bvo0dJ1tmXk7Hxf
u5WD8CvkfoGLlYEkKrneDI+vk4xCe42ZRpiNBCrJnaDct3yxWapq4D8EEny5e67S
Kysb/bjMnCr/fRQ1PEorRAjGSIO5Lv517LfNt9/5mItIPQz9q4PFuH8IhnTFGOfy
hnusXM4sDK84AD3sg6gT4gshhmi6z9YPpjFg5CAAcg+e5HtZ/3LnBM9nV0ZhhBKk
HDs0iYBVKqZHhNoVQkwnSLLrkUQDMnrkqrSy6RQ5fDx23vU5qKBniuYMnnPvQebV
o/oYt5m3d7KBlkfigtz5CH+7SS+ISbwQBwxhykmTpolwBG4deKIGUZ9EBe+PD55t
i8/Ww6Z1rY2KfhZXXoY2AS2OOuDzx+GK35fjSWBAT00r5PUuo8+aHpWp5+TjEhVR
GBYGHh+Xl+Hg24Z6X6/+THZuYys+tA4BW8Js3TnwBrw8MEYFnU4t38hw6BhnqFv5
ax5/656bUl6SejdBZeXNl8W1iw72RSkIsBcHx+ZZ8Dp561b7HY4WN720gslZDCX0
5tEJffKMCGguIodeM0Bg+4XjXQNhQSlQJXOA6ngAowNLuG6lQ9bdk4IhucuHH3i9
J5Rx+cKO8EqOtS9n/q6kJGuu1WF9hxY5ov75T3ukQAQ337UnnmFQENCcl1CzLSo/
t5fXlfTWXQmvCt3cDZ9sQWtKgyq76NiAaw6HwaZZpEHw1E2kX2VEjsnCfE8j/jTC
MUcFuGRMudoLErmwxjV2S4u6qUjvDABYZgNxvZRBwaNpm7JZ529d/APw5A3QOQ9Q
K61ytw258BlBQFA+4iW6/uV11rsRvBTaV9FwEF5DVea2IwbZEN7tB/IekL1Frznt
YzFc4iIXw8hmvIYWZoCdijHqQpvO3LK/q7s0ZHpLRmnVGAWz9dbvDQGlcIjMda5v
C1eMh3GDpce04Bns0+LYMIKOkxx0xMi5EbCjtEtoFFB38HWMR4+hjEdTReQmoK7I
xN/oG6RWg6vK51NXzCupKYgNC9CxaEdOpmya7st2uAQhagg4bSFWe++dSfciOO7+
uSTGAKM8ho6VXYEMQ02pyFqf81BEqM6h2IYNfHM3znqA6Tp9IaS0+CzUtj+yUpKT
Zcjj94DUcJgJO/i/9TcuyR3axUdrBGbXP/D9Qqm5PaQ3QRIn68A36GayxoBepntG
MWefus/X4R4T5H4J2giYVd2yq1My0tmzGkl4HpbzrjDKJQDZbJI/lp9c9tAr+DQJ
uaCps1je6OfqcaKX3Il7ruZpWvIdZ5BVY1lDzZTVSaC50ymAZMvm/CBc/zOTdbQR
S+dnwioR7q35an2M5SJCf+QiyvK6yHm12n/96RtuarXoWaMO91nUE1wgHyDbAzoN
xgaioawteHz6beU7xPAoGoxc3R6FFA4aMvJykb8wgysSpFOGddQGM6tWqm8lm9HH
H20z1aKEzveeLIKtCBEnkPHNBOu+WYScZB55qVGESBC9hseF//gFeVplIL5COWBd
hre4uzFR6MWX3Ucl0Bae2LS8gJTacM5Yrvauhy9E2bb4UPhZ22ONhzc3Ler3S98+
2G6Gc8yqNgoAYLLjRKFBp5y0IAfJDqfalkQHU5xSNAHL7l4/2fPUp7t6dBmmLpZC
/WCL1DW9/ZuN/c5o90j/Rr0n0oe0eBcV7vgH4TBnQoh0M0l7rGgEKIIipN8/lvKb
85cdsWCHt1SeLv5hGN26EjGEi5YsIwZ+F6iE14CkQsshHlv3L7/ZTZkzK06nREd3
7NUarVeOrZPqxSNfyOV0GBfvnnIuHqllABFrSmTvVr3mO4LjsGaqYeJrU9127wHb
xM8rieEA1KR5x6Ogi2PPJT6PoLrlffDTmfvjheKMKf2/hxgCcnaukyuNcuBIFOKE
Wcz38QBYSpv1+mbodi4D+YOUUoQ9eKrm12UAoIXR0WMixwn5Gm3pcTpmcBDG97t3
ZrF7EB6ov5Yf3KkrBpUPAmgk5xK54XTwF0NDktBi4tube4XzCnd2V0hjdyvzMIuo
cKIokT2etUZDhPela/7FgVxOtu8MFH4xU1i/3DtLHY1dAJT5bclPBTJYwIhxud7C
kdrf1NR7IK0SUTfAv717rtezA7wE3pPmyswvrmdWOOyszcqfvW0UbXQ2iTMN+A1f
zaPYKLQ/sGbjHot5Bcn49avnwC3Kc/S8VfecH7tnTekyNilciX/eLtaa1HsiuyUX
iesJOs7JV4k7cuojaoV1V/9S+ZrgXA34DcppOCO0sg0fRm+IJKpYUPpOur0URCNp
13OSUjQ5HxQYoOponHHXosPGXjOL5chwYe24dLYd/uZQnLjYakECzQV1PAIPmSxo
i6nseTQlzofkYACO9DH17CUzNrbimldbrjXu0j/tlguuUUx0dXiy/5FGzyDegzb2
ZiyHeuH0rk+Ff/hZYjtZ3d5QPOyKrUddafA1usqjwIWhjEiafAzVzkcVA8Sz/5xF
QgNGYmDtWe3DFgyRQHRpxeBqomMJAxfEvUQCC9jr4WruwwtISfJPlUjvK1YJC7V2
+n0IQcRz3JcEMCck/ckM4X8xKbQXWbJDB6CAIzuhDGHqCj53w2FXmClGQL6TMSdW
xxsUMhU/Vtyrzg+cL0mtEJDpuiSTzeoyL90cdtRk71yt7JXPVCPzZLtXHK8xFuxD
0gqr+1jhKYGUT7GnwGWXkilsy2sYH7v5GPAApRKXfrVzUp+/q+gdMjUaPDpQVNA5
Q+aaRyXGqAZ6sl9Pd0lTTkCChQ1D77cHrMhK96cnafz+MTLMVBHTJFY2/NRA12s3
5QA/xhb81JgVQL+5GWHITiN3GccMxxMC1yF8scLioiG3emwA8gW1h/8bU7tga5aj
o3I85BbX1Yha4SHXk6DUM9Ku9PLsJMw/sw7mhpKlYDDcavBHZD49Xb+4vWfJeJ/g
Hraq2eSdHRk7FASSJX1IbamBX2BdAU1P91xAXV/LumWqodJl37n0CXs4Zrsr6iq/
Z6wQgo+jcbS9huOs1qUVi/y65UngGPTRyM32SlhQbHaWIsle581OGjMf01aNW5t1
UELys3jbiwoz8Spx1FOAYLprBxy8y4ORFVfuwayrjlEnJ+jMfQ+eY+/cMSS9u+yn
qlk6qfmy/gRmHogL6b6zS9gR6HE/5/QdKMhOqXLLe85DSARhn10UgHias28xKC1L
uL8YIejctbtchYX+/vOb6gsElpCzM6QDecnt9W+0IJTRbf5j4LUeRObOra7qj3a4
n3CZkyUTy1Br/n/CkfR22KfaQKMVp5Ga9AzWkf+OoTDs9JE/pggTh9YEkhePWPd2
0xO2EJLHgalPT+mZ7zd+Yn2rFDR1eKN4FQITqt7qXPO4giuTLWowTcgOIfruUErZ
/7TFa0QfczGdNQ+vMtsJvwaPEn2XXZCFNqjDikHJ+z3kvERU1PM3clhX4fjDBg9q
odvFy5Op1VIzNRsR73QdNjFLKFTI9BsbcvPd0eLT7CRkAas4OTy2pRpnnwTBrpZJ
wCEZaLHm2ZWvUqhmqpHyck9+kRgC4vRM04E7eT0ejR91unWsOp+FukkDAUo988xN
PAu6F+wHtwugJnNo3gDR33JNbfQ6d4xLxGcPA81/T1AUp7R1DZ/2SJHFQqUZiHR2
yXMSQ2aBrwMB0m7uiaNpAjpHlkqtjnIiahs9HkIsV6JY1FqF2mxjnz7/oOqZt7zR
YHzpIpjCaxhinR+JoYm/X+tqIyiAKtcNazo8nqbSTKFszW8dsTMG8seS7h8zIdKJ
4+RWIMY7s0Rl4Q71gb/Jke26Qv68V+3dTPmJ8OMdVz5wRM/KAyp+AsL1X4rIYPsK
D/nDYcQWWbYFXReFI62YCzkCeiUyVwXFtGm/dzMvqOYBlG7/6Af21QedAsNslfUj
cX7Ml25uhEn//q42nYBI/a5e2qrqfgpiZzWJDj1T3sC8FBxqgVB7uw2nzyA8bkl9
yxL/F0ry70RmZyiYO7S/UxTaQsLCqbX3bjc/3xAlUyIzyPcAvOwxLXVNWwznyciB
ZJgohW2mpuYe5DDoHm1jmqTVi2YkhDRUaVSPSgYiBO7PJjQ16FuuBWiRKemJ404W
G18ajsZueJncBd2RZvHKaV1zQc85LpFFRgXfRsy8cADEKJRv4SephkHaSjTe/hBs
ZVaGvFE6J45XITygaRAiTP3/DbRiFoVSWE8Y94UPL2qp3DqioVtVy+BqT1AnGjLE
9u2sWI7lXvFBp/+Kqzp4jggHw/eXuigSzR9BGdhCIJoAwVZ1gGMHtYeG8sVUSVxm
fAAZ+NERXqwobvX5IY8WkvgvuH9gQGu3tt/gX8ls1cObBUThI/+4Etvs4uuGP+9B
fA9OiUo4yDrc/mo0XNe+VmIl6ArkGaKnJt1oYVrHrmE3J5oNM6KzgMBeAukfwLr3
qEimvTcI6Z+BvBp4Jvt2uyoa1O5EfEkjeVg5IA0Dg2+BqdTRDoOY0E1cmPQjxMTD
bt1hD1uKSX1QYnlrcM+wlV0ChVYvQQ5dLIS+MEKZKoR3vC+CmpvDHFuJFhb6Aalo
NFpi2GP1Zm/2Gp9WSKS91a6DFVJE5uEc6DZBLQ05bzt4kBEcyzVeAyqwwd7ExFCN
KdWgZllVcHRS9iPGJ8aazTrVpWhNq5VvmGhlKRsEigJODEyCarkGQYuwbxi2JQTP
ufx0c0XlyLHgi8LGbdPlj7rJBmGwe7cTRLfGjmAJlUn0GhyBy3XPZonkoWnMhJLr
YeFm9vz/dKqp/KwjfC4UEiNtFKa01DMVNQuxOA9JtTNl71B/8LVmWaZCB4peO07a
Z8fSWEgvRSufyWMfwm2kvMbxGcX06AthZeSz2r0lUsljMjmHY11Ao5e5R1GEYV3N
cjomBr94NatGenBW7vF/lmYo/8o+Y/JMeo8sUP2yYwijy6T+JofPTPdiNbvcAVOn
chcdylCkIN3XhnFnEml3a3RVCJxIDZoQZhZ70y+3/Zr4lurnLON5D3OFDFKUcx+C
0J3/5K3dsqhdq1/tuNhUzsGyrYDStNE7OHo5VMWCcMBKdklUxlcxCeI7ASVWjJz4
HOnCRtc+2YfzvKsuks/Rh/PwkBg4zu+1phA8j7s0pexNA1KcUqG7lKq9aKaeqjz6
thb82ef0Olwdjghd6aPHeCzZhifUxsJb1VJfBu219zvwNNteEJ2K+qDaG9BZT+G7
B4Em9ra6ych+mtVYh3i+YMFAHSevW/hVe7yQOAvFG0J6mHbqk1JwtLYEVv79QRo7
6CGa+h+Z4gmolunloAWSzw7dpg6XAuZ7B03gSHXLek7ZwVqu/N4gvAdSQpDaspwW
5AR82D0dYDIfnRJNPfe+s0WFKsmD7oJmJHA0c1coK51LtJlv3YzCBme407VsEVfK
6+7Ppz08CzwKSg1/vKIwPlvpuBlZv2WOx3+o1PYyxRlDOn5CT6dCGDw5Y8/lGpdn
JvNLKcPCen6mhgfR4VN1J0tWDbu0sVF44td68GFfSUla9YqW9sWvmlXRd6q9Lt9c
NHPPEZRE+KRMVPA19PtcK6PIS40C8cJwrUSLZWzrRtk/pYVACtg1v/Oos3nFqUI+
5UsdRYeQbGosgWXA+L12ZXZXkAo0i3djVOg2f5jzAZUPuiu8+C/ZeEZy1MH9uqto
M3aRQBU/BgPacJLUEpn77/CZ8+iAjdYlIsOwd3bGymWmW+AnVzoekjWSjH7yqm5v
bMRn9Wfs2nABEP/IHdsU72wWV1LNGjQNeFB0QVqKCQPYm5U+hg+gpGGnfRt+AeKi
401nvwX6vKlDmS6ePtPmSNasP5izr8iDOzYyci4C3Ww=
`pragma protect end_protected
