// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
pJWiUEpo7Z9xszJktkXCMfWv66YtEn/HG6eugEm6EsfmDtnLdRBVGkmH9YqjbP5z
83Xt7bZSnQ9OibouUvK470SLp/U9IeFsIq6Mawe9IHTmvsz29jodRdkEzuJxBA8n
1UUo2htnrGGu59K3ti2JYDogaPqXIJr3nwToEDI8eyc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11840)
3dIQBuV2jVPh8lUSyl81z8Dp7OjShjtrShVd6427p9LLJUA8B4b9kK9+zb8hu2PA
6U8meYssgFZHh7kp1L25uq+r7/DoiYc8qhOP4QW1HV71+zT7Ub5OgOjaa+GGQNSA
uagwI/qanxemVnBQL70PdkBeiSHNzK/a5L2VGCpJXnqXI+No0u1kEcXKTxSkBIbG
b4KlFfPNE68f45Yjzj5GW3BZLB75IswwKThJfw6AfjwzneO/8X6PHcFmvQ2ylftq
i65898se6dFHNV2wWF1rz3CSmX+tTOhv5vQQ3tt8NKhPFkzZe7EHsPuZ8J4dcS0b
xQ0AS97+WWDQWSd42zjBR4UgpmYWA587eEAwSJ4v/EoxlwJvO8pcWodhMYeu38Xq
uXG97wqa4OrNDqxUqVmxA85UTcv2iTSN3w8Fznvd8ZCCAmJbQsLAv2A6c8U/1kr7
hbG+MiPy2U0bMDAJA1WEkNewSMIB1b/MxSSjovHiVLD27qiA3bTRdzz2Lr1MPPYF
qBhrFb598dy4Sbqw7fT+uRvLMUGVV4UZzNmusb9wIt19CuuosPJ4pZ8kkakfkFRN
ruT6ZeH+ES3UO9fDJE44qTT26TLTSCCp9fGZIk+/+/w+MVyVOMTbvaU579FVPG6j
hGx5kKnJKKnE2+dYsgikd9Nu7IiSP2uuT/645eVGk/kM51lZyuEa6x7EVO6P9kVB
zC7/L5Z1y/Kv2lz/FRxw9nRR6bgaIZjKEObnOZAjnAyyQrp4azjerj/nsuTIPd6Z
7g8TYaF30orI96F2NYshRGJe3FkqVKJr4zeNqyVoAJxAvULodoPe+zMKG4dRXRxI
N6ewcA5a12jX3OR3eHQziFDJvzwaOlNwrpWZwuFd7uKbTVgKpbTWYqI6uQBYA524
IU8Y9XIEQKgW0S8NVTpZvyvsmcijZoD7purdgj7MberF4mIwTAJnCR4cOGZdXr45
suuIH3i9eIdu7YAYGSRbBEzdw8T5KTAmBBg+5v9Kqi7WB2IH3CHJVgEwAvoFlJOz
eQ1Bz12TZHhRYMCwGCp5EbyjT7cYzP+apfQ/8E8x7s53XCRpQQgoACgmbRjsrjAh
U6EgWE/hZBIsEPJB2wOPiwgFozhe/Wlf0HQa80W+yuUOAeMOBkVdYIhHZFygluyU
wsrtIFWdwMFfoZBWo01XqWNouLEQUPm+KM4GXGJVxNlPbhI6Z9Q6IxffRSQb/Kvu
l2U9LwpAj6hO/S7yqcu864f/mfi9zy7z3Sm8qCDTx4cN6bvOYAqUdJWDFPBevRZ1
KpAEkOUBK/l+t0Ljlk90TvEPo3Dn98fN5ghdjsRlH4DZ3UDnbr2kc4VWTgQ8I6u6
vG08eQPBm0lrxcnDQxjrWuVryDpgr+wTqEB2btQOhFB4WQoi6Q3HZvGd7a3p0Rgg
38eR8kbMhMU+JtTajmU2Jj3t7hbJFfB1zsEdBXIE84ICX0nW8crgnu0c5W1I3tAh
pqLCCCtd4WAjhYGJk1vfO+/WwvxmZDtWk/7b6GII+1Jfsy4mfRpdjb7jQ9t4CIBm
GWE84gaSwQjdFzJswqZj8JlHycsYsRLOMxb1GdN7A/Qb3QVaElIID1Yz6k8OzaXo
JMitgoyaPPbPc54Vzbck7qVP2SUixNIJvdPpbJuSgG+GnlOgAP3zCWh1moO815oA
fEIvbBik0ddafzIs6Cp1CVg6y5ixGTspW58vlowAxUGbWDApeLR//gC0NcLcRwQn
mMaQeQDxHJ6M0Rv37yWkXZ2oYJuFuR35xJoRn6fE0Ksh9rkTftbo0NQKgt/ud8Fq
JAXV08JszGPJt/Zvsg3cW7fr4wRpApSrDM093sFQ3qP8IuKS7KaCoWCr0fpG/VW7
ucipXo3Jvozob+tVRm8BTaF6709hu7Hi2QF140MvvbFq9rFjsOzAssuLM3a9cbP+
MsBu/N0d9vd1xsh4x3almxt0nPBlXchRebAlFs7NLuNozihsldb+dDPbtbxpCMfZ
YrX79x9nTQnbrTAXCm29QQtM9/gSYwBtc5k/ISQgiJMiPjJZ5EDXn9SAjKEQvjsL
IDSpr4Dr0KPtOXv6kjZYy9QgxuBm1hS+L4rpe01Dmizu1dEjbvEoD1szUCVleBo0
Db8Y69Byj5CtqTFC/1pP5tueCDJXERwBH7R5Lipm6RL31CDCi+FUWlnzVZRSSNLo
T3WTZNSSlw3aozwi7dHIcB5pLrIvTvyHrU1eBNCCQr//eXjN7qlVhiWurIwSW4wT
NqRhFeNUaSCZzBBGPRGRihxaofMV5atee6sZe61yxwzwIMViPbMe/BYppe2pJPdV
dES9wbXoYROu3ZDOAY1zjKt2HjRUW1ginoxJqO6kDk57lyls1jjDSVIi7dZ5JGjL
Mn93Ee4/LBWYcVOvv+zUvEjtLmfC2xMipVqkiTPpnaohP+3KpDjzdQm2GbHjU038
oDnrg8XWGiBKUjoVLbK0TBGrS4OwAZTxy1c+/dIjfJ5GTafKYfl5vSPqZVWivXKv
g1n15H+HPYNYVYtTGuUyQsskk5UV1laqv9qV2bKjiXcEq7wilSt6OgmOf3SqLlXX
vJ4jc5vL55k7+LZn0qY+ecxCT3T2psVEwG2uS/iGhCgtXmRSueiX/If8itbYxx/V
BoSNkYXVQw/rnBWfyles1XYaqKv3464Cm5Ybo8kV0RpqA5cs0np71kFDNcuh2X/f
VrwjtJp8bhcaHGmNUehlbCC/3MSOyMXF/aScas3oOIVLvIcFSFnmr1qaKgzHLYqt
QGcl/MMsUIBTxqzTOzXdepCr5eqw3yKEKRr79J7LwlZxFvEw83GvETZ2VXph41G9
LdwDM/v/Z0vAUE16O9x+oLUaKRdvnpz61Za4WpAQDduZx2NIq1Wi4/J6dGBMpLaV
azeNAWy/+Qme9tmi6CtSL7VI8JXjI4o1Bj2U4QH+v7JbuGl49PQeuotCUHTx+wKB
ohafYk1QG2ABum1oNl4a38Dn0nz7y6JPLC8PhK8/FaYbqJ+pKW/4ygetMVu28gQv
Hvtf2P8NSuSR5DN5ZwOF4QxyHTJIa4238QuOnqRNHhrxNo1KeBEoPCtkZxEK+4+A
ue6z4Nv+WW+uMelBI6eKtDQ+wrA9eBtej0rsweTDkpsCT1zjlC301GFgoajUlVo6
tk1occCXY1+mvv1IrALHAv3HpD1mNARaWzThoyOgfgjy69Dy5N1sUJj0T5pn/VmL
dvzAE0G2LeK5CypNdex0tFj6RV2oIuyYXO7eHrpnzUUycTtPDqOr9tuCUthVlmbh
RIVJBszrxLU7ujFisxupP2tiPc9GV4TuLDwZ492hXkruxVu78Fzhll46utlQ6QFH
iIt7cAvqUeX325FxaUBfvNMpXVDoBkXzOYJa3FN/uXSEEX8eIvUUGyaOBFEWBdvq
6hJBedyg/QlK0WGITHXcA49xfSp/Be10A/ksFpmMSMWlhNYz6Ax0YFHML25k0zqW
v8eHRZVAwLgxRhQXCtJnekwy+410xHZp47Um3J8wvvZ6wni7UNLzxvZhl0idJn10
lnULQbtp4RWyfofMXodKhQ6wnJMZKP21E5ErbsSnMyRlz16fH4ajmdW9vFxio2PA
5udieC7fPn+d3M3/EuCIPhBqZsON8IjJtlHIFyu2icrY2fMRuaVfNZCz/IFCj7rr
Bm8U36veZtTVUoDyXiKzxh5e9g1gQw1XsMWlHd/CMJVguXpNrP8UnDHE3xVOwGT6
dyjYYZcx4RZw8dy51HpWx7pW/cWqQ9XsdVDk2ZTJRYnjK72CDRvYvo6nEa9nJ0M3
D9QgCjwWMeb57TKwsCoXsQ2Cx16X9Z54BB4KqxZq1zKPlbnIRDTZDHfbIwwqnC9a
vGqupgRWDz9HJCQ64Xz0ZzI225BzdZQELuIVnXD/tCKA5hSqpumBnGcS0W0lZHI9
j+sJy1eXJWxI7fLE1QhorpUF06HoEtrSM/szhz9z3XXGk58eKdvZXIsg3oZVytU0
J68igJMT2oFyYqju3apVKelA5nbLgiC8v12lAd8JJTbmgT6vNvf/qh8COtauK6G5
CU/l7F+qTk2dp1DL6InVW+Fl1XO1ZGHt7FtvugLPcNWAktS8TKIU4AGixJhiN8j3
xjcpnp9n/B9OwfMZrr9FYxu/Ha8K2yvrKixp0PlR264ac/2vhIJplwbzCLqoVX+m
usY6YsA9kWYUDO39pRG1Du1P5AM8YLZYrMM8+sJxbtwOptAxZm+m7H+2JN1mKLV0
JB/CY/ZkvhKPREhSOaYzAJHh7FBg3crfiI5jTZGnRPxo77cYyG0bAdxNDT0PChgY
pa4huvLsRwIAkJjCZDHFP9m5gh2uP7cR3qC1S/Fhd8rV01paFcrVcYlbR8/Z9A5B
bT7epXI7CxWgbVvsTbV9MX5G6WZ/yUK4qgnOwctYmYNbAdubbttqYMX1MPRBekh1
2nIIenWyOojCSvmlnRcxi5xbzP3DUwQ9ZYu2LbhJrDgV79g0dq35zEu4DeGS8xpt
IoYbGAxU5ixsHYduR4gdZhoICzpXrUfiSP4aXVNTiMqf2WcX5rT4aCR3DZzFBtxO
Cc4SZEX13U65IWwSUHYe6k0hYAtjzY5Yvg3m2A+Ze36mkzAjSSlvkZ2GDy1eRAXL
m6cHz/z5vQboDIpw7h1HPNoriSr4VWO6u3AUb5wh8H4I5fVH2t6GUg3DfWEOPVdD
5hPQK7Z+eZJI6pAsu6YmrCVB2z8DjM2xWwU8tjxOTiFJj+1jrCneY9mN8yF7/Pzu
p5wBJsfIkyarZgM/xA8WPoeacb4bewAGIWTBfRiYxRw2uihnwJm2jYHOLa0ZEzLG
x0jjBo7OjFZLFej5Ai71Iq3cB1rY0pW+4EjTG6Vm/wpivkQgLqzE/RuHMhGhRDjf
W1xSzqoJvkw/81AxY0MzBY+ELJGkl2CGxfVIfxiCbVjl+8lEDlwzmst0+ywXVPDn
FOZcu4re39Xuv0KFbBcf4tzaX1dgWvDmlYbSRw2cmjza+CHb4gQt1z3N7SeQmy9O
q22Xdj/RhEW4e9UPsBBv/V3PZJ5IVpdTqTsWlz9E7fWC2mr7N5omnb5TdmKVlgEw
sZJPgdMoTQFmcIWVb+hRU9p6CdOsKAKZN24qOBWZp0u6miVYr33dgX/mcAb5DyFw
YQu+NE8wcgUxChAe2w0HK65NLzSV9mhFORS9VYfRRha/9Y0rtdQcbRRilkjWpr0G
pO27zn2be4f2flTKt0rQHIbehqvCIbvkS/KAQtibFqgET87qaYRtqSKbdtRZ/OqH
RGQOC5XAjRXfxWrfktv4+ZWSEv8S9aOWKLpaxAKm3ZXOGJrWtf80bIeGprpOstVh
JRRD+lwWCzw/rpEpz92OVz55859Yq9lTveC0M13WjU8PMtS/3uqKuNuwsLhSAPss
voRlXZ3CEn+/HKptr1lIeSZrwUACeoE0Fv9EyZfCcjFr+HEbWuan82g2X3gLIQY3
QMrifGUpGNCSxmFSfHXzPeyEKHYAa9S/hMJE8amTG/Qtrj3axGocNhBmO94sZ9Q0
IdOdvgrzuTW5TQ9f1mn1xIwdYNr1+06Vf1p2kEGJmH3oR/kChETWeczoElZlb1W0
gPiwHGnnjGtJVCZSIW78mdbYYSHhOQWPFZknphyKhxOJkEeCp+HJX9KPYZ7oQfBk
r78q5KlhxZIckGJNpRkYO8GYUwUOp5IaO9LaQKTwrpMYU/oxpoP27RK4UD4tI6rI
78u+d+qgHHYQbvzNu572uN4uIly0iyiwL5xGsbirh6jak7xyTJ9nZrBYTxiXYVB3
dee1zzpfbVFLmo47vaqtBVlt6Dh4AwSfXAwhaX8Md13vKVvQBZXxQZA1PyIqqnbb
3cKioM0gveB0S+f5ZjKymMFEi4X+B6MLd/DtoPhA9Oh/ogVFghcjlhQ4lJCvXu0Q
/itJSYL6eVCwZUwbB72dVIjGivU0vDQiBtwdXYpUEUww1+fE3U/2F0jXUjExYbwo
4gAlNkvsWmP0Z9Aixz6GfyCivjAt3APUj0mRL2sp1TYPMAXZhzE2yB5qlniV9UVo
dKNgpAo4rghlHXOs3h6f0BfW5ApJ2xoyd+4cd8fmUIcPrh+NjLwLIJ1GKUJnpQz6
Tz6CpawX+qIJfDudgdqmCPig68U8rRDl+Pcdq6J0Odsogy6zLaa+nZrJLZJegwst
C1TWqzJoma9N8zSqqwxvxbc0F45k/NVoBETYGOlwuHndgQqVJCD1qyNrDDrdxbnc
8pLioY+mthaQdksGcVCIVzPwYoqm1TOKRWunGB+lEK8eXv5exlGI1Go6dgdQOrEd
//fVfoSP5bJ/1PFX7bjbMORO6bRKBlR+E7H9fHc8PF/mZk8e+9W4OhT24yyatTKO
G4MoI0Yre6+GDODAHj1YbqSrwsCVhD/QMTRcDUhZ8bK+3Xb39EbKqG0wvTjEcLhS
X+Pe5FPmXVbfn6G3kVGY4QAUcv7kRiraVhjmYI6creqMSAMut326Qp2NuNq7b2kX
VBbSOrZsC2EvguFHXO4S5AheBqdJrA5tCrUc4fub7mJiBTCpBM7MSWZMDGcMyl5S
B24OMlJcSdfLJUoraP/tHqTPhT67cjuCIl3CVoj6RzLUTZlkHmgz2Zgt0ewhTcn2
peKWduF9YiiwKgUMaqzxq2mJqJDtTkHR3fX9VUFwcChi7wXjC/jDW6tgnjwwq7tL
KMVa1ANTpx4CFcCgVmLjJtE+7rfEfTN4ZZ5rd+hylafTE8yHD2f9TvLuWklZK74r
HkWpdqUuZifqEKwy/6+teF4rpWwGFoTI1tfdyz55U8eULPL25JmIYu9DaJE0nbQZ
I63Jnl46M3fg7DCiPDVUeF/PyitWbOfmGEW2RHlgm0Gn0W/5iWO24WMtiF9gGdAv
cKAF5vav6+2DtZq4S20U/kjlbG0rmYiM+h+b4TK3kknhUrHxCP4dlvDW6NG7K7tO
D0hMpq9DRCOciKfXC+hRo3uYC4IKDkRFGZl6jrWChGCqHorg0VsUtxn+7fUzVtS8
1lBR5GrbO46Qzx6I8LWrA0lVOeJXpnIvViwez1ACUGYVsr0Cq6QUnwhV2fjnoOJo
RHa9OYlPUm9StamVMhnnq2tS5qzVpaYZ4x8l55WlWUXEARpIv3JtxSSNfx0+6Rpf
xQAPXeKPg0/exwy1tmEAlytxi6WcmGnNcE7K9AfDjXGPLJGe5j6rVxDaZ5aqhwQ9
tQdznjra3fWLlyFjV7aoVew8oCbnLZSCfB2dvLN0Fs1C2Pz4ORCU4nQs5eb/YXtc
P7m7HgqVSWokBc248Jt76hf4A0qmcCJxwl8GYbF9BmVJ26VZ+3D7c2RrX5IXTzGb
cLhLlnKMp91oAVlRD5o+wvyBhJkGQfg6m3K/Sh/wUWgMvxTDFcqmlbxxCPepBi6X
yoVtu/Y5sn6QK8Nyf2qhdLCylFZ64/Lm/mXr7vMbl6mPZw218AFpF9au8t8gjBr+
eq9SiwThogN2muowGfKR3TYE+PurtbrjfzoIb9jSpGOfZ/RvxSC0wPRxUw1cuT8s
sy3wCgIsJ9dTwSKCHYUUIZ9FmXkExJ0p3HoqfPm/erGflwLhASCPWvGTd3XYLhgC
SFLsEbLOws/LjPjfdAK4sY6v5zocKqUhTjBA2So4x2bV5XPlOVoNDrcncOO85mTq
b4OdkarqomlSbDwb/Tzwj0VgBfrUTBbqIbCn2dOwjjDvVyFcHPddEF7PFSa9teqV
GY8E/34PJ/Uj5azGq4hTv6il5LcLTz6zp3aPB/iesMoilF3yJZgPAkCtRrwnh71k
hvNHfjH/ZjxvZNc2bvvkjPI7sh8p2BGmYfFKFByTYvECjm5se1pNtKzAd91qLiqc
CxD8/LuqqJHA06wD1LfTkUKBe9moSeAUHFgIp/9tVqI/1GYACRfpMzPK2k8zyvTs
1H0ucCztgLzvfhQER6a2VwpIkcZjKhwmRIRcNesmE1Y0n42sgEdsKIGVPJpiMEGU
wBCcWNPIeXEXfYoSmSckT/pUGDchCajzVn/GW2lntBlORrSJ315/v6QStwDzqp8j
08Xnjf1Oxdnr7b+P6qXOeRtQ+9yy+wDSgpij1fJc4EbBMoxFm5Gvcnjbv+dY9Xi5
C3UCOeOQHru+uLDu22dE7UHGMHjs64LAjxp9jyq/g9yqP1DOxrkHFUfOgYVxX4yw
9UIZcq9OrUc2WVwi9YLOZzr9zPnG53xjMVFlwabRzAVxx+lLB/XYa/aH7NpHbvw2
i7RSynw8EgX8GLShTjmROLaeyjmbmCVTKx/KnF7/O9WCdCInLuAtqVhi2kGBDCi4
4t4RwgS2QUU5fzOj5b7S3HSmLaEP/r6a4Cwj9LKRtX5FhgDbFvQU6mCD52ZGr6l1
akQDy4mxVfMlbEsOEyRQ3sNAfRTeUFd1uTbsdiJwVpaYjFlLXQjcOevjpWvVGG3j
vRmTqnP86sYkio7SQno8HoG9yCMi+hnkfqhVIkWkXp+bXTHGHizhJP4l+j79OrA3
Zrz69unxGUFqfdwLU4TvqKe5MXYESNx4KDFKZlxFmAL3fm4xcQ3xfH/2ys5TB4ti
6k8G9wyp3bfw6O3e8JMoJRDOeMax96IUlbHjpnKQl0lEfeQscdBliDHMhfXLur+y
2yiCENE/uDvwUdAodtS80VobgdmygawcpDlKByg9Org0XDBZyExY1/P/aUSKyFpb
Qw++dy0ZdcaAlX7+GYjG0N1E623UMoiTT5ovurfPsatmPvcpka5jF9bUPw74SmEj
t+CzDMvNCN/q6RGX7AceRyrrDkxSFaQuxsRAEHrCGy/MpV45cFNAQYjmuUDus4F1
jh2o3WcxD9pz00+mjixTM1wUv0r3YwgIqHzidscz0VeIxf2hqg/akAim92dbbP/n
SjvS1SIdNeqlnIEGCLWeRMsnx62HO5Ndf/fP6/TmCt28LpWlJ4GlChoH94gY7Xn5
kuRPw3m0p8tQ5hYKWqUXFIlWdNMzBswejTerSCRfTGcK9t2sI54x6m5XYf1o4vZq
gMJY6vxyWGuLFXGsGqIgWb24mx1k6bJIZmWFfg12wsZlJ0EPrxoK/bGQDw7recih
YdQM44kR7UR73SP6wfW8JyAaZYv6Nhi1IRS4TM5tuJjtJzW+/ahcQyzgBN8H5mPm
/7YPRpurj9txsL4IR75QazspsznBQdyYb92fK3KCJ8MZ0B5rpr4FhO7QpKL8JYYY
VFC4/P32yO41muKyakNraM5qfZGbRa68s9g0oAAQ62U+//5pRQW2gRRu5dhbY2oS
M2Sewg6nfH8soCyQRJzODVyV1iMhSjcZQVHYJYFRWerkV9Uo4C4znhztpEwmIXlQ
dtqfQ0uqPlFSAbSC1uSFZf3Bl0TQD4dCtb7PcE8EhHeDtoqQcFaN1RE6tig7LTn1
lwydyREh9qeQSy+YWYe9ptTl1M3mOTDBWWDaWc+9jQ58zRk2RaW/m1bnbZO44vzo
yAhgTve9HSIQ9aU0PP+J8Uy9a4TWYNwNcd7lhqAP8FLVTed92y6fuBeMkM3becuD
bJu4LOlyyN4pOg4ruvtEJaifSatZui1R0KcS64UQDNubc9X32215TTH9/Cso7itl
B752iEBsRV4nvRSNybErOUF0pHYoTeFyq20WqLv27imI5g8vFW7jMRjKlxIx2dJx
t0ibobMLIah4PQKcFdNPt1ZAi9qDzjCcCqR42RaKHhmy3qnzApepKQoSJvGbBfPg
zwM/fsLnROOvAouWeRbxafgg3aJAQzQXwZr34h8EY4FzX8qZvbJV9GcnuQsTixNh
E//+x+9J3rLRM3zKZ2tulEIx2eWchYh26Ta6mtBKe27j4WhDCeJ7o5gr7RRVFK63
yxRAHDX1ooLm896jzlGfPJPG2EcMMzKnAQoUMaLz9hmLvIG8m7irFp4D1ma4jTu/
404G+4uvR3pSLUmCbhux8rIkzDV3F54CtaHlj4DZpMSYKTw8tUxWMZ+S9P2BMF26
Z4oJegeeJgAPiVroIqDjx0mDQDjxTWCT06xcmWNwFPPBm9l5q4KdQQr74gIeWhUj
v38IRfEnZE5eAzd+y5qa4g6r5DESBZ3eh6vGx4ta1Lwh/e0obHj6rIzc2Yu4JQr2
S7dE4cTKl6AMAdlnV17hbK0/GcUssjlHkPBPNpFKAaQMvRqn6zA/WmeOmybmS5kO
q94w8iT3B+Hb+P9GGwtci1CAe6nue9n9tjaDsxDyk84nnWzltDI6owyO5jAZjO7S
4lNL/p/p3x93Lx8et5TLftx/JxFNaTufqnePXYLmbrdAnICTGMflaglHej9kv2XR
YEK4v7KjwAmFH+KFDbgy2/DE6PMvx/9kRZwRKBcgugP0ieQlUV/bnPKOqQKYHCEl
FepmaLbo+MaNy5T4YqA3/y79LwbqnPMFPc4L+CCCtPR+5RDMM8umOzA+vx26iUEp
T9JPM3F987EDsaURtZbdcvnKuiKt+LE99Ju+C/1IESZreoFIYMqZt8QTUylTX0SF
w+c8/wSJmMHBBLqZryLc4bDDBWQ20Ojie2p355x7P7gBceFmbg8xvWOaTrjp+Zl0
Ycx7pbnBKZbDVbYS/zLtMUCplW8QoE/KqZ1lntyxtnI0JL7yepWJaTNNwDINr1kv
sZyTMedG6PoKwV9O42jpiKbDwpre1xfLiT/uNnNgkwdjtRog6zntO6VJ/wVcwP1M
tWy7o/p1Kyc1HdypkSmR5Jk4SzFr3Fg/nz4v35knjOJAgzYUq/bSIp8pI3ZQbEVt
/svGq6FM6cwTkaE8Gjhh9zPnUnYM5RmW9o/XaLbBMOpmQTOVMHCgdlLQGQ0j9N71
j8Z1UaOQCAiMv8voWEsK41YI6RtUKjICVyE4NbzyBgdyKCrzdli/D5NaHdgrdIfF
ixp63xpg1tHOqlOHXevbglFKrZIi18yzeriSWynFWVC5EBsM0gRwFfs8SgNxENdm
oeTJUs6ySyvJB/FrnMbK5iJvNJCKhbMp5nLqR7FP0882doIEmTJTJ5v/CQUhF881
P0AFEnDlKIeHfI40ChQ+Bgttl2nVaRPbWwVrz+qHu+/D8SYG8HL4RKbLSe0EBnQW
mDypukCVDmI6ZsxGG0zNLViZq8RjhNW49/we6F7lHkv/y2QTDN62M4nTnT9JATqi
8cZaL2CakBasYAUqMRe9ViJne8NRxMRajW4gRo3lCfhJ5sWktAcy5dxGPnSE2RHP
kkV8Z67YsEDeISRUlEDcyLWPO89MeVWohtc2RUMdTGgK//1DB9ZvvNXxVm24C2bp
zdP2J6AFCQp5Lms3G9Lm65nIbkkDmScAo+1n3KJKQa7P4f51ofWU6y3ZVQXM80Nd
E7153YV+fBsBfAytast3bEwGsUgitvz+myL2/kT5GDmyu1gzNC9iuhDW/fAIn6NB
2PI4tXc6l1yMl0wUfun3+qw8Box/sLAMxgtgDidvQqTLfxnhoeMn/O/CBiXlmeqd
sqiOKc+V2FKVu/Ndh3k0W25KglLT7oRsf+5YvaiT41ccCdMwEAciIJJnBA0WVECN
zkaGc+yh4CY97Duq5M/LJIRSJElZGL6zTNiLcdoi0sE96lOjrrriJj7seCDSTElE
eBM0wthlXoBIk40i1x2DG+hs+QbJwAIsvkXRl9TcuvCV2u4OQlYHds6ypFk9NhZY
cG8BGrSTM4YsffMMYlP+O1UF1pFjYdYIejIlngPTv7jJy2CiWqLsMLrDmMYfrsLl
mDDPsX1AIOvB+9AUIvTDRfVSuvpMEzR0Vx0k9Pq1VEttfNdzaE/B51m+/DQ4W1qP
ee5QCrr5Cyq9kaq1+AkRMCS3kYD9ThA+lk14Be5SPG2Ork8QNYtNvhdzKviR3IQy
VGOp2s3OW0TaeHPZ1oun0MA0si+41i/AMI0kp5GWLJtZn8aRqXMIomsCfDOlgK9S
wg/SXngN/5xCH/84hbWZNPLV09ux//hY3I2M9xQAi0r5lUd3Ar3i2s+1GA19ILMP
BUVchu0nkkfoZMk3vJC/J8e9G9n7qQEckRknxCR0v6GyqPc/veM42N0DRnCYu6Zb
d9o/U3GGCVT7xwCvjZdr8A0xbtVROs5JOkoRA/yHS06FOMxykEDWHW5a6S+Tu0Ij
vmnPTcK7+jqFMWqMaR7PGnwwVbxYzaNXhdGQs/IpFkvDWC8S+EC6WkNfq9B31Vjn
1X/9OgrefeMi4VYz8vHHQG3TDYB20Fg/TM5Svuilk0u5Pe5WdBzdpR0suiiGynzy
VTchVbKf5MEFXhkHoH6bM/8442//heKiUmtOnG8erMwIJtTPSe92kQFJMqKs9Ox7
LBXKaPxbdWdwkMK9JvcqKAwC35K08ug87tPyU0lFirr0lIfePAaoBphxXwnN27rw
Rx6VCJgbV1AxhRU4vYQtlndPb7buW4spMkvLLfJ6aL0zn9NHhh9UmqUr19wlV9we
YU5b3uuobRKh7Cta5JEY3R996N5A50Jr6I6xT+uYJ+BvRL6XX1O9GegZn7fkzb/w
OJ4vVVhcaKUHe0L4RjNmz5bg3RA1gj7isBhGJmQchEtCPlPaj28LCZXN48ccWPOc
cPsju4dcRLGepftZTjs0S5PppAClE13xQ4gYzOEgoCMh0sHM2TNYGtHEHtdFhusb
armmrzjCkgDLlqZVtOfCpMZ6GrXu3gFqAxB70U/uwya/RarKK/0DOsryXm30p9bs
yLsBha81cx1W2l/P03/Tb6yLnVq9uLa/tugl4VVxS++TnF/zaOWH9YYgZFdEUOEt
V+SbrDZ1uH0Rfqvl4QD675JJ8ctze4qFIaVrXGpdKnfFq/iI0kCg9wf3zxH3VNT1
FCq4P4fAmt3+jgDHW6DM192bZI0972K27nvXIXh1fjzf0ceQg09qd/M/ZUaxmsof
TuyZDDvR9CJCvIf/UvzXX9CzkXMH/7QK+eP4clr4tzftoNKz+SP/NGJcSqsyJsd0
8XVbLvOCd4u07obUGR56/fUpFRSMDVM2avrABvjxU8LrNHAaAoO6InzzAJelZfYN
pkH5EdLPbBLY5e7ZT/J2Gf3l1YGHJST6avxQ4EOLuZE6mSwZD1AuShvUKha9wAn6
WBSjj8xA7d53BbAWETcjmMxhuaI+tWd+9JVckcCvMv39OUlDDPoXIzwU9Ync4Xgg
Sg4r63chXlagOKZA5SR5g/KStDvmD2VTff/3xRQxJIAOOt3EVrGAVgGJU/txj1DV
qwN9Hmk2s/gObH6BV6M7nLT4akgxhQALHwud5wLbl51D+L+0Fu/Ay6b8PSIxWrWP
225M2OWbVC5s0Y5K/FpI+LHMiCImOMCPS10suw866vprDe5AdqnLf4riR70GndY9
m/zQOc9b3igaAQMAbD6VZo+oKSPc5JiTbka0hBeaSj+1OkhDFPum1rWd/glY3Wta
R9LPOGrBrPhkM2A3bHKziMMBMzLaOfvAvbSOVd2ut9EwKZ6YVBNZUSeWfbOxfjta
f2hSu687z3CJNaD/x0VgcahRdGJH11+q1h6K2/L7Zsm92SeIOE2fT/LNOjizildj
JkBy+Inqab4Ch8LapDNOnZ6ZywWeyJORsl72hc6QsY93FZubRsPdNsCrxF2wDrHd
j40/V0y4hAJnlsWxWI6Um9oTQxTB4j2qU4JTD6HYgxUp2QOa9XEp6u7ZHLKlO8Z5
e2tEkDAY9A/ue1bdB9RDo5L6cRxPoUzVwZm12OL8ntLQ4fWRW534a5w6uamiwLeV
DJjPpGRU1Q05SM8u+51IUms3OCWZNQW5LHpxkl0KuMmiCdELP4a0g5EidKNAEbkr
brQnK3iieIxl6AzEy8+oDntJO+quKMUb89GWegZ+BfiWCj7UKASwEjMP8IdwyiK9
J7s/kbXTsVbSSXwGZ26n5EIBG+Vz7XSnsbyjvtgMwINEYsI2wte5SDxqYyf2mJLw
dXGknx+vSHVQ1ObPhZMgmGMHzCH0HJTGB8D26akARfMj7MpLupwljGQHqJ+sYlwb
W/5B+7J48Yw9F5gtd9roEYgZDslvkkwuqS58KF859CvtOtkMn6L3g9lKBcu2dzux
Pw8dD+36SVdjHL0BzgTWYkO4knQWcaQWmqEcvUmaIaG75Zzuj0dmKEBSkdfmlgp/
gKjxgVJr8D1sckJ6ivZZAzlzk64XgpOiSvDt8V4coPFfGzkgfJZnJ5+EFZ1GLt/W
2jKWTRXtoCV+/gUWf50HtQyocazS3roLEvWUoyqVXvyZXs/JHxlKxEngOhwY8V9i
3BFMYbMEzohCB9v/RkFD3Tbx76goYxrJCQ95aXzdnWktXahNZzentXqcgmPC0w7B
gR4WZhDpRKy2DjzMQ7xBWkaazR6UsbjuxlhJdq8Xcl18EBm1xWmmdgUScfnQLTmM
NarEI1L+SINrYC2luPle9D/CEky1fBdWDuqgTPIvRIt6pmHaIHwZ1aO3JmMkQOx0
8jYuQfZ199B6r8tIQPZH4NbG2mZXQZB9ynvBQIr1bIjrmi+R7JGj2PY7vLTX7Coj
6X2ccN5Rnd8Xd6OIAm9gL8HSCVTTu/LVrqcmQ/ASp5rjfmn+0+iuWKuq+CzK6UD7
e5z2IWTOP5o5S7I50nu3NpEyA3c9lSPq88YQGMztEqWwpcsxxV66ghwzNLdgUsiL
CAhirTMLaVxI2se2n7Yl+PQh91xXgx62tL9lAH+2xYk99awokJyP8aHqCg1hvTrc
S2sYG1hvyG/xY5pi9ivCeeRw4BQBYIIc7J9eZFlAVYIbOT+BXILOCIfTKu+qCs/R
EB0xltGYYsKteEcU88zYd+6jQfP+hM43Hpc11PLyes+E0IFgTY8K48KprzwI5O1N
88UUWsTICKFs79zR0My1xO+UHPYjS2DdDNLlLugzou1bRGTOswuRVx8lDMrknCc+
TTHWUiUrwDJYZZyNqHJaAv3vy14dHGY9ibiylTbwJA0UXfy7RIeMSHkc/+MVSgCA
osAFyNZkQ4vtV3OSYeb2UP5HFYrZRGmriZKDSk6zXRKH0L7jgDL61HIx8IXdL9BS
cnPXc+0YfKIOI42OQ6RykYL7RvBnPpcYxMsluMBMWLRO1kV0KAF7kO/FsWFVlQos
sRBhUaej9VEVaA2thA/L94JQaj2Q/4PH/QMcSrDpY4j1Nn0tIZ9WXNUgQzrpVF4w
4Clgaqw3ymWEz8+uAvGImVVHbPw5r9mxs4PHULSU9YuSdnUyTMbUWjvgMKGsCx8k
IeQK8dBRmVzc7LP4mNyMA2jbAcnZjCxfgXcAwn+3ntew7jbO/rTHnsf8qcUVbond
qnoEaJSr61LvT4KGogsSZWlv8cA7tunGpa5KuOG3i3mdUD6N9F7JGzGqzPe2tHHB
WZ/hnf/M5TR6sZzatNsxNr/upL+krBuNA1uBtqxZ5xDSxIxwokhaBks0z98A70tF
NKUlTxwXQx0GryV7ZKjesXLQRuN/yZAWLlHLDvmt/x6TBnFsLUTciX7rYpcaqqv5
5ROaS5NdAh9HMcWPq1B5Mdsdg1HTy3gO64jgPS+NBLI23wgzobYN6EBLlP1fosxp
XGI10nCR8N42skDcZgwUe4MG3fsMbZVWjHBlVhkUpb2If8xjZe8kMnktufJdENpK
fa1stpIbPCUboxaPzbR0W1tOj4kuLDwfNJbGnj0ov/uFeiaIenWfXe/VB6dV0sWo
Kbhjrje1Heym6+F2GEcxBEdc/VVeu6zC36o49oTF93Yz4aiWda2UQnAO+MpjH3us
wbeLWMWK6rXWp0uajQQWzXPfj/f8ttiyMqqNJWAIIkpbkvX0v8GmsUH0TF1IWlXG
I3BsD+PiYAsDujCwpFZEmFDHhUiyz6EHe5K3nVFXT8pey0q+US73w56aTJNYa1JB
cZhrcmL3QBFEY35zCBMG/lP1PUXbS8ojufz8aaaw9nw=
`pragma protect end_protected
