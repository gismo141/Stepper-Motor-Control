��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�>	��h��H~,
�z�*�M(�b	������LV�laD=tp8F�6�!�~�\@NQzB5�1�kR8�W��7�����e6� �����ْ����5�}܇��M� f�/�_�p���Y۪�^�ow��PS�*'��,e�/�W^j��������ք��ݜQRiZ�-
�}u�d�|"4�����fTD~e{�I��ks�W�oKG��]��6Du������V���r@�Wcle5�t��"��a�ǎ����"b:ٯ��O�A���k���֩y
�^P��}cC5	,R�W)��ɑ"�C��Wh9U�sɕ�B{�T��'���Ч�k/Ƭ��7�kֳ�q��	�c8Y�&s�mCM���lZ�~>�f7@��(�a�JL/��������Ly���C�2g�& ;���ս�\w���Hu���4J4Y���!P*Z_|޼��1xA�/���m�������/&���Cʿ(
��,@�d܈�K����~?8�d���s�s��c�8܂��l���SX��G2�`�<Tt5iP&JP�2�8|�1*�)юa��А�t������p���������7?}�s�{��־���l����M}�)� _
�o��&pPW>���X+R�T��<�V������4�\-N�����U�g H3$#6
�q�֕�,Wz}��E��ۅ��Zdc��(���f�6 "4����a�O̀�R�mrM��?��Cgh��7L�����43K�ե��Ƈ���3ylc���}�Ū�`O��b��R�|t�����.���!�F#�0�}.*:"���|�����Z:E�\�d�I�\Q0����v�֯w�j����Ć,{�+b�Q~�X0�h�(D���p;蜁�!p+~MP�O��X#-t��f}Ɏo��`R>V>�����^��]W�X$�7ˀ����KҚڥ�}��7�����*�דyRQ��#[�H"Q+���A�ÿD{�@�
��LH=֜B_�,g�B@P�S*�[f�y�1�+b������N��l�e(<B��R����(�yu�)��?����O]��EW���(jʄ��t��G���K��EӮf��_�E��vQO�e�ƻ��mՀe��L$�$�=���dr�:�Ru��lJ�]��Ʃ+Q#F�o����X,�'do;���1�~����-|����Z/^�(�͒������B��[�d3�+��EO>�/�'����H�q[�lF*@jA�o�P��y%s������y1�x���֫T ��2B3����9�T ��'�9Y`�s�r�3V�l:|��,cX�(����t��2w�osG�q�U'� ���j�wM,6$K���.zsh�G�1Q��a����H���l����x;��\��b�\���7��[��=��g�茬@X����|��K�cg
�0~;J�쉫E��c�@��dK���NW9iZ&��������rdy��D�$��'}@Gq��C��W%��O@�ʙ�"[�L�]UI�k� q�u{�q��
v���\M2�3�ZqL�<�ݵF�r���M�k���4�+��Vq�ㆌ�d��o���`�b4҉�uq&w�!�Yr��v8 �9e<����b�����5I���g���N#}�:�1����Qdᷗ���-��:WT��d����ϻU=��	=�E]�����։�F�)��>*�^�e!-���'&&�p����� ��5'�_SL�1/i&�( ����`�	��OX���/4�P5u]���Sr�Y��?�P��Q���d�W��+���m�X��`�Вxۧ�,ݪ�AeV0�R	�k���pܜ
�*Pb�m��Mt�>�.�������ދi����P��EX�m��^\!d����=z��t�4�M�r��?x ��ـ �6�.��Jz�[����_� �ՊK_K�h9SB�\����\\\A@e�Cm}؞�du6q���m��S֘;��2%(���&�=\�kmh @��rs1�<�i8qC�	��;n����Xm6@n8i�,P�� ���`𸦅V8�殠��eE�p���_���W+�ƭl��u�E�ɻS=�{p�>p�H��E��m����D���/Y�#L��ovH�r�x�X˖o>Ժ�Ir|�&�����2�\s����)��e�pE��=|���RؓN�4j�V�~�1��O?�I� I�'x�r��`=>Y���^!�
��|���ٴ)���Ly�sT9�I�m����(P���z(f*�<*̈́��3��������jv/���ȷ`��PST�bSӠR!��v��_���(�h�����j����}A��%�g?�w��d�B0���j|�|=���7��dp� �7�����%�" ���g�)�j!g>��^ ���9W�q�*��w�g{�&���[]R����bX��o<�dː���2ǖ��aW��]�K����Cu�mřy�V��V>R�Sev��}�]�����)�,b�`�	��V�D��sS��<�Ƙ}�Za§�~�7��-w���_C~h����ވ�������Dࡰ��=U�ԣ��h-)�G(��xw���呚N�WG(�.��f���ʸc���S�������'��!�����V��/G�9�]0�E�v�տ/�V�L��9e�	I�y�h�2]{£�&�Ê0�N�i��� �ϐp�(
\0�5M�A:7�v�������.�]��ce=��� �"B��@����L%�s���J��F��aY�_���x>�� ��&�����N{ݷВ���e.PaeЗ�8۫��d���*��&�g�žX��~L����y���/)R��X��D�=�d���X���ԏ�uo�΍u��Y�
��Xf�-������~��O{2I0X��ES�mo��	yA���[�N�~+T���/~H����Oz�
[�j�ȞD���d�8El���r8+aR��3u��6$�KX� �� /�k;g�,/�j�:6T������C�QP[�O�Τ��ld����W�'>]o �c�Dy��x��R�3G�����Ī�f+�"'ƦN�(���>B�g?�R|���*;4t��Ł����(ͽ|�ݓ>8i4�Q�c���U�-)+UN�c�H+�90��HY���F�Hj��D��
�O0��p�ls��h`/��2$�	N*�~&yTa�ߔ��(���W���t��%e-�}��6��u`�=���T���U5���T����Y�|�e�X��4�I=���_���v�j��ǢQ]D}��<ER�z��R������tmMB��9�
1��SFsUMz��)����/��H�bm^�kv�K�J;�1c�m�c����,��i���(�9MW2�L3���wōfiq?�Sw}��A���8�8D�taҳ�u�a����*n�@���W�s¾���)}W�r/&$�R֘�G��V!B78G�����~&z�^dFh7��Fs��qH�ge�5�jѷ������OD��S�n��!�zI��8СwM�������/h����ޖ��}�G�K�|��m&aJ>���E�=�%�#y�4E
'	7�΁��@ A�z��4��ǡ�ȍ����a���''6P"(+����B�pHk��DW��b�x��#��_Bܝ��,?�j*F�[�`go4������&�.��[q>��0\��:�QOm�%�Fճ�.;�߿#V�*�0����e�%[��,������{7f�7I;��	�ef'f���[u��$V_U��	�3"��_'��>i��<H\��`�v	���&25v�Q�M�-��/]H�,���PC��3�Jh�=PGAl���-��=Xp�]>�s��� �^����S2�y�)�r^M�]N.��lO{G��Vs���H}D��y�N�sj�b<nD��0 b����i��t�e4E�V5����L�F�Yi�]6�ڴ� ��iHYٽ�T[��7'R�]Y{�:��l0�_�]���*��������Yb�M�A/�3n��n�e?���pU+��۠�;`;���	�gD�Ȟa��Ny_�X$�^�����
�N��)\���R�������on���p��)�^��9�����-�zY\�˩�<�'ȥ;k��J_0�emf� �4.F��?�ߚ�3B/���xc��95x1s����f���w�^���ϏX��2�:j��ծ�\����e��#�f�XyB�1����/PO
��@41T6��U�-\Ovf�W-��N��ơ@����bƪ!W����g��q�� ����J�
�+����7p��/^[�
TOg[F����8mts66l�5 ����h!���?\R=h�A=�Y�C����[cS6F��7��k�5�M|���������=zLV�nD(�]Ü_�F��$ͱH��
��S��#/G���L����]��V1�M=KDUۭ�#��B
�۰�̶�=�ÿ�{�ny��A-b�gp�����Q��1�3��
2�Z��ckag���d���3c�ˊ�@`ay/��od[Z{D (e�=�z�ƀ�<�� �k��̍��SFS�3H�5�߽���QJj�xͭ?�oj	s�y|�e�z�&E�Ў},�LN�G �_B[�'9��`U��s�}��0P�쪨`?��G�)z¼NjYw�ȁ���0҈��Ch�T#��bE��-8X�j��j
�-�t	`@z��gJYj�Ɩ��I����gL�41��;+B����E�C��^ker$�{52U&	�� UX��z�����.$�f�����%=k�\��c�	�s�$�z�*Aι�
;�Vg{{Tvm�ԁh6:3`��Ta^���s�*���EQ����x� �H�!{'<L�*0�5�969X/�0���9�hK��2 lF�4���m�gY�U��)=�M��	�9����Y��L�)W�7ӭ$$a)��b���Ђs��-��@��� �,L����J��!h"߳��hW�+):��k�0s��r~�pı2L�1��[e�<+S�y;��Y���Xۋ��dn��$=Hw����ۏ�,TKC�F�B���ѐ�5�]͒�YR>op{�%�;��æ^�E���
�@3�ka�$Tqa����䊄�<Ԁ;�k�낟��VN��˒�_&��7ҖP��N��� ~4��m7�츺��q�p���ز�I�����'�;�"�4vO��^��ٔs��SvɪWd�=�ܛ㡮�d�j�f�F�B��0!�6��R^�O#+Nw\7Gn�3�Wqp<�?'^�d���)�{�x��Vŷ�Ydg;�L*�����׎��K��a��^S	�z"����n}vBs�Sj<dӋ���)Y��̴��5\�y�1ydB��("q��ĩ���(EJ����R�L]�%>OZ'�}����'t�7!��_#5۠Q�O����(��9"�ә���ඌ�DӬ�ա}6L@�W����xtĉ�Q��p�ȁ��^�jq��P��w;���\��(�����J����ǜ�`�e�_�M�uf7�2��Y� ����{��V�� Y��H��V�)3�[	���a���|���t)_����4pZ��_Yc^���soR�?��5T���a��	[��h��/���3�A�c_0��X��\SV���(�fO�1gu8�/�M:,��ޠ��4����[��{cg�����fm3��iI��؀
r���%�U���/_��0m���[�jz�k�Az����39�^	�D����:���b/۳�
v�]l������ŐG*��7A����;��.B_�=���џZ-��n�گk�񋹋��xO3nc˫?�$@9�G�Ћp}��8���%�~���f"s˱<k/�:U� |}bB/�ߢC���>F�V��g����N���Y���l�4x5ت\»���v�r�.Z�]��,�g���T�ɞ ������GS`�	���� c�=El�g��d��u|7��H.J�f���A��:т�k��+��Kc9r��v A`�a�1�-x�Q�Q�<���9��jۣ��#�<o�` 4��ƶJwS�a��-w��T/�&ݶ��G�r4���
f�����!l平���8�F��N$S�+
����g��g5[�)|Ǝ�/��c	mQ��o)�?:�q�[(���� �B|��ݱ����^d������R��,~&oO)�fG��Yv�d���ӽ��k�����#Kˮ�F���l*CcY��J4'�H�� `��b�����@��eB+J��@�
!�X���:]>5�'5>dem��w}qt.����z�>G��'��Bm�p��-!P��]2<A\+�+(��;��햛c/�0<``���9�D�հ���~≋������@}�E��pܮw�p^���D]�2b�i�?�����$5�9���#R��9��$� ����#_�F�(�O���?3�M*���c��OC�mt�/{UF�ސ�����V&|J59p诓�,b��X���}�v$��Y~X�vؼ���7:�Y��Q�	��q�~L &);��]�+6��D6�`��J[f5�/�P�S4*�D2P��������V��*����{���S;�����*�9�#R���&Z�n��}� ��t���o�R->G|ǩ���p<6�@�z�P�D��gó2�J�y�����t��gn)�����ȕ"��8��/�7�:�Û�jC����*��)�)���������_~#s�y�O���/�׿��m���d�Oc�/]+$�{�Ծ��7uJ���#�<��Lդ���w�Yu�����N�� Q���{��BEtTwhW
��,���w�4�H)F������:[�{K�8���Yųy�7p��MF׏�<S�#�J&�-�_�
n1s#����Rz�Wjɔ��ӯiٝ(��DSC_�
'�d65H%�Z���I��[Ke����}����Zv@��RV	��s7j���$�	<��J��i �8��dFbx&!��5��ջ��@�k�BƼ{E��[:�@�������K��&�.�u�u�J�Uagp7{i����J8����,�L��w���vEC�'-�S�>^(�0���M�/c�����@q�?��q����(�5�&=���)2?~�.����[ɦ���*#u�pw������ȟq�l�c`p>�?�8�OԴ&{��x��mJ /�w�F3#����~�Q�u	���H�����X���]��q�y]�)o���w&�4J���g[,t���MYi[�;��P+@Of��1Jf���O��$�I^a�X�1Y�O�	X�7$b6�`�g56����+V�p��������ʷZ�w5�=���d���a�b��p�d�x]�WR���r1v��׉ :{��xSyaPDwԲ�3�$mZ�-:��G?2H΍���<c�x��uc�(��n�u't4��&���7-3A-�o.f(Z��R�3�/��Jש�Rd`�ǇT��	ċ2k�T�8�J_��c-6����k��`���1�ݷ֖�i�p^}z,����e��|����+aP�����j���;���p[�od��E#�v�zڈ1?�x��RǿZ!_��:߷~�z�2`��� ���n>��Ė�MSz}X����
Y1�-�UX+�8�MH <��?�Z/+9X7S��1-�-�^N�C֋/_Qv�ֱ��GKS�-��<>I]�k�]�7��{+o�	�[�{T:�@!�zx���hz�%�jOg=�<��*�*M� ��6v]�r�3c����e�����z�m�z�q�yR�]�˟5��Y	�ݸS�N-�0�a�]!�4}C�tE+�`
�V��K�ǮD2���v\��S�_�:�^�#"m�����P=V��WX��޵x�������Pi�&����0"�f���a�J�Ѩ�2�a��.J��>���ucY;���l�R��5>�N6�n���j|8��/��+��Q�I�n��{���FR:�R��0�����ga�;Ck<����1�b+�FK%�i������tj������T7��K�j�(A��5/?s֓��`0	]�0��?z���\5�[�K�E��g ��5��DnU��QT��95��s�oOi�w��5�հ��ap$`kk2�
2b���c�Srj/y�
�����>�hOبy:S{�G�S�J��@��v�}�$�ST�A�D5�)�� �3wQ�)�n�񌵨o�k��sr��1"�H%��4�Id.�C����۔�XO�6з��4Y��nK�gLV����O<z������^�4�_B^o�&�E-Ma�I׆[^�,��q�ag����Eu5�R�du����e�4���4�t[,���Z�q�G����p�f *5q8���7�E��O�IR��B���(�+�ĂJ�p�6~��>rG���d�&^y���S�k@�r��uV�R� {��죌~�p�\O)�%۲���^?~z�[��@�3
���>�dmտK�:r��;�t��������b5$�F�,��ojս$N�&ŗ[�"�����7�)ý�u7UxJu��ؘ�)*M)N�R�[�!V)�{�,Q�ma��u�<qXa]�I�����w�V u�2h;d@K��
{ ����It�㏩�ݞPUC� Q�I ��
a�Nٚ�OW�x	@{��|���ɦ>���������_#9Ԕ�&p�xȩ��dpvv���iS��&�(5�� �������I�j�~�;�kԕ�,Z���N<��o��ہ"qa^	���@�:�A2R|$���`�sf2�Z��M(f��2����\Y��L{i�ᰛ����r�.�/�Y]�s(͖S��5w~Q�P�5v�oB��x�C��G�����H�@7Z��.�WĆ7��WhC�����DS$o�������������,5 ����3��0�����|5Poc�����=����R�4}�e�ꁗo�eW�Jr�*�`��}ł�o�!�W6�7>xU���/}�L��3�;�ðY�3�B���9_��żl@�'��>f-�כf)JllGb����HSy��E��j��؜(�_�*a��a�I�ڜh�Ǘ?�*-�P��#&��9e��[ ?�7m}OkO��W��CA6�}�%qp�!?[e�E�<,`����y�5v�b0-�U��J{�\)T��bk�n
��UoE`r�j�~(O��u v5�c&f�"W��C��Qߨ*��E�
ϓ�sǯj���sO.(��0�I��.Ɇ�4��#�sӰϛg�����ԭ�	󄭀6�t�)������Y�C�cF�������U�C�<�)t��P�4��;�1o��5q�����8Ƈ�zX���` 6�sbZ���?Ӫ�[<�i��Йw�7I�Y����š�G;��&h�;��)۞�_�c��������B+�m���~��H�ں����$�P�6��#@�r�^�s,�8��xS-c�E���*'�jU����Zx��s�	� ;��e��B�Gk��S���x ���\s�0m��"��c�k�x��t����t�Xw��a/�̝լ��m�/~9�9���F��qUȵ�a�rJm�+G��F!��M��*b3��R�d��ʷò2~:�hA�b*�~|(���S�Lf�h�S��w�O;�|]>�{� �Y�=�i+���y�`�65��Lg�,�M'L���w�'��>��j*�z,C��v����mP܀�?O�_�� f���f��>�I�/sI~��)eZ�!%2�E�>y��vڎ"�E��d�ao�5�\]k�]\�Y��uP2>�h%��o?��*������G��� �ׄ)]��bi�V�*ߣ��.G�9���9�R�h>�-�{aew�v��v�P�����y��RD�|ހԅ-���YsR���N;p`��e�R��D���5%�^� I�Ax>�Q}F���Ԅ��'9���u*(
.%t{&�����e���!�D�k]�P�<����}j�F�ʜ���1Ւ<|��(p�8\��^rm��O]Y��=5���~�ΰ�'�u5�Ǩ��%A>����$��M>�`�Z�=88����^�%y��@bG��A�#B���RMk+$�=�|���^!hl%Ό�,r���.R��ڿ�H
P
�tZ%e���{
�v:�^;hd�mh�ߑ�3�@�@7�� @�R��~2l�.�d+����L8\�������
Q\��.2��J�L�F��k��u�Ɣ����W|X�!=��b���i�]Z���\7~�F��_������=w���\��n��.��t��NK����z;Z��O9K�cW��Yʏ��-i�x&�FL�\#�s��j��}��e�1��Hv�`=!3[g=Z�n%m�N/D/΂��@�_	ru�����H�6J�Y�:�HIe���. �٨��������Ȩ��GѴ�,m��Z���kpt���c^��N΋�=Ѣ��R�� �2I���;XϤDD+k������Q�� !�T��ړJcIH�fkYM�r,��j�t5����S�4�Ώ_�С��`	�y���/G�0�����֨���=&}U���Hf��ag���-�Uf1ea"�jVF\�_p�	���Xf�V��1	mF����g�p��S>Ub�Y@S����]Q�U��J���c�fMK|H4śZ���S�5�xcu����s�co��_l�Zp>�=�ۭ�c}ܳ;U�TJ��]��V���@���e}o^�I��w�~Bp���ӸQ��Fl��!�B ��+'=��x+��h���4�����GjIx�9jb(��[��J��$I�8�L9X�sI�k��v�.G/�~5���..2ך�@I_�Դ"Q�����k!�u7%�-u���:]��ٜD!�bg���n���^"5e9��K�Y��<L��$��-��)U����S1S��u�����Ä�6<��u=��_�AT�	@ٖ~�8J����g.��bN�JL���[���B������Ժ9W�B/��7�ۘQӿ�y�^<	�_�{�#@�[�.�q�e���7$uw�b";��k��u�px�6|+�$�JNԓ� 5:����@qBe�'��پ0?V�$��vBvfWQ֬�b�2.����9۾�Aҟ7���Lʁ:��7 i��X~2�a*�g�����>�]�Ⱦ���(��7J�d��+���"�m�!,��_T������+� y��x���NE��2�o���u������.��5�SЂ��d�s�g��>��J%���= �Z���D��Em��f�/�9x;��B�Iy���9#(d�����Z*6��L�]�R�9�1�f�N�=�y��q�A�w�8��tu��v�O���$�$G�܎����YEaL˒+Ҡ�^�)��}H
�{�Q%��^��`8�"�'+��Gv;���0����xo�ao�sQn\���+H�s��s
�G��Og~�����o��u�iͭX+)3��Y�Mߧ� ���V��i�@��! ����B�X�7�o
����SgF([ͣ��>�x�
ܱ�(�kO�f���H�g��`k}����4��F8���t�'��/��Ԯ�o��YOen�#KcݼW�:=�V@mجX�j��l�W�ǑC���Q#������b/�*}��d�E>[3P���5|�S����S���:- �8�M���<8�-{"}�nnD"�%TƧ<�M�&\�&�й��ɩǛ������$�N;5F0k�`�.&�%��6�Y%V����������ө��4�v�J�H��ԑ��lu:y��^`��4yK�������X��w{$����a�nX��!�k`�hS-,$6�J92Z��>̕�N}bE�T�k�Զd<�2�����.盔(pÜӪX�4H�����Rr��k���ơ��Z�~*��ƨ�RIT���'~U{˨#�O�s�r����=l�3�;wW�c�J�` -���]��O���-e��ϭ�]�E���w�lw`,%e��}��b�t�KH��]@2:BE��%x��\�)�@�2� �2��|�`�����Φy|)�s�%r�d�S ��4�X$<�(��Sm�ڳ�����:�gb��*�'�{�[�C�	9�5�vGy��O�d��U��D{u7�@{��=�%�PY[��<�s$S� ��B	n�=Q��@�e�x0]N~-���d�]�1c���,�O<C�J���|��+�ͽ�-��J)�C���e�Q��HǠFo��������"p��X(�lm�	�jS���y��A���Κ�`��}��M����%j�K����(kTS���V�m.p3�N�,�dF¹i|�?�jm���Vx�.��h$_��x��˃�u��H*\foُlŏ�AP)����o`��ǥ���~o\V���0t��q2�D%/"x�s�M���΀(q�9ꏰY�!w�Xy_��DsYM��(j��S��2�s��&��ErCS�!��+�/y(�A�au�Mgd[5c5KV��-�d�s����b�|{:��µ	�y���>$�D��T���PvSl�e�K�	eq�s�b2Y�Gr�4���gB'�z�g��$3��4ȂO�
���N>pTₚ>L�� ��`�n>FJ%j�y,��J]�3?�#�B���.$��^q�
A]�Z֗G��#a���,�(�t&?T+漭�o/�Wq�`j��c��1��n�ب(�������7�n�W^�}�;������
�y�l��ڒ��~rG�{������kY�F�B��i{d��WO�JMj����_o(t���53~�{|�(�Ш���L[����dIN�;�sb���(��Ie_�xr,<�aE��N2	��`'�%�������؀�z!!P�"n���d�5�A�g^�I�����Աsu^
�sD�v�d���%�h3֭�¸�2c���gG�=G���0����Ԙ���	�����vb�Ư��=C�w��B�=�E;�rMD�
�����nL~Y�ɔXX��H�;�Wɺb?``u�zNQ[��j	!�����:��|Ĥ�k͆ ��Q��y�l�ׇ���Y����od����LyN@~-��K5I_2c��W�Ċyk�H-�`�Q�sָ{���^Ԭi��(F�7���̾����bsn7���'��[ �qpO:F�$�l�t䙔w�-*sE��+�6_]�)?2��,?E����U��~��G�cf��r0��"�&�*��ϢX|����Y�Lg��DeQ(�9���	X^A���m5���F��n]���`E"}q��a޼���5�;�u��t����R����%7��d���vdT�Ud�"��EC���8 BU%����9�bʿ���H$��&u9��4W
+��M�uF,��&����0TYgE"5���&�P\�&\?J{)���%��6��f��	s3m�:u���XE����\�%@�F��{X�n׵-K����e�XY�)�%��#���<}2
ވ3[-dc��si��]�Hkʞ]o ���'�>�C؄ҟ���)�6�ۤ`���nk(�֡�є��� ���O����>jy�٪8�{�AL�[
3���H��H�6[��vy=��'�*��P�H���oVA��O��?��f�ܐ2�g7�[ė��֭0�B`�-�ć*���/ʓ	F�̇�T����Å-4��ç,�C�4�ժh!ԏZ�-bi�4��q������J���܏fm��=�[��'d{�<2Y$!'����گV��:3{�Ԓ�m�V�/�x6��ń��� I4q�%�Q������#8{-f���N:��B\�;@��kJ��>��MDy�w�DO&��KMc\���B�������,��7��[��=�~7�	ߐR��Ė'q�V��B�#�ƃӜ����|ja�v�uG��_�������G��Z��*	y�c� �V�i�7JʃB��Z�!LB�q~tT\�����+��if�E�(v �bG���]�_����T_Z��9�rP�]x��ќ)'7�Z�7=$�7�J��f7�I!nT�\ ��L(~߬2����1t7����E$_@���A���G��6�1f1$�8'`� }�S{��p��������{���yv��Qǋ��bp.�gN�JiD��i���W����{Kz�$v`�J@�[v�9wP��2�����V��������4{!3b4a%���m�W��Pǣ�~�O�̍Z��}������.��4*��q��s..�:ڟ2]��7(���pS�U}��r�E*�e���)y�H�=l���d��o�|�� �l*�kP+�D#�/���]�-�Vi6OG��5ԍYM��m�0SA.�rCF�.IAP�����m�JWB�x
;��N�&\���=0��i�������H����x�k3h'���(X�hN1���i������Z�-���0ncz���b�ACi�GA�����mn�+��Q���]��!���	E��Dާ)8t��8��瑍�B��'}Ia�����[	:�+���Q?�.䢟��o��;���6�T�k)$��{վ�3ۑl%lu�̢"X�0���]	�]�1�;�^#�>�e�NP�%|�F87����r�_���v�#�d-7��I\��g۝]��H��ϐ�<3aЗ���f7��H��@�^!�-@���*��i��n�Dp���.z�>!Q_�툚� X��ߺ�%1�M� _���S�T��n�3<��%&8��õ�(|t �-�Z����ɵ����}�@/6����zC��w���@�6�E���&s�ծ�5&a�㕷ܵ��PW��)�8�g�5
�H��9�@b�z��8�*���^&۟����4�W�" �<���Ͼu��N�8��7��.����o3y��Tׂ����fD����[+�&���`{!��2N�F�u��5�&��Ӽ��gFE�5eDw{B�`	-�	ܿ�(b��a@,��s@���8cS/��v�.!��iX�[~4�m.I�r*ц�h��/�қ�P%9�k.<U���@=r�l3���Ì��VY!;�y��n�r�8ݹv��d�x�g�Y���U�"�;�g��=�`/U��du����L=���X3�Uq�ev*X��Dꐹ3}@+��Y�8菭,�t�GD`.s�`���� �Q������D�&��©��AG{��N�GD�K���>��T����F��s��jy'�z1���Hd0b�SuY��r8M$+��}и[�>����y՞7JS�j��B�S�c?�c�^�,[#��i�jR���o[��i�h&l�o(�!�2�3#�f	Ea�+���D�&��i����1k|EkߡL89��8c��m	����-�L��H���udhr�&����ڭ��F|^d��7��(��rp����Ѐ\��zy�7����n���ZQN�l�C+t���s�X��7��굽������G����S�:#�������γP5��s�)��������Ѵ����߯{AN�p\����<��{���������i��ʸ�x���+-J0�Ѻ֨[��7���B @!²P[S�z�a�`��0�ܘ���(���6R��J~F�\BW�+7�3��T��u��t�U�{���<����
Jhs%C �a-R@�wM�1���2bA<K0�P�����/8�(8��5��(V��P�5�\�n��lKC!�r��u3#��?mI��V�L��(G��1����d%�8�y��:K���"��/��Z��%sk{���<���o�E+nnҬ�x*I���O�VC��_����Q��l�H�SO�M�ch�l�М�E���}HG�����jm����<�D	መ�,Y�1ާ��jد[����!��|�.0�~:��k0���1fԻaX9wF�
�+��Ф��������� �*Z�mP�wL7$p��3�c�MYT�|ۭbl��YO�94�RV0���![��������_�E~Y��/�ٜ=�Pm�}��2���r�WL־�B��� lF���Z\���2JT ��1��H�R���S_�X�@��y��8�*�lb��W޸^� �h�cn�N���Q��&-N��ȫ���L	�w#��8��U���C�l�I�9�{�uxj4��N�MB�����v��\W9�uP��Х1�8 r���$�ޙ�3"�oXE�)N��_w���8V�6s��1.]��r`�����U�.�o�c|��ȯ��K��U���b/���qX^��1�K�7�Fr����f�`�j�w�E�Ux�@m�JtկHv��k�T��-��kr�xdz* 1�"�u�Ex�;�,3i-R���3SKm�cOR���?I�j@��ZJ���>�YRD"���3�,���$�b7S�/�!���	��s7g.���u#�T�1Q����*5�~IO�ک�^)p�� p�JQ�3��o��c���ir��7,)R�o�v�t>�W�Zu��i.������ߧ|�u,c��p����)0����( �J+�+�;jv Qs�`�ބ�^@&�q��oFOp��v�Œ���4	�����FS�W"�+L�SMU�k�:��e�'Z�qh�wX̒�"q�^{��M�Zs�HFX�-��HF:O�m�D�^���rS�k��Uw���&�j���7��B�e,�b9^�3M���5���z4�T9k�μ._ J�HE��t)�O|�����`JtA�y�Рj�1NB�X��"��\g�K@⪄w���L2�T����=�#��<��Ӊ|	�;վ���7���]�9��a�g0�5j�]�Ϲ�������z��@C0�`��>�����Q7?�2h��[b{���D"�*��X���C5k)�γd�T�� ��]e!U�A�zw�V�Q j�o�(R]��
�2�~�s�����%��*��g�5�M�����ac������C���IZt3\ϲ~\�VNrN����=R�BÞ �݋���=3�a^a��=���uJ7#�=Y���J5�� %�*Z�G;��{-l,�.C�����P���U��������Xc�Y�z��;��O(�HjZ���1j]�<��a8;�!�������JD�p_ɒC�&d��C��E6N����cA �U����Ne���U)Zcl�D�B!N��o2�U)�����$q���/�o����<`⡘�M��=�?n�ucf��7�T�{�"�)�ͫ���T�I}hJS1g*G�� H�`+���T���_n�|1}�c+�-�W-�>mn"�X�`�T��^շ徸�D\��".��<����V^gP������_L��Nљ�}��c	1���l�Rt�f2�to	@u����.�m!]�M�~�*�u[��0(W��y������!ߧ[�k�ŉ�����I�r��P���q��r�4��X��&د�|/d2�4��)�F�AWyu�OK���D�:��b�e
^b"��c�*J�a�f*�T`��Ȉ���Ͻ�y�"�A��x��N�M3ْ�6���Ś��fn�7. �1>������>#G�(h�sU��G%��C�#���*`�O�G�٘�����^�Е�;T'y���� G�s�/�����F��r"�8�����|��j�_�5�������e�4=�C����$���I�����8ڌ�#l��rYm,S�%#�2ٽߦ}��X�c}�$,�9��;�W�:��1<��p� �>�	AM�Z�2S���͂��M�v��f�'S7����l���D�;�e�xw��M\�����Ĝ���jb�'/j��_U�;ߵ?��w�va�����Q�􈻰Q�eT\���ZE��ɀ��`�P~��-c-0��{�6Xn�/��;�~�~�>4� 1�\*�9�_Ld'<�JHɿ�J[6�����X�eZef��B��E-��LοB��9����%Hj�U��$�&�O&�o����?B����ŏ�-Ư� ��:x鄆}k�����B�C,]�'�6֕�� �M��Iy�}��������lG���JUu������;Q�Mg���vd�D�6������Yَ�9�%��f���L�� i�����G`�Ar�f�}%
>�.B&i� qX���a|>���i��2j��e�1o��G|C���D��U��4���o�O%54���"����K������\-�:$^jQXK���b� (���#H�S@��[lu?�wE{�B��`d��ԇ5��q�>�e@p���y��	/ӧޒc�*��C�T������o�c�	�����|v9��v�F�<�E/����{s�6�T��@��uY_m�гj��0�f�����FtIU��Vt*���_��'_U���yR��Z�/��gS�՚��r��V�ؔ�����������۟W�[�%�?U���I%`(�/}�`7���$7�up�D$�:q��ek���K^L,~�AFS���J���b���ct�2���
��GdM�.�,�0Ȫ�D����i&����J=��؂-�?��6�וYF�Ȅ��3, 
����Ck޷[���A(�9\k�q��~ڤ���T�c�L2���Nx݈�J��s�v����&]S�r	����$��^�顩g�TXQ�ck_J�y�'��%U��B��]Ss/}�,Ԛ6��	�ǨA���݄�b)J5�u�Jz$n�cw�/í���&ƨ ����黙�p:P�>5�9T���Sl�'S��ni���@���h
B�h�xħS�.�I��T��Diy������g��^�B��oOAx�_��=��@���Zg��@1���b!֍࿵�p�};X����F,��,7tɲrˏ[��1��l�����k�(���!\�@�4�����;^�F�ԥ�+��U�?Ƃ�ZIʀī_� �D�ţhhUfJu9*��?��^R�M�&yx){b�ѾK3aD�7�qqU��X��zE��G�C�W�ءj،�t�b|�,�Дӈ�kM����C�T2�[�.d��t#o�BFl?�@�`~{	�يf$F̞	[D� ��
J�yD�՛Xl�2���Hp�]p�\�)��N��u�vRL����X�2�͹I~& ��ې�q�r���`�_p`V��O�ƦzV%��H��4&Ւ�v�)8I�ÒjO��6�k���T�V�D�4۵>D=j���k�hC�_z�!N�܆G��
v_Ӌ~	��M�Ղ����6�#!�V1�lg\�Ӈ�':dn�O&���mf��
܎��x����ɍ�BK�T��!q�5���&ZV�wo j0��<��9���C´_3�z_i8�{3�)z+b���0B�u@#�ws����2�4 ����Ҏ��^j�K� ��;;���L�9D�	�J����8��h��M|#@	�9*E���E��M�Uk���+��]V�L�qHy�|�]��; g$��ϵ��h�i���p}�s�ϼx˒@�����@[X��DI�Nl�0�6�̪����E��x$�oW��ۤh�, ��I����q����ho�G�zO�HB�)sun�-�˵�Vy1�J+�d�`|�[��l~<BP�-�a�T3�C�����>��G�΂3'+\;p�+����Z�)Z�,�X�WN��N��/x�8
��N .����m�pz$ !t��m�󾉜�a?�*H���f���H�u�%�f71;�/��T')+�2�d����I��9�Ԟ���*����ɯ��ֳ�������ɽ)���B����ֶܲ0$��MI�@5��;��Z��i��HX��F�t�߬��4lx,O�o�0_���o�M]b?%C�&��}y5���m��{xx)	��F���E�L�/
nz)Ms��T�+������Z���<�'4}�<�`Мp�����:q�,����ݪ5LWRq�:�^,=F 0���NW�U��5P����������|���j���0[�w#��Ax~�:�m�RH������PZ�J��@W�Z�fR�Z���jy�����ｎ�&�Xt2�O����8���Y���`O�:np������J����%?�G���*z��E[�
��[T���F99"���
����Ѯ�a�u�ܷ�5�na�G{��m���f��:�kp�_	R1�OJ>��k��ĚW��lv�L��F$����3@�L���͐�LV>q����6o�}]�xZs��܈=��Λ��[�a3���
�}zJ�,lh�t����	��k�d<�y��W�J�ߤ&�n�~��	��Eq�>L����m9��r��2�oӃ���n-P���;��6��76Q�X���aY�o�Vȝ��A��:4X���3�\�+Ȯ�����+��6���+^��6�8����d���r���|��in�U�QS�qκ*�,1����*7��4��(�3�.XeY*h�=��p��> W�f���	8�u����+,��Փ�?���O��:��~�Gi�V��bA2x��1�� <q��p]Ц`�DYH��rH}8X��^���k�P ����IC��I�=�C_Z��"Fl�R�%C��B+�w��� ���#��܇�u�J��B�}�0���Թ/8�7��	��ﷳY|zoQ���Ž���D�̐����'�c��v�Fi^��fC��
K���Q*�z�d��vi�_����������2.�\�4&G����K�P���\�jn�5�2挥��9{QK��<�+XU�&�l�ӷI>E@�}g��2'[_�4�u*��>��Hu0oE� �a[G�/ؤ2�)�\���0�)��׫r��m�*�ʹ'g��k����e"��r[��!:'��QM�7����F3�@h'C������K-'(Q9ڏ�BV,�4�=F�g?D��rP�;�;�oڳ4,c�--ǔ�j��X[�#��<ۯK]p/ʁ<�kW� ��~��$5o���IE1�hGJS���FĂ�=�7R6��^�,�4�_��U���M)��ʥE�7��t0ɇ�T��-ַwih]	� W��I�y.��z�ݹ�\|	7o��MU2���;B�=�y�9"̇��R�6�Z�Q;����֕��Y��dItq� ����^'V��dt����<)��$qH�`㳏@b��[YrIE>"x%��v�<B�%"�!*��ً��L�+�Ռ���	x@�,\���Ak�V�.�KM2��*���^�~	�b�K%�U���������BT�io�⊯xjY�9�3O�"�7ǌ1������Uy>�/�
hQf$?�eb,���h��Jn�P�cMk��q/�M;Q��]�0o
Q��$��
�ܲ�6��- "�(��`|�0�h�������l!Z���W�����cj������a(�n�{7j� �qH)Y���a�����J;X��w�����������#7������Q1���(���O�j�'�`����$�T �P�Sl6o�f-�3�r�^p��G�B������+�tP)k�/CP��:?�B�������>Tf�[�7�/�BBf�����)m[��
�S�OW!��Ϝ����ȡD j���)q��D����_�Uo�nc��E.�5&�@N*2�3����l�Z,�/RO�D���O`,b�\ƫ��᧓Խ�uI����N�@����E�%�u�$�dI��,!����4:���0����`�+}�u�ǁv>J9�9��x����:돩ī[�|���WdT�%�K�L>w��~����@>���FYU��/�?�ύ�L��| ��Cp-0$Z��V�kx9��\[^P��'%�E]7fc��SdLGϗ��~�� ~I�c{�ި(R��q��D�m����@m���I.���oz&� ��e�ĮK�j����������A��=[Y��C� �,�~ lG̃�����/��O�����:��3�V��J/4�W��ۦI"�z��1"k�"l�A~?��{G[x��s<j�Y���F�������l�+����������j�[�*�{MSԛ ���,I�`=aFL١]S��ݒ�d�d^�>����`Z��4��M��j�dxP��K��;�M�\���;'��>F��[`�u���28*�+�\�X�p��ɯVZ�[��5#S۟33��5�}���]X�����9YL���U	�y-4��Ѷ��m�"s���@;6�7�i�D�ͥRO�P�x�ֱҥ³,C\���h;%���Φ02ubZ<���2ƚ1��֯׭( ��wW_���?�9l���V�g��ȏTKs���^��5�>���R��nG��H���[���Q�|ݖ���S�)6o�<\�=�~��;��NK����34n(	l,�n�d 誨<��
�7�XJ�_�.�)�T����nǅَa�
��R�u�C��+�����H #���归� �,֧�d$���*e���V�w=��b�b�pa�,��i}#KWr�6�����<	?@ ��`[%͍in39�K� u�W�Q�~�GY�D&�@���T��r�y�+t����н������5�r�O�ʙM���L�����<�����'��,�[�:i�y�Ձ��4��]����<��J�(�����F���������X�r�xf��T�����HY�8����\B��cxף��H��8�rX��kH�&�bW
�y�q���x�� �4�jZ��9�W��(����^�s����@�����/Ų׮8Dc��*�+]��*_1`��'�4���u����HM���v��\Ƴ>�t�z�'07����9ˊ�qO�|w�K��h{7Q�S�:F�x���D���ۡ�vl���4S8�}ù.���%��[Y��ҙ� �T�ܱ�*������T|5�D��]d��26��H��	�	}���|ȃ:Wm8S
"�0 �_6f%(�����j����-�v%گw��bU�HU������NG�P�z1M5o��><@��E-ҾO���pp4���6�6�.�h+h��X�]�菀E����%��k��ͦ�$c��X�h/ȉ���8�N�����zh�o�uv������p�gʚ�eN喋^�A��or�`^�I��3�OG�]":��������w���#���߸�9�pb/J`�
f^��O��Z�}��.�F��Nm~DJ�'�L��π�U&�j�C�7]���٢fY��_�¿�P�L��	Z5���=������v���m�jXRR����{����qY�,M9=�%+�jrfV��Q@��d	����������}�#�ܢ3���IPٝ:����=
|�Y;�tH���%/�H��W���h����t)Õ�c�xo�	�>HP�^͑�jbj�Չ��.{p��v�~h���}2�������n����Ts�t�p��/���o�IPo��X�y��K ���hB����88�M������ �3H"�V� ��X-,-9���C��[�k�s^�Y�����	:4UIݲ�%�_ׁ�
X��
C@�+b)k;���Xd4g�˄�ͯ��B��\���x���d7���_\p�����۰�/���&1z��ǺNwf?���Y�-(�&��`U+2����^��w���9�;$X�Yj�*�M�@��%q��0a�:���$�K�8�}I^���Eb~�[�9���u���������z��E�7���`cL��S��uPΎ��Y�<�j2K�¾�ϓT�{68�b^������P��nE�+���B��2ls���$�	�h�sGr�c��	]��\D�Ak+�]��C�
Bk�����G5�2����	��T�)�~9��ƣ<SaWQ��M/������?��)���<0�:ݱػ��R\��4��a*|2�(��yOc���	�����u]��l��E��m���ν�~x��3Č����.7}=��V�i�E$8s���%\�4\ )�q`��̯*�˔��	�ð�^��ְ䡳r�E���n�(ϥ�0�pf�ۦ�������	y ���[&��JXZA�n�|ӗ8L�	���p����i��������&A&d:��J�[O�
�j;���\�k�i���Cȥq'n�	�;�qJ���&v��*��ȕw[9���}�<'	���q���Ϛ�k��pZ�OD�}#<i."�\�_R�۩�ߒ;���0z�B�\�h�5������P�ʥ���,�A�H��P+���������QkB�е!P�nF\o��Il�T�#q�5Gi�����q$�U���C��2������r}�d��a��hT���uq��-	�)m��J��;>W�:�B���5��hG^�UJ�*ID�OG��X����`t��vGPM#���0W0Yz<���eCi�����~6��bmev���`��os7u(�M1=RU�h��Wuj$ܼ��7�5a���s2���7E���ǇĿ[8V�Z�1�1(YL�BN/��v=4s�	����y�YN�?~M.�\+΄ؗg)�@�#��s�ق�k;''�ӡ|�n@�Rk/�Z�u!��m���!޻��N7M�l��'�H���j!+�d� c2�->Cm��V�-G���|�Ϊ������Q���ʇC��E����C|`D�)�;�m �l�X@�T�w��� !��ww��V�WV�,B�$i1ט�<A+my�>���yr�R��dw����3�lFJ�����HV�����\��l5%�Z�����_����k�@6P�!3��#'����}�
*�p�Ғ|1i�7��¸�ad�6���ㄹ����.���H�d2�7]M�G 2aj�'l�:�iS�d<�C�qou�,l`� ����}����i�U�;�X:���Ȇb�k+��ݲ/-Ѿ8�G�ɶ"IY�o��MS�}�Fŕ��~�����Zњ�� V���CM��R���('��Na��X�F0s�W��{EP��`G�M���}%~6T���j���%]�%�]n�##�[�������J8�M]��Y���PZ.,H��OϪ� �m�J7E����iu�g�~l��T���8SC����e�P��߯ѰY��;ۆa�ӵ>`J��G�f�ۤll�?ܲ��p�~D�=JJ�7�;&�hu�o'A��O���S�FĴ��;gG�2z'5S�E��"�2��Q;�(ӟлgZd��@B*��r���~B��q#u�#����7��i�@(\q�*�t^����PC���F�'��V������ha+|���R ��p4�h���Y�Lz9�8�����&!�꩚�O&�9���WN��h�c����k�+KA�Њz4M7��6��W�F���Ŕ��D�e��`����p���'��2�=�,�Y�R=⛮��ur{���~D�G������l�����)7��a#�C�Au_�>^�R�"K.G�fp�Z4*g�v$��������\f��K1�6�;T%�m_w:z�b�z�)�z�%�s2��tR��˄��.�d4�ԭehۑ�\�����T�����G�u���H`.{�h�ZH�	��qv��{�L|Ӊ�m���,$��g�c^Q��Ӛx���b|nf�����Β�)�GY�{ -��3�JV�ʟW]##�:�@�"P�cϠ���)E�
վf��7q�'���A!��9-��Bj�vF@R�e�<���S/X]��fLp�8�r���*T9.!�U����z�yt�1l|̑����b��E���z.���O)8���k�<��|24����h�;��Wv��	�h�U�e�"u��(�o�EK���n)��S��lT��s�w�֦��"]��*r��n���8�����p���z����4'Si7�f�^���#��؝�ل���p���?З:�y��4V�>�g��Y{J};�1�z�n�0���Yc;���n����^L�8Q�!��/k�o�8[LY�U�}%Q��(
N[�z�s��4_O��e�s�S�@�)�g_3j?}��r���_�.��>u�'g~p��(�u� |����Ln7��Z�GX5DsB�<),hnDsȄ��)!��� 6	F3#�d�xrd��G���������-�|�f�<���x|��}�]�������J��:?�K�a���U�8�F��T�7��/E�����чk��{�cf$�d=��6�+�!GymF������:\���e���1�ل����톤E\�g�8���y|t�D����3��"'�OEn�D�@)���; ���|�����S�)!�ՆF�Ç���Jz_6��F6�*i���1:<@;SWM���{���b�v���-#gX��&@��nf�X}oJ�@��"%tu

n�H�Ui�����)�S^��s[>W��bЃ���c���
)���Y�x�b0��ǚ�9w%+9��gr���PSa�CL�/|�� �tʽ�����[���>�+����c�Vx�B�m����'�4={A�{��ڔ�h�VcBY����9W�Z�k���;E`�zHy|Kִd$ Nh���c5�u]&;U?p9k��c�I#��bA�{�
�O�z�a��#���v J<0�Sro����]�%�(��18Q8ɗo� ��P��h�3�OLov�lY��] ,)���cP�Lye5׋���鞶�E��#\F�Eψ���7��W�'V�ҭǧ����c8o{�ۈL�.��君i����<��Ħ���k�s���+{�l1�>�y��S7+΋�/�� �Z��7,�pZ�G�HS�!���M���N3Z4Dd�l���I�\��O(I�ҭ��uo�=�Q)fU���� ��92�V��~A�<�3���x��p������&b]!�l�{|��Y�<��7/2�y��rG1�\�L���F�o��3c�Gy�5q�"+u偏�V�Z�����#��:��-ڄĬ��(v�� �wl�)F�T���_eG�Y�e~�������B�v0W7P��">��#җ����^��a��=\�=��rо��~a����!��5�s֬�ؾ�|��he�$O�� _§ݷ5��	nSτ`���g��F5���P$��*�_�X��f��U۳�Z��6�u��F��*��f#7t��*�pʅp�QEӁ�oi�oI��b2�����^CrS��]�)>N�YWr�9;ThuLpe�;��CV=�%��t�%��7� �5��c�L�?r8���')Da?���ޫ�a?9$��ᛝ��(��}��L�da���t�y�	�D� ֝NBu����43�I!�H+��N�SY<��� =P��k��V���Zo ;Ȉ��̣$n�d�j�b0�!�0f\P�n³���˂@�:�h�X����{����]s�/��#��O���ǘh�z�	�1��"0)Tl&�Q�OX��
�3�@����$,r|���v�����E�,Y�_� �%FQ-S�S\t�XzT2.�?
��Dd�����ŷ
P��#$`Ր;��[������;���t;yL+�˖��%)������������e($�˕�@Ύ�y�>��ʨfw�C�b����C����xP�6} �Ǳ%�'�L���Z���D>3���8��!z(�ҩ@\�_�f+��{
�qZ��Ţ����g������%~�29T���F(5:�ޚ
�ԃ;��[���-0v}�i6LXo=wu],���L�{ �k[�jh���(��ݎ��9K���}eIdQ�����Mv/��)�T�6j��F��ܵ8�u�۾�����8_�羦��" ���2������d�p`wKת1�yn�`]��9m����Th��J�P���$�<P�gCx`@W�Z_�#('t�~'�Μ������?!!��d<��;mɌ�`t��tk4��ǝ/����A�t�I9�ۋZP���� ���D�D?	����i��<oM��W)t�:��֊u3�0 ��3߂EW�� u��ƴ/��a�H�^;4���;� �Q�]���UEi"��3͓��Nh��|J�t0c��"�,-�e��_ �\%w.چ���]�P��h8d�@3a�V]��y:)�����%ގ?5�6��1�F$�/|ȯD��)@&l�J�B �ũ>��c���`�f�U7�h�2d��/��¬�X��]�_��AƬa���W�g�(3��7'Ά;�̏�"�C;1��I��#��Dr�	Y��F��wF��_I��@�uΌ��iR�`���@[oԃ�lY)�iV�BQ��^]d�R��˷�K�Ҥ�m��ļ���(|�=��@y�"R�k�#X�in~K�H�ֲ�N��Kx�e`�֏)O�T{`�(B��ݥT:h� ю�v��#�Yz`Sr��T�2��$ԧ"��	܏��OI�װ�W������U֦	H��ާи�I��7y DÀ8»��y�d�IeR�����ī
s:�L$�٬š*_���r�jwCB���W����O�?/����&~�--��GUO��u!�3_1��M�g�����!q�����g�VfL�L��DcxN���tr�-I=w�Mk6�!{{4��{��ީe����5����2��E�|����9�?;����B�׏m�^�VM�S�Kr��ͺoyY��8.z8a�g2���3S?��5��3gLH��2�{D���񣛑x,J��e;yh"�� �i�F-�GC�a|��L�<���+<�'X���϶��R�(��+�ȓ�Y��B�*�l�T�.~�n�a�}�	:�D����8u����:\o��Ƭ|:����6�$5��jO�F�"QP��bO4v��|��}��tmk���n����$��3���3
��+�i*1��u��cF��z6�Ш��y�`��:9�E�(��7q��]&�l�aJ�#6�@�.�j�\eU#��j;���K������Z�_Ms��{��Cb����SږD�a-q�擆s�Hj������&vgF�����:N�1I8X�Jmǔy������������=,Ԥ��x�OL�P�eQض��*y�h5��	�b��֓5�k��zKdm��'����cIìX�4�X���f;Ķ2f�w�=�s^#��Md�E<2{�g��"���o�ƷZ�A�����>��l���灩MtQ�����5�Ee��n�dV�����.=�^�>�ԭ)���dL7I򗽵�B`�a�>Z�we���Z��dF�w.�%V��Q�G]�̃x���Ҁ8��i�I�u?�i��6���4���}���p2���Z ����Z;������!�4��y8���u8y+q�*�+=_� �c1��sl���̎�'�/s����&U^�ei���]:���aI����Yp_i�����j��Y����k
���̮��oH��:��J!�>�\*_���ZV����R��"��6EwtYU����;�wC���^H��[�}����J)��w��|]m�������������6�X�\��g��է�����,��}�u2��WS*_�a4HgO�Y�c��v�bc��+���f��ig�a����)�p���N{a�DR]��Jǵ�D��m����=�B��qwln_%�o^<����@��ͧ
��ι�72�W���i�{zǬw�v�me4�~�x��%�[�L�Ä���9	��W�~�w�k�T�>h.�[x���H�J{p��n�0����P-���|J�_���1k���l�($�U1W~��:�K'K�D��gp�ݛO���%Q?���g
F=�1�����.+0X���Z���v����&��٧�� !s��,l�W����(�n����v�����v�����8��;�Ą�i�F�/�����E�~����-!���A�O�_�f�$~��DTͳ����R�U�Sأ�v��Wh��'pU+���@�L���^g��Y�W7#ۓ#C�Y/6O)	-���E4��z� �;QϨ��Ҁ�.r#��d�����iH�t�E�.��f�$��`m e�Q�Mr	<���>�D`o�Ȇ4�X�|���Ĉ�?���Ҙg�P�MMo���xܝ�:]IG#��2�Pg�W%��Xa�&=�{IO+�=�B�[g�M烳`ۜc�W����]9��X�u_�4��4�����|�ק�a��x�]셟TY!DqX�ў]�G��:��c��� R�\�A�\���?������`��o���e�E���u�/4%��C�����g/&L��Z^�r�I��b�|P9�%"�N�]vS�ɢzxGBp5]-� �SP�~�g�|��N�Xz)�9Ռ �����ߘz,f�"�6Ѡ�U�e��	������e��h"���|���G��;]d�f,D�#gJ��ܻ�I�sP*<���� �ٝ��VSo��Fa�����5A�yO��%SLf�8�_95g�E�������ｲ?fnѲ�P;����ǧ&n!����7����^���߱�on�J�P1Y�0�ǆ�m���V`S��(b���Wm�i��Ɯ�vC��%MՋ�M%] �� �+���ߙ�7;���`�v�3X��]7�T��y��TA4�@+����qO7�ާ�0��[Z���O<@��gT7�4��Wj�qV=����:��'��X���#�+��#�GB>BSD�gG�[�X�Ř��ȑ�4�U�+v���@�}�I�B���x���l�7<�5����ľ�Q�	�Db���h������f=��8h�L<K���ϊMϟ�-�Z��zG�{�:�R+:u^�<A�*��b,�2��hÒk3ET�"�F�T�/�t��X��.��X#�BQ㆟*��}�ͷP�}�,/�y%X���}�|)��H@F��=���ڕׄ�8����ň�eY?�X�"Cl �T9��y��U���`������BY�����ϗp&�0���i�VG�\��,��ᶇԮ�`]6��R�8"���h�4֙�ޑ_����\�%���.m�A>�3�3	U�qk�K�`�Oe�9��h��)i��9{��K����гh��s��~����[�Ϫ��o��n�<��Í׈����_|G�>O3����~{"uʆ�2ِ������N�(w�W�N��O�N}N���?_q�!�bJ6�Ք�Ԣ��*,Ozj_�P;�PM�����3u���rq�����F��ل@��;?�$��*��sP(��w,���0ʑ5�p^���C�����|�I����NW��(gٿX�� 6!�5淁3q 7����nWlArj��Aw��gl��[]Sn�gM��2.SK��j��jwd�;JK`Y,���~�wp�^!���3��L�5����Ii��� h]��N^�<�y��Ζ���X��_1�B�8b��@��<VE�4_2&|D��:k�����27��9��4me�ٜ?��$@x�d0�����8�T}#ظr��߂zTj�IB�� u:��lR(ex��'�\7mC<.�a��%�Em�R9� �H�	U�w�tV��C���Yb,�}��O��fYNKB�,��Σ�\w`Y��@5��}��|Ɋ�t�����u$D�V��tzd��7�ѕaW:,R���3WQՋ������|�m����}}�߷��$�V�ir�ԝ^@�̔�+z�!'
���,g����E��Cl�6f�l�>����uE>� ~�@�<�hD��DVV�m�n��тQ ��_ͯMl�P������f6��6��t,v���TJa��0��6�cIR	��˽P���
:fP0���7�����k-�j�qQS�p�h�V�Nlg����tkT�Sk��Qw���T�ƟEڝ\�q��T��K\t���Y��#��W:�&�����8ˉ��{>kV4�]���X\��t n^���X�N��xLי�Z��wK��ס曊N�����_�V ���9��pBn���=�H��"��Lџ�g�7W �K�׵aA��<P��4v>R�m;�?�/*_1Wo���]�U�ױ@���h��e�~`w�c4�L�T.Zݎ�W�Rb�c���n~�vw͖,��@G͎UԤp�>5o���cU����4���U�H��x�=��2gI�\H5V��1��%��]�v�n�0��������byتa�����j1�Ub+�j�)����f�	W�����C��kOZ���7�����,Hc����d�Y�S�tl[��0�Dw��A�rA��3=SqR/8T�>�2���P9�Ż�`�W%���=���-i?�V�����P��>C���}i��F�����.�+����;��($��q�G�~�_�B�p�$PԲ���_�e�%0F55/���d��T�e�H1�6][�#lfo��+�?(�
%�"@��S���劀P���`��I��V��p) }��&lȝ1�s�F4�'|MI�.9�($���{*�#{�N0�]�A��X��ѡ�����ί��Јe���3�X\��&�D�!;N��ΐq�,��檦�]�F������_/���[�X�az��}R'�&ȷ�r+��\��y~�j��Co��q���^��y�p\c�1��J�����z��0ɹƢ�����kt�7�G3]�J;j�w�W/����"��J�Jj�i.������t��I:�f�A�6���ww�Vڠ����]�;�L�,~�	�v5����1E��.��.A�,��{�/�������;�<�OX�&��?�K�
AWo�m�~��e�v�su<��0TR��� zCr�{<,��$����s�ٗ�K���=A���;r��ζ5��v�y�j-|=��\���.x:�;��@�i [�Nj3�	�( ԯUD��i����g����x#�"�S��G���9�ݑ������;��xfǾ�[>/�bvt젥�L�����#��,e(�	�U�m�P��B�b��y����L�ael�I�z�/R"�o�['��`0�ϭ$�����"SH{�q�hUno~���G^Gxh��v�PR�HL@_�� O��8p�+����ހ�Nm@�|���/��������-�k�>�xx����,�C^�c�!�I�,)0�:�����}�gHqI
k�#_Y�%(���$�%d�����F}t�WI�%��v�Y�9=կ==;�<���6j���\�����( ��`bZ�|9J�%V������q�ke�}̲5֟5w>�t����������Q�� �|3p���%�q���c�����q��O4 )w*���/�G磨(�I]�� ɠ%���Ʋ��	�ج�#`�8O���p��nM�3��K�U���� �!��(����j��ј9�?���P�4{ե����Tk�fO��#�I�ζV���I�(�ɫ�J E[����k ,�#!����s[��nP��UbZr���q�j-܉�����lH�p�;tkߠ��IC���c�2����@�$b��"����yA
�e�8hտUx�a�:<s� |F팎j���������L�2Z�R�i��q`���̙���P�Z���l�O�5Q@���H�`����"J����*/ene���Ŏ�r�P&�<3�0I�fy)��m���u;��i.���eD��	/N�����'�A��ꌨH(���"֢�}���YWRf�VɌC��qs�B�q�tsڊ���F���_օ��zʽ�9q:b$�� [e7&��~�Wvk�i��2��@�J��߷�Yp���p���ȠJi߂X�%G��ۜ5@�;�▇����=��v4�(�ؒ����]����t�A.8�E�F���������c��LU�bp�x�t#���xB��W�W#��u�����ē���
��vmX4��H�B+� v�������V�,R�����`5P~�T��zK�LQ�ǖ?*����>+�ii�#׉"�#��+��`�Mn��E+�v���/�q['�t:���i\T��&=5�Hدf��jd��#�6���x��?�'='��"�ϨN�/�y��K4�'s���|I��&�a�@�*`n�]L��i${A��
��T��uI�[��*�a��=,�Vgԍ%���1"̏|mΜ���~��m��D�;|�0�����q���0�<A��#1Pa�}��^H��Jҽ�K9���Ֆ��^�N?Iy3t��D-�TqDx�d���K��F@>U0D.~"g�<0aL�6,�.�Z�?�����55�i5`>*lwʅtv+��Fȇ'H�57O��Q���	�)�`E6ZzZ}8�X0��޻t�B�yB��|C^X���%��!�_��(\��G�p�xy��]�^�T���,�z�VQyf�Ӳ��ʡ�Y.���V6x�'JTEC��/,q`v�H��-݀O��Հ�T�7�Ǚ���3��b2B��u)��T��Ȗ��Q�N��������3R�h [כ�#}�!��8yS	i���"��8�\-��M-Ɣ4�1�o �ԅGS�&p�ȇ�u�_{p:[�B�IBu
�
�ڢ��@!B�'�"��yzk?Ƴ���_q��-��R �(�{�*l��󱘔Ώ��Y(���,xf7&'rzi�M���LճVc�����:q)�[-2�����v��k}@=��v�b�?��pf����IpYw�)����b�F��\��WA�ԧP���u&�#u�6�u:ӎ��,+��uc�ЫW�>�u@�B؋�����k��\�������j
�?@��=/Ǩ͢i��s���m���� ��F��8h���	{*yv�ݱ���d�Lk�ao;#�L�&�A5����Os`���'EYEzO|�����qA���ȇ�o�B~{�ȇ�iTm��K��C����p�����(|U�ZoHv����WI\�>�2^|�Iy��Ԙ�5le��ٯ���M��D�.U�?e}�8�6³����ܭ>��L�^MN�����U/~s����rQ�;~��qG_%*���c�}R��|�C��ߦ��V~S$�.�\��l���]�ݛ����Tit���l[h_��>ң$��FN���/&K�l˃y`�|C����([�h��.<Z���Q�FLu���fG����Q���@ �r�o�dw;�œ�+G�E����woZ�I�]��k�_R�X9����(�܉�,��� �G拏^>\Yq�Nrk��}�[P!.��3z]ή����f�J�Y��<�i��ݙ��8������D����w!��"�9�	菩�R�[��G��?�vQ�MĵX����մ����oz��ׇԔ�,I��2ŋ_��ߟ�[Cĭ.�V��jO�<q�4�ۛ��m���Z�T�4@潮 9r/{zg,d^a4���~���6��B��J���43��4Ka5��͐R�]�"D�s�mcrI�~�+Mh�6i�0r��a�D*�D?M�����$��tK�+{!������Nl�����*�Ū#z�@�K�Xcw�n���:����0Ʌ� ��p�� ?�0	 ,-��p@a�y\�S����eg�P� >�uŧ�|�l��l�2�3I��1<�$�9�aT�DBcظ�4@
_���9�wЬe�Q�c�q�,я��x��(�&���J&�צ�A�e��4uc4����p���'�W�#l|�Y�*(��E�/l�=��.s�b,�����c�>���)<r�qW������s���aF���/@Iqr8�Ϣ������Z��Z�4Nў����C߭�@)�<Tgr�d��V��QQ[K�~�1��`�b({�ռ�g*\��I��w,~����6��#�U��t��O:]Rh�i�@�<_�X��PQD|�E�Z|p�h�����w��!�Bq���>�|�1եfa55viz�s/�磯C��jv����.��{�y8`p�3��&�h���S�ل�<���֛G�i����p�G$Q��[�4���zE�j�"L�#V:tc&��rF�qqʁ��i�Z#������vbOL���:r%��UZ����p&�ã≡�2�
�x2U�J.g����c���Q)Oa#�׬[��>��3���e�I%�����'~����]]��P|*1T�%�8,AgbM��Jl}�j��'��J!�H�
�E��֮��p�xf�Taf��v5.@
�늌�"�>h�T�c9�!N��#��JRY2KK�#Y+�ۑ���K��ՠ
�c���
h��a
L�}�}��s�E���Hٗr0<F����hYM�M��.�PO�4�����4b�*�R��������TZH���{��V����� P4F�뀭��</!v�|�*JD��0�P4���(�Hw���4�z��E�H�F�����!%t�(��>yc��Y{QR`M�˄�1�҈{1�E޾ۡ����M�*yZ��ީ�1}+dZ-j��m��A�!溦y^��|8��� �p�6�?�H#�R?��y�
o�Y���>+%�_ E`�&��N%SD����dMmM+F�o*t$�-L��O�T��|9H̓Oԕ*�D������Z)!`G6ڃ)�����=��um���rhQ	�v2�;}�k�AhaߏW���ǒ}#f�9� ��mY12[ �|4ލ6#u���ZU��6��>S^Φ�uwP��AA?!4�l@�|���ؤ�ƞv;!%��j]�v�ڽ�����vV�jl�*C�4�u��1I��33K�h�Bt���I�z�~Mr��cwi��˲�0IG�����Ќ=)/�z(2��/��Z�����y��t�[wX�y���PrC����Y�1�6�,ȥ�e���h��=:�����Ӧҋ�H�y��zs���̔D���1���7�5I������a�5��%UM0���yR�|�8D�v�������N�3��w���)�����O�L������4HT>�b�/j6]F�����O?h�D��4�I{1lH������q��	��N#ų�cϖ��ߚ�(t�qF�4_��b���Q�b�,���
ѣz���Ua�/�y��	�غC�KoD�f�T~,�6Uu�,Q�2/i%?`����4����t<���/��� �hq���{]�%`eV�)5/�Y�49�B��u�-޽��k�oG�K�#�lk�����2���Dlȗ�l��}�ґ�|���
���Ս�+�DM��\/|�]U��鞰1M�h�x�LG\z�:n�\���(�;�o��Nf������Q�?��=�7�p�GM�����*��S�^��:%�-�M7K`���b
I`	� � D��mo\��n�4QL���:�2!��4�lJ��� $6�_����0�ab�؃4@%���TPcj�����$	�]�G -�G���Zo0L��"OM�[T�U�At���g�Sh�Ȥ�ny�<ǡ�� �˖Ĭ$��	�,��w7ѱR���C2I)�oN���" ���-�le	p�J�O�ր^�^����_�L�� .a���Nƽ�4�v|�|��,��F�C�D�h}�B���č{�C��D���N����%�Í�Ц�
��&�cgBnٷLtK�F�F\8�����m�-�xm��P�:�X�We�=.���+Rb?����w�ۭ�ܓ�y�7p�÷�0�QRj&T܄��`�����.Lڰ��Y/͏c�,��ye��B�F:��.e��
B{[e
�8�=dji�d��2�()��&�j�ە���(��%'�·n�~f�w<čJ	�/�����]�h��� �R?��$�+VS $	L3Oq�����j�*��g�"r�:ͳWp��"O��ݓI �Y3_�L$j�V�-�c5�vUV�����:����z�c�9����
o���V��J�Cc{y�q�٥#�F��	����݌�s�^F�
 2m�Z"gD�m˼�LH��e���9�{/��H�Q�&�$G4���q�|���`��-��Ub��D�h>e����a��"�[�wI�����F1ћ�����>_t$((�x��l,�=|�o��T�FA8�m���W�����)D�q6{m_p�4�i�l|}]Rr�� �k�������6g]��$�I�������Ѭ��[�p�C��]~��(��sC�sāQh�=��G�K.�h�������Z_c?l���[�mzZ��H�)�IE!L�C.��V-�ej�o�PU��̉54�Ep�f��0Q���m�rm���A|--�*�l��5����(�h��J��5#���F���6�r8�z S�39��$p}�FT��JgAِ'B$��N���gG5�P:�(��q��,�!h3�Z�f�[��/����~��q��>��E����vGf���a�2$��<�D��v/h#����͹���~���#y���tΜk�S��#�wи�@�A�b�g�T��y0.��Q?�,��Xa!/j���]kd�۴/�^F�!��-�G�{�Fx�-��;�H���*�9ӑt�� ������=��U�CbЩ�'�u��&��i[eG:j��Н��W�	4�x1��. R���*Eb�F��W�ұ�0�4���f���,���iP��7;��f����ZϽ!^W&�0$s�q�ޏ�88hO��!S1z��:��{aC$�����1zT�c�(o�I�� 9�V�+ݢ7w���.�a����戨7[X�|�FK͟�^���Woy
�����n�d����&��}S�$ٞ�ߑ��=J����9���:����k*Y*�w�}z%e��L�&��_b���������Wn�'��B�s��@� ��1d���yڔƈ�&�Y�5"0�Ӣ��Br5L���嵦��^�p#m��	p|G��B��Eá �
�렵�=f%���8�ކ�N�6�����n(�_�B�߶k�D�5�BD� ��̫���S��҄3�x�=�7�7x&��~;���0��1�ѫ�Ӳ�@��~i'���6�m��a��������˙��rDP���]@m�����&�d���y��}/T~lǎĭ>�TE�����uz-fy��7��i�yT[I��+j]��Y� �p����P*ֱ���چ�{U3��i�/m|�!XRr"M����@$�^ �������:2^���%�j�v���ju�h�8(lf��X��)}jI����gF(@���l� �R� ��#X|��b�eՠ�	
��S�VF�^t�m`3��p��j�b���$
�`��׎.���9Wy�!RRz���Vk{U�jr���O��3i�VS��3�,.}n�4��E
�	�uPW@=S��g��q�S�r_���y"�+9�X�����l�*���4m�D�#g��>	�,���pKnU�%]�x��#򕟦�_gVE�n�RB�&v�UB�����y`����۬A�� +��Õ%�v΢Wٰ�曒��?K��\-�=��$���/j�w	2�rM�������O����!�E���-�ą�� �
��u�Iq�dZߟ��_B�}�����P�L3�d� ���0��X�#�[sR7M>Z���!��a �5�}\"5�!���Ԃ�\��;a�b��i7G���n&��~�Xy�'�Ь
�}��Vab�]�+��0�)g�Mھ�x�]ݔ8�.JS���S����ѻ�3�Kg#��CC�a}�_���	��G�UkR)	,���X]������(��� �H72��M�^R���n+��@d����0������YT�7+~ElkǸ���>�9ĉvڏ:�M��iz�(�)��v������PC�o�� v�g���3�
�y�ZګI��x�<����Qq9�CH&��ޥ�_u�j�2`�!N,�]_.y�[E���~#:hi˚^��ۢ�2� G��D�h洐����Ue�O����ܨ,C�i������͸�z�$�Ti�ZX��9u��Vs,���a��AQᡍ���u_����q�
���''(fcV_��L�X��;Y?�Iv��f���Zx'�i�l�{��܆�d��A�{#%��t���\ji'鯓�x\�*��x���Ƨ_q� �0Xmq�1�_���S�e\�x
��#�6�������L6)/�WA��~����jT�Q�[�1����
��sR�E��=���e���Y7-�gQ�g��V��Z�X8t4^�n����Y��G�������YX�׶���H��А�R��kpv�|B�ˑC�]� ��8�95���z��@&���'E�z�ݽZ���kBh5��e-�T ͟6Ӻ%��-�=.11)ќ�>��A�xLp�h# ��07�[�1�ɪWiZ������g�V�d���/z�'z�Jb���s��[�bxʈ�Qc ��?�i�iIޖ�������[���f,�#�i�+˂͊v�����DO�
ˍ7�l�>�_��X��+d2�C܁�iGo`!�5�zqT� �~jb�O�g³+������G�Ȯ]{�Ofxx�?�2!�������v"�D�Vˎ���d?
�6?�Z�[׳�@�7��ehپ�����������xt���"��`���uQ[�:o���`Ͻ���W�c�����L˿�|�-�}r~}��D�]�Pjy^u�~�Fe� ��M{� ⪝����p�*��a �w����Z[��5y�ᄱ?
���5[4A׺q1����lnAB�CƁC��1�aK�������x��?�bO�����ޱr)׳�{�ߕ�l�.5.��Ȑo����j2hؑ�r�pNG��G�Uq*��6���-���%L�3lH0��`������������W�d�	�CLy��b&���n$�/\�/N	�>w���V+�Vr�X9�S�<�p�jL����^�*�%�2f}7#�"����W2b�1���͗Ƃ�8hp&�iP:Y�>x��f<�Ph ��y���52w%�u?�hX�@�?�e��tr�p[N��l��K�3�����xu�d�pLD
\���Q��%=­�Ĵ)l�L�h��N&�p���bjc�&�A'�@�ũ<���ם_�`x�����I~Օ>��L�Y��d;c>
��n҇��� �E�����5zz.�27GU�o)��ڲ�Fܲ
/i��*��]�����7%2	��6��O��c�92A+A����8�Cf,^��؈��[���wds�I��bwS��x��mC��oTx�6`&jU��i[f��u����A)�*����t�V��I�\a���E���S[��L<rʩ�k����oPG����+B�Z��2Y�>~�͡�C�Z��Cq.w���u�j�ۃ�s��u"\�UK̠5�J��>�����G"A�L�����MW�^�.�橭iC �}�����婿�fLu{`��+�\P҈.�)��%C�$���Z{1J�h���e��u����A��@�FL�3l͠�
X@V�>vr�����,[� ��2�r�0�rM[�H[:�S�����=b�������PCޖ��O�;�!�-���+zi<ZQG��E��^�6�fg�ǝ�y؞#����=��9�dp���؝n������S5�2O,\T������p{7f����\⒩�'��$�@R�@2d�Pv���-��b�9��VizX2q`~��6�#|�O���h:99F�Ґ�G'��p[�S�X���Ԅ �C�yB��,��5^L�><_�:��

$��akIן4 �tև9�J��T��ez��XN�X��ir,+���mp��f$���:T"����`eP jqJ�2iN�Ďe~��_A��XM��pM�^MO0WI��=���k�SK��0������Ő[����ɺӊ�蘢.G� ��TX��v���H_�k�¹B;	�`Uh����Z���
�<���V�]W*�N��i�1Ss�E��4^Cs6�'��8�y����Gs�V��(�!���6��*� ��������o;��ռu�(,�w�-3�g)�SͲ���s��NnS[��_��O�H�����jKĆn�9�_�T[k�:l�7_h ҵ��nB�x�^h��,�0�@(�La�)z+���G��?^�|P�K�[y����,3lTh��$P�m�V-��ޢ�:-]��a��kҝh�<_��3BjIv����>£��{O�)�<�56�����w�D+�L�4eܜ��"�L`���f��N�{��:hBcS��/~� ��"x�}�T��w��^���&�0�!,�b����	~���[��'s��=|ҧt�)�c�oG tT��2r���>�i?�Rn�/h<���	�,֓��D�{������A�c���Ek�6hC���3K���c{e����ϬFG+O��ô���'���)�A�Ⱥa5
{���H�0ˊ�~���RS��n#n"�Bz
�h��
�u�_�Nٞ���3ZB~f��U��1��V�8l��o>��!:��!О��0��YA��qvVFlԕ��ۀg����V���O�-��.����R|�E�`��8��Mj���+#���6i%�<W.ƷP(������>F�vf����K�������vf���M��g��»/�����}���N��$v�������ǘ���tN��{��p'Ug��m6/G����I/������Z/ia��l4È<T���g��Q����o�:v7 b�J��O£{�;A�@\����6)���@TQb�Ț~���k����}�}��u\電���X�Q�] �Oe���� ��g	1���h ���LM�V��a�P٤��$L��l���osɚ��FF97������Nb���Z�r�Q�{Z�2�SN�;ʖM ���<�jު�o��2��L�6�r�2t-�^:T�'/��	s��#�/W�� |�6�I���4��vB�D٢�5�� �wV/�/��@��;g]yB>�͍�E��
Q�E�Z$��jVc�1^?�GD�1o�	�p������bj{�+Y�p
u�ca�N�:���ւ����R���U�P^�ހx1y�0����Y6;�_�~�`���9�p�i�왡���,�"#���*2�a�K��)r��I���'�+n ���"5��g�P����>iQ|2I.+�_�ھun�ЫV �;��'Y��λ�N��5X����>�[з�L��y������>)w� ��ul��\���]J|X_���F��ĚGx��HK�]���*w�u����.Lcj3��IYZa�c͏�a��M���Z@&?aH�1!�� ��`y�I��X�����rNZo*�g�+�g�����z~���e/�Lj��t:o:�x�(U��h��`�~J�F�4m�n+��懋����RO�o�:)�D�߹��Us50�r�����e�L.�M;If�g���/Q�۾�JU�8|˾5%���2����t��V=�w����t�>]���z��E��Y�P�D�3c�*rm*�'w@��hz笓���Rn��PA��sM�)�A__�g»t�ͨo&n}z�M��|�-�	���1-G����)U�م�����see��,���z<Ys�*�L��aR��AX�!�j�	k��b%�g���u��`s��0�H�+��|�Cu��X��O[�)@u��Ҟ������%{����1�7�g[Ɇ����k�1�{���F�5��H28�;`�@j~F��R�!��&=�Y^�.��$Y����M�m�b�����o�{U'��� E�+\�`��o$,����J<_�����l�(��V�P�K|�&v��z�6��tA:�[�z}6_yr�!C�x@4�*��o�j.�n�8J�0A�{T�y�J���BZ�'1����
o,`[��ԫ�-U�K�SQhC;)]�h���	{��:��'�l�Ρաk���1��_��޶�ǔ4ӑ(�s&�g\x�dV�	m ���S)Ye��RD�M����;�N�4���.|���AQeLO�)�2��PV��Ҵ�W��6����e�Isf\P.ð�k{�$!5U+�i�m���]R����x ��oHwL'�S	!1\wxe�k�?�� ��� 0��%.C�j"x���=�k�����C5�c̅�b�k��9Y:�&<�����VՂ&ys�Vg���2@�%NYѶ��YFd�L`i��]��	u��x���.s
��V�8*�L�aatz�e��"�:��-�i���U!זs'D��4�zW�ۚ�������3A��2�Z��k�vό�����ѥo/��6�x��0����y>��p*��pl;l��[�� )���J�?��E����QS���R�p-�5qnk5S���aF�������0�.�+pO��s��V�]�f_���Wlg�A����[�'~ռk��a��h��h�LL��� �ag��Y;� k����w����h��pW=����`#z?�:�xj��2��K����{^��t���V���� �	y5U{�� �74��2;9�8�����s���j�k%敉���Z$�0�T
�c2���0䒧�,�7�ף�Ey�k�l�����W��B��h"��E-���@-7����+�$~�i��OK�yC[�?����U�	� � <*�nA&:����W|�l/4'v֛�"_���?*����*2)E��B*�+��adu[[�7왋��j����⻨��L��"�4�/�~������&��F�R�����	y��Yw�GG��B����G����W3_e�S8Ka�R�󻩋�P�y<s��z�|9n��"�еjy7���k�R,%7�%D�b���mf?�7�#���>��ӽv�β��9�	��EZFҡ�E�C�r��%�Co��U��_��xZ iah%�/BǘG^��L�&�ˠ+"�󃯏yZ#t�I��EE���`���U)A-(�!�L*����oK�&ԭ�i�vJz��o#ǆ/��'�7�?}ġ��o���!�*Z�\��k`�W6�3���'Cʛ�VW4R��pV���Ž58�������T�r����A����ڵ��<�������6�g���o]J�����fơY*�݁�إ�G].�P:?���_�Iz��@W�v*L��Z�g�#r���D7�C�wm��A��Xog0��|W�@����C�W��bb��71w�]���d���FX7�B$",T)��{����P&�����>�y�!_o�j/��M�u�W|q�JA�d��;�� ���bYG�?Z!!tP�5mj�B�p&{'�/\P�@��gu|��Z17B�UI	<��}��,�D so���P]tЎdY!__ ��W��_[�n�^r�Mr�t��uV=�l�`5����*��|��J����u��=�W��}Wx-�l*8����(d<w�̨J�!�$��>��:=/U��`=��l�)�;���3�Bb�+^���D��o�d���E�3*i-H�H�{�_��2�Y,>^g�ɔ�F���^�4�L	T��I���2�8�O2a��kQT��N;�Bq?��Tl���S�3�V�_Ax��-�	)m�&=
P�c�lm>��dɹ����ݵP$Y��<_	B������\��,m���`���q]#�}�0��UU0�Tj����fb��y�Ή�zw�{�z���zB�AB��J2���E�(�s_�eɗqp���\%�k�$bʮŃ<&X%W�\w�2Z~�t)W�(�c���,X����x*Hۀ"UQ�p���c�sI�8�~�qN�F�35��l�i�Y�/>rVf/����.���,�!���i��'�YGh5�$,2�F��;ƶL��
�($��*&�|�	����;,�n��� � �6��ߤ��,Fv2n�ت��N\�x9$����v��g�|�=q���� pʗ�d��%�}�b����UP�mk�LYN���:�Ժ�A"Uw�:����<<���x�z�r�O�*���cW�HH�~!�1��p�ߛ��8���= �����H.��͍Ló�L_�0AqNU����C�E��8���%���ƶM׎��fڹ�i�(���Q��E� "�׸�)���h�%��KJr�m�ڀ9�ٱDf���(���H�f��"ݓ�?���9��璦���$׷Z�Rl2��O�O�Oj�;�ѵ�� /�	%`+���l]Z`�D�-Z���_�ʡK�S���c�F���a&(c�:b��)z9Ԣ�>uS��AWFiVz0���?kḪێ6|٫������b�����ܻk.!�߶6Q��+*�"D�y��x�V���y������ॄ�%��C�=	1E�܌���Q�P���cO��b(�f�)��d�*/��X��4u�|�\�2��(��d[��4$� L%2S�!c�����|�j\���pp���*� ����Xk�rV����׶��*�u��Ԓ�� =�z�2����J�e���^x��u�oYa��/j:v�"}-[��ɢ�z/�
�ٻ�5ء6�(���+�zD�Ӣ�`���c���7g�g�h�b%'�6���H��<����8I�	I�P�cAϻ	��7��Ot�tcc��Vy���ܓ�x�{0�N��v�o��
坝�LS�`���we�^�i���"N�����>)�~Y����9�s˝�7E�q�X�x�3ƿ�e�&.i�rj��-�:���K8�
�"�Q��ô��#��K�]�F�3����in�$�%"c*Im�w�;�>:�o��f��ut�BzE�����	x�+�0�6�Yæ�Qډ��.v�i���֒�����
�1Ve�q�m�&d.��K&�?�K�6�4�s`w�1
�"�=g��z��z��z���[���7�"�G�}��;{��Y���/�?!�%�R���E_"fY<�c�PF���n��3�̔�̶j��&�vg�zq7��d�{��P.��E-�iy$,}-����7M�DV��R���+o߄X{����^��d��s��/�km�r8!�N�i�J���e��,�) -逶A�ΓP�&�u�<���R0a4dV))�S՟��u�y�SQ8a�Ґ��������fX������u�K �6v���q[h0u�;�6�Z�*!�KMd
"�Y֤��Q0�QX�n��kO��.�I��i����u�����}�@ic�OH��������j���8��y���N���D�����P���0}��v�����3y����X��6p-�)!��h��n��`cr�0����n{3���4W�lX�%����}�ͪ��(�y�%��3n�5�j`�Z�c�-��/���G���7Z�{V�hD���W�T�0�a3�o��ӯw�9��n9~�ׄ�J%5dE�?.�F)U���T��,i�;��6�k���Y�|hV*N��4I֋Aa$(��`���2�3h"��G��u}�.q٦xJa!�>��Hpt�ʲ�ўF/�S���@�4}��+��3���m���i/�*���a��M���7va�+�h������)�aj�j�ְ	ɇ�0�K�tD���K����oO����mWKCv��6����$
��.����2�5.�]�Y��yչ|�r( ������Yo���6�f��D�J���/���Iq�t��?D�����Io�}荮��UH +0X�@v�㽴����j�~�0Qp)Y�a�U���	X�@�sȫ�-B��̨ҝ	k�M�KUۉ/���&�ș
�UT*�s��:I ��h�,w�%�)����neK/��3{�G�n�C�}yV��*�Ծ���F��Þ���\������6,����v��u��koxa�����Y��0�������h{ŵQ-��߇��v���]����vm�:�䧁�5�&��iP�KC�G���f����0�dД�p�k�+�c�͒#�j�W���s����Uu0~� JiT)�{9��O-�v\Zܑ���L��h�@ɠd�u��l�5��s��_���ߺ>�=�����sש�����Zd΀��h�����Mh9��E,�$P/��r�>c"����yJ��M4~E�0��2��eY+v�.Ц�w/P���s�޹ů:H��`j}%����'$�S������� Y����A2��_�R�L5�4L��;q(^y�)b�,����1=��F�&�	�4L3��ܚ�=��qcح݄��'f	�V�/��־��Q\�YN���:NP��̫[z�כ&���5�V���B��(�
�O�Ò*�RnE�o����J�C���As�O��a��M÷���x���H��Q�qK��tU����M~�Pk�}U�*�;?���!�h�^�ee��-�חX��AV���y�8���'M����~�!X]X��=nL���E#����'n�
B��0Pu��~঩��:FMWf�lv����]� ' ן���);gi��١�=z�Fh�2�b��MmPKC�q��p�\�~ ���q��Y,z�����]~�%M`]�q_\���`��6��Մ:�p��!��B~܋b��,�Ǎ����~L����Qvc%f�Qo�,�8�5f�i8��mW�6*I5T�<�g��!(?N�`���L���(��v��r/{#ZȝUF��}�R�6fR�φa���.hVd�]'u�cC���9Vܯ���J�w�5C[:��u��WU�M��1���LN p���4��\�ݩ]��M���.
��~�ϔ�#��E�ձ�M��N��Տ�4k�	�T��E�|j�2{�����=�?�.��xv�62_]������3���p���V3l38k�;��8���F������ /Ӎy�^���$M���c�'$c�u���K/!���_4kvP&�j�:���7�`�1�u� ���j_��t<T��e���6��@mQ43_d�wt$�o_Y�p�ǵ�����j�<Q�G1�]���T� �	#�5�Q�1��.= �dv�M�����2;;n�Y�`J<TQQKxSb�����J�gl��3
~SnK��↬(�B�Lׁ�ˊ{nV,�6�|TzF�}��g����am<&42z·%�_v�N��Dm9��5r0��Ҽ������^d��/x6"j��Iù��Qg���ͭB~mDa�H2�8�>,u�-\l�h�(&؞	~��S�"��3O�nq�U+�>5�t���r&lRK����.�j-_k�	�A!IHW�W��EQ�������5�5}����K�󣰕�*��C���4��3��������7h�T����{˳N�gQ)�:3��M��
oQwZ,�f �_��H{�ADy �i�Vƴ́��r��2�)����ū�ݪB"���P�ܫ<B�������Ed�I*�W�;9;��9`FkUF�����Vp��-��η���6E|�&�<�Z�j��$��C����K�,�y'�L6C�
�A�z�)����Ծ�䦝�=3�<s�~<,��2��;NX҉�����j��`�S�:�7`���Qb�DU}t�@AIz������4��?����lL�F��@O0�)��w ��|jBu;M�쐪.�rP)6��]�V˵�64$��i�Q��m�MG��D�F��3�P(��JD�'���g��jV%Hl�"M�JC)W�ù����&�+G�X���۬�X��S����	O�$
���Z��a��}ST�x��*�"\�=�W0���-��pn�4����/�3;}��j6V��1����6�Ma7�KUTz!�ѣZ�f�$���J��.�Wڮ0�~Z����\SS��/������#?QIݴ:�xS0��C�N��>�^QQ�0x~���u��W�g3 ���cY���H�A��vɆ��g��Ud"0b�����毵�ӳ�9�(��$W��x0���#�cЕ��;���U��f>�]i�-��C[�j%�l«6-�~�,9�-��ؼK�\8"�NzеjG_}�q��[a�Kh�F��r1�TK����A���[PM�@���U�;�M�ɐǮ:��M���A&+�����$v�p2 �~��#�%|���\��`�N�n�~�!tc6�+ޔ�.*Q;�uȓ��[�A�5�?���1[�F�sp�t�|c:#�m�kZ@�o�,�/�q�i��g���=����(��:K�cvO=�$6�A�|9���ݢy=h~%�s�c�B蝅��V�Zo����A��18�lx�ݘ-�Q��P}�X�PUw�س�skt�4頩�c����~=��?���n�U쉧�������a�r�K���q8�d�R�2����d_f�)�b*��8)f��{K�N� �6������}�>�kޟ�����<��q+Q�׾�&����_5u��/��9?'��'�������-��6N�����-��E由a�xױ&X�&s��:�7�� �INU0Qʁ�;�^�>.���H;*)�p:V3j�P~ol�
��ض�i��\q��������<旄�l�B�[�B��5�.0���3v�-<���hko���T!E��yp��+f���-xF�����t[�ap�_���CiWVZTU^���i��B�u@ASNw���(H��)D4�w.f����!�?�L�x��n�MRSDa�4������X��)s������&��\L��WV�*=���y�f3��˙.����:E\jt׳_�p�X�8��ܓ�)������������sh�G�M���.�V�sY�Up�n��u��"/�����$��f�]�l �l?$8��|L��Iu���{3Z�6��t����;_���HA&ޟ��0I���3��}.�>nx�#��^{^lG��w*�	H��Q����	���x!�ʕ�X�)rB� /�$�Q��ռ^ª���9d�IHţl[|6��-���RL�n�v����W&�}6�}i�Ǜ�����[aS	s��p����n"$���SP>��A��"o]��b_;�Գ$f�_6>U���W,^�Z7Q���n�
�x�Xe�\���?i��
�����/D2vk��i�-y��kǓ��{�v��b�P������d{p���m�Z������V���U^���y'2��Y���z�z� ?W(���ygT��m�e@E�Lx>��&#ȃ�|�f/s�y?G�ǽ�z;�w���#��X^x�`'��5;�<�t���������j/��mm�x�4R~k����c�۫��f�+�H��Hk��Jf�I�J�ŏb.Tۉ"4�b�B���\=��`[x�G�����ѻ�/���H�wǦ}����o�6~<�TAƭ��3q}5����M��w�$�������a5�*�Qc�ҁ|`�LQ��o���Ġv�a=�/��\kã��z��葥�@�bz �Lx
~�16���Rb��h,.���UĲ():�R����FJ�����U#��8��*}�O���LZZǚ��&Qim�y�˕�6�"��f�]�H����
��U�w�ƣm��Կk��Y�|�y��u��tNkc��_���T�D4қ�H7Xc��zP��߻֪T[goN��pq�!i:�d����e����[�!]2����ޓ�6kv�o|@�h@�T�"��x&��CkQ�D�
��_m�{u�O��,Bɮ	y�	$p.A}?}2�u.�7��t�l���G��4�(�#<ݣ�/��d�;���ȴr��f�<}�^.��� G�_3�Oj2�v�M�����$@U����VEV�
U^�&�۶�Ms�D�HM��Ր�}�}��xY�j�ܹ�i);_�����Pi�^Agk_�)��J�O������jl�K^�<,*�\�E���T����a}�u���n9���|D��-���` �G�#fHomf1��)(x$N�c�$���Y�d2 Ivd�ȿ��)�$�q~A�-�{�i��i�þBa�q��-��\��'����L�Flz�'{�]p��|�����U�� �hK�ÞQ���%�lp�����+,u�do�L�=J�h���Ka!���X�T�S��O���	�F� �V�oJ���E(x
��jI�:���qL�<O��:��E�#]�J�4ۮEJ�Y��<�:]]di�����o�@$�"�jW�0+��$��	�Y`X�?���N�o\� ����$�����!��4	��Z�
\�L_KT�#���r�Sm�uF�a�F��	!�� #��a��Ua��q1g]Kt\3�X�A^�7�̧A��\�ߋX���X�C�՛.�.��t(e����b4�,��mȍ.������~�u�7+c,��r����_ho�]��FE1Vs.p^��i@����frmX��`�}��nQq1��D������J�ReߊS�l<D28y�ލ�����c��������7jƁ�W=^.t�ñ"y� �׾������d�{����~r���E3TQ+ �I�.ȮǤ�&� �_~2��J�M(���X�(˕�!l�Ɣ��Eٛ%%\�W���_�
>�J?���Kk�D�Jsg!������.�� ��k��p�c���a�7��3r~�6��9���:?鱤�KZ��ʣ����غ����t�p ��p��Nd�$�2�ed]
	��a �H!�,B,���R� �%sx�0��pl,��k\�Y��I��h����T�)�91y��u0m���e��RZ���%��oQ-}[+�P � h����gCO&�Eeܬ��(2Κ*�Ы�v37ڻi~�q%�a�R;��g�،�~M'=�j� v�7%��t(�B ���Y�>���MS�LF�G�@��ݐw [�ѱ��$X��T<�UJ�]ũ��_r�Ǣx��ϝ��d�}�JY�����i��A�A��L2Y���Acj�Ne����m��iЅ��\/$�%Q�y��S������qۓ�L�<}{����О2������Qx����>h����w)c,����ٿ\`�}FVF���ƨG�N��Zv7o�&셴h>�MLV��܉��<g��a�I�i���|@f[����O��p��K��#��C;����=����Y��~4�cQ��M~�q��M_����^4��-oT�G��bg�W�C��&I�+��I&�L����@�s)��nȠ�^c$SUE�O<����}B�ؑ9Z*���ɯ�?�Q�C[�Z�Y�%E8�uH�C$�� G�%2d��*�d%��S[�mѿ!��6�����즹���M�&d��Į
���DʓéA��<�J���`��׾]���~F7_v[�U(i���p��D*��h������1FխZ�[�ʝ�}�%i�=9��]��S3�W��[/*��ߏo��be4H����M�	f�[�h~Ȭ#�>�/�_�0��"�2H#�"�j����*��Z����0H��6�(v�ÔF��#�4E��7:�(�ET��L���*��r�A�79IY���^$X��ulh����g�V(�)o��r�v_���d��ӓ�A�@���߶��R37����f���l�0��!j6����t}W+ְ^�J����.�R�~|C�|�~�;v�z��~y�ʪ��I^
'S�5M��x�,m"�/���κ�'�# B!�08��{�,<��ͅ�޴����'9�k��B��?U������ft$��%�d����ξ�Ԁ)P�� ����HKͬ n���`^	}U�Q�R�݃~�k,o��.����ue=[Y�qb, A�x@�e�V�w�P��9/�!���h�b����u<�BM�!����5C�?,9�/���f{�e��[������B�zuŐR;�ӬE1#�,t>[a~� ���k���;y<��qN+=�R�zo�Ң$�^xc\5�ǵR��*�!k���x�'"d̸��x�_�?@mc#`����m�n^4��W����%�`P/M��m@��J������6�}�M٦J����@�-�"�q��7���BW�ě���vy�0��"��HP�2���^K����/�c��}�b��*ռ1;f�!�|.�|��2��-`9����^�K�Q~�Q
a$8����pv���A�����5�
�Yq�����&ƈ������A���𧙰n�fB�}��o�6�d�A@C�jBhi�[��L�k��i��������f4z���=���g�BrH�&�A2&2�&jw��y�xs��Pk&�F�$�D�?��J��!醬Z��g��B�5}B5e���qI�ok��Bn���+S���q7�`Zh=�D�C�R�Ƚ��w(�Q�Mj���1~H�B'm�ۿk'����#���/�o$���$:��f+#!Н�v,�^���$�0��"���������D�'�ϿY��0�
�('�c2�!�|�6�HH̝4?{Ya�f3i,�.��LPL�-�)�vJ�����=0B/>�����(���i�f��I���;���Ӹ��%��T����t,�<�}y]]�������C��q#�9`1��Y�a��RN	��2q5��:}�2�IO^�`�A�PqK���[�b��!�	kq0�"��s��8�ow�I���u�v��!!v��"�H;��&�o��}��e�*]�����u��.0S���9�r+����rT}8��/7���mu�Jp�O8��}F���<�K�ވ"��������=\
�H��L�K��s}$0�P��~�~��Q� ����1�)�o��3�,�$ �Qj[�	�������4z�M�A��.}13�	���ޗ�<@h~���U�	����R�,*>t=ܘ��=h<�O�|�o=*��1�20-oc�j~=��W/���M�W�Q���ו�E^6q��������R��=O
N�g���g:�˻(aǆ��
F��L�}sTO�rj�� �\��Y�gJ�݂R^�VC��}��Oѫ�Q�gYԗ�C�<��u��x�"�������`@��|�PMİ!������^v���Cg�x -�^�N^��4�6w�H-~K�a�H��o��!�Q��G�R���J�b�Y�[+7Yl4���?���u�v����I¤N����2v3�u��W!�Q��2 Q^������i&Yh�R��z*|J�1wv�tTbKJ�J���rj�WZ���6��oF���^�CtQ ���Y]!z~�΍��R�׌��sط{2����kz��fU�a���������y�#,[���Q��=q ���Z]���nW�����"T�w�P�-�����>��.MA�+3��T.�ܞd���ҺZ��T9c�%s%
},-š� r�E�ף�"�
�7A1*ȼ^���!ေ����+a�ӏ��`$nN�Y�ʧ��yع/�t����~�*����QW��5��,�-v����N �K]�w�i��Hʽn�.��cT�H��Z��ts����<���&��X�d�m���3�沣AE�{��{$2*Y�ó�X<�q��ǥ ,��:�����[^�6[���e���`ܠ�n��F:��n����շ;������C�A%U�������C��(�x�m�z.o�˳��?~�K؃Á��j��� ���c�����������UtN2���1�Lx��W�Ev~ܐ�@�m2�,�F�(x��t���t����2��q��<�_1�ܣW�-��>���w��I@5��*{���Xa���Uq�=Q�H�'����֏Y��LR�V�6�P� &���w9މ$EIL�(�j�ٖ>4�UQ2�Q�-���G�h9�_�(	0�e�T�
3I��s���{�&��3�O ,_�g�/�3|�ێ
led��������9x��O�ߧW�h�o�|�K��_?�;�VPd���0�Я�R���qօ���~\O�94�������(��9L������p���u�a�S�qE]9�b`�QA���/@#[h��D��g��{<�> i��g�i����o��+J, ��!�X>�'ArOwpeq�>�b�t��Y�ҵ\ޓ�·�̤H��%-6�D�Yr�BfG����(Ң��-�S�������*vM�i�����ޅ`������4����D:��������F���b��G9IiS�����ҕ &��d05N�w��*��t��c�� �T_d���6#���\.:a�X��_� P�
oqEM���0�pEV�Sq�^m[��o�IJ��e�('��?#��,���prs?��q���y��m��.�0��BF�^k>��Y�΢#.h9n�o �:[�*bu�Mҩ�\��"��8����gѼy\E�Yx�N�G��ɬFY�=����Y�>puWɄ��n�j�}�f�V�kƳ�{��g1Ӕ�OU)d��A��z���e=�B�5��{N�����t0�x�
{A=���W������!,x86Kk	DMsx�(b~3�ͣ~afj��Bϸm$MyBϿ��v;�;�'��>��#����U00�VPN�`+U��)va[L5�/4sxFس8�:�{X�k
wq)�J���3�mVr޿N���)�5nUH<u����`-���*�;�+����v����9�.ۉ"����H��r�w��mɔ��d����H�O���`��D���/�sS复��:d+����*�
�D���v�
C�ofpJ Ă@��q�KID�
��>6x1h��:?c��7�v��)b��JeD,������?���"q3J�6��v�G`!66n�<�2k�=!�5��H	2*�y�A�������t��aMh�*�<Ϧ�MT���N����/�+��S�i`��5(�,#B<��?�7���q=H�aMm�F�	��q7~���V�22%W ֧1e�D7�@�*j��I�م�FĹ~E�)����Yn-K�K�����ڴ��͕xB�YY�O ��t'{��d�y����RA�1��)�"��"w_r��[���W/P�3"Fx�m,�����c(�o���+���d�e�:�����jB��r�v�������6]ʮ���^��/�P~Bh�����2 ��D&��$���4���>u����%�s��D9ȍd.|�wM�v��2|]����@_}�ߢ�Y�F/��Yց��6
8!�$)S�Q�(���=/�N����o���PLM.P��;r*��R��TT���Ҽ.#\MV��_�9N)�n����G���@�D*��P�z�x9-�䝜ȉK�\pP�-e���!mt:�`��\��`���ˣ�� �1XGN�NzV�V�΁Ô�����'9�|��ħ�E���[KWp�_���I�.�7�g�P�i��?��`�j+ڔ�R�hB�[R+�3,�m���s�C����w|��6
ӕQ)��q���"��\=p��Ϫ����P���1�(p�L���5�@*��&L����+]')9F�,��vf�$@-���E��xTk��g��h$pV~s�ә��@MVJ���C,��I^�|n���%�g>�� ��[yX�.&q7�ZJ|�q2a��*A7T7A=&h]�5��m�P�@_��3��q�}�`�8�����d	���cJ�%�6�C����N
vu �.����`%����1ѯ}
C?�<�3ܗ�ҷuY].Y�w�6Foӓ;���qE����#�{3�BPÑ�k*�R������؉WsNaFu���B�У ����d4f�N�Bf��}E��3V�H��H8]�oہw��q<YTV��/S:��T�EQ��D��U^]Ҡ�bϹ�UiieC�l�X��ŉ��b��o��Z��;Z���dmx̽�GLg$�Q�p7%W�{���6S�y_z|mnM����')۸4pm�k����f�%E��]&q�d�(^�r��|�����E
�CH��C�b��1�ۺk@7�^44���-���t�҂Ie�?;�F``췃�C��4Z��{�����@3ee�b9�}�Y�5�`�-����u���Ƃ���Ĺ�vbjVHT�\$F����1�&��]�]p�5�ӛ=���iZ��-�|PnFx"������51Oۡf�StB���#��$���nNo�ь�Ya������N[���~dR4�~���W�Q��3�f-��ݟBv�{��'m�(�ܲy�����e#,��.�z���p������<��u����ag�M"��/LG�3��ޙ���B��qRJ���.�����ŃU��1����X�˲QEfu�0��RM��~ :��~��>��RV�`�k-=+4���O�r�ӷ�<?x��ί�����[AS�!��=�٢Dj���_r�T�v��X�m �t�{s+��e^Qkn�����)�ɔb� �^�q4M�K�o��(�;�����^S;��+��ۦS�.�[i�Qm�9L6�`�Z���߾�JKks�"8`eD�f��B8<r:06��t̱�/s_���8q0��������mː��T���P�D��A�	�,,�J��/��P�E~@�Ũ��;YN��%��N�j����=�	�!R�i���?N��Rf���t�_��أţB@�4'"� #���77 �s9��D��֖E���2��0�4�/=�F�~�>�����E!��.-T��B��D���0EAd@fm���kQ���#[��U��J�ic�,q?w~��I��zY�9��%�t�f����`��:&`�F
�AA}�_r1w<=AQQ����L\����z�������{�6�x�rc�}�Y�M�<�Ͱ<��V��_?��He�iq:�	Ʃ�����R(�os|�ӈQ}��T%(�<?\J%b���w��z�D������ ��9�����X'mP�i>�+�g=O��ɒB��2E�$(M���G���$�H/y.B�Ԝ�`�F�(F�q"d�� �ՙC^fB���*�FJ�����I
�\W.����6>R���Hܩ]��Vb�d�0MYr,�����ȗ�AȉTL�����E����Y�ŭe�x�6����Z)�I��>�^F>�r���&�s ���(�/!H��T<������IF������\�$ E���Z�������-_����1u8�҂��J���0��<��LQ��c�W~t|�Ppہc_���.�!�Ũ	��C�kl��<��6�	�f�yJv�5@�>�����mφ��xBR�|�]��B�GZA
��O�E�rhV�U�>_���5^I��I�L�-Y�:p��|�J�AL��KS��X���^.�w*3�}MV� �%�!&�-Ii4Q�� �3N�]���U�IQY���H�e���YWLF��ŏo���LЧ'�fp��;/x��$*�:h��\�,c]i�߲.�zӳ�]�/��D��q+F{%�FxN.�B�_�7���B�0�p=I8�>'�i�2"E��j�Tj��QPZ숝��l�lqj�����a@?��u��6�ؖ�P��S�a�w�e�|t��P�A��7��=���� �%@��y��q�Ca��v�o88�q�k�5��j�M�k��F�8��J�2�Mt(T��s�m7.54,L�Y]��$Z`�	���񟿼��f{���X���+Q�ƥ��y���+t�'��E
�Z�R�V��2?�;��mE���k����;R)�9T����ϟ�����(�
}O<.��M������Ǒwy�{���gm����
e�n�vl��"�j�6_+���+R�y��i���!�$�M6!�D'U\��Ä��iD�C�1�w~K]��&��C�ԡ�Ȃ�n�"���hz�;��~:�i�l�=���dL���Cl�%�˗�<�th�T��՟��`�䳤�S���Ue�+G��1�S�S�+�a�Z�m_U���r��w$�i�����3�k�(q��TS���]��4cq��Mf(��[8��se�H�g��8M�KPj�<�YB�1�K!f�+�f���ͮA,J����0�l�PO &�l��n��T��q���>��V{��$�!;/ٌ��QQ��yB�4S·n+��g�5@Ib��%��"4l�!�8,�m1��<d���WP0��ߋ-ǩ(G�B�3�,��D|��0�o��[�C�=�L�)��b���y�ìT�~E�R1p^pKg��)�;�(�K��m�ڙ�B2h�e�:���b�a�d,WH�C��Oj��=����\>Yo*�L;��קI;�[m-��=�D��'Ȩ����Œ���:���?��a�$K�ò�5.WZUΕEC!-q���	(|���_�}w�N�L��v8�<-�����![>�-��"�'�eΰ ��Z��0�e�H��ss��a��}�/�M�˥�ʚ����;��}����c���4�D��2�5��M�wP�h.���DL,�ń�0'|�wa���=g
�����7�ߤ���F�=}	GK}�jD2�4q���^�Ɂ�С�Eo3p�>�4�Y퇮��?�=�:,��Sɮ�1ջ����&�EWdO�+��$.�PT���2& ��uC57���Y��-���9{�XF���9%�qn]8��Y{<Q�}�{�x�Y���b,��.�u�f���/*F���*�>&�T�۶瓣Y��6�Ӊ���&��#�D�\i]թ���Jro���w�&U-�������*BwY��Y(�/NV����9�[s=�o�ef�
�)9\IM�H�eʕ+q�V�.}�/�)2j���2A?&�,���[�c�Y����9���`͖��)�=�ĲR f�S�\7��E��u ��!� �m�]�,#_���WwK;�< g�w���:]X��	��9J�?���C�?��V0�G�
��6��=b�U����~Óe'�w}	��]X6�7Ld��u_!ش���A��R��b�ͤ�UH�i����d1�s�KX����X�T���K[��>O�����&F���
d8{
�;�N��
#�'D���8����ď����� x7K��ݾ�d"���j����u��w��2�~'7�(u��U)m�	*_:��i����$դ�����g�)�N{���raP�����G%#�l�ƻ\5Z�vL+�m�_~�zy{��[T7�j���[�KpݛkDJ���y��	Η.zӪV�.H��z~�#FU���Z��L�!�K_c�b�`
��m#6
B�v�PO����S�eq�^w8���Ahr�C����~�^^i��B��(%�=�Ԡ,��@xF%�q,[��<��my�T��nG�=I�c�����s��څWw�8U�ӑ��q�IzVK���ɗ`	#�T�%)��ane�4F�Ү��4�˶r�|0�'=���4�'3[#�8������+���I��_n>�b�<�;�:��a~Hߓ��~�I�8��S��1�nų*PH�BE��VU�s���PFUm�CP� ���c��%Wo�~���_ŽP���� ��AM��� �1^��,���.Å%�a^S+�ǓQ,� � &���?'0blBL���;E4Ǵ�&�L˽q_�9�S��;�E�g����l=�"{��?�C�^{���W��EV(�Q�{͒��ϔ�ѥ���C�<sPby�SZ�m�̴���g�1D�����d5����W>�A�ڃ'��Vڠ�%" 9o����=�r-��˜pac�.vW} ��e �O��ac���&��3���R+LF�8D��ˀ�I �.�r���d ��8�Q	��XsE3j1GrY��*�r�I�b!R�Q1�/�����uFO�E�L�g��\:��t��T���q_��O���m�����Gԭ(aF{$ 5�"+����s�Pp���$�G�ԇgĉ�Sw��ٷN6z��t
!�i����-˴x{+���:��@�Xג�g!�#�@ �Q��wN������e�\ݨZ�8gz%�i��r�#�&@1*��_^�Vg���·�h��Kco�|<iu�jQh;�
�t�8Ah�[j6�i��2J3�嬍q�^��+����kOF���Q�_�ܗ@����WZ!�*G-!粧[�f�ѧ���������mh~I�<�٦�Hm� �H�*h�'At��_�
T���V�V�HU�1�W/�����)*U��� �&	k
�����.��R��a��C�*�JQ#>dpOp^Y��p�w���kw��A5�j]���c��iSj<� ;��W��]V@������5V2�0c�p� �~�C֫»��?�؃�;~�r仡"��j����/a�ļC
����?��� "�K-H��t
���[_�%�:.|�p0Jhz�䥺R����Ԁ'���[e6� �Y�ׇTMe~�g��uܡ�A���㸍^��^�gz܀��ޜ������٪ȞV���,�"h(�=@T��0���=�����oV��`)	F�a�9�y��=}�*��I��5A�Ӹ����=�(~���#�fX#{�>A�m��A���^�H�l����?d�'J$���6�籲jj�AgJ\ A1��{�un;��=j�|�~��tף�,{��3�f:�T�
��@�͆hR'V�"*�x�Y���ׂAŏ���^ܵA~�I��!��������}�A��%�VYp$�guަ�!a������\(�Ӿ���ǰz�H�c�Ic��Z�������*���өyn�nU�(%⛼�~�'zPG�����Х3�5�qT��|s�@#����NH@(�ΦJ��Aa�����8J�6�o�W�X�%r����/e]��6����@!�	3��&��s���o��R���`Ѡ+��/J�_X�T D��_��ܚ<���M)���ɷ/��>\�㥂H�ɩ^Bu�r��r��E�DQ��Ģk�(U:��G�������m��I�d<�L��8f_�D�t��M�M��;�qI*��_$�����B!D�*�9~)/"*�Z����9R9�',��M�ߋ���N�s^��q������r��8SW���l��>Y��A�p
n�Șz���TG��%jdY������co��A���O��rJ�n�����1�owy�JMu�tG�[)�$�[����(���B�z��]�V����8�:��L�n�;��*�ސW3��<�����)f���B�t�'���Ũ�Sϧ�<�P�`Ǻܒ�ӌ(A��=�d��A�7T���7w�6u�6JV�{)����Z1Y������F-e�e�e
bZ����jj�f6
���z�Z��3�Ǧ۹�?e����~v����S���IVM���Ѐb	I���F"��@wi�l/{+����*�,���ә�����o��P��eȹ��m���Nl���,��ا�wd���m`E"��GU�1_7��k �#l[�b5���"W�2�l�{ *8Y�I~�v� 
��p5�p3�O�F�5D�F��s�o�ۗC��֩*��l�N*v�$A���OF����?��J�j���&��q�k˯���f��km����ZD�_�1�PGj��L���u&@��N����$1):&���:[Myc���c��>~X$t������
�3�͚�C��m-pqT��^}���ʶ�C��$RC	��kV��.h�5=` C�J�A���U	1`�N�(���z�c!���d����?.w"E`�����[� &	?z�W1Ůc�W�7�D�ώ]�9�����r�%���(5�C�f�7ۃh�d-.-��V����ǂ��'�Ɯ�T�G��	(EY�,���`�(�$V���xP�4e��%��X�M.Q�Z�#���2}D�4|e�?]s@)	��8(-�����ꧬ���l|���v[^�8����� ��t�X�9���\զ������B]�ȵJ�-�Y����i�
0�����7nJ(HN���s��H���s�<�Dr�rs-x�؉�%���q\�=e�\ܵ&�O�R�>'�`��F�aaA�%���I�Z�.>�����z����1�+xo�t~�c7�R%�+���.~�=]<�_��Q���f�s��a]������M&d��#[:�JvH��IPQ*�.�lyQ��+�g��6.��g���ܫ�#u��� Q�Y\X!Z��
��:�P�k�Tu]��u�����⁢��T^��U�ZO�|*�ëU�������(]#�ah��Z-{�dJ�U�,m{iG5*��6B���9�o���w��/�X���+�;�]U��.Z(�&'�=�vxo��:�pL�"�IV�`���U�����D|o2�q�^�:y�"�v٪n�Y��"��.X@^�E^A�����[]���|��F�f�7�2� jnH&�e�/.�:��v@�CC9cxt<�m�-�6�%�Ń{������������ɋn7�|����y���|�<oR�IdOy.Ӎ14� 4���CNȎ����Rڷ�Lnb-�5^@�u�|�:�m��(���Әý�N5&_j���I�l��>+&���O���,��T�E#I����Sr$(xg�&���÷�
ո}�m�0*(,i:��A*�l���.eJ�k��`t�46Ş{er���ːV|N\/�����9s��rqX�"�n/�����_�����*��a �Y.?B},���� ZNP[V�?�����!le�[��]�`b�V���	��+��#	�䡍]�=ЎG˝��`���"�/}����yTy5J0F��F�g~�+��KGܜ���x�z9�Zk����B�ؖv`I���b�Zv�V���K���)&ؤ��͡��5�Ĥ�B~�X��6k�$���O����$`Kn1���a|�|�ƌ�wIf��f���2)�{/�^!(3�&G�ϑ�N\�����u��ݷ�1�h^��띤��=� ���_*g���h'O�#�@��0���Q$���X�����<��zNmX�O|�����X :܅v���i4O��X��&�^�)4�[	qL�l"m�-�4�N����Zt�Nz���3�J�>ު8b�����.OZZKީROη
x7�l�z��5�F9�Iy���XL�{��8/
}�}���O���_�є@6�ف78�#��D7D��E���ߐ��0���.1��N]=3cD�A,�O}|�/[�@/nRg��₷��,	YS��ޅd��-�����v�=�I�<S��=�+��	cz1�+�p7�z7�ԙ�A�6$d8(̤��ӛ�Y��I�?�ϱ ��������#���Eh�M(�#\e��g���Wo��=����h寉gۊ���22���=��j9�2u�:��|Y�ҹB?�� �*�a�̟�U��c��fڥ��X��Ğ'�T8�-�w-�����j$�
a�@ޅJ�i��Y�~n���(.;�0�+����o�i�mr8�H�MCe�����y�*�HۏAW"I���4�u#��"�'LM�V�z܌Y�A5yyOO/��lʍ��eT>H�j�Vˌtm��#Б�^�"�R/�ᨶ�R��F��-$*tA�P̤\ z8P>.�'&U�q��b���u��o�&jj)��\�#)��"Dx+�/ ���IG)2�C����𻺴I�a��=�i%H����I��޸Z��1o5��,�Wů6y�r�g'C�'�������
lnu�v�����AT<�d�wE���������U Wy� +g�vdCtcs�������d��Z�Q�B�x�7�JG��m���y]V�g�]�عXw�D2g���/+(.���IZ��8�$c��{�d#���vN��0D1���c;˩* L��3'c����	��~�d��.u
2H�㘺��fȁ$T;�6kTa���E��9�-J��^�"$f$	��L� ���k5>��-�%l,��6�~�)��)p,?�p��OT��ob�$����&�+�(����1�d$�D��-=�:n���u�)�8��'���ae��,dk�&*���4���߄��рg�}���?�0�Ѝ��k�D��d�E���.[����^R�g�B��o���G����b-�ٝ~'�
�)A^<����Fئ��b�R3{� V�o�m2A����_F��]��CӳLݺ<�8Q�>��VX��BV_����ld|���Yp�,5�@cߘ�MQ�=�������$w��p���F�+��2A�ذ^�/��w��C���[Y��Ӭ�B��_��en�á^��>��z9܎H�X���6ѐ6��f��k�S-��Da�����O2N�8�һMF{���1�� ���0G{���Y}[�rN�����4\=r�� gy��tB`{�ϛ%
�lfn]	i�Q ,���2�*�1�uTd��Q�,�#�L�t�?����K���9R�8�?�A�J~��5�A[�H��Ч��/����f߽��ź={~�:��N^<o%^����$�9 �U�k%>�ǰ�""b�,Fq�X�+�)�F�0��}a��b��u߻-�_�pcp���Ms�d�3pk�1��C.��A�T`�����$�����?3�F�e�K{x�;�b�L<|�$ 	�{,u[/}-�2N1bt�_��x����� �֍��e�,te�v�-����bQeU	���4(��reJD2X�V��}��'y�er���`����@�+ѫ�S$�i_���q�q�P%�9��X�b���ɣ8@p!�*�
���UkT0s��f��އP�ҝ�n������\�*B�:�6�"�}��N���������(��g��Π�?�?�!��L{�@=;ŦV	1^�*�\n��5�����4���"�*i��%��=�/2�&�;$�i������F���ȅWZ;��.�B�7�>2���c"�,7P����,P��Ҷ���c�⣣��h����o�b���3�w@5���ߔ���Q������J���;Z��Lx?��8z`����o�p ���!��4��O�w�!K�y_[1���)ǌ��6�Ӛ�N��`V��A�mzg�M��X�3N��G
�-Mِ�	5.z��XB0j�묒0q�P73��Z��i�ZU����I�#���Ofl�k�� A�4� �Gn�6+���ܴ����I�[գ:M(<�dU���G+���d�.B��8j�U��l���%��V]�឴7gw�,��I;g�J3r�򛮵?�5�Ք27�l|R ���m��K�*�\:�i��0n	$7j	�c̕K�v4����%;����o�x�����D1?n�����l�}�r533U���=��Q�|�7]���R̗V�#�3�h<�g ��: 3q�l�~���{���O�,Z]@,|�e;��3mR�ȿ���I��M0V�3��N��XrUM�o-�<e�Io��tD��!�e���z��dʩI�.�e�hz܉S��V�e� Fr�n&��I�H9�g�02:7�[hٟ�V�j��W^���{�b�s������Օ��ٚw���+ԋ��x�S>�#[������q�:�?�5ww�C��r��N-��o_�<�cF��=Ǹ�^�����c����ϑ��L�D��:�Е�*	�H��}%R�"�n���nP��v�O��E WAE>Z���n���ku(���
���"����^b�`M?���!B[��,v�^Z�=֪n�VŽ�*��m�.9���uy�- 	�x��W�M?}$��+��V*�!�M���x♹p��o�fР�m�����$gf�T�j�WAb>�O+	F�w�.�u������J�mñ��B�GWU%C����j������k4�h&��͘岴�\�$����&�'��w�Ib�1sT���^�oY�E�A]�MqV��*����� ���}N)Q~�~9=��l�9���Zy���5����t��c���<�����貺nS;��t�;�=�W����ދLk/@�;������ʠB��NGW�IB�1���B,�m��|Z�S�}&l��Pj��g���i$b:�Y�`VZ�wф>+�*T��<'7IpB��AHL�m���0�v���H���\���ao���_4�Mk¹9�
7�6�#h.�Pf�r�:�h9����g�L��؇U/"��ٰl-���oe�PdTQ��Ǆ�\��z�勛���Q��6�\�� A@��W�fT�b�ͫk����Z�]������*�$��3��^�6׊z	n���;��VɌ�uI��}�He�R.���=|���m�'إ��������Ɉ2�i��B%�����k4�$rk�����K���]�9�XQ%���ڲ̉Hf����5��)�M���\�]�q��П�%�� �s�eXz�v'�Ж���0�<J�[�G����f��>��p:�cu�>�ȯ�f��>��?1��}��֩�C�̠��0���/�>F �/\q	��)�T=������ݢ��	���O��:J�ka9z����@�q�(�W�dc�A�r*%" �oz�ޑ$p����3x%��sz���0�ӟ��Ղ�ѻZ�]�j�CsҚ�����a�%��ǒ��s��D0ؐP]a��O"�.CҴ����`8�L��mc��P+�3҂;����UT�Ɔ�yL_q]_�jI�V�i�Нl��@�q��Z'����v�UZ�U$+$� X<c;Ie�cu�%n�i@'�Qh��*��	n$�?��3��b�j��V�����1�s�}V-���1;m_�<,�����'�O�t���i4��<>�γ���F�=0�X��\{^=����]���7bG�J��R�Q��P�3'����T��L}�����ޗ����IM�Uxm��x�����B<�f�qI�+:�WO.�u�)�����f�����n �>���m7&S���Q�t�;Q��+(�f����#��1�e��������|�2M�h�>�~ⳃd3f�6����8l6+�$�V����%�����"A�%�/���[�Gyo4ahH��*sy,�C��� o�>.+�|C���0Ѵ�U�,T/� �
VY�!�[>�r��51J�ܐ�Sn�d�4���!����H�bkm4��riw��'����GA�G�<�N�5�0R����rd�wz/@m�3j X�}pu
5:��m���ާ�W�Vc��YY���Ѕ�2�ԋ�d�J���V����f�u
���t4���~�γI��@���MT
�4"c�)�T��gZ��
�j숪�*?~�Sqf\�K<I9�WQ�w�����,o�aةCi�1�T�6؛R<�� �����3Yyz�z��)Uz�͆B��V�+�!Y����?�����	���]�(�ė ���Dv�hR#~�YR�E���, \�ਞ3䱩��!]��b?��N -�;R��`wv�6W��ኞb��F�� ��͊��p�$Ppc�6�ω���:v����Q��%��3����-���ٮL��,���$t�]ԯ��u���^��l@��u����� �#��}~�|7�j�uoz�l�������W��&ً�{7�����>�P����^���0"�Pmӡ�X���<A9d��Wm"� �w�����C�9�ū�_|�k�<XZF�+(](:�4�����*Y�2�S����ʎ[蟦~���B��ra��ք��ڟEݻ��^}�~dtƊ����Z�[$����[�5����k�-�U-9$���y��^L�/B�}�H^֫;��~�?��.�)3�G~��	�;���ސ���8��ײ�i�wq��.sD���7���TDlW�ꖢMD��,&�+��v��|��A<{05ߚQI:��|]��_��������lq����'	>؎�A��U2DBj�/m�+d�ܙg,�0��67�hi�7��Q_��>�9�y�H��ة�cv�P��Ϝmي���/��Nb�-r�'gE�w=�h^I���R(ޒ�:����l8x��G�j�7���`�ٻC���a�]x	�,� ���uF�44:��":�y9���-�u�S�\�ɾQX�CT�Υw�/t��7��B$ità��a�8� x���r�LC��ʗ��!�m��=�������.���C�=��$u�-׉�V�V�v�==(�n@B� �?U"D%����}X�	�����Y�ek��X�o]q'��+�>��Ă{!E�X:�?o����Տ��s�pI�gJ��~΢j2u�H{e�R �G�''��f(��%9^�_�J�$�:|�䧱�5��nu�.]ͼ�*�(���LS`���D���|��}o��+k9i�Z�b��S/�9����z2k�[���(ġP.�i;5g�<�tP�X�x�$Z��)��=�0�_�Y�+d�%R�u�ܪ��N8��m�][��^�K����I���#��c"%N�u:I�6���[6[>���~DRwwΊ^���n[�ٔbV&s�"/eX����Tj*#WyN�	;�2."ry�, d�,���ȴ���>zB�D_\T�T�q ٧O֠�{��<����Y�{ӟU���hW�K���Э���� ���y>LM���pC��t[Rb��۲����q��\҆k3✑��cz��Z쑔���w���j�Ѕ�:ôՒ7H��-�nf�6��1��h2,�q��ա(��U��Y~h� ܄1j����V7�W��ݡ&%y�r�F����5�u`��a3�L"���;�a�_<���0:��Cƫ?���v���4�'�"\ko�n��G�3�>ؤF��Z+��v�?1G�?H�4X��9(�H����lqM�٫Р�<��tH{�G؁����;�AlZ�t$Q��3|{�U�ȅ1������Fd 0�JVd��]]�Hϩ$F{n��'���9�y��#"Q���°�k�Qˤ��p���5a��ڀG~���m�rGv��2ݟс� vT��g�5	�_��C�	���]!XI��_����A�룜��RbW`9�Rn#'�zm�Lu|�O�~6��B�/�8e��"���O �
ȞȪ}ޝY �	����yb�K�9�.����5 ���#�6pn�a�k�Q��b�/����>ƽ���n��� ���	H 1�i�+g�}a���c]?���r�J��ٝͻ�����3տ6�B+!�ա��py�*�Ɩ�Z�D��[qu�/EwG��+�:8��TP�:�I�r]�i6*��}�ཤ<5��(���d�3p �>��%W'N+���B	Ô��3*Ү�ϵ�5�9Y9Z� 7R��-XD�
�$�`��(��v6&I���+�DF�E,V�Vz�6����,܁҂}0^2���AX�7��:�Mh���L�{A�ʼ�$U����^����j����O$6*s[���n�A{Z/]"� ���`u��0kI%�9Z�Ȥ���B���s�m�_u�뤬C�� 1�[}���Ű�^$ې���-S����:̏�|����@U%��Z��.�\��͢�#�'�:C��ΕQT������3Y����T!�|B>^t=��}����Uw�j�L�i
���:S*̰C�r�q�)Q�*�aG�%� a�0_J��x�'���k�)C��2�_/2�~3*���xl����FF��kp\�
�f���r�{�A#*?�ܧQF���q$5�6~p|�$a��x�K���K���JD=�$j�<�T��B�;��E��2Ce���*C��+@;�0h�P�dߜ*���4���;��dx6�DK� P���B�:=;�K�sSl&R��]t��T�)����K�5��2\���	�u�� �	���F�f_�<�{>DjaC�a���b�O
������&�Eb�|��c����y��z�4)�'�y��:hIu�^�p�}�*#�o���^��h�7e��X��*-D��agb�5쑚�i�[��&6�z��2ݻQ����#�.��x(�����9�'1��1C��K��m��a	}G�a�&����՟a�_L G���H�i�s��&)�TcEA���MP�(fB ��U"XzX�=ҏ�]Nr�\O,�$��{��R����_[)�� Ix%L�1��q�&X���G���)�<.+)�F��>h�݆�j�� k�ٳ0y1�x:�Q1)�X��3��2��k�A'PG����t>A)�M���ZS h��dO]"bFk'�E/o�ӑ���mTJ�����F��c��+`ƫ����W46Ժ����B��	Z#, ��eb��XIi\Vt20�=���c�;|�t֥M�\|Y�z�9D����A�R��ɴ9 e:��e�Le�G�_a�|�~����
)(6�̔H�ͯ?�
]Jʁa�˔��]�c��C �9�`vhS]#q�^��}��-�x
m��p���c��;j5dX� �4�t�x�cR����9W�k6��@ ,�?巻�]O��z��<1c@և�P�w#W�V3���S���=�1�Y��@$��<BI���4��*�{��q�X���sN2��a>�ģ�Pa՟���l>����rp����ɎR^-��\�|\`��xO2�q�9]�� �b7����/��0@j�A6�`�	�q���|f��F����֙�zs�z��#�<��)�*.���p���f����vw-�������\g	*��$c��-D�>�A9�u/�z RCFg���}�ѭ X��$b06��#��N�k[�U�i�t�ǀ�z��Y���k�E���e�$T�.�4����;e�J��Ʃ���	���D����>�����mQɏl@7W;�ը�d|>��<m�-_�cl��b�<��X�}F���0ո�\��N@x��J���ϗ�?Át�z��n-�;X����E��5ε�f�h���G���ְ�������.�v&�!H��0p�o��-�`_�T��D��2��-T�5=8���Wz�þ��]M�JR���M��z��T�QтV��"�9*#7+/���O�y�^q�L��; SJ�gz���&�5��u�1A�}W|R�w�Nu�]f�wma���D�"�B���q�3��qALD�%�@[�^@�B	.�����C�l��}��EfvNo�9�Z����z�(���R��x�_����en��1�|O�Yge��Mn
�;��\r(jP��T�D�����2�x�Su�Gw����֋����C�ӎ:�|"I2-��|�����׶�o���1�.�{���ӿ�daz�K�,�����r�s�4�J�X�4��#���*�e�̟�m��ۿpH����6S��o�:=ӱ���b�t�:���Ԩϣ��e����".���-�Шf:���+(���\m]�A#�G��~<Ђ��`"Ń��/>��B��C�q��8�|(ֶ���s�&������B^��H�v�tNp?ykU�4A,�g7#����`!��=��+ƻn�*dϐ��ј�1g�X�X�9�k��r����T7E�<�#����N{f�j�����)-����:��[|iD�$^�`���/��x�J�o��q�?��5����Q���+�	�����	��ɀ�R�<+��-�E�v_13����iHț+?�낭i�R����q-W+~��q*~R�S�UFmG���29��6޻ӱ�u#�;D�=������YZH�p�[��	�����0����y9�������P�t^�G����?���lK8��Ƀ�8\4q�%{	����t#�rX��o�Kv��C�����U{{��&r(^�Q�Ha���~a����l�/��1ް]�97��<�j��	�,���V��������&�����(f��@
���Z���
0'�Kq��@Ԭ��%�P�o��"������)��w��!���ib�s����T}8��T?±Y�:��%�'|� �:/�ϊ𘽏ם�ǭW|��u���k�(�L���[{^��*v7u)i��i�"?�j|��Ȍ^����D�hjeT��~8>���Խ�Kb'[�)ƌ�Z�G�[դ���S���s��L������	�D���V&�ܤn�ѩJ[�_�/B�<:!Ak6s�^���V,�t��FxqC{_u��3�37�J�&�uU'��7��i��a~~�#w$[a��2B����.��3�<tӳ�����ٴ���|4��n�����w3�Q9h	��Z9F���|r���D�B�H�0�,��t=�����K`��)a�|�񸭿�d�֓�3�G��r(Lr*R�������.Z�h�e�jrM9�����6MYz����������@�_�2�
��q�t��=�XOVI߃B�x^`7�0��%*�0��n����T�m@� �e4 �9��&O�ɦ�3�ZCcS�0�ZjA��.��������[��X�ޥ��b5�;��|�
M��:V�d?�΁r[?i�7c)�`��>}�Ĳ��Y`29c�q �}9�@���R8t'y�Kw��OQ��-f=ܠ���oxn�Fx���,��dC�CY?������[J����=�^��W�R�O�����Sq�0D} ����#��Bh�z�
�VN�ݍ&�9������[y��}�l �n=��#����=�/o����xP0q�."P�魺��'��網��΂vX�R�}ō�����dzA�"���D�k����4Z��WXa��X# \�4�@-h�^S��B+����w��P�8� e�����L1ֹS���2]#�ȍ�J�xmh�@�~�G�����+)�����`������ADZp���T��l��K�QPd����gn�0Qc2�1ޙ��@B3�m�{�`�����[j~p�ÐB�J]_�eNn��J���=vMql�l��m�-M��0�o���(��d��1d��� e]����'y(�\a�̔�.g���	�tQ**7d#���Z��_��,��y�8��W��1*�Kܒ.����u����t7E�	o�8��M  7ǟ&�����y�g|��V�K0cE$�B����,� �=����O���)�@� ��ɚ�4�㒐u+�i�iʟ4À^^U����f��� :KHD��O�:n�⭁��տ�2�$o�'�LHT�R��׃��m�l!��N/�0;��M��+�9'=���ǈ��;B@и6�勘�24J�z�8:�k�,�3EU�'=U��գ��E!�oAާķu8H�S�r?���q~�	�� �ja��S��~,�TF�T/�R�@Y{ȝ-���9W�%_m���Œt�v�Q2�$2T�9��¦)z��N�򶏖F�0N�cj�w���Q��ɳ��>=##�1��}�������[
f2����-�����7����Ǿ��dVwK�2d0����I���� ���L�"q�����ROP�p����O��]á�l�xk�>61�+�y�>��%�S]c�\� �f�J�Վ���j��5��o�j�_��x{� ���{�r�<�%.�8ࡘ�7���4\<=i���Hiv�����?�C��pZ&#z_��< K:�v���Q����ݙ�{�c�EhT�Ee�f�?�����֙!�(�H�n��AQhi����_/��f ���Z
ރQf�Y��e����~	�rx)�J�媃��i3&*�`��a�Q�ƌӪ�9�s�ݣ����%���E�m1g��(�7�z�	�X]2l�h�ti�~o�uA�=��h�u�j|"|�=(�HoH��x��N������2<d?c	
��B�a�#�v�@�v2LнAV��P��_�-��M�tȪaU΍��O<���jQS���'{�TrX������)����dQ��hN�9�ff��tG��&��md�
�efU�����(�V	@����zXa�_�R���g�� lq�x�S4��	/�ɷ��Wۢ��9� D=ɥ�fx��>{�� �6��i{n��}aO�j0U���)2�����vj--��7�(8�0Q��g%^y�1�D�g4�9�O��,�(	%=����%�ͭ�#�t�q����>,���JK��b/N�_�{��W�؃��pN_�5�՗���3��r��`#㼤y�/���=}j*ױ�C��1沁����2�W�ɣS·'����m�7P�04I�D�u=�	��S���K�����UM<�d�[i�3�B�2������B�ol��ϲB�%���#_��	8��1�%`g�#<~�[ZE�� 2�d�@�2�>��~��4Ɉ� ]��H��{2�S\��7&CF7S��y��M�c��
/M��%�G�yಚWF1�=Н�����5��<����b1v���؃����n��w�\�r!J�.ppM�^�?ʊ�K����^Ԏ�սq5�|k���X3�7:���F�m�G� +bn�A�i�<��җ��/dc}�mYC߀��f��+�}�0stRW�,,��GOLx#;���ܿ��P��KCP2� �VJNC5�/��� 5Be����".�|��l�~VV78�J�b��Vd�Bӻ��mf��{ͻ����TP��4���e{��MG]�-1����(�=8��B�ITFp��: f��A��p�}���Z�����l�v㪒J��&أCx��vY�_Z�0�j�4G�����U�K�����((��nJ��T�ߕtZ�+���1w�Ƚ�Z���X$O�Uѓ�r��"�\�$i�� �Z�����Y�˧�tK�Ȅ��L����)���s<����jX��N��SF9�dU� v8� e�X���&�}����N7б�N�)ϼϱM)�h���|Z(��y�W�q�"F�Z��;��*#)i]��;��by�|f���r���97h��4p��Zȧ�b�A���C5��zF���P*�M������\,/ G�Bġ��k4�x������E�WLB��߮.k�D����HO�	�{y�c�\�s����g�צ�����	�+��0<�<xFn���8t��h6bfH�9S苠EF��^�������i�ӆI$��� ~}_�RL��ټ�)�CE�& �W�M�/�$Ү�s��:��͆�]�n5L���h��y$G;��\���W�cFz#0���|�9��:�1����tuU�����W��
�(���
,�"H @^(�K�:}̯!�.�и��V�8Z?���E�Ff}�I뒴c���l}F���14�e�jK�+t�,��?�<x����,Ѣ���x^F��d͸��}�=�,X3NҨ���O�f��]���X|�Q�<�#`af[i��$[���c������p�'Fi��ĥս�̠q���xi��c	���V���Clui�GrW3*��dl!��q���n>|O:��W(���7�X�I#8��H���<>��a��.�#`�Ze���6�U��g�O�Pĵ���V�r���*i��,ޟ7��9�=Q���ϫ��Rd�r�
�ׄ[�M���ay|��~�.���
ۮ�1���3V/�����A�}�f�v�"�l  w֓7�ˢ4�7����ug�R�2𵧵�9Y�
�^HwpT~�L&�L��+�W�п��Y3Ȥ	G���<�$M��������X���*�O�h�i�z�/��N���j���xCS�5�x��bM�|i:�V���ǵ�_~������`q�a�b��p�cLm
��Q����mΫ�i`|��N,�=ml�����,j��.Fgc���� ����Cv��`����lc��b��m
`��*js=V��8á"��@����c#G= ==�^8�I�`�
Gb�V�CL�!sZܰ�\��wktR���Ҡ��e*�r��������]|0p�w*2���(���U�*x���r��k������Ux��C� a����TJf��/��w���1�0~��{j����Ъ�����G�=�p+8W*��sm�u�|���oZ�M��&�w�+��	�cv�.������*���&u�$z*,��MkF�Ь-J�iYy �q7H#�EI�ti�J�&re���Si�Q�1c��2(���|=�`Uݛ��Z���j-'1  ���u6����?8�BⓌf��'�!?�G䷤9��X]BJ�݅;L�>�B�Tw�8\:�i�QS���9�����VRk:F D�6X�w�.����G�I'��q�va�Mr���S[Lw�Ļ`{t�[`�:4n�
�` C�mK��h����>��N�6)Stj��dzP���û����{+f��,�i��>�@��Y����ѷpNz���)C�oQF�I���S0�U��q)�G]��{����;��%b��M����Q������4��#$��q��^�N����R"�_���5���gg41�ŗ�\��Q8���c�J� �}�#"�LC����,%�Ij�ݡ�Ec��<�Cjˉ�䦳Vr�Q���(7.���,�'y�>.�b��̤�3��S��a5tTxJ��{���,8GZ�����k�v�\.�,��.�y�:*��)��j�j9���+~�Ca���~�g�a������ZM�e-��Uڱ�i�;/�2��Q��ǝ�~��=�a[�1൫�^��X.���*��Ҁ,e
���o�[��:�����_��;�7��q����)��Q�"�$q��+���O�f�-@�Kt���$�6Z�c�Z1��#)y�w�H宫�;}�\,Pfy]Ze��j��\�Oh�6��'���#;�ㄧ�|ОS�C�!�2�nL��y��������6�~��e��L���+ּ)�6cq	����J�^?-�_��j}��3N�3��>��Őp�2�]�����l(�򖾤���\*XW���YU�d�/V��Ɏ�����RN[}q�G[�[J1�v���b�1��moc;}gqpS�(�6Q����ߝ<Ҧ��Fo:����No���-���!C�mۗCo<��3~�AfD`��3�D)N�e�AN�����_�7\tl	�}��i�I�Փ.p�c�h���_�	�� �7���BLs=����ϭ5��і�|����$/�G!¾�y ��G/O�n&O�����+�~��ۇ�pV?ud�v�	��tʙ@�is�wu��e5`���:�i�T���L+��?��\Fn���P��}�F^<c���JwK���!d�a�������1$$�I���)\^��.(��cMB���:�n/]��HݭT�P��6�|4�6�u�J�oz��%�A�>���̉��=62����I��XH)C0�!��:��Y��U�������y	�o�r��!����"�v��cU�"Df͸&� w�C`�97oѿ��Ϊ�O��&��?�xZ�e<
��b����#bp���󬨵k�(i�Ӊ3F�k"4�0��k*{�h/".iY�<��w� =�|��<����|���$}W"+i� ��x���u�V	n��T[~B"���W�o����s������lBT0"h�~��bh~����Q�vS���4F�w�tM��B�Y]�D�P�EX����j��]�42f�}��VA?tO�rl�%�U�l��vt�~]�:8"\q�${��j�Zx����D�8|�搢b��� ���H�r������2��W�/@�'�2�ȃ�<1�Ӧ�x��J|}�M0�e��H����^Q���B݂�W�`������y�H��jv��n۷���xT·>�F7�dK���<C���J,ʆ7��-��>D�夃3�y�D��ǆ\�ˢ�v��YkO$z��1��-�;�|-j6D4<��N�&�Q��Ů[ɗ�	��������:�%?A -+����0�진w�;�(�,x��I����넅�`��LO� 	c��7�$���i8!\�a*6����g]#���9��5oN��)&W�)��
�Fd��%6\�'�[�O�M=�jl��[�.�hDgqu����zBb��5_�`X�|��3vuRFE�L�z��+F�v,"姈��C�ǧhUg�C*1-���PQ���ƍ�TG���m��Q2��H_P����?�9��i͹���=���鷕�f���6ܩ�<R���Ľ$N)+,e-��ڠ������<Cu�M���G���`w�8��K�ڙ�tCb8=9R��]L{�9���دK��`ֲ����j�6�X�|So�6$m&~�����
��O�A�O��Y�|�ml�NS��o$�޾Zb{�bGܿi��g�'5#�� �d�T8�|-�$F@�x(.�u��W�͟��O��^�.�9Gm�f���!u��1��y��N��?(!"���l�r�%�1����ߜ8p:;�t� ���B���e��~Z!��x"�ѷd n�ǿ�5r	��i�����c�g��h͉X[~���Ku��L��]��|,t�U�C%I�^L=�ɏO=������������Կ��[�m͎�Y��̷h����Z�y(Ժ��\���'���f7U����W��`%��H��x�����d~���RM�j�E!7��C��
̾�v~��&�}2(u
�V
��$N#�b�\�\i"�f+e����h$>]�WJ\&���V_�d廆U�S�Kq��&����/I���~;����Վl�*++��H�Tj�qǹ,�׍����	�d�P(S�V��Z��{�|+(KƂ�ME������L�ۦ��(���9b@�Z�	؞`�� E�q��Vܟy���j=���rɲ�$���侀���^�E�7^��^�8��1Kh�~�9h�!ʺ�X��b%�Д�t��ࣥ������]Ǿ�k읾�h!�e`6�{Z�� $�7�Ԛ'9����fL�t��у�DBâ��| ����NP`��b ]�����n��'��u[:_�'.�o�~(5���9�Z?!�Rwn�<���qSp�.աi�^��g��t�^VfG���K	ޏ��a�S�����k�씦a���h���RKH�$��H�|��H�H���60<Qz4�޼�źxA���
:���sB�+^���f�A�a������1������Z����� X�FA�ͣ���?��H��=q�5p���-����[�������@{�p�3��J�|�N�["�v��GȤp_�7�#\
j���dWk&4JJ�x3
)t?��,��6���1s��(�C$��2�ǮFN�Z��ϟ�Ҧ��А�M8
V#%ר���ܑ`���w��*+?�@y1oX"�k�݃M*D���@D�N����L7�-�rm^Z�wb�0�>S$H���]�ϔs'f��A���Y���"��I�ϛh�+(C*�M=��@��}n�i�T��v��TN^4�-8Z�Ϳz�R��(gri���Dq�"�J�Mc�	Ě�f:+�a�EB�+I:�~�8n�XA����8������q< P�O��A�s,�8����Y���O�zX��Ȓ{\�>��r��H�	IJ��"Ά��;�	$c|���EO��Xݟ���a��_�m��bAmݜ��aũ�4��(�F��e�l�Wp�ȶU�06�����s�J�=�ű�`⢐����?����������c�iy��1��e��!��rˆ�)�}�z¡.�N�{ǿ��γV���_U�.�сv����_�κ�.@�<��:�4]]&�{3
n@�h�3���
�w�G���Qo�!n�.3�G7�!��j��	U9oߍy��}帖�<d���&�n��v=x�`���l#��b4�+t5�
��������d�%�7��{������h���ލek�>�{2��3��&���m�sqJk��`���s:RÔ��L� ����W<�_5M",w^� ��x��;�V�먀~���م����:N�jND�d�+G�}a9�A��]o�n�CX���萝?���&�NkU���m?�׃�A�����Բ�=��)��L0�"/�2�_������o�};L���b���7�"��R�(�ג:��G��K)2�H[�؆���Z�ƶ6�$����x�W%�&�Ggw"s�&=�R���O�/"4�{<�x~Y�j�Z0C>�M�,(J�}����$	����VҊZH������U�~E�N��H�ov�O�ߌ�yʫ��ӹ6�k�HY҅���BK����c�ͯ�����-w, ��P}������Q+��m���2/*�~_�}:�Ï�_��^1�1�0�X�IK!w|+�^P��.(.JX�t�~}�Z�����f�rf�i��_Y������I�n$;�C���� �;�B�qֹd�_����s@�)�5��q6|��XRD70u�"��}�gR8��s�u98꒦Óƣ�(1)����>�u�U2Jx1�6���1W��FR�&=�@�����}@�p�&���Ւ�.)�O��]�L>��?��2���>v������z8����1\`�z	����o��0��>$��^/���/����s�&�+�����	I���U�EU0(zb'��J��nJ3�r�Q�"�Lp�F"��i��(�(n���7y
�`�߬ƥ��؆Wt^F�7@O�Ed^"#7lo#J��Ѵ�L-�~J�\S��wF��f��I� tH�H��+����@�$�A]ew�i6�׷���� 0i���
K��~ʃ���Z�>
�J�"��i���B`�mT����!��LWS�\G	�e�fNtY�i\�6�4��4�(A�����~�5]�Y3�m	�c��q�%@#M{Oz���zP�8����hNo�IP%k@Z��p��O%`�YeyS|�h5߼X߲F��Q�vhk��)���tg�,)���~�a�wCf]��U6��� zŘk�P	ЧM��Єf�ϳ�3��j�.��h��w/��:����:�]�� ���@+�Eh�!���0vV��)3�c��b����d���S���0!e����}G�0���|�Y���vZ�3�t�߉+s�����ء|��H���si����Y�ie:������V�!����5d)�lx0�6�P�����hhG�gb`¦����"r�IC�B�}�����*CME����FaOK�����o1���*pC����.cWTu��S6�6��>Җ������9��ҁ�;���Α�1R{ю������~Zpf�)e[׀���H�h�[�T#�yt�5��Ң;D���e{��kT}q�ܮ�f�#�w	4k�f����x�սrB�U�l���nH�����N��F��U6Û����g4��R���)���]C����`%�ȴ��1e�����d,*�@T�%!��U R����T5d5(RW��yo������ʙnI|;�m@Aj���!��B}����]0[��	H��>����Ȋ�\��Q���f������DU�=C~���f���Y6���D��lH�W�����7RPx��c�7g�$�Z9�M`zl����z꿌I�H&p�P��܋�� �|9��^f�g�"I�U�=��U�%��]\EUqy�L>=>����: ������|�ʸ&|/������b�s���q{L�/ �����4��V\�J�w�#5xz�~G��w�*?�����7If�
������/`]����h.�#��3w['6��������QB@�O�O�T�_y�?���?�>�e�.�a�wH�I�="'NW���/��WP;*�3��S�S��ng�=5�?�}溺Z�VO��bߤ�oA�A���dߺb�J�F�"m����T���J�� �r��ĺ���.�tA�Y��RbI�
�'����Q*�K>����gGiZ�5O��9����yD��D0v�ܥPҨ��BU�u ��A/i|Y»!T㖀lC��^�d�82��Լ��=��_4�r��p}n?I>ܯ��0hv��oY���:�L��!��Wb�?�{�S���:b�u35��~�$�'OzO0��H9�]}Lr��$��O�I8�"������;��3��3d�
�R<L3�3�I;�ae[��~�X^��z��`����Oi���S/�,nW�ԏ_�m�|Vnbq��r�P���N��~��k�Z&ʮgsV�}���'��q�9x�~�)�G���S).�#[!|[����?��Lz�(��9�I�Z����k�F�W�=����8� y/�|aJ��jP������Ca�E���&�H��5WQ��濙���%�������X��O~)3�d}��Rnv�������b���1E'ׯ�lІ+�P����3VX/m}U]�z�t�I�I��VNM�,���07���&��TP�|SaDo��\Vd� U�1�6��?�م�e�������f�}����[�t-�K�v��}� =!!�����T���4�"������ ����H�r-���Ķ���>����\o衣��=�^Obl��h$|��;��!n�eK�s�5�45%jŹk�	�~.�Bo��L粠�Rqq�j�-��`<�':3��`��칐syY?E^����ä�y(��<0Jm���j�x�5��h-/Ym����Ɲ���O��N��u1�L��h���4|d�9_ ��֍ܥ�����,�?��ċjf4`���^�a_��i���z��k���m!����@yf��KcC}��Is��G_P��k�(����N!+SLz=���@fMBZ"�z��Wߺ��(���	:/_�S�1r�!�!ޘ�ވ��Q8�޶�H'�ႈgd�Ȃ-y�c7ʎ�{��)���ߩ�*�q���$Q�J��fSdh�y=%��le��l��*�k�2�@G�eݜ1�wvZ�%9�f@w���Ť`Y2�����������b.����]|��%/�=O��H�Q|�s,��,<���r�+�b���7f�D�з�Z�j�K�����!w67o:(��u_�`�O���W"�i"H.���Zg�9<. ��?�SD,�s1R����f&p�(-ߠ7�V*|�d�5*$�����x��n��s|MH�F�d$�(�-����{��� _�XcC��=�aO'�����k�gGU/:X�{��kb�izi�Ss�wj�iX���%cw�x��gG!��a�O�~�PMx��l��2tۙ�x�����ڔ����yʽ���ip��a��jU��	��.gGk�'�
=Ycn7��/G"=�>�m%������酧i��9N��RS	)̞HW�0�ќf��l3�|����ӬRļu%e�=J`��}�S�϶���������^��*��S�/���P��Jf�PZ��lA��/8�����Rp�>����	L<u>�S{�(���~�-j)̏�:�`1�?ҝ�,N���ݯ��k($���X����3E�
�:��3�u8R *kKW* ��R���[�W9U[q$�I��ۅS$2�co�?�5f�Cգ�-֊I�� וh���E�O�PzGf� [���pbwK\!¸���(f��2�P�S�y�f��lE	 ���2A^8o��j�-�>��	��-�xnl�Х/��"�l���()����!	���˖96ye��Wg��S&��c$=����s{\��2e�������ߢ(%f�Ȁ�{8hC��'����eb4��oa�U&�:k�� ���"Tg��������=|@�롛�f�wm��9���D������fe��ʼ�H�}��Inn���m&�����n2w.��2�06���q{�Z*zx��H:W+�_ ��s�b����z��AD����P�q%�jԣy��k.�\��R�����x8h\%d����8	�7���ғ����X�U�����ģ�U.��mK�ru8����~@�-H�*Vp��@��9�$������&t$������E 7 �w/�i�L�-\MU�JXUi%��]X>-�Bs*�6��t<`�	��YWwt&�yS��8u������*#����H�6�:ǡ�H:�J���b�5:a�#uo�S�M�q���Y#	ܐ�ftP�{PU��g=<g�ϼ�	UeA_�5澬pvB�AW�6�L��~{t�`G߾O��� QZY�ku�q�?|��m��I�J}}.f4�&���.�<������;��59c ��"�ۧ�����})��Ǽ�hUG�!ɵJ`U)q�S���NH�8��0�.��`"�97���X��w%tb[1=���@�`�
6��M�z��Ќ��}�Б�=Q����H:i�"������t:*�5�Bo���~a�!?��_��NM>&?�F�|@��q�oU(����[�� �K��j�1����*mΥ�0�)N�2���VY���O�=*���kmЊe��N&r(_F��d�M˛�zN��P��'��|&gLa[qH���QЬqpq���<t�1��O(�$��m�$��>� :&�s#a�xn���jRt���Ms�B�lH��Rqz[.���g�+��n���wb�&\�ִ®�eZ*d{�K��HV�ǩ��[	y%R��]v=bKSR����`F��������4l�B|�Oر�My��)mK��l��~I\B+e��y^;��}��h�et��V�,���R�xݣM�آ}c4��#���3ڠ�Q�5������s�7�Hȩ;F}7c���>���S����C�^��,B�C�7�HvM2�m a�*����&Z��|F�<-��o�C�5��%V�r�"p�"~��xy�5�����̭�I�ޜ�Y��.	��Ek��,��^�Ui�s�U�(��E~�h܉��+�Ib�h��OЎ�����i�� �nN�/�R[���!Z���p7�Ș�̮���9��/$\�VQ�N�����*B)�7)0"���V�}�8����M9{T�OA�ߩ-.�
����p��C!X8	�5�)Q'XX2߆�%���s"�7�4v:w���&�����d\��wP|@"��L�n͝��h� �����,m���+�tXKIt�)��ڣ�?�.*�]���	ij��0�7X�ҹ��
RU
�������N��;'@Gl��FUS���p:����`@�	����4 ch:�{��SaPv���g��An����J��E��3��'sgJ�
ި�)c9����i;��Pc�Jn��X�98>}�d;��G��g�P�%$�(`�^�e� ���h�|&}�~'׫rD���<e�Y�tT'��g8��V:�c-p��a30w�����՘$���:bw D)^��7��y�%d�/چ�m�c3��S�'W���J�&��vԍe7k�F��D�W�Oa�_��N-�em�^��0ҕ,k��6�Fʊ2���<E�O�V�l��žY̋�������BN� m��v�iD��gE���m�}YC��C�1��%#�B�Jk�^U�4��9���ӆT�+�?)W����b#�y^l��0IQm���$v��I�����zϧ�0���"�A��~��9 p!v�U�2�e��u�1��'	a1c��$z�ء@6΁ն`| 6�܂��J�4.g�2�`T�������cYe	|�b*���2E�V�j:�N��<3�O���R�$0K��x1���X�L|܉2���F��K����8�O�xiJ�*c(�կ��H����,(���|k�L�.��F"��Q��b_
��l!�N8EL���,���­TӰw.�����(2����8�{q4?2���0u ��u4���d�tѶ�Dn�j!-#y#�f�bL��Ga���p�7�>�.t�$�a������y�f#��=������Z�^i�{r�$P�f7� �2��ȌF=���m`ڶ��L���*s�w�C�}eO=����W��lm䷿�U�O>5Ԣ��ǘ9��w������]��vV|R@�a�.2)|6��0/��#�d}��M=��)
�bS�7ȁ��8��ap�e�b���{`qĶ�rX�KhѪ/t��|Vr퇇�9L<d���o���&o�=��A6cJH`) \�O����ޅ c�K/I��'�K���[�U4;R�Y(����r����(�J�_������X�E�r���U5^�4��y��n�Yz�m���f^�δ�|�|dK��(}Tk+���,�k��#�ߤg�Ef��р$c�PV����l�;��"M\Y�"t��Z$<֑��,CH:�a��y�c�# ��U�ine�gM�XƇR��Ӿ�`eh�[�u)��v�?�0q5Y�Q���
؃�3;�+k�%���W�ЅD=
�2S������G������*8?ǍU�6j4���ʭ��F�epéT���r����6���q�ILwf��i���D��u��>?�7Cz'�~P-��������z)d��s}�&� ��#fe0ba��$��.B�y� ܠ�r@G`����q_��������u��s
��T��yV�cOZj�X"S���1uȸ&��=�Xwc��l��F��\��S��=��ǹw�J�@yb~�� ��0�~�.�v���_C�H�9��)��(��f���B��_�,oY��j�t��Y��{Ym$nx�sz���c��-��#Bì���͞�1��S����7*Lf������:'��{IҎC�P��@:����v�5��>�ؕf�b�A��/��&M_�s��:9��?�`P�S0.�FX�4�u�%�ÁcsK���=�'��^�R(�����tfa)5Eq�
�$Z�-��^��m�r�y��ǲt���164���D�����|S{zϢQ1_D�G���bè���XdMj$�v�٫%^pS�f��B�k��T��q ����N_m��0fw��u�n��u9۴҄���ހ/DH1�s�B�b�g��̂���&✝+v�|�wTD�@��Th^������h�
��E�p�3�r�W{�#�=�Y�H���Ȩ��c��'�%Iy²c&3����^4"b�ꮇZ���\�'��Ǡ$�=˔�P����,�=�Q�7�L
��g���*�0���Z�Q
y��5r�oK������+�gn�����8|6+�{�x�|+S���&��f�zp�Z/1}�2!���t�wE%��R1S>d�%���dM!���`�i���X=�����n����Rۏ�}$AY�X���[W>qh��.W�=Z�����������Ů^D���)~�n�c�+�~�c�EP����P�K���B���0�����Xv�;	�s�߼�J&���c��#�n���Ƹ��al��`,?l6��1^��#�'M�������n���Ùj�?e� �b3�q�ՉsN�`�N�	=U�S���{��Џ��I��R *�>˧�&c'�j�F�7`,�J'�)뿻���U}���b�^�p׵����<t��&���`1
�ǽ�=��G?����(���I�]oBo����v��~�'7�¦Ho�gS�5�h��	����28g�B�魴�Q��Rws@
�	w�ȯ���f5{_��Ƒ8��9�&_Ե��H��o`����<�mj��%+V���¹f�=�l�άa��p\��d^ٸʺ���*��i�d�±y9 ��u6SY͇��`C��t�?z�
��[B����~���LU��@p�ųѝ
'���6�
0�����U.�w���٧������C}�
ׇpS��6��t��#��,?�	�ѥU'��8T �C!�2o�?ނ$�\w�5]������Tf�]��Hi5�1)��$��,�W
�馽���������Zn�`K����������c)X�u��[��t_ϒ8o}�������̴��{�(|Jidn+�P='�����xd�Wx-/�d2M�U�H�0����ȁ`TL��|�"ULA�������1�C�y�ݯ@Z\Я��|S6t�f�.�LMP����}S�g����������;;x�u�>�>�8MNR�����	�8=����Ȟ��������lP�9�.ʞ�F�ŊLIRn&�Fr~X=v(��pڂ|��KRC�v>NTݱ*d��IM7��8���������$8;ۘ��0�������:�I��95x��!H=�\p?{sY�;�eq��DϯET��ÑUy��)p6��ר���wKڹ�K>�w2�).��S7�/�o[��ј��;�%��f��b��o��q��_��G)>�"+(�aq;-���"<�L8f�����䢧���*ヾc�Jը���N��ʓ�<�_�2&���b�*^����l ���=yf���X�h����bB���cs� w��d���C*�Ô�zB)/s���.CZPJ�FҦ0T�t��g��Էhtyz�@�H�빡�*>�E�.Kl��׊��Sh��?)?]�`��������k���2j��z��,��R�K��D�m���-r�ϝ��	婭5�')��
�r�]���D�j{�8���5���cਙ�t_t����\��*s�	�R����f�c���Eu�'v��t���:
Ͱiw�x���:a*cտ�Yg�.�e�G2�|F�֒�m�n�v$��:[0&�Y�]1e{44�֚�1���[���:��Þk���f��Q��G%���t[�ؿ�PeG^�]����U�6d�E�F_^v���kI�;�_����f"u2���L��+3v�O$(�i�T����Ό+��qN�WV�w��m�1=+s_O�V�F(�������ɷ�QKDYy�3C���T��i*#�溒��dl����l.��-@��"ͫu��r�|hW�����݃g��?��i�8f�ݟ������;
����N�&�9�$Z�zK�-/g�y�⹎ù� /�B�<w��tK8GcT��я/aSQ1�r?G��(�O�$x�8f�NW��l�3��}��Q��2��E�g,k{f���#��f�-����w�:���^,���_����dQf�9�8-�OrV�'�h� ,[�ȐT��B��A
�_s˂axm �܃�k\���[�tV)6��{�t�:jQ��Dd��AM��&��&n��p�o�6����Sc�j��BΗ�P���Xq�k�?�[V;[�1@�Ss�h܍�ud�8Aس��WTm\�?�`��S�;,���|2��N��8"ת�߉ϲy4$M���ϩ�<���o��ɔ��B��y��x{f�{��l�N�sH�<�Дd0[3�v�A��X4�'د*h b|�컳�j3�˶��	����0%�e�b��e��?zX�ߝ�-u?��V���{���d��d��e��{̇>�NQ�F=�����yZ�߅0L�Ou�*g���+g��F�	W��T�Ӌ4��֓�1c+���=��t�B����{�=�����ꒁ=x�]�&9�̟>�UL��a�4R��	�Wb]�#&���ĸ^�9pBԃ�B!�}��׳�y��H�S�CЍ�J�\��^��h�5N�)H�'���q�&�cR����%�O��nl����fƹ�&�qBϯ�[�MS2�t�pk�ؠ��u�Ѭ%�=b��d��E�ǭ���;��p_��?ǦQ�q1���NZf��7�t�Ӎ�7I�W*���>(^�uTiA�î���)�	��kN��I���� a�p�H�7o����>��5+FV��A]Ԃ2q��n0(�Ӆ&	bK~����V9G�?%���v}̧#6��$�&�5c�+R��T�m9�(��Q��۽�`XJ)�&޶��X��Z��I�)N���m��U|_2��x ��׫i2��%����2?���_a9$cB�eg�	\�v� ;�l��/�~��,J�V�I��Y��s�JN�,!~sȿ��S�_".Q]�g�ȲKR����eh�	�%dQT��˞ .��>&-�l-T�Vs;!q�4eT�p��<���Y�C 1�f*+[���~?����<�Hiry2�5Ǯ:�|��"'��z��",�[� 5;0�C�u*1Bb�8-�[���!��6��vB�R�B����[דX�C o)�,/��'���7'u����K%��S$�t�"��st�hR�nΣ�`���
	E�&S�AI�_F�$��>w����G��9��nb�7ږ���F���"wr'yE�_j�qH�f ��Ա�j'2[4��m���s�U �c��a�H��S�j�}[3�S�3�����������?aE�ޅ�&4�i�\	�4��RZ~vj��|a� �E%�(���Ho��,~�=��D[�;�}�-�� t�h���QA
��Y�����Fd>b�J�Ne�>�Fځb)ޫA��C�R���ࠥ�C�����χ�=�G-rH���������Q�����%%Az�H��Qv��`DR��-�~��[�9��E/�&O�f�������a%��K�=K��E-��S�ç��nT2Ԕ'+�����$��	3]�&EhA?X�:�࿚�4���v�'�^��1��wa�$C>����|K'�y�"���V!�GU�#��z{�A��b1}���p\"�2fa�6W�{��`�&s{��J[�a�2M�Z����p7?��z�x�/�mW1��{�xM���|H5[����x��������'�����hm{���~0��P�O�"ތ@��S?	~�O��I��C��%sX����菷����atӿ*5�މb`.����'�o�{��1urr�t�!W&�d��YO��ѝ}]�����.����J�D�C�@�s��"+=�8���+( f窤RV�B�UfP�i�k���j�!)� �
��=uˈο�5�_�����PFD4�Kqa7s���D�P�!��f��!Ҙ��4=r�.�퟽��Ub�q	 ���̹7����d�aV�ks��ǯ��hI�Z-Z]d:�����0�g�Φ{�㡺�C�߭z�>&'Y��l'��V.�5���6,�`�xo-����5��4�a|o2�( ��6����ϼ�W��fhk���uoǨ����L�a��������$=3[���'8�����#ߊw�$W�u_Wy��xf��#Q^��E^z�}G�#i��Ə5��I��	�7�y4u�k[��?"
���7���$4w�G���Ǐ�.����$7n��"��d?��4���TH�=���b����6�ܩ�~^�F�T�x�L�X(ŇO�ⱕ	�I�W^�F�T6yEQ�� �E�bq���\�r�Ù�_��,S���R�S�Ǚ��Y�$!������T5[��+S�>Z~P�������b���o`�I��}��J��+�8-��q6���#��إh�%8�*O��?�JC�]�%���nǙ�5�1iƩ��Zp����L�K��BJ,T���ݺ��(�3��6u��*[�h2��~/��F���H��ǘG�;W�!.kʜ��X��(��K�$��$r%Gar�8��X�z]dyr��M�i<�����ۗ�uq��-@@뛁n����R c+N������%R�%�k�"/�-����vZ�v���`�Uo ��Δ|$�K,E�0���$�@��B.�/�3�3�nF����WO�o�%��S� �1�<؟��6�����襼|�d�RR�:� 	'"�Ôލ	yk�+xk}�ܔ��q�6[H�ʬ�2�%�4��5����r}������	�F&XF�'|kCаA��{��e/6�=�٨�&	��p�"_�>�,FܿJOԬ	M홀(~bL��r\��l�l��i�L=m��cJ-~B��(o��<(��&\���吗��H��a�،g��b��p��3HKl�jux�ǌ��c�����0sNwr��||�6��ъ�*��L�a�Q�Xw�=�m�ǵ_���xy�@,~��j��ǫ���[�O������2��!I�%g����J�fYu͞]W\|EWջ�,��h:�J��j�!$�2SQ����hY�ħ��4@�"������=��QJp@ő�}�����m��+t��T��;����R�1ZW;�t5�ԣ��W����|
�废�y������Oeƥ���:U�{!R�ˈ��Ӿ�y����-�$�M h�RE8������,��x^�zi�6�-�b4�]���K�xչ�I���p��&�&l�#�>��@p+a$��!�O�&�jk9��j��G��kp�"���2z9��||JY4�x�bt�B��k�U���/�«:�
8R�H�Av,q�C�Mk��xw���v��k��0�SZcn8��M���i�ҏ��䗄�����tع�&<��u�py��g���.*��X<����#�����)��Y��-$U��fC`�P��eKU�!&��g�Yv'���&�+������5��h�Wޣ�0�yEF{eH��i��]�T��
(���Tz��ж�#p?;��p�h��Hu5�8��a�"��]�_���FCC.�i�5��˹F����4ʾ_�N�t=����O"A�,4�Ҵ�g�kt"O-F����&8|��o�J�Kmt:���3饅־�����������v������P��A��Ih7��؀
�2"�!텠�_Vnަ�-O�|�ζGo�-P��v�O�Z�p�n�_�����f~�� �cS��K�EG��^|	��b���fAҕd��}�W�V:Fw�F�I�E�Nlt+���R���R�����.M��:����#t�����@�����{�d�d�f�t�q�p��۸�]�ů�e®���=�+O;?S�0�<�+�y���XE\0v����s�͟� �ږ/��P7�C���� ~2ߥ3!딭�oC��x�;���Y��ˍ^���vw�ջ?���BF� ���s,|��C��%��;�J%�kX!	�tPC݉vPx���If:�#���Ӧ��G���A��~��
���\4��hO�F]. /�w��3vN�;`��F�4� ���Y=����XO�rKC�ٝ����/agZB*��
��`��ѯ�6	���U4L��!�w�L���J/�w��ED^:L��p��0�
L��[����=:nN^�KXSj���8��V&���[�w�a�}���7yΪȡ���=%�\��!��0S7�m�MvUT�5��!q���t�R�j�ԍ��W�4�5�������>K�V�Jn�7�䐪'UC�nɾ�͠e�V��>����x�m��Uc�Du����Â�Mn�B�� f��)��*Jy���b�"KSt���n�M�AM��@��4p;�ڃ�������F?���ɣ���Q�ԋC����..�2����"�G���v��]�y��狾�l�n����y+��~t�O�a�4ӑ�(�o�,˷>�v0��'%���n�l�՟�������l7��5��Ǣ�ƖS�2JHM��]�+��j-�$�O�^�T�U[ق�@��lx���1�Ru�J��~9��F�,�8E�=�ź��lZXfd�2p�
�o����!Q���޽5� ՗��g�B}�`�P� [�<,͛'���*�����,�ZW�yB_�Hto�;�Z�St�3�i>�k�]bXJ}	 :^���VS��ʚ4GD|�G(�m�:B}�L��Vuź�v](�!/"F_����%�����x� 01`���	�/��9�J^ɩUb�G\�;�?�k1�y�����Q�6twi�N�*#�P�yE���mG�,9&����Y��C<K�M�q'���о�4b�)���҈�ø5Է��M(��o�.[��fV2D�̸��Z� '���J�戛>l�yA����.XYw�݈��gu�jM�+d�h��d�XC@�1\׺w��]��R��i$��y?�ߧ��t{:���[�Q���M�ug������>����R�#�*�\z�9�e�K��Y������Fygz�f��dP���l���C�X��w�Z�,�,���ٰ�^X�5���[k;s��x�U'�<:�|�ϯk�fd~�]V4��!�M�uv)����y�B&I�`����	��m���+!n}xo��Ͽ\���$"�ï�����jt�p�V��xJ��4t�q�y��{G�������Qr71�0�SX�o]�5vO��%��j�_9ZL�9�Λ,�"Qm,��kj�ߣ�z4��N�y'��|T*�z���,Ŧ�u��m'�o���V�8x�S��Ěj��11�|@P0���M_nt�o�s/��L��FSw��+Ϝ����=�ʶ�X�`5}���I�O���͵z��O��_�,`ߦ'��EO�p�Vc���3>�YG��9,�;���V\�o����n���>G�S_�Qr�Q}d������5Ucj;��� � �]W,�o�d��?!"��v�;����0fgQLX��u���q �\<��(�h⨗�2�x��Ƿ���lQ�T��w���-�ߧ�������]��)���<{5���5u�4��]s0�A�L�Ӎ�)@t�ݸ�/f�y -�ey"�l#;>������ʢ�cy y�1�.!KRͽ�n����.�:�Nd`�����ލ+۪�z�B�.	-	�z���	�	��X�Y��v��Q�uw؇.�Y��9�乷�/�S��r��X�`���ZT�����4�BE��
Ԟ�U�	E��~
�R��2������S�]�P�� �z��&A�6p�K���1�Q�H�%j���ֲ�*�m��5����غ���m��7�oǤ���:�[�_#&D����B��rm"��@H+M��l�_�EOc�Ĳ��V�f7��iKJ�(���B2l�eV��a�no=��T�zʐ��'3 ����ۄvO�뙾�M����@��u0!�:�5�C��<i�}Ŕ������c1�ϖ)T+��G~I�JE˔�"v 0y����'�A��^s^�@7n�hD�_��u,	r�d0?�1 %2��~#��̣�>d��5t�'�i6�S����(G����I� ��ŗȩ
�s�2=����a=G���U���>_זxL"�b.����O����$����7�>F�m8k�e��F��#|�6s��	�L���GYE"��<��ܻ��%��g��o�"J�������[@�4�:.!���xc�ň@}��*ݯej��� <	�!~t��E4mj-��Gv4<�3R]"jEv29,�n�&ҵ�,�;	8q��$$��t�� �v���.�g4�����g����*�H%��Ċ���ś�(�]y��4��90ܬ���=��K̘l���鉭�fQ4q����`�|\�WC�k_��{Oc�goCΐ-/��mfh+�E�]�UOR��=UNy`p�
c�s��U��i�F33�:J����.�ӏ��ԏ�t#�4��f������I]����k(�]�v>��Db�u��-�vp`*Vd	�������Cz�n��ȩ
6f���
�>�)��{Ǫ*OtP[(V��Z���Ym�@�F��I���3K�2��!�޽&=�ʞc�F����ҽ��֞X�xuB1J�H�S���PbK��c�R⅊nf��f0�r6�v˧YO�N	"٥c�Z���#�v�|B4�62�v5���PL0�^{z��T�1n�E����A��_������Q����(��/�	@4�c~�Qmsn˃�9&%��O/��w�_��7p-���5����SK��t����J@j�h�<�5�[9c�^xƦ\�,����eЮDrKn�O�i@M7$S�-i���u�8�V0�{�O��j�r|��.�Ũ9-�$���$*��aD�3Sٌ��Q{�$��w�������3hBC����fU��s󿪷��F�vi���J�q4Ǒʥ�5�H�:����cg�ڸx��ȥ�,ӫ�L>��CAiQ�@�v��|�{�$�WP���0�*������'�F����@oܩ���\J>�s١im�n��kf n�<��j�U��ݚ:4@F\�?�	Q�T�䆀Mo�Fm���E+����0]e�ٵ�L��L���,zGw�MF �������r�����-�XIW�Kŵ�`��R�+��������ͣ�����ȼ�+���[|0&�� ��7̯-,�&T�	����p;������q�ꋙ-��	�Y��8���N�U��l�=�gBؑ��D WJ�k�nʆ� �hI�Ǖ�aH��\
���0L�v�!QfL�\pm��rQu�>�\���~�Atp���j�[�>x����o�����^�B��+wQ����0n��.4okr4�����(R����{1���E������y.�3w՞��v5ߨ������kB�= �2:���ƥ���u�>�F�	������l6j�$�3����~�x � -o%A�������v ��j���j�m���D��RmO�[07	�@�z�F)� .W���{Z��E�r��y���)�>g�v�w�!a��n��L�ة��eI�4G�$[اt�i�|��e3_o��b������o7����_�� ��c0:9�Ԑ8M5�ly�k[����4 t����� G�s�>|��w���+��w��ѓ'"�@�5R>��O�s
&w������"���2A�`(�B0T�N� o�$�~���&�D�V��<b�yP1Cq����Sr�,��jzt�net'���'�;�
��D��C�g
��LʒbƧ4�[��R-^�����ݤB����(�P�s��g53���42�d"�1&A']�Wz�[G[�]��uxc�pQ��g����]�D�+�f��T�K3�@�f�C�� ���P������ߡe	�i����G�/���gta�P)<�����b��<�r���ѲE��1����!��B͡�/�>퍣6�aՉ��c�#b� �M�'N:�m*�K�6s=�v�A��hq*!'
��e�g��H�k�{Qa9f<!SϨ�6v�r,����R��u$�`��X�/�7hZ���r��R��<��E�����Z��N�R�W��s�����?7D��
�.yER�T�/���A��>�sA�Ǭ�S��9����}�7;ˠ�@� �tq�>hə��f���nV� 9j�A-+�ޫ@�����\\.�"��A:�����1k�u$9y�m@���x������z�^��9�X b��r��܄�q�����i�v�����73��v����;].�FHx9��ҵz}��F8k7_��O�����Y��R�ʚ�|!Q�n��|6�~{�ه�9j]�r`�CRJxW�t	T��P�U�2-�H]8~n�+���Η��/���+^e�
��Cq��j%�J���x��M�O��Id�������i�������>@I� ;�\t%:�,Y��6}��Û�����YexA��G���-���f�F�Ί��wi�+H��2)U���s�,.4�At���~�����i_'\���wT�s�CX0�M�(�m��׾V�a�<?����kGP�ý��﹁��AE=J0�HӸ{����蘤��#:��F��YgI��
�$^L#Zg 콗{i�z�Ay�"��yr��D�����Y��m2mZ���iy�����Hڸi!�^m8k�z�!�O��gc@��Di������Kt &m �QI����/�?��{ڞ�5�~�jD����ESD��o����#��vH�<�R�i��R���v1��Q±�p��3	��G/o�+X0 ��%%��ȏ�`o��/b�-L�e�k�d7��= FP�e}m�i�2���&j���ۤA��3:�/�g�9
�nB�Ul���y�c���Q2�챘��F;j��ru|���D��ś��
�M�
Q+n�a�0�A��'��5����:���ޗbu׼�i����Չ�ELm_F<�Bw>S���V�V���U]��9]o,T,=ff�ESy%F��{)�����~���,�O\���뻫Zl��h��/W ����*������p�hj+��IV��!mL���)��S�<n��rI�u�O �2�{l��V�3�X�%�V�C2xaDT��u�v���+ꏮR#ʹb���J�kM$���ű�M�a��p�(Cb{�Te��
F�YW�;РnE��}�ڹ���4�`��p�\�+̉0'��	�t�5�*$[��?n��M}�\�����m6�Ѭ�l�[��A�0B��%~_�ۆ�L4�(a`'�$p���NK�.|��O��Q-l��3Ǒ� L��n�zݓ��	�~z�Sݻ��� ��X�P�J����-����.nO\�m:��L�:���tQc�[�U,�>J��)�Ӱ���[�B���+�24�;�j/�*�?l�\��B�E���ZXh��{�>���!�0d2��-�7T3ڄ`���Ev�0z����u��l{�]��bz�c�a��"��{	[���{i�[6��z�Ï���
$���|RȈ�:~l�2]o����X���oT;��0�?NQ`h6?��@���f�䭼�b��{��n��������-�u�`�O]�B����:"A��-�e���P�y��v��]Z�����E^RG�Y��W$+��A��cH���`U��{�z���ʧo��K���Z-CL� ��;r~v��HG�T㻌 �G<f6�<�_�@�w��z����ǮXdgPqC�g[� B���v�/9MWK���oE7C�z��g��rrc����ۂ��;A�%�>U����fP�z����	$E�E���l��_4��b�<y����J����ì��^$�4�|�̘���:=���^��� �P��kL�W�D�?�Ǻ��2�v�0��, *���Hm"Q�ar��v�S����E�	ř^e+AL
n��k�F��^�^����W���S����?|��|}l���a��֣.4յHGq�U�(-�oI�����Pm�Ƒ�����B?��u��K�i-/���a8��9J��� T�c��#�B1���� ��`pV�w@Y:2�ɀ�`�ۯo
DI���q��v�YQ�����t��vƾό�0̔˚2�C��p���"F��a�fB�V��Y�r��O_�A����?������L ��Ω:�+{{��nD\N�*�
#�h���6�:	̉����"�F)�)��z�PyU��_�{0c_�2"9���@�8���EpM�G��GN�\�{Ǘ+zKt~�a�mᑷ�"�nk��/2E''�`$�dD	k�����)�%bB�b�����Ktf=��I�a5���G��t0���͸� �Wj�"�y�6$U�t���뻄c���Rſ,6��6�ok���&(��i�8�)���+�����2�b��0ߘx͋�-e�P�4~���*&ǖ�T�;��i�Gj_]�?c�ky�ӓ�6�S�#d��m�J��(�k��\�3����dc!ʤ����4�J�~qݼRoH:uo0�Ra��'�d�|z��Y�{hˏ�oO����L���� @s)z�	հU䢢���^%+��q�W���X���(����}�	��O!X�hO��bn5�"��S�, �*��MR�̛g�;�<B�
�m���� j��.��:�D�h�?ھG;�@��M�ƅ,�"����=�s����W�o=�������ɭhN��S5e��;�.�~8C=w~d@sO���1�R���{ �}7�r(V���/7}�V5�\cPQ�
֖_=��FP{FE=J�	�8��a�E��6����
��~G���E�5��]�ۘ��������j��2�,	L�U��MX��ֿ:%��#+S�ÏU�i��oJ;��޿}|� �dN�r�ۜz�����;�g���̼�>O�2$���ًP���̉Y�'��$7��V*&Y�i�ٟ����pVl���Y��ﳊ'RBL��GyD>2-y&�l�Y�*������Q̇�A�d�[Y͛�'��qTS`��
k����`R�\{��{�e�ގ��#�?��Ͳ�~{��앃Q�"�jٲ��>0\�o,*诃J�`�Q���tZ斈�{\��ڙ/w��B��G-�+7���a|$Z���~g�[m�Lr�,mމ��Ue��)��)iɔ��P����đ�w���?�PX���Щ����,��I�O�{,K�΢34��{�)T�k-w���%�v�����6ˋ���L2��#I��%|�H#��so1�kk	����}AbT�34������W��m�m�����k�AQe�Mf�l<����:��íCf�RSN
�`�uѮ���u���逡.�S�ՏQ��0��������~ �i�,��v�Z����R�MMd�����22�W]]��$S��� >q��ψɄ�K7��U�3��F��-n�zΧ�N���.�9�[lDt������wuD�Fq��r��F��_Zr�_��*��FM��X� 5���
{��{��],��r@;�f���_o��|"�u��a��X�"s�����Nzb��"`4]�g[��cO�'�z��p�^�
׃�s��x��e*��!a��jL&�����=翯=�����2CA�v�����)���<1�M��8��.)^�䣭ӯ�ӓ����︌��K���Q�ծ+H5�:ǃ���	�����,�^�f�(��<"�YͭD�]�N�o��<��.�PX}Jkk���D �F��y�d�T�R�^O�M��7���0u�+%G������2���V5����Wrl��5��>'	P�ciL\Y_�a��e�� <�Ù��3{����#0�p��ꫂ߷m�|ێ/ظ?�̷/��C	v�6�V�f����L)�bd���8xqc�x�� ���NL>-x6��Vs�]-�X�׍���9�s�Ӵ�mi��/��:�%���6�fpC�n*F���'��w�g#�'Ӭ�J�(?�_p��|�m�i�sAD����R3�E�b���g�b��T!�#L@2x�I%��̰���,�#I��
��c�f��$��j*����:9cJ;��������$������t��ezJc��=k�^+����	2��D�aº�_W�&	��5�kW��ˊ#��$+}���W��M�c�=K��v���8u�m�8�>���E`�2xx�>�
Ex�B]g]R"U�����f����ι��~�=Hu�B�
���Ѣ<��x�?�����c�B�&��Oַ�Hp���͏*�V�2B,�M�< o��P`G/20��d�ƀM���i�Bk�cӕq.$D�W�Տ+D����yА�k�ؤL�w3�k�$q�Wz�/��-+��(8����S@���/�	J� �(4�$��O�*	t��Y�)�e|�-�x���8�7�)}̛^�5��+�U:�f@W��m�*u�v;;~S�~X=Բ�
��D:B)�繲q�.���!�;���.^��e ��� ��>�Pb�H�"��}����/�7 u���&��l1}��Lݸ&���7-I�$6S�17������l�Q��;�F�G_G<2� �����}�96y��i�#b��]Bn��r𡭑�G�H��ࡷs;�'�e��A�c�/۠���Y/*���_2~�v���)ۘ�ŗ(\Ce�#t%P �����R�f=�j������\�=�W�����e�4@&����F����c�z "YIS�SZ�0X\�Ò+���u�����%n3�j��7Z������g�*�� �e1�X�=n��������y@�����=7,	+]��[�$�`Op�w[�9�Q�v�A<�5�T�xE��P����(
�ı�ۊ��6A�S1%}�G[�a��t�7�Z��ˆ�]U�k��C{ز�Yxd�C��V�����fdK���`���S���4�sÚ�șd��%��aYg�]X���Tҥ��Ʊq���f��b�Khc"�1�.T��2�����Oj�1
;X�pV8��sb�n����������԰����z�[X)oK�S��%-�8�2�bLs�/�F�X�QB��(���QN���x�]�eA]��Z�����&BG��r,�Ws4��Dr�lD��y��Q��6�:�+[�\��Η0��)Dpbǋ7bxu89�y9��@r����>J`�L�.6ѝ��k<&����{�E�Y��a����H��:�XTD����c^�	��[�$���̾�͑s��M�&�^�r��y\ݱ��U4��A�Ņc����t��n�uO�8ٽ�Kg�Q����x�MRlA 
�p��~��W$�}�:F�'�jܩTI�}E�,>kS�.YHcHA.)�=uPf����`)}��g�=�٘-�LGU�v��tM���-���J��iہ~su�7{�E�pݾ_��׋�A/-�H5�Τe+x\�2%�؟���q�SV���)@���C�}P@ 1jf��P$ɹX�;8�@�!D*�Nm�u�'�M�-�Ѵ�j��Ǚ_DfvR���G؞&�3>�AX%�Xm�Y��S*<���榲�p��1�)��|@�J��,-���>ϒX�6�{�b;"���:���� �Ct>A�yӾ�ޢ'7��I>�
]l:��:�uQ'��f����>��?����!"����u��j����H8�y~����0���EF��7�X�V��|����IE��A�X���wF���N���g+��9�;�+P���B�R�۴dp�NR�Т��V���*TD<&�w����b����fw�4�O��;�I#�Ϻu	�+���2��	��%U(��f.J�1W?�YJE߿����|�v���K��&������+S����ƛ�-!x�r����F���3E��Q�y�^I����v�ig�6ϸ�/��XY��Dw�+�*��2��>������j�y����ԗj��yy&u�R�f$#�vM�~��*l���P��ޔɈ�8�tr�?LU���ɖ����vB"3i�5���|�Q�h�8��sqg�h����}����p)��eH�Y�ۗB5�����xsl���7���P�����W���e1�y��
��y�乒��M����Xe���b%����N~H]�T2���nl�����eP��:��Q4�9Ѿ�H镫�����%�H���hQ��l�6"�0�qN��+�JP�Mݟ*����7�aʚ-ạ=��@�"-������`����Aqڝ��i����AGe�Nus�PE��@�6/�p��$��~i�S�6�v����&���������j�hJ�u�����,U��� �e�������[�wa������d.�u����z��MN���a;�	%�չ���*�0X�8v�ݥ�
����5(]���U!#��jJ�!��=��a"w{W��%�,�s��p,nDA��&'��c�����g5�w�+�`h������3�3���0�诵��`���5�y?h?"AB0����e�;9K;@�v~�=XI�Ҫ��+⺭ g&����8�S�2��q�
tȹa�zP�^�o�1��8��h��y���nϻ�j�WƲ$�����s���*�y�IG����ē�k���I�����y����qVs ������3?��:Ա�WaQ���ēІY[��k�����w<��UG�%�	s��JH����YӲgY�$Cd�`ڌ��1��̅ ��!�KO����uZ�C�lV�ae�z�6E���y� ��:�TR�^׾�eÂ�.�B����&q`�:u�5B9�@[#Iw�"1s-�����n�X<ƄH̷�@�E��wSM�gNQ�0����9����:������^�ͷ�2� �uyOY��{�S	���Z��0�z���^��t�`���*���מ]ڢ�rd~K04�Cj���O1*�v�1�L����N.%(��OM��d=���S$C���aP ~$pF��@���-������z�?�����⹢��Y�ے8N��ϰ�����
�2�Db`2�ظ(!_�<�-��'�ZQ���]��J(�	��Z��?Mj��[Dx֝ʱ�%/R�? �m���B�^ �B ���n�
6������Zm�t�[C=��#M���!���ه�a��r�a*���5v��OV��I@��ۑ��1`��aQ�,\-���4!�_�1�γ��_�w����B�6�w�~l;�>�h����Zg�q���KF+��='X�'T���/�t�;�a �M����	#�<���	��z� �֊���۳�s���z��5�!ݮ������ʅ�"��2vއ���%�D:y6�tVg����`�+��CD�G�ߞ--P�|(�{_��/D31v�¹n�c[f^#��.ΉU�QJ�t���ٹ�5s9e�pz����C)S�S*��"���[b��� �0P	D��6������Y�b
|���a�UVM��+��)dG�����3�<զ��7��QC�g��t>��֔m�J/��s����ߎ�uNª���� 3̹���F��S�G>.�����zm$D�S'CI>ߪ�}�ʇ�2~�z�a>,%y�	���:0��4�ΧD�%Q@ ��Y�3��ڀ�A�Lj_��u�l��SF=�Q�e�!!�v��J�N#���*jƲ��|����O�[����U4��[,BM�|�a☔m�2I��Uу��M�2�_Ѳk�B��
pa��+�ǵ���8[�'�|=<sF��nԟ%]��?����(�93e�YC'd�^����C�"aX��������#D�0��Ν��K,�uJ[���%}g�V��+{;�P}[y�Fv�ɉ-z��q���?�m%V*GY�b�{ǝ�+�Z�V:$R�oH$�
n,������A"ذU�q>Sdo��n���^��ō�B�������R��[��dr�jC�9���c��2����j}��<�T�1�?P̎������BA�L<A��o���3vٍŊ���!rD��]u�9	)wj�Ȩ-pӥρ4�0��8���dejT�"�\<�L���g��6i�˶1���!�ćy�JkR!IϊŅh�;��'���TaX���+�8��ĨD�M�1�%J����y3��������!�|>����Jʆ�F�M�r�'�����D@&=Ǧ����"�{�����k�iP��w'�Go�d�_q$2��!%�N�gV�/H����<��0����wY�ޤ�~�̐�7�kFwk��G�,l27:��S�c��C[�E@�X���ݓڞ�{@S�݈rv���$��+�ؼ���%�Q��{��@� �r�mn���&g�Aܦ	�d��� [�����u[����Fࠎw0��T����}UWt�Z?g$���88�OX�fU�d���h��k8�ƕ��E�)h�����Z����|N�ר��`���pcC"�ho�F��;7�8  �/H��J�y�w��{k�$L���{	� ��;oӄئ=��ԕ�����}(�:�[�D�j�hw`�Rqx8a��w%�L+�:�èp`�_Sұ���ewP�aj4�����3�C�<�~V�z@���v\�Z�ޔ��K�K�8�8�Vh&���1��n`4qL	�^��^D	�T��Y� �k�kk�3ʹb��S�+��z�����z'�����������w��zٷ�
t�� M�VȾFy�}���0�p�� |�d�q�ұb̚�>��q�ǃ�*�?�x�	�BCF�k,wp_pB˶ƞ H����y/��?S�[m�c�U�A]!^�M���	Y>�������8u!�B�Ҥ�7a29-�"��[�୊k�Z����3�Ӌzs���0��p��f��䢆�x)��)�S6t�3d� /�Uҿ_Z��#�65��$O+R �Y�P���Z&q0~A�Z�yhq���<{{:�� )
���9�pHl�Uq������:������K{����ye���PVUd�i�=�K>��bZ��Z^s�(�Oy�ߎ��9�XX� �oZ����Z�[� ��8��<�-�U�J��E�DCd�w���rLQT�ˉ��~��y�r�����ϝ�s�Wn,��(lx�!��h�_�����L��/�Bk���z7�����Nãn4Ctr)�����~%Qw!tXB�Wk��9��,�0M��h�\XR�}��Z�4�ϜuD�6b�� /%4Aτ��$�
/���D���n��� �����k��\8m����0x'�#�B�s��Z�@��n	^♘�um�x�x�8�OMԓ���Mn�^St8����B ��a>K!�n5�l�A!��@���Ɍ��Vc�����OW���.�?Qpׇj�ؽY=��� �0;�t�x��Qv[��0�T�q_����`Eh\Mspp�F�x�*Wc�GZ*�����`����B�XԎ���Oɩ�|5ydI�$�xj��5<�A��(' �n����14��_�*-i�`��3%��`B=��88$�~	@Gç̰�*<9����J��eN�H����i�Ȧe�gc-��H1����}M��G�ܯ�h�VL���~8�O��	f�N �F�_kNV�t78���O�O�Vé��aOڻĄ N�;HUS��BpM�UN"U�c��/S\�Z|�
w¡$)��AC˺�������,	��*�m�+L��d� �����vIď��~�H���;�@���$_N"�1l�[Eb$�c��X<��3�F��ѡ�ƥsQ��`!#�b������MwK�OX����?��]!������u���g��Ei,��zaI*�e�W;��}�F}y�;��d�I,�l/��؈�� ��e6yi���KR�lV������n8;��qv�8�ܖ���O8u�]����?=J3F�C�v�~�"��缺7L�s48�a�.����r���\�~`��4�wq��,v���s�����9�u��n�\�)k`���m/����O֏��R۬�'b�E�AN�!bN]�����a��&S�f�&O[��	���d��0��p
�C�(b�פ��㮠�"�v��CŰ'h��#PU���z*pc���̰�s���`P ��w��g���J$fW��bi���V<�բuR�ϷgU�|���
�Tf0{�_���z%w�(�眯�Yɮc�U�[�������t�k�<:�3�_	����Jo@��z�؊�Sq5��K�2vf��tL�����O�G͔�l�V�����x8*��U}&|E�]��z����;�&�0
+u�
�wc��H�	��H��8�}�כ7����@���L?u	ҽ�|Fetz�r丆j���4���X�I��xK!��Nohq�ز|���ҿ�':j�����-��h��)ey���Ck�@s�y�8D+ (�1o8��W�`t���n>�|����'�v��>8��s�Dd��ӷ(y��%g�Ak��+�aPd�w%7�%Ո��$�.�!e�,d,�,�b���a>�-�ă�f�����|�R�,�-�o���ɦmǁ�늀�,�����t]��م8ϟ��~]H��	�� '����l����3H��l�9�!�^�c���L�M�e9�+��m�S����I��v�������2�
����dޕ^W@�"���&)�
aWbPLb=�)�5�]���ؖl�qmIK���.,ϵ?������_.~ö��]Q�^��0���@��G��{ ��U���%ұ�e�B�rX_x�v�y�!,d���7[S�'e�����1ě�CZ֍Pj�C[vj/U._`��A���9*�I5�IдP���B��Z�=r�2ٍۯM������o:8�$�~K��d@F�O�|5�Hm�]�Y��ʀh����C�T�CV��^�d���t�qx�Sm��ŕX���8��}�d� f7��k.��j�g]7Q-Y���ƾ��b^������h�j�[�f]�5����X���t��k����A�x�a���-��/,�F�5��>e�}X����vu����z1mȗ>�F��k����s&�_�` ��#3x%5�҇�B+88$� ��i7�uV_� ��J;���Z�%pWЇ���մ��o��z{���SdG��C�58+�)����
a�$囂i1����vi� �^�MG!����"�'���M�פ?�!�L��<~k�Y� =�5��7����~~��b�d ,�"q(i��phm02�[
��OeS�K�n�1�#N0���h
�z-����3
1p͞�SP����H���WH��s��b��V���Vc�yu�i6Њ`�������S�1F�)���^�A�sc��"�ڨ[�Y��L�ţ�
�!�Lc*��5%�X@��)*pܭ���k�n&ϥ� Y!?|�q�R�;��)��ps�������es�|젌O"fS��hI~LE<���#�4���5E���_!�a���b8�7P{VɆ��hmL�<\�����86������T��#�S驅G\��1�顬a�k���3H�7ܒ5�kO��V��/K����{b8��㣾�B|4�+�����4b�Y���;�?7찎��߅HX���8�^;R��Q��2�I�0fh���!ZQ������2�����ĤO>j<�e1H0���Q���p1��"f4�+)A��v}��B����36�^J�i%G�K+�kjcg�X����ʊ �X%�4N3;x˧�Ҙ����~,Pp���]�K`cDQ��h��b�֋�����^(i��[$!��j*i�@+����P�ql�L����|L0	�`�oY�4��:W��E�<>�;,��GB�=KJP��c��4��ҡX�+$D�FE�$h���,0Y@ʸ�$���=���E&D�7��nS��e��I|�>��aC*w^��i�Y��X	A�O]�G��?B�cV�t�7Wj�E��3n��u��)�_mr�\|���1��oZ+�K2t��S\�!
I��a������&*��k��;���,�It�K��Q�Q`�ͅ�ӊ���$��R���D���f8)3�֩暎��$�#��`f�<f:��FWGyiø���\2��^�
��C�ϓB��4�ӕ�j�kV�|t�Z��J��c6/b#�r3��0�rf}���P�ϐFj��z�c�hD�nSB�,�=��>��|C ���'G�_����8~�E1�N��l;U��Se���v�{��#�#h�f#D+E%���N�[�0e;��J�B�坖2����*M�~��ځR-K�8���/�al�Ev]�]<�����l�Tf|.&�3��-�8*
�x: �Z�;�ٟx$�a�ɒ��w������YQWa�y��AT�Ę1��n?���%��J)܋�MTMI7�������I�1E:Zi���j�'Ǳ�@����˛�8\
Α^���Oy4m�I5��>���$��IuE룫�?�	6�`�@>d�\��r��M'Y+��~rCa_�V=�M�U��d�xP�Pr�u�u�|U��#�W%5��ڠ����E�}1JP������
;��	&	jM�~#�a{�wJ�ϋ�v �$��(���t�βE�I�H8�7#{J��-n�&�O�`�*��\��QX�@7���^j���5{��2ˡ�����g%��P��ì���p1��,��aMP�a;���u"��\jǺC�3􂵌��aoх�= T��[�I�_9�Z1}��&R�t�w�p��:��.}E�s��ڮ���Xk������NI�b�I��G��IdA��_R�YoDx��Ƌ�(�ꢛ"����T���z23�?�$~��ȏ��Tx0 ���)�4*D6���r $?q3�G&�p�H^���8j��_HU����*rw�,��I����l=�	v�7�T�;c����1a,Ú��3ClM��,kU�f2@.��SF�7��s4ƈ���'|f-� ����� G�V�G�M��]|!k��i�d�:)�3�s3wŇ�%=+k�44�3{�Op��6=;��b���C�.�OH�����A���`��-ԁ�������,D��!���8�E�k14b��s��j8.�)eg�?�Of:8�]Kx;5��3%v�ֆ���{N�b��$N<g��S�I��h�	�U�n�"q`'�7�7�߼9���4�m�����וx�8�Ou�>�N��j��m���{���,3�9��h6U~�&�JB�w��=Ex��Ѐ)�s[����{ �&�8�KAgڦ.����RH�{�_��i [��0^�r괤<l�Y��7�`,�lVԜ��H8�6�Պ�����	��L�e�W��ig!Vz�\�k�O�K3������EU\�J	����|����d�@�"[8�f6�+`�C2�.\��t�0�%�Y�� wl�;�|�Pg۰��b"�L�H)<�����N�I�ъ�-�>d�[ʚ�@ G���>`�}��D膏
�3�w�������Jm�ےΓj�YkW{�\�p揩0rR�'���Q���D�H�gR��m��E�O*�*����[�d���\B��O3жj�����$^���s����"WЌ�E��j�zT�[�/��r��t�o8���MP�ݐ ���*x`�D�mP���iBߋ��mz�(�����x<&��B'ބ�9p��.
���ٞ�k$P �����[D����v
Ň�������(l����\$ ���,�~����뺛$�]�9�UL�d��ۣ��^y�<���fƕ��á�4|�<%.��0k[5'v{0�aJ�^��?�d �l/�_;��.��ޥ�
j^���!`glz��_�!j��\ @�`a�ph�q�⦯�����W��Р�-G���z� �����94q�⃸�<���{�����z�*���`Pn����^>�`"��掕�?ԇ�:Ô�����Z�:��5�j�����O���L��<\d^m���YgJ�3LG�%�i7т��V�'�Z�M���I��/��Y��gԐwY��|!�w�d����Eə ��~��R6����ۜ0֧wCTׄ���/�B�R��P}��J�^X�%w6��z9���!�ё�R�2�%�CgS�JZ�N�	"WV�2�J�cz0k�q�}�����/e3�R�*s��Hj=��e+��Y$*�{Ms������I�0lG�O���T+�Zh��$	��V �R� o*�Y�,�p�}2��&�Xdw�oa�n�~�����ݧ� ���>�*|s$s��#�r�Q�k��D*�\�aM^�,�$�t�e:� �6s�K�h.T䯄$~I�����}�8v�K���QR�y���b�lG��{u��g��i (h�Mwl�
@w�S{`�1H�IV�m3N0���h/�����[N�pU�'R�2����W�Ll�j�p��.a��A��0���M�̾u,����B0U�hP�oԤ��j�1a��Ey��P\��R������*.tĮ ���� �t������U�
m�wJ��x�k��v�ū��3���ｴt�*x���gCV"����x"��u�]�I��[��~��u�����I--����.�T���)���W��Ad=-�������Z>)��֖��P�Q�m@�;�A?	�b�����>�Hӂ*�7:�?�����gZ!���/\����Eu/��\aC՛b���j����h����d ���%�Z�u�e�:,r9K��g��ً`�����h����e�{�<C�
��f4l0��Q�f�4��Mz]}G�$H�g���&	�Q]�JP�x��	�V&���XN��d�� ���Sx;6D�2gV>Iǂ�a)4����R52�M���M�t��|�:/%c�4�cX)?v8���a���(4�>�� 'B�o�'��Ȥ�w���ZĂ�+�Ŕ*�CI����?%m=�<<���>!���P%/��ܦ`�R��7.� rs�䯄?a���n��O�z��#�sگ�+���k�ʪ}�Ko�fp�
��ђ�'��=���E��"D�	�Q����Q��Ȉ�,Ȁt�or�$}�0P�df�D|�T��\���)i�wy�g��@ǩ�%�V|~}�K���$��#��W�Q��w����n<��,�q6��9�C޲@�P��8ՠ��� �0���S�\qI����<��R�~�z�6������n	-�^b�/��2E�����㐼p�e�ڻj�Pm��f17f��cs��\�r{��H3���8��1Ф��z&��� ��ES?�黄�:ɃV�ϗ)���=aOW\��4WȊ�u|Vޤ8�w�PrO��{:���#^�i��*�m=�C�+5|N��=!L1������9�0��SN6�$�w\0:LRs��=�8�@-�>��N���JZs�m����t��dܭ{l�Ŭt""A�+�&�|'�|X�����b���̕8b���+���uk�|p����Ks��86m��nT�x�mKhKMuԠȳǩ�W�I�J�[�N�XO�]�4d�O4$�|P����2e���wr�snH��tN4����Rڝl�`���-o�>��~GԗZ�9e��
���Iw�6,Y)�?�X�$�"��3g�3!�u6�(�󐗥[���t��>�P�����42�@���/%4\��W�4�uF����Յ���Ph���^�3'K���
s��H�����g��%�GnJ����k����h�Q5e>�K�F��p|����xI�&K��SL������;��'KX�n����]R���h����c7}��l�������^ ��e���˽�����//;~���d�	�KN�&.��A7���bnX	Z�zV��k*���RTPqB�G�x�H�ë&zh �|� T��N,�_�:���I�ڋ�M�o.ԝ/쵦�֌�,��]ӕ�����+���]���W���gt�O>WJ��`OڹZ\FjR6{<��_v�T�mL���V6B�;My�Ԫd�;$�N��\����(��Z�D_>�4&�Ŀ�٬�~�'�F��i��on�?k��9�8�Y��&�-ĵe��&V��b�,��+ř;^�̌r���y^㘙I���
1�1�G��-F��(B�'7fI&����D=s;`� s%?���1K����ꔇ�!2����81٪�m�q���v���(C��=;38�=i�;��O�{�/�X�`pқ)3�<*h�ъ�B~���6&lQ�[=������57���yP=��-��)�n���_�V��3�ﰢ��3�HZ\��X��Gp�r�^����=�3tB��֓�����=r�I�`6b��a����}��v����M�O��߽I>�Сb֚Ѻ�W"�od��/jO3�d��Hp�Ep���lœ�4ݻD��l���5�*3��%G����7��|��(��t'߸�t#�k1�k�Q'� ��]S<'_�����m:���|�(K{s�pd���?���,�G	Է}��O	S��|�j}���G�����B��R6��,����K��V�Gu~��^�͓��k��ֺ<g��d����J�g���A�6B�#�a���wKe��:y��ɯGm����C�(<�<�s�}��}[N��I>�7� ~]����G`�K�j��s���^�����j���}ѐ1p�e1�7�Z���5]D�~����ǋ�,��r�"��L�P ���;2E:Z\�-k�p�"*��R�%�G���,)^wE��!�(�$�;�$�E;ɰH#��Vq��(�3�.fR����>���_���}*!�V�-l	���rî�����Rќ�čPG�TI�$l���;@��$���sL8"�N¯��j�Z��b�D�}��$e={zo��I���tB�~��vK��2��ÏD���c�����	v��)}sr��v���"�4��">$�S>#�� �J'����s��X�ZZ����2J`f^Q5�	��zff$��p���*H����tVNBX�P���r�B����>��#��߉	���>�[!K7�p�����|�#�]!�.#j��D��-{����n�-�!�pQ�;!���0p�	�ALG�
�]���,ǵ	R3�[�$��"���M��f�`��{@�+�'k.� n%��.��o�Ͳ�1er2�tD1V~b>���/����k�Ae�T��B�wL��)��K��e�1��k�7��lW�̀ˋ �cH|Q���)ڄ>��k4.ۣ�Y��֧�X�Ir�����O������Xb�:lZL[2X�G*wĜ�0�`ؠ(@,&޿�S�ʆ7��H�g曔uJ��?H��5��K�����{v& V��p�/���Ř�E)�x�E�*�ye
�W�=��k01���ʆ����	�P�q	�[P
*C
�f[&~�_1I���zU"z2��:�S>���- �ﱥrmC����R���gT���s��攧��$8�΅2����*i`����sP�S�c:�@�@�l�X���E��i��ǿ�`�7�r����8��w?��_-Z���" �U\N�u.���I_aM��_t��E.��n�f���R��l9���T�T��=�p@���+�T��0�bô��WB7�!hcԌ��r�[D��|%��E]�j�|W�b�$��l�Z!�v��ΏP���1�pt�2�,�=�&���\�ţ��!��������C�D�"�N��&��\N��E�*�ov�R���04��S��|Du��u���@�L��0��=�G��O$���Ϯ� (�D��,|��>db'�wK�-Ո&��.x]�e��@Φ}Sy�m�/�$����2��[����-b��F�����<�N��i]Q��u*��v�lEp�G�Yo^���$��45�1℈$J�eś�c�Dȸ%͟�Ej���N��R���U�� ���	\Du�627��P�;㳀�c���?ȱ,������(�#�� ��g�>�dw�Pƕ�ʉ�Ԅs�R�p�?v� ax݄&gp�iǾͅǚ��~���Kl,�G�Y %!Иm�M���K��Ê:�;����T0Kן6����ReE��J$�L��<K��|�Z����/S}�1S�z���<pG��6��J�9��8h�"��X�~��,Dς+{�׫d9m�K� ~���[̶C�vadAyZC|�9�w'(������ƅ
7'G[�{UTou|���g��?�YQ��t>GdS�wM�Gu���¦�f}8	3�R	���.�ky��]��Y�6*�E�/�k����.!�iF��>�Ə�m���_�p�9^��:��v��Y�F i`à�A'�bw�,��9�	k�l��W�������C��$����9�r=v'��"6���H��b��L�X�f�*"�v�OO�"�pg�M}�]��)�n�h���8���!�𗉌��}�V��d�H�Zm0��������ͼ鏧�Ƃ�v���/��9���nC��=�1����x�����c�Y���f{P��6�/�Y���nl�Q)�Z?5Y�m�ɽ��y"q���}=��S�]�o��V屲�Z�77�\]P����?�))�#T1U9$�_?���}��A]0\Ύ��"#�I�й�l���?-���;ny�;��<����� QO���1P�;��� �;ى����:䬋�;sʳl񼑒q�;w��2���8���<����d)��i��!��RH�c�H�6�-J*c��y)kԗ'ޔ���J�q��FY���衒�.�S.����1RJ?f}�0v�dH����"������Qޚog���*	#C�j%�ox�g���SSc��!���2��e^��&@�V�v)z!�o���:7X�e �^��le����FX��hXoЈ��ZgPOe����
&n��Zɓ4c���28�Tt/������윙��o���[hr���(��g#�3��G��p3'�0�O����;�_��0�?�ݘ:���̳r���f�y��%�D�O}n�[.x^�!=����t
��2��yD�Q�u����Xd�X.��R�#ѧ���>k s�e�{�6��[���ۂc��֋�3�1�m��f����r?� h>�Hc�=V݄�A���U1�H��_�"����c��O���`��mL���=�U �g
��^�����F�.����i��/o&T헻(Q��+92�o���}���!o�$8�T�9h����`Χ9��u_P��R�oE��	3=,�ㄾ�\������+$=$���]�zJZ��`�c�H8���9q�l�µ�T_��2��BgUv�P'���!]���E>>B��{*���Ճ�@����oZ�N���}	��~��*W�
]� ��H��ߴ*$ ��++�����E�cÝ�<{N�Et�v_��N���l���3Cn*ia7?i�)m�Tc$2�Z$�U���%P=�ai�s�����'ߢ��Xr��R��;��r���S��y{?�y�:<��m[�?D�I�QJ����WD�&�:w�w2Jgt��2��|�xD 4#�\Yp�~��Ǜ��
u�Vރ�ꄪ�o��V���J�N��[�_��B��Q��A��p���z�q;��_aZ��8��������XP9�M�5P�	|z��j�K`$g-���2樬����|�=l�La�e��KMu�ZI�B3+n7��y���.�t�!����:�0��C����H�#����+�^2������&�[�Џ+�3��Lo�������f�C��f� ��B(9�hգ��!���Q�Y�a��U� ��8�.Yhc��g�݈vp��ɲw���=�����̯��i�k�7����������}|�I,ҙ0��~H>3E@��[M���ymm5{Z�@'�x����;\��ժ>WeK���1��~�u���Q��d5� q��T{��e�����R7Z�]r#��._��w��L��U�b&1�ۚ����@��7?�?N�[��W����Ɇ;�۳:0���E~�������A*�O"��x��?ь�E���9�zF��z�d�r���w�T$��� &�t�Ա},M����=�>Uf�WU���v�H �č*�M]P]��~�S$/K�/i�~��}rT#��|��y�B�#��P�E�4e���<[+
t�r��*�㈇�I�1��uB���f��:0�i��c���{mJ����,����¸���yl�S���Y�'$E����?�B���,�� �!������°X��.�����|�^ѥ�_Rk�����Z|�}��_K�T�r��Rk��&�H���-�D�q��Dqmq:8���E��]f��R}R:s$fG�	�E���'��)�P�1�k�����
J��x�ׇ|����ό1h	�Z��[:SW�p�M5��s�P����S��1R���Mv���n��mŷW��:$���`%��o�!���͹`��4��<�T�)��\�Qati�K�٪���]���I=�������>���T	N�j��Ĩ`l\,�z�*���L��R;�x�?�s�2fx9�h�K�,�����HK�`�S����d�.w� =�v�����jnZkI�G��J��y[�%�uXP����Y#Sr	vN{��_d���)���3~32��$/~������ ���O�,_��Um�Ai`�5�J��٫�	�=+���:�R��#W��lF���'�@7E`��Y!�B��~�����\�K�p�\��6�rO�KvM	)_�j�_ۘA�ķe�9���}Z=l7[z׋�>a�-�v+OĦ�s4r�"�w���g�O�|���8!��4���ىYZ	8��Y~�<����|=g��6�1� �Ɏ16�N�QLi)�vz���P���T�'Y������>מQ�?����[	�����
i�	���,����4�����E9�V�����5]�C�I��my�BvI6b��@��X�9����s��\��E��Jڤ�B)�'t��IZx2U�as��6�8�����C�"���IL4���\���H��ʬ�s�WS����h�Ɨ٧~;��dM��T�`�A��Q\"d�tl}��s��=2�a�l����ҸGJ'6�m(�}�A�ٚ.��D���x.3hYq��8<6`�����"V��h�2T��(�bW]�M���i�4�+���U�5̣
:Pm�>4��c�]�+��@%���
(*_�_ƌ��΁������;�.1�E��j�a��0�ı,oD�(�aT����L[�FLN�Y�s6�)�g�0*�3�G���kV�J�Z����D�Zҟeg���t�
'2��?,~��W&�/�M�~�����z#T?�Su�,Y��Lw\|J�u摂9w�oQ�NT�M�g��*����>�*N�۴�X{�`�F�k`��.�q۝��?�^��^9����s��<@YU[��cdk����r��%���L��J�u��{��##���L5 ���5,`����%d��w]ǉ��C7���bhh1����AZ�|=�e��c���;b����r8��O�@%f��HJ5�!�����M<�^���ii;x�Y�f"��G�Sbo3�����_�����=���6�1�����8n�c��I��)֙���Ū��9��!�D(��PF�M=�a����Y�v�n��N큝�G%6د�	1�m��u"�>�����!P��Ns���N�Q=�����5��oC�q����)�[���5s ~	0���jr`G�xO'���%��|�p�g���%�k�p�P���@�������n�WS>V�6>ҏϰ]#�+��Y���}af�X�;�w���M�A_� M�A�f�OS�R�Y-��==2�Tof�l��i�V�����*τ�ȰYհ�)+Uf�c&P=�r}Z����L�t��Qr�S��Ĉ0x�����~����Q!�V�в�jͯ��<�P�/�K�{k��K�;"b����c��ʾJ����l�E$-�%��<:/��Q$�L�D��x�[�����/W�1�T�p�ZJ6��'8�hz��D�:�^G���=>wr�+x��u��T�WoO�ϴilGY�/ks�J��S�5ht�ܕ}�p�b�p�o�6|��A�"¥�L��J��y@C����;�ތ��[�3
��T��^���x�n
id(����@k��\����%)��;�1�'́H�6(��������r�ʖ�;���6U>I�Q�P*6q���ʟ����1G?47CKݰha;���	���@�LS
��[/s�t[,r��J�قN�RZ��+%������|����� }w��K�7�~FT2|3�U������z�=��������U�JX�W�T���پ+7�^v1��:�Ey��ǁS��̮L/Ԃ�6p��eU8�tA��j�5��71^׮��ң:��B����a�s�XצZh�;� ,�%�g��p�f�bh�S>�'�,��:��z�`�a�+�T�a��> (gUG�iI�i��u!�\3���οml8�$HE.�,���%����ޟ���N�K8�����NY�_�%<u{�����۸@z8�ע�X�zO�&������<�	Q�^�BH��z%��6lr�]+J�/v0o�E�'7���j��#?7�a�R&H�ADwL��CF� !���3�4NË��Rp���K���XH�[&��F�1y���IVi�X��%гv֝}nb�Jj���3h�vx�PT�JS �t�<���ᩢ;Rc%_�Y�b�JmH��6����U6�����JtzZ���SDUZ�����D�>Jh���� <Me��S�$f\h���@�&�9���M"�dP `���p��*$��$9>(����(�UK�/�2O�]c��beR�h�2$���
w�S9�AC�^� 3P�7��̡��W]��0i���D,߮��n$��:��&˔;³���;X�t���"3�0��I�"ҕ��X����t4�b���Ky�6��#m�d�?�T�M�k�ψ��g�����&c���zz������65��)��tXZ#����^|T�e<UplMκ8�=���fJ3*D"� !/?�a	����K�8M� S��a6�J��k��$��J�T���𧌷�^�����$��;�8$���O.E�6�zF7o#���5l���&E��'�0�,e�-�>��@Z�E��X�r�߄�� �@�����!��@`� (�w�r0Ocv��M��/�I]Ӕ�ǚ�9�Jw7.G��pУ̵�/Rh��Xq�ͪ�,�ԙ�A\�,�@ϱ���"ځ��ME��/������~,�K��3R�fP\7�3��	�Ѽ�-[�O�!�>�URr���q�A��GM	@���[����=��>O�D���O90�2H� ضF�P	�u�T���^M���]��n�n%\:2�k�C��/~ڽ�+����:k���p�#�C�x�� �(�T6Ac-3ޥt&�m�9��ob��Y+��d���A��]�7(�<�i�G	�-���@�Pn�7'U<����)��]ٱp��tx�[�`ya��z�J���m��-�$Ij\z�c�|�f�b�$�&?s/�Ra� ��g$1v��>�3	wtWb?����u�S���W�S9��d��v�c�����d��o�\?�Q_���w3��h��5�8���z�=C�xnBa��p��W���R����U�;¼��]4$5�6�j�!i�8�|]��i�p̐����~�y�J��MJ��o-����5��;U-Ɉ8��2_EF�&I/��/{�v��6��G��0Ws��tH����sp�p-HɉpU�n�>���$�2��F�8AK:�|���44��S	B(l1N��G��ʴ��U�d��Y��ӱ���T���n��B�����y�� �KĎJ�<O]uFv��lPl�L{E}6�1�}$1'��Oty<s����V�@�|����\�:ZV��fk�gV�w�R�^�3����nD���\4fN���1���Xih]�r��0&Zea������S�Z���|���M\�:µ1^�
�)��JM� �B�~�i� l�ɇ��^�x�J[�v����8�5Mk�7ou���Q��4���4C-��,p0}���!p�Z�P�Ŕr=�u󿒘���A��%�l�W����(	�Dz��F0t�����
������=P�q���E	���U�U�_���x�||�Yz��ᩒ�����k;���쓠k����O��>y��D�!��_�B���M���_Z����JX��T���}{M9���J��"�vO����(��}G6�hU�%h��޶��1�}����Q�r���o��nƤ��Oݖϵ�Qe������?)@Y\?�6��qJ�FǇ��<�r�\x^�	Б�����P��������נ�$DΟ�E\?�سڝ�m��{b�{���ox��#�p��Nl�~KE�VY^9���i�d�͹�ㅊpj!��I����*{<���XL���������?�j���,&˺z'[Sт�PV�/��Ƿo��Y[�
=zk
s��Z��̝b&��#�!�`= E�jk7 ��1[ӷ�DlD�v����X���_���qK33m�F�Xpm|�ޑ6W�ɪ�b	y�����y���I���W�ǈ�.��Z:�'5�e.f�1�ڼ�@	F���<�?�X(Z���,g㹇Q��JP��}�I��V_ׇ�B}�%0gXF�P�	rzl�C��C��������gJ>b�(�_j��6Ebw�3��ϳ��(=b�&�A���A���/������2��mr(ǨA��3yv'��,/*����g}Æ��9]����,�	�]���wb�W��98�������?��G^š�T���H�_*T�y9��z(��|e:���?��E*H���p�5DEm0�+ô}^Z|rJ-吩J�$����!O.�ҥ;��"��6<�0Xw�@/��:� ��{צ%h��h���!_���)t�3��rM:B�~i����z��1mO��fgS�p��ΝB�/[�H*����=iO�[9US��+	��3����4ݡ̃C!�H�%�J��y��[b.�]�䑜R��u�F(<B�X��E�24����1�4Cu���/�h���͵h�!����x ;l�R�h �1��ߞ��:
�|��:V,Ǭ��)���T�Lv���-ܬ���"u�����Z�1��?ș�g�S�!ĠQof��'���^��#� ��]��$��&�oaCI�x5�xKz!T�Pa�~�"��9�eQ�L���=�$2���)˾f��`P�:-!��̓���!m��Z�W1����3��.�}��h���$�{�H��p0��ɳk�$��7��|�1ל9�AA\\�xW�V������\�N!��3���x�?���Ǧ�Ps�N��"�;8�Ky�w��dM����;�=�g���(w.�:�{�����8��;4�kab��b�m�y},Pl X��eƨ	ݏgR2�(�U����<����l&_ ��+?u�v%3����W�7ߣO�2ߊ�Z�
֭2�ƌ5J����͞oOnQ���Mt����L��txAʃ�8ږ;���\�@�M0�M�㙴�Q�]0�(P*�9��p�<�n��џXs�-��-k�bx�N8��2��@*�I��!�ؠ�k,�+É~��T�bED�����TQ���݋�*$�]��qY����� �N��W�5�U��u���ܺ�I$�� �7B��~`6��$r��y߬��'"���`��2q�_f�|��~NZ��ÔO
�	H���n-�X�W�& ���Z���u�g�H�rN�J��	�kM�Rl������	�ݯ����J$N���	��<�_wZ��Z�aWTAyx�\�T��ڪ���w��_�m���p��)'#/�Y�
L�~'NQU�� �QI_X�)n�-�ɐpغ��s(&�{Y���Ɠ�f-���/�g�F}[�ƪ%����)tJ'��h�c����%�c%�e���I82b������Tt��p�N ��fԇצ��O�E8@v����Q�]�p�Xf�mRͬ.>��d�z\�`��X,���׮��e��Q+��~ ٗ3=��>�C+e���7�Ʉ��$8�$?[M�NP>�tV�k����(���p�Wnدހ~ ��B�븿\�A�4O5�T��rӤ���j:�<����*���bűD�F�<�xX;�L>!�9M3�9�Y�^8�!��&"^"62շ�����fq�S�A�!Yu�ǁ�oY]��~Ecih��S'�D��tdJv��f���b�>���>xO����D���2'�8�їn͵p��A��aYR�U�}�\���j^�y͔0��5\v���M�<���ۑ:�% �K�+��1��������,�f�q*-��p�b�k�M�D�a�Wl�DT�hK��~6�b�R��p~WI<��:�c>��&7��r��X�vx\�f�Xv ����~���HX�Ǡ>��a�w(o	/P�;��N}1�p�}l0����a"MZ���p��>(B�Q[�ZQ��\=�C��m!�Ԋ��\��X�l �2����sgւ8,E�Zk�s��X���HL��D�U�alQ)V�R3 ����o\���eE;^Q��3��3� �&U�w�`���Ew���*��[Ebj�.�BS!WVkr�}���%Lgi�S�2&���b�c�R)^��#Ǖ9�ɑ**�;�`�:�Z��x�|GŤhj���I��L0i:�;�%����u����P�?���J-�W�N��]�R( ���^�R~�J�zŠ��2�ޔG�N��rc�s<ޤy��;E|9��"��,�L~�PJ��:ׂ&���XM&����^pܲ�L���� Z�I����wL���e�n%�����Bi�XP���}��6��C#s4�ґJD��Q�l>>s;L{��_�jQv� �Za��m��v@�cL=��g�x��m.�%�m��Ҟ���m�htAN4�/^P��ݏ'�p9�f����I����3*���C�7"8g�kx
j�)|X?��(�dP�*�F��	}Q���$��:G�:��r�d^�8�,7��U�q��Ė^Qe�M`ܒz�֧�6�q� ٕށ��')ܝ�>���lb�纰+�(�Y�w�e�v?���&�� �/'|]._�������P���G�G� `�i��{��lk
}\��L����G;	V�i�����ZT�+s�L̑;_8@)��!�S9I%��/'L ȿc�Ԭ���r�4�ց�
�{�:���YR�/y>e>j��
���@Ǣ	�ڧ^�s��_k}��֮=6�YC���Ɩ��~C��'��Ќd���w�U'�����`0/ư3r�������Տ����H�;��h�Ć����&%�::X��"Flx�,��_���VH|����_�7����d���d�ݲ[�����DZhm$�|=�c��P�o������e�Y�Q �bzV�&�ܽ���X�{��B�O���h-kE$c���h�!ܦ}/s��*7���It��@�x<���P�g'���i��{+���6u���۳UL�eS2��o���n�1e�<»�c\�%C�46�%Mu���l������ςj`���|W�Z�fR#�!�<	3�j�WGM2u�t��P��".Dm���%ղN|QXG&����K&�.����1\����s7��ٔ��J�F����e,݄4Ԫ,H����y�]�Қe0�]��Ͳ�v�Y�kmޙhwA}�#�� 2�Q0��L�O͠(7�׏�?4����g�L��4vM�gRξ���t=#U2$��<��i�g�W���}�e7��C?ķ;���?����6�$,�N�jb�,pB.J[K�/��3�Q�J�w(�Ʌ�N�Rd��g�#�>�y*<�5^\2����񣹷�fDf_~��v���t-���w���֙�'a�໲��bC|���$��'c��o�
B�1D��s�ic#�;�s�hc��5ެ@R!C����{յD8�:_���-a�[���^�)ucw��*��`���Q �ۈ-]��ݱ��,��j��@����X*b�����k(����'�"��OՈ�B;*`�<-Ȩԣ�G�b�^�ː,�G{�?=�$��(��^5�+��p�z_�97�@
����E��k��:��=��at�f�4:B�kj>n��+·�p-N�%E��¶(�A/����<���<�Y��%XH���XA��T�4�wwb��@�{�o����<���q�0���@�[ǨQY8+��EaG��䭡�Y;�@F-�gZ��v��'�2.*�~(�$l�({�������?^��M�$����2~��
Leغ������ϙ>zx�?D�=��n��UD����?������7R#	Fފ�ۛ9:aR�̮��8˞#5�L~^��O�a�-^�#��T����p��(؅U�E�2����N6�� y��%ѫ�^�Q��9\͑�Y[���d�ڑ	w}�`��p�<3R���F�cMi��@��
5�tq^�GeY/�?�73[A�r����'GD�$u��>��X/3�ab���_�Q.�xG�.�/y,]��e��0�E\��B�{x�t�"�fe�=��Z�q�@�5�TW���L�Cge�~�X,h?*���̘�,=����<�O1���V$V?����a�
#�T��6�x0�>�^�4����s��0"ny1K��� �#��&H��'$@P��w[�Z�wH��N.r�UZ�kK��do��(��"Fi����jk���}��fX��J�3o�ScyiNW��8"`qS�)������w1�od}��Qh L"������jV�*i?G?I���!�����u�=��MǷ��N/��z
�mH�Q�9�TT~�������܈���&��&�l"�[-U�K��i�wt^I��afq��i_�U�u� ( �g.\b�=���v��k�!q���$��nFh�|X؜�9u��۞�٬�	��(
~Ϙ�R�!��p\?�4u��-ӱ���I~}���G;�'�|�����5���&�fz,�Q��ݮm�@B}���R��`��+��w#�,/g��aZ�50��R��l'X%��'r��Yqa݂dθ���,!�+ɢ\�/V~���{�W{����t����r
h(�n;��V71DU:�L_9 ��֘zr;��jxI{���Yq`ӿ<��p�ބ�E�e5~�ҍE��� �B.X(F8��C?;n�y�Z��C�/C��u����]z ���6�	H��5\�����Q��	p;����� z��IS�	�!�I����-�<�@N[绔ԙ!�5�4�E�>N�HV%h,Cl�m�g���sO�vځ2�,��JgP��GI8��b΀���1'?�*�k�0\P����~�z�{^� �@��ٳ�n.!o!�s��d��3��[3U�h:��08�szSGlf�h��M ����� 5_�!_n�r,�ލ{�������8�yy��b��y���wɵ� �lis2�k'��g���]	k�f��y�O%�mk�I�_^_�������ǳ��]y�3Q!`g� T�S��� ZiyP��B�ʣxpЧ�[�<5z�����y��aq���� t%;�!��S�n���Y��~ΔT��|/���^ie[�����h�S�T)An�%wKe=���׈���y���VE���wz���� �|7?2PL���9�w�m!�:��ƀ��������N4�LЛ�C[���L% N����9Uz���,��0�a�*����]/zU�o��,��н��	(T4h���l�͏_�eSW����9���%Uy�lj����np�e���k��!u���¯�r��a�����uQ��T�+�4���M�~���7ڬSbyق��}j�tn-�N���{�l���,��:�zZ��]L8?����b�!�0<�p�%O,�jԀ!ѯt�)������I�7	�+�	5���T_h�/�k��4�C^�p������p�Ŝ�j�]A5��y&����ݔ2�Q�?����������B֏�hEW�G�o�#�>�?cL����M�<��Q��-I�V{�1n����$jﵭ�������1��I�o��t]�%B��>��[HO��;�L��P_�l^2�T����wW������K����E´$E�"�Q��^(m����pzu��,.�*�c�?��ahD�����	�~W"�.�tn��.�J�4ނ�/)��������mcO�:+%��i��\y��0.㋗�~��qP���$���I4�b0�٘�9� � ��hL�X��]}�!d���e��u)J{�pc����@ e3���Q1c�J�?�Kΐs�.�l��9ǚ�%�yD�f)���q�ؗI@��'^dڑ
і���3��y����sg+3K
�*v�#��B��vFZ�!���h�Ƕ��j��,)|�0��0�a�Y|s����.7�C��V�PC������:�Z5?#�5�v���gM29�]�˅�&����`~ZUg����.�vi�&����6AD���Y<�F�_�O��Y���iM��x�l����LHG���s��ـ��-�7M⟾��rS;V��?|00���_���
�)�� c{���X�Hj��Ԅ������
~At�a`��U�Z7N�z�XGr�t������FQ?�s��q�_�i{�"��|�/��7��D���}[�g<JW��\/�W�n�8�{���9�Q�~��j��"#|��j�ܻ9e ��H�j�X���[n�J^V�k�>�DH��ډ$d������A��%X��-�^�̇UY������0���3� �k���t�	�پ�]�t:xFD�L:�<��J���ڴ�2XZc��Ȑ,��@�oI�j܃3!��0�q�i�Z�Ɉ��6$��-��`�2�m xe�����C�:=������G���VBcm�����Ã�w��6�M�&le�ۦ�x��#J)�R�٪�Rp�� ��#�	�)��!
<�9��
`c��cn=�w2�]��?�+�݋��y��*Կ����F�7W)��ۻ��5bk�#m���hr���`�$����H��ຜ �ˤ<��~��u�}��<�)I��k��	��\��{�Nd�I<u�9�G���˖� _67���ç
��56��R'ڜ�6iӐ��pu��:=��^�0��<P�1�3��d���������ܮ-B.�jS@aP�9�p�ʷ�;�5�V�ɟ�EȹX�k����NX��zr��T��[�r��[�B;|Ж(����jR 3�a�0��T>���֨8^��wz�X����[e��OV�����D��9ru�H
�j�Ci#.2�RΟ2].i¥�΅#�{���a��<�wV0)��儰��1��#�Y���V��u"3������fi�\"�2�a���A1<MB�x�0 �7�n���Z��Ql���r»��㩹��S���k(�1��>��l�k�D�6��ly�5�A��HT�_w���x�� 8�>�����aK��hi=����9n|��쬣��n���b�] �Uљ_�úS#?� ��j9�N���K`>Խ��T��[�ĨU'����ң*v��x�Nh �k/e�*����K���Ed��a�ҟfܜ LVk�t1{����x���6@�
'�E�������r{��HR`��Azd�!BG�E�@�ζ����=q��:1�	dV��?dڒ� �\��e��G��S3GI�_NT�ȓ%��"���u���6�+��q5�kG���ʳ�9#lW"�2�Ư�c��Z�u������qנ�Afp��Г�u�_N��v�HWbӏGmQa��#�1�k]�YC )�oDZX��ݜ2lm��!�3�w�K��ԭ�st�z36\K1�J+��m���s >
6�32�-LO�T��q1u j����B4���;ݾ<��{�=V�$v��fV�����.��i�dL�jS@dҋd�����I�S��GWP�S��7�>�t�:�*��o�&�?����Q � K���-e��=�Gk2x��w?�q�#5;��xjt/$�7�0����x\��]-Z��tU��������k�-����Gqk��$5��߅ø�7�n���v=��-@d��4l�PA�T����+�D(+��f���v�L"�М�bĉtA�7^ }2��l�o�����s��,�M��	D�U �uFa��:Ii��_O{��4�z�4�I�~���E��?��e�l�d�}���0�UC:���A�Y~�?9	�Srn��/�Ͻ�9o���{�%�"ց<|!P �ɍ��ISN<7�N,�3��WfԻ�Y�g�WoMJ�t6�Z��S��1q������q�v�Et����;��i3���a�l�]Q������S��ip�?O�ly8�bz2���,�~�5�fW0�촍t�W)Ԩ7����=P���G���&�Z�~�~0�,%6�kǖ+Û̲��P�:��� P�;=��\B�c �" +VȾ�⹘L!��db�o.p,��,UI����j�]�Vs�J�>T!j�	�Ԙ �v8����"6IC֊��/�Wv�-� �s��c�#Q�DB�d�.��� �Y�n5cRcKfp�%� N���q�L ����E�癧]��S�^ٮ &7���jNN:�!z� /(��fM04��*/�ł�2��Mi��@�&TR _���-N�H��8�[f�LLf
�L~MϘ��Y��go-5�"!��bl��&�+(�,����
]c���?,j�����șyS:ϗ,sD��a��-7f�؈��4����u�Pv�卋���s�)�W���M1���ʒ��݄d�t*�c�mU�L����x����,څ��w��[�o����U��Ag��ǟ���m�W�f{F�]�ʿ��%j�	�s���+ݣ݁�)�Gca��C9HV,`{��`㉩����ߎ�C����ۛV��>g�]�s�}ɿh��L��p��r��n=�H�-T��,�bP��2	@�0
�%g�JWQ��S��*I}@FJ.�L}>6���6�hz�3�V�ѯ��)~�<��3`�Z�K���M3oG���hc�S�'����QF3�w�|�'7�
Y <��i�-Kh�E{%�����!yD܄�dgo��i^딳�h|�Dۗ��ٲ����x��� t�$#�-w��X��p�836��n+R#����|��-KTIةc%��Wv����^a�7�"�YE����J� �f.`N�����}h͗H��yX7�M�o��!�H��;��Z�aY�!��E��g<��y�7����A׫4ʐL=��ؤ@:�yu�\p�&�[���[��2�2Vb�dWe,�ݩ^)�b���a.oY�)䆙%��b�U�I�GX�Bf�+~�i��n^���k}�f&���t\?����"�^޷��yOGq����k�c'䮥�&ޏ~$��th��װw&��G���EH����N�[��2,^ǩe�<�d痗��'|Ú�X���*U4	���E��#934ObK�|]򟑱�B���EY �O!�r����@'@�Z͇��%rW�tNf7P�˦�yM�� ���	��"�{��,$���^H?���LB�i�ȗ�0��2�N�5�0�7�(���g�.^Ox�`G��g��5i�\+9������%�u�i��=�ܼO~i��3��E���������HV���N�Mw\ �7R#D�S�D�݉H'��'���H�,��O�^1B"��N0�^%�?��
�,��r=�Alx.?�C�#�T���W�Ua�(f�k�SIgڲ�4��v��t�'�D4�DV�s+"!L�C3Λ���	��{/󂏥O�HdQ�$<ڼM�D	�=(��Z�j:���MG$ɞM���/�P��9|���8�.�=�Άo��W\�U!k(#��\%.�|�:4C��[��n� ��-ZbZ�_fĴq^a"�	��e�n	�~�J���z_�E��]����۵��;a���:��>��͡AP�ҡƢc:�~�DiD�c�,�xQy�_4m�&��.�a!r��ɸ�˪�
hmi��R�B-j�n�/��%ݟ�&�ϸ���dve2 :��%�${1��+j�>g�B&��3��Aw�,�^�?�G��ל�L|Y�Ww���N#`�踻��E�р��
� ��`�
���n-���z,��L)͟'��Ъ�n2P,>�bq5�L�d+A���o��ޥG[G��X�2�mӷ䂹؋�wW@LP���B����y� !�`�>#����-�c���@���\�̙���o�gDn{���6��"������_�=3+��-Ho�������v<�����ʶE!N��Yq����LҍX��X��W� S�b��C��ު ��s�ր�_|�� ��R:{�G'zc�U����h*ȴ�92�"�������})L)?)F�tS��nu��j�E�3E׀�Z2�a��p��&����٣:|�m��u�Z^�Q4�eM� ^#�:Ags��5�颖E�tZcA���Sx�;���9��̦+���<��Tu�'�e�Y����,���Sc7~~�3�q�D��#���&E�h~L�킂(䘔�u��Ol�*9���upU�G1U���r�����[i���?���V_1���Dv!S�=��}dh�ܯ�&�%W.bQ��Q�v�ޕ������~�sy�%ޖ<��o| Y$:�<	�Vn���N^�È��Y��U�aZ��Pi����h�|�{l�����Rk�������l�^.Z	smdG�yD��Y��F�5�ࠁS�,���DL�b���:!GL��_�W򄈑f���G�B*�p����Θ�1��uY�<q�4�M?�%̪��& �ǲ��3r�U�8������G�ݩ�����pT�#.��H�&ge�t9�%6π/ͦp�Ї�|/c�W)�;~-�svU��}��L��}|�B|�����L�2�>9������'�,�0�0���jK��ON�Ҷ4�)L����t���cb!/�i|�|������h�:�x1M}FY�=��-&ն�Yc�|�o�NU �����Le/}��!ɐ�૿��Nh�Z���@Cd!�VTp�&��q$_@>wh�_th��W��q�^V-��<c�J!;�i���A�j4!^�v"������}��X�	M��}����a >3Һ����[ܛƊ��*��_wv��5�(v��Nm�h�;М��oQ*���k�B�B�,KQr�0($}�G0�mOL���)�Uh��A�����J���߶�� Er�?�H�����f�q�箅�_��[�Q�K���f6(�������و�mz5 mm #İ�4�s^�v	� ��+����jIC(��G����EB�z��ŸτD��m����#9�,�e3f��i)��`K��2���9�������`�O��َ��|U-+��z�|ݍ!'�_厒*ri:rd��<�Awݢ}�V�!$'h�[�|&��%���N��/�b];�f�v�A�o�BɊ-u��J�z7��MDp ���^b�R�zљi�c3�h�Դ�<<���3��y �ƕ�����TRLPH�W�;�PHTq����	&�)A���,�u͗��0�+�f��(7�׀Mھ.�g:���+��#����Z��*y�8�V��ج6�i9x���	��h�� ��^�0��C8� �S��,f� �u�K%������f�v@��
��)�O�z@�g�x�}J��or�JV��}��_�4�5�/P�����8&o�!���V�}�8��O��1� �E7u�چ�-�1a����>�d�z5��Z�s��F}��χ�Uǽ�IF�;2z�����M\U�Z�(��;<ŬD��T�qLQz��&a8����������n��Z'5�R���C�.��V�I�y2�Ո��5�8�:�V*OS�]%��1�[(�Lˑm#]�˨���&xk�D���� ��҉�K�M���\bm+D�	���x�$�2��맔޸] �\h1�Fe��wHE;���'�����<��VT�d!whn���� k��$F��U���ը�W]�p�;2F�Rf5͎Y�g��>�����.�J����<��F�?vA�xW 4j�P�3<��6;���-Q��}��׿���E��Ԓ����:s�F�Wb7R�k��6�͙�	!�ړ)Ao�½ "�]`#t8��8��Ⱝ��	��|!��f��1�BNh�(ؓt:�{�)�̫�ܩ�Wh�*��zb�+�8��§��e�'��l�&k+�v��!�}�$�@����4E�5��@uH%�1�k!ݏ=t���	PW'>8F�CC�Kg�]X�ء��,�*��v	^���N�]��Ɂ�F9k5�N	���ͅ=N���� gw�@`�˺L�f^�g�4�
�_	9��7���!��X"a_-J�A���x�7H��nt���{).��(o�wBUW�P]����fѫUXL�)�bD.�B��):���֖3�c�D|�b6I�߮�����Jk�؄�I�.���%��O;������ejf�52b����p[�꿖O�L۩(#.�3���� S5�@��D8�1��sЏBu���~�!m5��ӹ	�[4��,�1���%��<�m��
��� ?��k>�����!,��H�;��WTR��9@�_�;=�k�F���C���d�3uP0��?CU�d�MaUy�>_8�6�'�됴2��!���'o�p�(����5��)�U?��()�q�6&�z�����.�D��0�A���ne����2�02��?:u� H�}
XrE��i�v1��$��̊�x�r[dG�0P�CV7	۷~��FI��%Y��7>��y//��z�lp��YS&��7��y��d^�m��~e%9<��v���:���)�O o�T��jެ>PEҢ���%cW9d��O������7 (��h�qg���Ԣ\wX&��#yV�.w��ۊ�=�w�-��]�jܓ��kU���{pE��Rsx[��󊍮!l�����Cc�w]���E�ɡ���1��)
����Z��u���^s�����A��G�ޥS������o�;׿3�_�|��~�Q1�[�|�Q���_�����?�&���p�wHf��[��~c,H�`��C��/���9|����X� �{	��t���E�W�-�A/�O��g;/X� �2�G��	f��p�&���k��>,�y����^�����T�l<vm�����9J�Cazyj�����ݘf���9�Ep�(�$lA~��J4�>�ZI��(���*��w����	B�����{��+�n����:%J��ٞ�U�ׅ�l<�-�c<����d�'Z�"��$:��~�-�m��{x����P�
qC~3Xz4�gۗoӾ�
�O++CE:%v��+'4�S_�Tt�(��Y@�C�sU�F�������;����M@���N�N�iQ��>Ì�˼E��r������@u �4��#<I��j^U�v3p�-���*����`�z_� ����%��/)^Ncj	���0�{?,�G�v��DT���@�˨���F��?��m���T��濗�[�����0+k/��Rwʘ���w'��@�+y����S��b�T� �6��-8²-��Ȁ�ƃ�H\�0��l��hT�{Q�3�m��N�\�9��-&��ʣmD��Pjq�+�%����/�
D_�{�x�ӮĎL0p ��q�4ѯ�,�p��T�<�ٙ2_�C�~B�1��ҭ'R.4�0=!�����j�����&�@�$p'l��Vl���|�5	^�V�Q���Ƹŕ�uW>L*�L�>_��CS-����[��l܊���m���$)ʛ%�
�*���H._�X��~�T��u��Rh�7�=�.���j�j���\h�n�"�-*�	�p`�
�]��V(�����Q��]����OߔqG=���4��6�v���WA�����$i3��S��T3�*����"+(/�uH fC{��9�#5]�a����{ce��G��9�ih�:�hg��k��1��x���k��]�QM��\�؋����nȗ��k��՟ñ+vL�Т��c��J���2���/��i����{��3�X�$AES�z�S{�Y2�,H��B�w�������ۑS}z��c�2!�_S2���!��)��X}�	m�@U���� 9ۍ��DԎZ�Bd�8�\l�@ ��5ށ��ĞCG4��ٴ_%juP����Zv=�]�p�l25}+s�<�[M���Ɨ�Ty<ް�|����C'K�z��A�7ʷhfv���r3�Ȭ��A�y�0��UwRQh��t
T���w��������0V	�����h���1�1U?oG2�Ak���ƃ)Iu\|-Ɩ�����;<g��r!�]:e��� �*�0�_x]b\�98#���c����,Z���e�@e�U���H�*l�R�#�`�dmlX�4Xe�|,�!���] ٹ[�&#�+_m�`7�4��>��7�n�Xz�$�l(��Uٚ�+PtM�ƖD2�s���K��� ��5̨�o�p��^���z-V�-���F�u������t�p���H5c,uC�.�Rq	>��E����?|'��"��A�7���S{Q���˜��\x,�a��mb:���!8�%\ҋL�fW��J4"�A'�h�@���Y��~LϚ.ި���w��mn��r��zɰ��q�a���Ūve�� `t��
��a�ޡ
�~(��H����`���d9O(�^�y��j�4�!�8o��Ƹ!��4���y9~�/6�ޗ����{mք���&�)�i��e��z�=���.|������,E1P��v�o�A�nrO�e�3��l�"�b�8�4m��JJ_̈́��z>u9����(?���a�ܢ�(h�=�U�SƮ�i��#)/h���^cq��e��,���}g���kƍ�\����p�6�ܱ�'���G�����J<���40X��^�]_�-��֌�v�K�g7ځ�ۗ��Y���2�l'`|]/́��]Io (Z����~�`Qm��ww�B# ��چ��N�S��;@�(��鼟J�>�O`>�Ґ�T�,�\O�z0�!ޏT���}���HQ�z}ؘ�F~���d�g���dK�!����d�hCF:�W�W%-D��O�6�{ s,��폏[U�u���K�/|���p�B	R;�X+�:*�N  �E�S1���@�ݖ��cz���da���Ȕ����.w�	�U�,NY�6����~}1���G~*����3D�
k������ҪR`��\x��&79=O�2L��Xݸ�N|ȷ��A�.�N�w�DL��7]ƷX�]0>��@�[���Cm��ޖ��P�>��ݜ��?�%~bJ㶱i]:��=T��y?�v�6�4��:�Q�M�%����v��zM��J��x��9O��@���S��n�0���G�B���D�����tݜ.����qC��Bc�~G��퉽�ib�3GFA�j\�/7�-��AJ�ظ/)�|);���V.j8=�ނ�Sy)��fC�)J}�Y>'h�xa=��MX��J_'���D��IEl#ʠtD����fC��8��N,����#I�͂��`�u��I�9�=��5"����]�H������:�}�r�t*5�S�ŝ�Q�P�Lv�O�l=w����v7"6��˸;�	���Ӎ㶛�sE�y�ҔI ��zC�V�!��ƫ���/E�-�3E/��*�}���
�����eR![�nɖ����0aW���ض/�B�<�q��9�������)��i��,��Bm$�?C�0���Z�Ȧ��YF��������_�$����J����/��lW���b�l����7�ǭ"�z�V-z��_p�x��cD�1^"�Zha�p�SY�_���ya;.x0��}9f����?�.lG,3�["����f4��-��z���������όd�V݈^�{�z���<���+9հ<�{���6:3�N<T"{S�b3�����Ʌez��a{������bR�6D �����r.�
QiV����݈X��+M�z�X~P�"��|��T��I5�[��[�h�Dv���$��5�.�lv��O|SGRdߊ�Sy�Ki,� H�W7L�ޞq���b���D���C��Y<��\P'@��l՛�{d���5tTX��������n�/k/+����#3�o�SX��A5Q�g1�y0���Y��;�K�ׁ��+kkl��#;��Z�H!-Z#�yaͤ��KnvO�E{E���>)ga:7p/���,$��EB磲wʙ�Go3�+C`�iKD�e�G͎�n�T�3f"9	�c/�_�g�����	w�yi'L~Q>��.�:F���F:�3��vA}O�R57&��� ��F�dC\�(����u�h��ne?�m���G\�2M�5�<���:X�����!��rn��H"w�g��>�����x�W�E*��_~fa����k���^����&F�;3٩��4�Ӷ���8n����C���?0RUd;�V%�Z�h���oN�}@�f�\���-�;p�m�i�P�;h0�{Ǻz����P`���&�ǲв���=��l��,�%C-����V�.r{SA��}��_{�^KfA�=�����4N�<��2��3wF�|��&���J�RU �(�C�q���p��Vv(˿�G⚄��fi\3�$����j���������@jJ`�_SEDh����?�th" �A�^'��C�nɴ��
Z��������/��>�p��&��4K��3J9���l+QV�q�+UG��Ϡ��p�7���4v�H�'2�*u�`�ů�K�2ơ�@��^yৣ�b��"�_rA�=#{��n����[8���gڃ�؊��(@�&�Dc{+T�!�3���Q�lޜjsf����4(�F9�]��m�����G�z��z�(;h�Z#�x�Qa��
��ګ��5΍��s��@D�`���m��v�%(�0��􇷮:Q+���o\�2|z,=W��4k�Lֳ(�]j� a&�K^ǟ1�	����2�1�s���#�/��-b��5��K���	�;υ��^�g|MC��Σx6	:q�/����FƝ������u|__Z�A�p	�p����������x>/@���Fl������ �������V�������tVG��q�����")D3����~QF'3pt9�4k��C�r������R �	mL�8B��j�72AD��UBY\�
όa빹.�c�¯u��/)�
�V�	�/��`m秨f7o����D��c��o8H�(?�/�9��c^��h�9p������aqO�
vD��^�	U�#Յ������'��m�]��Ǎaۢ$��p���G3I��U��;D���9���V�_���c���b��|�k��V��?/�	�-�5\�0I령@;�_�)wr��	�(� ݍ����c�4���=�"����w����2��q�pH=mq��L���ԲiLE�Xw�2K�-^% �X7�����A^ؗ�Z�̄��Ǩ_��U�bX�����Y,{:�)(����/uaLj���*�S2�BM�n
���I�]\p��T��I�kk<����r4	ĹpWW:=�UW�GG�nZZ�)iy��5&<n�:sG��L����f%�@���s^��Ug�� MlB|�y�"Zz���'0��[�N��m�z��W�Qٛ��mae#O5�YW��"M���x4<��є����9V����ZD���Y.�V��)��r�

��J�n��c#�Z?7�?Щgܗ�_Fb��1]I%�W��w��O�|ܣ�Ah�)� ��\��4�%\���5�t�TM�c��'4�t�o�]�G.�Z�f83���?�.=�ѸX����J@L���!q����n��F��Í[����'��е��z.J���0l�i���?���]��&��Oj�a�K	y��a:�- *z_pŃ-]|r���-�=1- 1O���|��^��i�,mU #�&�Ó�* �Nk܅LY+��yI�NeS�>�19���Ȏ�a�N�8Fl�r�cp��o�f<IU]�6\7��Mq���wf�t;�C�����k.�K|X-���eص]���`�:�J������.�u��y_�$����Q�5���+�����6p�̯�2ժ��^`�:CU'�'��g(T���H��ǯxI["�a�}�ىd�mM��,ϧ�����M�/�S������q7���4����y��k{7��_��p	��$���i(����;��h��D�a7��vxM-�
��;����-�r�|<�����;0'����D�H���(�A�(cϻ*_ݱ�f����|���z'>�@
"��X��QO��Y�CYW��ۘB�/�k3�K=����L^�H:� �%o
v�.^�hn&i'����jV�IԵ��Ү<��J*��M0����M�Vԟ𖯰,o�$[ZQg�h�IJ��]%��hr~Q^��]�b��x{�j��������~OD# �<O|�u.��U����'"g��:�j0�P�k7�[�G�L	�F�HZ�8WZj�Q�N�@tD�}���]��MȨ}ff[�2�=lړ߀������e���BC�����l���H�#�6�9�
�@p�L�+����d�t&C_�gH��TË�?���!�x�<�`N�\�7��sEm.��l,{|y>` �@=~�^�+� �v��i�na=��r�ּf�����Dma�#p{��'�c�Y�c�	����M���6�h}a�gZ�=� ��.i���N�'�	�����p�]mՎ7%�.Ӹy�,��B�7P $�
r4��`�Z�j��qFg�0-��\F*o;����q
�`�K[D�m�E��o�9�-�g@x嗝M6���6�L�	9�<�L�S��CXxX���Y�.�.r�R8��-�����'��� ��`,��cl����� Ey��P�"����/X�$Sʁ¸�i��]3}��3ņj6i�`��2��@&�Ǝ,	6o�N�߀���x��^/�ã{j��KN�/h͠+CB/��D���~BLU-�}:�P���777U���;�y�Ŀ��:�v�t��ad��f��1�L���.yf���d�<��/�
�ݯ�>�\*t�xl���Q3o0��~��]䘶�g��������l��QlT�,��V�T|��/�m�n�"G��%t��a�8���`�c���3�j��{킍�ѧC7$�YSXŨ뜪uʇ}�W�6����_C�A^�SI^��Ř�~W~u\M�.��<�8��W��W�*���x���
(��XEB{@_���T.�ɂ��1����������* xo������W�����P}��D~d��d��N��]^�So`�+�E�(왞w���Q��f�?P��Y꧷��1���'�C�*�S��A��0�*�n�O��0@�HR��G��4%W�����%�kl̦�xd�{��
n',��%uaw��f�mKm��*-&�`�P��/�#�=7�[�����_��|㸟s�h���͕��t��P#yd/�|O�όZm��M�����������eq�.fz9غzAgE���2l�<�<l(�9��߆퉱�+09g��SV�����B�8����Ϡ�2>b�QL���|t�*E�Bqӌ���y���ص��ᒣ���q#�1���
��p�U>-*u���l�t��$b\h�R��_ksI���S~?��7hO�$��?�����k�Ⱦ7	��M�ϰ���xvZzX��7�|��ڡnٖ�83h���s3Y�0����Ϫ�Q��`AE�#�Dn�FE�1Th��(��Ϟ �c��0%����JA����16���t �g1'��P$�.n��ܔ`��=�n�-s�Ji��	5t����y���=y�Z�'�R}�)^�<�&7>@����=*^���|� ]KO~?�6�����*A�ķv�b�s��_.�B�u�x�3�����D����d��b�5���:�6ͺ��J��oe漠�q$���P�t�3�cy�fC/�#i!�7T�0�ثj�$����ya�^���0t�B0TF{.JƖ�죚e+b`�ᛏ�1`F���A�f3S��¤'Q��a2�$
7M}��Q Oƙ0��G1�C?e
�G˝����V�=�ްЪo�uщ�����i`f����(�-���
=���Ӽa��"�3�X/A�T=���IU�6?k!���L��Ԟ��'2?
*�Ydu��N��L�n��`�S;�i6~�3�7|#�Ue�O7F���<���i%Z����crdc�FS�t%hA���y�E���/��s7�$�4l����wc��n:GV��Vhd��t!��WT�$���Bb*P��������fR�nk�ԅ�|3�2�7�V��{Y�����-J͸^�2L��(7ݥ)��B^o�0uU��2H���!l��AqI{�\�Z#�Ԩ�Ȋ/1�)�9_�?�<�kI��]���B���̵���d�i'�c&#Γ����gQ�P|����)��Z/~W҆J�_�8����:s� ��,؃FA������mG���ն9S#�4&�b�lg���U�\�l�A���@<hD6Q�q�����ˡ���ӣ�(]񴘜6� ����A��$�:�3��
lY�����A�U�aYI+Lj����(Q{vN ��*ܒ��?Z�i��w%_�Xm&�5�B��
�\��D�Y��|ga�h����Д��}������'�u|�p&�pW����`�Ƅ.��EB�U�{TwC������bt�3�Q�sw�ܐ�y�[�`���PhQ�0\_�e##���+M��k���=/��:=|
���Y.;��V2.x��+KY�fbt��[����nѾM'Bv��R~���X᾵,8�>��]�=�?� ���������p�O#{�D捘�gZ�&��eV�-���D��85��\�W*7𦉙!�<W"�]Č~��d�R oY���.������I@|�c<wG��l��j򆼎ܪI�(�xdo�r@R3�Dݹ�ׄ��@fuB�:��!ض6�<�`g�o�d�����Н��3���V�-|)w�$r[x�I#�-��3b�Ǖ��@k!�(�mb�V�V�.K�%zG.w���hqN���c��8�)CΰR���k���>�,iͬജ�DƑꏽ��wb��c�HP�R��?�@��I�xZ�ջ��K�8���� �UY�+��@n4"��c\��[��x����ɍ����{v�J�uBp����y�+�l	��1ě�_L�c}ʸ��>؃qV���V��H-.�|̻�� ���C�k�9iK�n�[����F�H���f�jtCp͓�� ���+1��������W�ۨi�J��p��
K����$�.Z��۩�,,�y��X�%���#�DC[��
��M� v�+��v٣���u2�vOQv�p2Z�e�s����0V������ơ{l+����1�z�#� 	�	�t��U�~\�'Z�f�&sO�?>��d_L7��w>�3�!y� ȖI��cW��ϥ�7����Q�3���(
�m����}����X�
�;�(9�BP��7A�zf��Շ[�ceۜd|x�:I�Q�cp�fZm�c�ZHբ<����N�D��w���鮿dS�O5�3D!!��{��\!�Oh�k>Xm�N�}���)����)�wφ0u�<�������:��j�s�-�ZS��s(-�L�	��?���,9����o�0�$�����
�i�Q`r���Ɉf�&+�����Lx���K%.%¡Ŧ������@�lK�j^ю*kL0�D�G� ���Y\P�w�=�u���]�s���A���%�B^)�F�������h��`c{���V���� ��&S>�?�7u��k}�)��Hh	����L�����c{�^�|kȔjoun�2!q��R�����+XLw	�%�x�Ԅo���4{_��H-��	T5�����$��j����.uK ���ŕ�����k���!���=	�����_9՗�Լi��9ٛ��E�^���g۳���&�-
��މ�;���m��"�a綍���7WJ�0���Dt�&���8�#�!;p@��8��}�����O\
�d�4+���SQ���/������~Io���+�s����s���U%��K�˥�i�Nhxݤ�JJ��&a��[&�.��^�QzU�=��oT�j��qԘ.^�^�fm1��ᾂ?0�M^�Z2��u��ZAM�)^�t��n��^����VːzN�i������2�G��'Q=9��K�bW��)>���鿋��P��	P'�L����� �j�
�8���8�	��ԢQ��Ŝ��H�q���=�|=��1߆{�ZLx`�@X>��\�	�8�y+d�?�����R}�_�j���ytW֑��P�Y���Ib54b��<�� ^�]{���g����m=�!��&���so7N������O5'�eo��&]����'����0т����Rĕ+�@-D�Y�lW�3����25��:U�F�+��2��rJ�D��HF*B`��wS7����.�߳�;����E	����g75�qJs�H[��5�=�����a�pU��_��k���hg�q�^*pL
��2�@�e ��C�f�Yo�%�qbSz��2^]C0����04M�������k7�EКu�1#�׿�bڍ|짴m�[U�3ÄL�(�:�I����]�`:�� YR����\+���,��C��zѓ�N����o&{h5z����)���WQ\�^W�o]OĝB�̴�n�n(�3���c>��MlB��~�C5V>�Z�tbr�h��[�=dW��E�m�6���n��Ķ�{MU��g��xǎ�2g2��όưs���/��nfK&�#t���b[H�C	�1@���R�9�����FR	m�&�%�G��� ��Io/Hװ�K��;�o�S���"4g�c���)�5m��]��B�f4�序�L�:SI��� W�}�&iTeejƬvr��7��/|�W|���o�� juN�N�l�΃�1����i������&ʥ��x5�-C�)"cu	I9���LE_%)Ç:\��r}Z[��g2�݈�
��%�B>h<�ũ,#���]Lw��n�^m�w)�_��֖.��ςW��wO�U��u��wC�wC�8���Pl�yQ&1��\���u�V!/O�FH��M?E�zk��BǊn��yF&��_�����o�k�Of������VS�yb�H�lR`U��`�����3�b��p�R�v�߫& R�Slt
�QB�pǝ�HdXW*CmX�8|]�!��.&�%U�H�w���O��D�2�9�uN����N7]����ճ�"P1��1!4�Cz���\�?ߕ�-�m~����>?�'��yj�m�n���H1���1�;��,�}�=��ᜒu�6b��g\�N���Ւ�`�J
$��Y��)E��W�\_u�2pxjl���Y�?��4���Ԛ���9|Җ	I��������!q�ɜv,�s�<�:5�s-���BTh�H��F�U�V����׫ݺ�`=�D̒@��w���v��7�ޡ�#j�n�3����<�Z�H�k�˸ُ[��Yb��������NT�Z��l$��*Ҵ��j�]$�W���;�n�"	�w�Բ�A�"Y���d:p����:��hP(�B%�R��!���Q&�R-��i{{���xP�z�<:�c1ͯ�BV.icڋy�l#-㩌u	��"��\E�������I�z���F?���O��ͯ_v�O�9�Ŀ�'��zU�ڜ��Ճ�{�
)h����G�^�*���_��8	��q����ع�HB��L��s����Ȉk��&_��ٺā���~�S�������b�ƿ��$2�%<��6W7�Ӹ��_��@kI��>�1%E�%���\��_76��}ȗ�n��8C���);:��w����U/�#�������ιbɈ���q�⾟��]��wm.�D��<ae
U��l�l�K��l6���z�WU��fT�� `�W-a�[�u���g&�+nӗ;C�%#b|g�X�:i	!R�#D�4h������HzD)����l� ^18f��G���)_������{�݇��j�����E���y̻ȥ����g'X�{�b���;�����-��'�� L㍋I�
Y`���P�P2*�+c/�Qt�3��'H�))ۃ� �yl�"�`Lrg=� ٖ��	̲8ؼb;�)�EB����n ���M�%P���>#�E�	v��p��0�C�]�����i��d��O�B@�At����K�Y��b���IQܗ��t	��%o����Y s�vP�T���OΑRX}��eP�%�
�����Z"=V�h�7���Yp�xkyk��a����}�e�:�g��<f�p���!֠@]ԃ�D�o~<Xfa�=��b6{	T�����H��^�4%y��]=�3�ЉAz������1/�k�X���٠d�b�*�}�}�Bq_�`�1�"'�9����^�6ى�G����c�R[�������è��ɜ�T�����Z���Ǆzq�v�n��"�v-�{�H��p[m�ė���o�����/)ۇY��E�ʺ#�}�_A�yr}*���4�z��f96d�D�bF4O�T���}���!`�"�xy�Hr�_-~R�M��% �C-��8�>\@��G��e�ӏMM?fα��_
s^R�Z�`�:�7dяx��$V��S]'r�BL'5��sRH����I�����e����[��x����D���.�o?-����_�L.t���E���zg|L����n����39 �+}`�k#�p�����E�����2X��_*Dܬ0�=�L�7��n+a��i�v�%_7�B��IT0b�H�� 2iZФǟ&��8�{��tAo��<�<����M�m�dbAZ�c�e�{�a��"$s�N��,:���y�q�9s����2@��f�q�Ԉ޴��z��3 C4�`���������؋[E��⎮��Ķ�:�\��b ��9����FNiuM%z�s���Nt�z���2���Ӥ=��%)����"�.�v��� ze���HS��&*o#��zcgq1:F;�D�<�3bF�B�P�C%�����M�TQ��G���w2���&������;�$��cϿǺ}�)��4G����zra��3Y	 W��*��RW���!Npr�0����d�F�!��T�Ĥ�����m�#��N���1��"yG�r���}�qޡr"
dv<���^44����9���цj����5EΌ}��Y��.�1�L���K��"!�o��G]��C�q	>�#M�Ϩ�jp��>�L�&<MQ	�=�aǍK%ul�JI��
�[�t����v��W�������U�F,�)$i�d��'���T�S�j[�^�R�Ț�-*�}E2�G$� m�f�Q�D!�}��}R�yՀ��4�C @����� �/�D�l=bw����M��G��,a���B���WP����Y����&��Ǵ��'��	�ρ/'u�_�嵩�Մ��
�LO�L�0�Q����������(B��!������"�nŢ9��[bˍ���5�_ ��p���'.���p��}EU}�vs������</J��y~r�/�J�#�7#���U̔��qTn�
�k1�0'�X��4���_8�[0-��X[� k� �.;"d;>}@�|�]BY?k��s�l�;���OH��%
Gۧ�+�H5B�����:�˓��i��X�AZ�p�2d�P+J���xy����W;[Z50'�蘦���Q<� �q̧H�~�m3+����V�%���cFV�v�k|�hߠ0�جo��Я&��5g���|��su�o�F���|�C�t-��"Ԍ�\��C�WD��-�/��[A{�tiPŴRH�{��"�����)�J��ʾΎ��JJx�ڋ*､Bq��2I�G��A�f~��¾;~�� �(���.��x
����U����Mt���ե��v��Ff�z*�rL�L��S�i���.��bT
���d�?��}�+����	��-c!pt�5:"��x��1���_W	�=�8<��Ȧ�� �V�]ff� ���lLI�0��0��5D���qY��^�Dڌ)/TǕ�]�Grj��p�f��a?��	(c�ls�����쭒���'�	�1^�@�@M�Q+��ѵSg½ d���<-�|�_��]$6����i�����`�l`�ܸ�6�5�~,�s.5M;z֘��/4觰s�.����}���ʤ�Br����as� :���ඕV�����E8co����΢D���Nq$͉J>����S�ao > SQOL�+H
��Ε��#ʱ����n�ygj$��b?d�J�;ĉ�|n��(�[o(+�- q)�=��tQ��IQЅ����(HL��ϕp�ȵa�L�;�<��2xS�}��������_Yם1�ƛ��}z�J)�0L%��+��^�<���;xO+�i+i�._��1�&��&����y�/݄��a�� �M�/�WMV��4۶����>��D/���8���� �ۑ�,/�!^D�=���A�:���a���3��T�G�"k�8@:e<'�b }���j^'��m���Y3����U��@?�gV�ȝ��	�ڄ2X��7��	��a7��'n�3pc2�L���%��g����j�\5H���"�3���wC�l�ƶP%榉wb�20�����J��.f��z�u�.r�k%�x��Lw�~��#�7���o�����V��=�4�a�RK�$�j��� rr1ͻ��/�$V�3���̱�/��+��;�����M�I��B��cn�w�H�)1x(���;�����oyϷ����%9j���dq���^ԡrJ���km�k� $��-�u��0癷Rl≠y��ƳL|��Yu���5!�,sс��� �T��(�x
�3!�^�P*�y�/&VɃ��!�BmQ1��%Ll_P�1�IߤyH��:��ΐ��ad<f�$���;Y�����b�R-�K<xF�
v+�}�E̮ʩ�9X�E��{Yh�ͭ0�*0�w��p�?j�O����l7U��D+�zѮl�.���;*�����ss�բ������W�$�d�	���ӗ輇�Hثۘ��0��}V�daP[�x�����fk'�k��h�*|���_��
T����]�,�{"o�n�uѽ�"��rs�@(�	��t+�{�(IlV:[pP��l�+���C�o��b� &��Ѐ�
U{x�������X�1Xǭ���Q���C����|ZY�w{ "�/{��Y-����X'���<T�RA��8�c��p�p�_OT�#��D���EHt��6!
1\*�J��P?���zæ�5�[o��$^��E ���)c�B�������Q\E:6�S-��}�?�*��gր35dO�)(���cx�I澲	��+�̼���m@���\�;uSǮ��%N��s555��Ù�e;�m����������LU#�C�&l���FtJ�	:�礃σ�V�D��P ��L�v�^���Ӛ7�Ɔ���H:��D��V]0|J��;ïmS�y*��zT|���俟�Qm��,���X$CD�Ha�Ȗx����c���2K�d����ky��`�������Q
4s��}0����9Ai߱S>\��X4P��\�9F��#�ϣ�3
�?稡���qp>�)<K!�Z ���p��bO~c֚����Z���d�5�AH�d�a�s#�ǂ��77�CzaI��<��(i�B�=[7^@�$�,b�Yn���9<P�Y��E����s<����.ל��V�rܽ�|7b�J4a�]	�@�کd�(�L�%����M{r�뮁��Y����+=Td�ࡓY��ϲ-�	},�/�&��S�H��W��%Ą��ZJ����J�Ǫ�T/�gJ�5ݭl��P^��fH�:a^����a�x��K���G+�[|��+Vk�����b �{�=D�$u�CW�AV�5�.�"�3�C����:���������k��9��:=UU2��Ⱥu5B
��q�gC:.��L�bG�����a� %\���~�IFC'�ǻ�����?�1]�x�~�tR���X/�>���dg�R�gRĿ��Vɖ��E��!AF���=��t���*de:K�)W�B���&2�z��^N1�mQ����+���Pfa��cYvzE�xZJђ�q*��	�فM�KC����۱F7Da�ew=���I�]܍�+�dd�4�}���3�Б��L$�qW�o��@ ��x��£w�e[�4��J67$�����S}mw����	e��-�`�Yg��]�q�p�RPO ����{�ɹB�N�'��2��K�-h�)l��h%Ca�9*_��yl_$E��ܧFM���9]�࣎E��$��;(93��(����XFn��`�6�>�;�K.�K��z�f.�s:m+��3��}�3�,DƧ<k���o�����H!��h~vع�zQo�\/%	�tYq��>�N���	��N�� }����F ��.�/��ݱ�Qfz�]䧨?��k-�Iܖ"1��
��a=�>Z�c���-��:�ځ?J���z��6���������6��CV+��m����B�7s�?S�e5�`�x!J<eQv�$<MYQ���[)�Ay��S�U�����ýX��IF��9a_��U$ȡx]2-�di6�fāς����p��p2oJ����D
����=�3l��#�0(���($�]<ձ�GJZX7�D�S0���+y���A�W˼HW�Fw
	$H�4U�w.��60	�O<�0� @���Y�=%\q2�ӏ4��x�X�?���C8�Rr-:x*h@t�����W'�1�Q��1Z��jkۙ�|��ښ��\Ia?=g�i�J!!�po��"���I�5��&�9�[W�!�3�ĂW3(�n��;ɟd�d���j�)B,�9�>�9XR���Xu[p����M�ݺ��-.���9����=jd�?�":a�Z����o����S	:��f	��/��a����j�"�(��t�:����0�Z�KO7)(�:	�)�=M�KnmH���Z���9��鹆�����A�ׯ�$>?���\u�
�#��������couRUr�If�ִ����7>���r�+���p𠺉
	B{@?}�m�$�Ed�*̍�����h׬�Ȁ6��ϣ4�?M�貈`�ȃ
i�Ҫ��wO��9)�b%nc�ݔ ��~�[y��6�������?A[�l�*�?ql�9ʂ�^�q'�=���uR�,6R� v_b�d�Pn=�T�TCHd�T����"@�wW�u�C��֑�p�7Pk�r�&e����3�b�,�(���T��}f����׍r��'�g$����
b5C�5�z���o�jo2v�����l��������!�e+{�r����pd ��%̚f�\)
��.h�uÍ�Wu��fLBAUJ���9|��q��ՔZ���e2���a|>�OZ��ê�+*��JV�<�I���o7�#k���>L����� ��:��9�a��J+�H�,:��{��,����i��|@4p:Ř���1ԨP=����H�ɯ�ٞ�"���Q~-�z��I~q`�v�I|XU�9/5W�á�����}�j��Z(�)����pq�����g�ͳ0��Π�{�+e��ȃ�7�T�Ĺ�����/^J�>�qe�
�4i|X��=$����ԁX����_���?7T��!o=PXf#m �443���#ڪ
vn��o뛬z����f^WE~�+�~�(lfBW_��T����a}{�iA�۬|�y
W�3J�O���gR�A�Ds��?��I�t3o�!���(����A�5��ΐ��W�9��.����Ju�d0��޾'?&` X̊3��
�KGש�UP���N`ϡ6�9��'���D��|�E���h�<��pKpb
��i�4���!T=�ZyVV�1��8������b�2�jc�|#���էp�ˑ�uɷJ~dK�O�6�櫪BX7�¼��ku���^/�)b>�rm�X��e9���z��ٗ�n[���~��(3d�0A�J��l3}�,c���c�őہ>q��Dߥ�u���&zfq��I�g�`�mv�\zUDٖ~xAtF�k�����3H�����C����hN��f�[ﾜ|-="2�y�̑$� �>V/��;YN�G5v�W`ݸW�߬D���L_xw0�]���"3/�)��WTS��>�i�M�2��ҟ�08�5�F�?H|��z��G�h;���]�5�	G? l�u��ԑ��t��a�}F,}2+�^Q�w6���eغx����Ul�Un|2�2�R�?�|K�1�[��ڹ�ĒX�iI�� ���D�q9pb�v�	���c����)T	�SΤ��f��-�N(��N�W�j���k��֘��O�4j��lB&}b�3=���.<��FD�&���7���%�/�3�
Z/���/]!����Mf���6�1t�&�Me{��krۭ���}ԛ��{H2��z��5��{����I~��	-�Ny�_�=�z��(����Q���NW����M�*�?��������&�<I��@��"�P,��o{�0j�26Y�Uc��q-6b2�+$�Yebr��R,r�>�^v������Ɵ>��f� [�,��G��!Q*y�#fMQ�.� �&&��п�<˓����	�a�M�0��܎�ܙm(���d����Ǆ|�x_v�X5"�G��S*���G�(�ꎱ�SxB�v4�&�db뫬$��=7��7"����T]��!ϒ�R R3�XA����w��:���Ā��Yh��=�b&��/�0��fn�����:�2Fʓ���o���7Qz���IA�hgm�7�&�x\���5�����b�u�N����cY�;�/;�X�篦X���>COr<ym��b�N1��ߺ���w5�泥�[D�<'��B�A��_�	
y�qЧ��
���4��}�k@�ų.�
���}t��!�|�`�^�J���2M�ș��D��"�s��op�|�[,R����,�������"�j?��a�(��n�ÿp����t�E������@R�iO����<!���K���U�AP�C�/)�'���fVl�<V^�d��ha��^:��X�xO�D�-��=�^&�@��1�L�s]U�������V)��+�'Md*��Y ��N���@^ҤVo��hӸT�B��)�4B�>���%��b��օ<��,�
܂I��+M#��Ѱ�$���Z��(�r�=lrv%6�]���.�ޗEl��B
?�A�m��e����U���]V�O��n��c�҅�ˋz���a��!��Gj�;�ک%_��!�o�T���~N�Ma8T�Q�	�[:s��������0������մKP^P��d�&��� W'ͱ�~z޿Q����n�q��4��	����W�YH�^�U��:�`��<�����3L�H�>���ĵ�9����4cP�M�8S<d�K�%x�%� �S�:�xQ��T��xR�F^F���-΁~���@PX�y
�gZ�2hRj:n*K���M7��}�����А�`4��=���T'mSS��������)��0r,U�\7�wЅ����c���C>���?tt�9YY��5�H� +	���|�f5�F}J>������r��c`L���fљ�(���+�1z���b�G��X�U/��2�]QQ|3����r�h8YX��;�f(� '�L�P�+��/*�9�?�3Ǿ��Y �����V#�F%=vIz2��NuαǺ{����%�j��쳳�^�,�T�J���;<�K�:��	��h�By���Kf�G��/�̶�n��8�=�MV�����!��cS����P��]�)��q���߽+��ي��xWM��2}�4����i�nQ��UlAe��IG��Wmȸ��#o-�,�}6��B�Yۇ��7�w�ҫ�q�&���:,3_Ùfժs��9Z�U�r9,���:O�G�:���Ͷ �;�;���>���q���{1R�`�?����l:�~u�]���"Oy=O�NKDφ�=N���:�ҍ��*�ϯ�~�f�=��ι}	�vb_��il�V�tvp��*�:;��.Ի�f�R��W~N���ؚ 6�=⦚����0��p��:(�7q�.��Ȣ3���z����0�l&Ao�8}��L��[jT��g�5�&�q�T����-Ȁ&�+~vu3S��ip0x��Y�<��%�7i	�h�Uj���%�U�&��Ǌ~q[N��F����B����3-K���2��W�������l��6+��S����FlI�w>c����Yܿ��B��<�(x�?��o�E�CU;�
0�_���ϔXly��s;�D�
��c��QN�F��e\���uS^��j���eƷgz\x�,�����ľ�"`]h�!������c�ʠ pF�k���e�h����}~��@4�ad<`q��w�ᛧ;ͥPx���J�|a�E�9��܏6YۧT�ծ�KB�Vnh�C0[��Wêǽe��rDV���Q�7\�.��ms���A)M{q�"�d�����h@�r��
�¨S�&�t�� ��
C,��T˫�	����?3	:�ٙA2�+�n/&�X�;h͕-�;��TO����Z���g�@�y�.�]�  d�?]�o��Ƽ�-ӲX�,�T�炑
(iQYx��<���[,.�b���5���NSӆ����	1��$�j�H�w�uN]AYy��~�1�/l�`ߘ�$�ٙ	��郦K���4 �wQb�qD+�lUH�N��\+��Ȥ<a���.��K�*~޽g�y�z ޠ�Ny���4NO���Zʏ�>2�pK�����fh�}K�H���Ȳ�ёh�E��n��x
*�ue�.i?�Ѧ�����3(�������eB��)�: �]��J �T�Qw/Z��\���,&.un�%���H]L-.�i��,��<-�A%)%D��J�*�8�S?yӂ˵#.�iz��9��R�@�DX������S���}�s�-%�������l�q�4>Q;Q<�a�����(�����̚1z�h�cԂ��J��!����;m�_�.�v�5��F����/�p4-!���W3��[���:�׵U�r؄���:i��*���#ЁA�����0���H_�7�C�Q���z�hQ]:�ЧJ/D��g���q:@nO-�Z�|=el��b6�^B�݁p��Ѐo��Yģ��:!B���ܜ��������Ӝ��YY�j6q9-�K{� ����KL�Z
���z.z�����Y���c��gk���8cU�Ak�;�ƭ��Ich���sH��Id�rң� kb#&�f���,U6�fqh���6PK���Pk���f�s
��Y�Čݛ�(	���')js����e��i�"]��0&�fIQ��Z��i���B���r��ƾ��]�ڴ�[M��ۮaL{��F7�։�%% Wo���Ok�g����`�}���&U#��8�v3c�@��	��|��*�xی�"��H�Ssl����K�z�W �����|sض~���~�{I��)��qI]Ȧ�!��C�u@,���[m?�k�<H�ttAɽ<��z�R9B��ħ����ϑ��>h���:��l��D��s���[ŌS�8��v�l��[ ����o'�p�]��!�ޫ�G4��]40u��:����}���P0>�*.ȡڬ��L#�Ds5���� ��s~)g��H�E�EB*�C%x=ZgKq�\o�
��G�qR�y�7��8*�2ϣ�wI�J��5�V;<� SX�TJ��+���Ҥ��$���B2�rK�Z�38Uu^@eh�	M��l��yK�L��LBU�"�TZ�<說���'B��D�
����y�w�h� Rg̺� ���x���NG8F&��HgX�kK��P�6/�׾�#�=+���HZi�s?�ͩ�Ë�)����-���0�Q;�43���ԭ&-���F�>�7�O|����j�h��}QSP ,���O�m��˾g�L�3Ap#qͦ-�w�(��J.�Km
���X��ܑ
8�[���c�D\U��E���E�!*C3�#(���x� O��ѱ�O,���+�Vr����+�!1��&ĵ3|*x}7
�����I����nӆ8b�2+��B r*?��?e�'�]�x0��� ��^�X�\�LHVY�3��4�zh�\ta#򟮣�hA*l�R���~��'�k�d�<�M��B�ц�m�mp(?~���ح5�@I\�7���j������y��U���6�7���V8�'�Y�_*��	�g'4d
$V-Z�!ŀ�j?#��*��l%�<�]�^ݥl�i��,pyVKnk��3�'.�o��u�|�l̼�'�(�9�R��57y������h��}���p��l�T��(�Gi�L�q��	H�Q@��ɐ�F�E(G["v�0s�U�'S�nPe�q��6ʓЯ/H.��~�UE0_���*�2��ǒzG�X��p�6���Z�a���"d||W�Ʉeaq`aab��"7/�u�x���@E�T���4���9弥�ry�w0Wu53�GS8�u����%�SvT��n*#S;�r����ң�};�@��m��&|y-?��Bﺬ�]"#T�@�@��m���n���+�`ky��MGV�V���i�H/���j�j~;@k��Ӡ�";<(	s3� ��|�)������k]Jb|��eEAc�*bs�Q��עF;�C	m���{?}�J����P�x�Gͻ��3N�݌�t��`�L3�ZU�e�_�҂RI"�4����|�t!71�E�e�3fu��R�zy�����A�b�hiݍU�E���U,��*�� �(��M�uGc�ł�����p�5�AN>��e����ɔ����L�)��R�z\�Z���e���.��@���f�?K���b�����E�*_b��$���>�%���x��)ADu��u�|�A�ZB'�M�?	��,(�m���Օ��ce; ��ͭ�\A$���+��:���$Rq|O�Q5خ�q��% ]}Z�c!/TJgiUNr�}�=�:�W ݚӍnO��!��XG	�P�c�?dD�w%3�L��C�fl.D���y6��,�dB���)�;{�������>;�rsU�[;�
�j��1�mN*r���������n���wFѶ\�4&��a�"@fy�xu�A���_A5��Dļ�Vpd�T﹘�Ԫ�}8as�t�<=݇CSy�1���Qѻ4�y"�6��XH��:�0�qA3�i3�jZ��+*eJ�A�ȩO�v�6���S��+k ��O@�Ac
����34�����$�f6��z%��];���0H�9�0�Ȯ
`R�M)�Ot)�Z� c`�,��w_L&t���4����Fr` �T>ն�-'QZ]�&�r!��j�:�/5����VOP�O�jgpvI{� ��\ZZ��SĞ%���7+~��=0;M�?�\(ߗ�%ߗ����ѷ���Zqquy Qg@#�S'�����°?���R�x$X3�Sz�/���	��Q����!�g�#D+� ��u-x���청3�;�ÂQ�X��k)��>��s��Ds'α�<�����},��&�A�z�j.�ܐ�~��m�L��τW�]�M�&���bfH̦]$s7�A��"ɉv�2"#U�$;6%��(K�:�.���͇CY��C��1XdҞ��^ t�6���n�L/��oJ��h�}�	�[�}�'y>��O���l�E�8���������~�ɼz_����$ D�G��7
�eۤ;��|3)hĹE9����04q�QZ��A�Ud"�ދ�`D�)R��e�@$A��I^}H�)���~�Wטx|HQ�tS��Zb���Y��m�h�EJ7t��t*OF �U�YkOMJ��M��*�|��DdO*7�[� �����7 /2QɡzW�Y�o�7�[�/[���s^���,����P�ra��5��#I�t�z�C�ַ�XU�yڻ����\�s	b��K���c,Y�c�ˑ�A�Z�k/�y�c~���UM�n�p<�E�����\��8�sRLY�] C(_`��j�QݴF0L�z�=��@��1��}}��úƶ5��J�.e����Y���t'aW��e�A�
�40�0>��I<�}W��NQg�Y�#��΄�����Kf�WU�f�#+w>��N*��O(�ͣ	ZGMF1z-�x�����}�A�7f�VX%k�zI�˥p�;�܅f�w��\z=5���_���ꌺ�1���GV�XH�F�~������"��Q���Gz���ը���|~7����2���E�SŬ�X���5vg��T�����F�n�ۣ|N5A����iL�@R�WD.����Fn�>m,"���
�Ru����"R�	�cǵڐļ
�T��yx�%�D �i�O��C��b�g*�SP��>_b�C�Ā�	er�V�H�[���_�|�~��*�����!::�{H�=6��|��(y:���V�*N���E	~��qw��;�kRg(�Q"N���bvo�xZo43f��5}#H(�q?љ�7���<��g<ČصD������ �ߴ�l�TS�1E�Z���@1��|��kT9��t�Q�hfĄC7����U:࿅�|��4���l��T��\d�W�Q<t$�NnH����n�$���-zJЇg<>�����]DEf}@��:�f��2�1��dX���G&���G�PA�&6b'd%���!�X������"���r7��v?���b,G��q�����GXzE�� o���r��`e�/Zq#i��4��N����F���+�4p����
 ���3����p�-��|���d��D��,�^ݽ��n����I�^�h�-ܓ��)��ָ�k�a�����&�z�������X��'Uf��6o��MDp�I�6:�z�9�)Q����q�Kؕh�`%q��[�z���(����QM��-���{�-�q"�w��Z𗝊�Á�t�M�[۝͖=��|2WU�^��Մ.�q#ju�����,,�Q��::l�}�1��U->>�ȥ���'�[�
Qp3#
���EK�h��>�Խ�q��s�~n�q�nӂ]v�%KH�9��#���X��r|l�i���F25���p7U�O+�|h����\�v���L�����_�G���ZdJ�p}��x�5��TwΨ<���Ӝ}?UF�D�|���Ѵ�ī�l����Ҽ���N��B�b �<Y��o.��,	�?��S�`MLb�U�)��qG�����@��Ö̧�&���%����_Z\i[$#��	�\KP���+�
�o�ԃ��S�_��$9��᧡�$��l�V���d�30��o�i;�\#��]�L���mi@�&�Kf�b�#��>�.{��
���Զ���kk��x�j��y�C�ij��;�M%���)�K����H¦����uG	!֮�gț2N׊�~x�'q��}3�ʷLN�'>٥T6K���̼�yB��dA�����'�_�fȚ���� c�C3���1�n\F�Bʑ�)���#�n�d���U�;� ��5�'Vd巀����������w��y�
�%��P8*�aJ����nh�'��F3���Ǥ�Ay.�Z���?� 
��P�����Y,��#��hI�ft�/��!��koʖ�ܔ��,�UatZ�x��N��9B�(�a�VƢKqG1�Ι���"o�f���`Qг"��JS�.�\��B$d�	�E��m.�u���3�SP�@*;λ3!ֲ�5PД�S(�\��B�@�F�F�E���e��#���,�2cʜ�*;�5}�P�sm!)�*Y��F@DT�J�+y�#��
-0ed��b��s*D��{e�C/)naU����U�p�G������];N��y* 2O�'�p���kQ�Q��3�i��l�WJӧ�`7֪J�?��4F��F�^oW��3d�}���O?^y�{���nt%)f���r:�*�H�:@b���r�{�cTs�g�V�����s~�0��kc�9����o>N���M�^Y�X�i�
g����L0���#����.��R�-}�o�U�WU!�5�~�e7���f��G.(����Y,u0�9�������ڥ�(��$���I�ytq`��|*��R��E�kώMv�L�P؂�A4�����_}��g�pçq�/O��&�FyX#o~(������P��h
��y3��?� �"Ӛ
���F)����+�֝�n���mH��T���"��a�s�:Ւ��}�h���f�p��X|���wqt�tx��'D;~����Qo�^6�+<�<b�E��J�¶�P�e����臆��ITdǙ�z�x�W��]��JU`6"��P4o}!ߟ���J���Y��ݏ]PL�c��AugF`���h�&����.�:�54�����!xպƳ�'/dN��JN��p���9�_�~=�CǼ�Mk�.:@	x٠|�z�<�i��;�VA�V��07�'.��ah����qp�V����R)x�,��am���'�$�PF�A�� Ŧ���LtO}�:�V'�^�{C5�̫��:�>��G��Pwc�q +�TV��EP�~�s���-�&�(���6��&܀�X���wt;��*a�}*|��	l/��f��R�3������Zlp��#�����Ç]U}~7S�q���Jb��]���4NQ�{S�z���͝N��f�49֎����j���rMyni�,:������E�M�4t������DY���!8��н�NN�m��H��B߿�ZI�ʖȀ��E�;��.�"L�ӑ"��<j3��-8��������A"	ve����բ���uAӨl�6����Nؾ�*z��8��1d8�`�M�W�jn�Ϗ@�pǙ�Ԏr�I:��yB��>���q+d���֚f�?�u����'�tV.�--�#)�p�^�Br'b����K�� �����%|'�[�]�p5Z�����go�\������/<`Cc#�(TU���3a�h��Al��D�h�5N�&܁*��?V�ђZ(�%� K��I�� ��FI���#�W�=�y��X+��OZ'R�>����.� 㵄�z�~��,K� ��JteWi[�P��{8��.a�8s|��"k���뾣��x�M�7R�����b0�]�!�2A����qju�PHQD���a�֪L���:t=�_�����L�L>g�����o�?
�Q!Bƭ�X*'�EY̳�`���@Aq��U���o����JW3��J+�Yt���տ��_J0os�!��UX���S6�"����h5���V�c�VG�;ۇ�[聬�n�_��Ƣ�z���L����Ib	\R@�)v�hy�ܖj��mTó=$��i�=7�Kv�԰և�KdY�wB)����@�Hݮ/g'�/��?�Z@�����|LЙ�gH��l� ��*��nyl@&ȯ���w���[�gO$�ls��(��z�y0z�ދ:fG�.}�#֊
�⯇Z�0���F/�~�a�RƍЄgD��d��VF��L8�Wh\J��L����P�?
�)��W�ip�j@d�]F�ܟ�����:Ԡ�������x�w�������1M�v�+�l�zj[�y,�&o�Ct�n!��,f;Q��
�WIb\��Lr.�Za�6�Du�7R�4�4
5���¡�7>l�IrQC����s��"�t���F��m`L^���r�v���ۨ@��Z���Hm�h�ܯ�� hB���ŕ��&�ު��۹_�'\{�8���DX��v���3>r��8P@�y�*�
#��{�4ɚK�;}@,�hAGTi!�Ƒg�Z����=��(p�g����&G`>��Lt���|�ƹ�HYu ��z�l�sEj������t��ِ59�=.e��#���������茞�-6��#52�`��}#-:�!�j��Z����x��ȸ��e�VH�i���hI��Ag#>�ihւ�����O�W���l$tIf<#O��̄��\�Z������7z�!��kІ%L��p���Џ�^�'>gflpl��{ǿ|��"����,���x<ՄS����k�`�w����X��ѡl�ˎO}�pnnY:�m&L�R#~R>w8Ơ�j@1I��'�Hx�֡��fS���(DwKё _����'n�$�#������F��Z'Pִn�થ�NHC�'e��T�$�K�;�K�>I�Z���5�F�E]�c���o;BY���/)��P��@IAf��F�	���a�Y(�͌/�
�|V��c�휮�>纨6K,kx{��A�'m�m`U��ߤ���/��:��(N>��)>|�gJ��qf=��W_����v�fIt'���4���G`�j��!l9�Z
.� b�������X������n�H�D�(�vz�#Vvi&��Q��Q�[n2l�	�ɻJw�DH��Ok���B*�̶F/I�CS�crW��ĹC�c0C���C�<����o�A�C���EK'��A�_lte�	�L��	-��}���ke�0_���F��.��\�圇��3����n�)��uz� �i��X��wP�7��k1�S=������LԒ;���T�j��u�M�ȍky�%��O[�Al������k#�I�T��7LG&��0����:`����2k��|�PZ�vF���UR�a���1�_7s��A!���m7�{)�L�ܛ>�Yy�J�āY�IkL�h�R�@�]x����,�s��3_[�oK���D^�T������E��g�X��Lf7T3�Ò7�� gcMrٙ+rG#c�.�Y�D��Ŵ�:���@fKT�$��Z�mj���pُ��GdE6rW��Թ����/,�IK*+����NDCJ�[��@��f3� Eг���٫�N\�^�|^�涣�v��Dq-���S7&:E�g9���).��j��Q���%]�N�`i\��h�#�Qru�(:��]&7�Wxfi�7��+��6����Db<�e�.���;z'Y�},fU���u�!�,��#v����FJ��~`���aG�~��}�G���OL4]���`�}��oH�6~u���,q��� �A��evg��A),@N�er��2X�׻��
tq��f����v�\~1#��K��} Gi���k�g����΢o!]�d�dζ,]
�~��W��,YF���eHeZ�{$|=c�.Q��L���R�ځ�w`���	:�!4��4�_�Vy���K=�P��Z�U-�\���$k�A��ت��73�N�߉9ͣa��zO��c��!鲱o��L[���QGT �	��䀝<�;bBB��p}�2!��A
����y<�~��0������>N��%xɚ{ڥ�3#(��ܻ��(����}xf1��׮ڨ�#F��5��{x�5��v��1�\�T��D�������s�%sO��t�дւ��̿`!�O�����ʦ�H�pa��bU(Zr�5����O	|0���u[��d ��Ü�>�>�eH��G�G��#Mځ��`�?���Z���"�Yf��H?�}q?Ԃ"J���nDż"�{�+��A�D֜p����	���Ǩ5WTĻ�R,н�0�Y��_�}6�.�9�S(Q�6b�1�!.o���2������&c��>S��� d�;���َ4*i/��[@�s,j��kRs�d �gl}��*ӷ?vBŭ���Lȋ4�ǧ4(!\7�P\>#�nk����\�ҞaQ򮪷`f����*:���Ut�dϤO�Ԅ�҅ֆWy"�nߋ7�Q
�P<-�L�r�� {M���������)�j��pu�+7B���j�t�ȶ���y �^��`�.H8�#���̚�c'�[\Efݠ~��܉Y��}��ǵ?m��� m��C�_k��x!��C;�'��;>#�婹��2�o.J�[�I����l���� ���,C+��3���q��
����Kp4)T�&�t��"�DV�$fr��i��X)C�2c]G������`��=U��������p�)�.���_����T\��z�M�-�X�t��������ty���M1� �V�r��B�((ȗI	j9<yj�?Γ
jV��4�6?@��B�"i�h��:z(��t��<\ E��-�֛�'��:U�=����F�zIĐ�.J�5��`��f6�N'B�O(�K�#��i�6���b�{��_��4D�bSUxE��0�<>=v�~w'�T-@�j��A	�����%|��э�T<鿠UR�f��f�	��Z!%V�+�>�W�!���R�d���^Q3P���ںĎ�m?��{��zN��^�'/���GP�>;b���dl(�B�w.	q]��7��V�����������-�1h1�F!"��\�ȸ4����:�1R�f!��2l��y[���/X��Y���ed�T��� SȄR��F�-�b/�e�䰾���ʹ\��9�tl�j�k���g|p1��T�TJ���A��1������ 
o\g^,���БqOf�z��P����3ʴ�C�&9R�
�M�_�̷.�g"��7,O��v�1��ok�W"	^ŭ�.�IZc�Xb�G%�5�S��oNX�K���j����y,��&��)�%��+\A�h#���ߔHG\&��z����!��ت�/T�[�������k�V�10���QEΙo���7�Zk�[8��)�KO����Yf����ݰGm&�FzAϗN��Lwv����	�V���E�hW��A��ߝ��J暴4^����g�[�u�e?���g��yy9P�	t�UbSe��xѻG��AA
�����j��7e�}F�ü`�����-&p�Q��'�J�"�%��y˰��0qF�����^��y�!�W�����(�u�;��|A�UL�5�}v�nI��g	d`KsX^b��ܸ..�Ј�A#� \� �v�6��5G���W�U֫6�������/J갥Ng�� ��3�Ui�- H�Z����~���6^i;S�D�r��`��P��|�
��?�d��:�{!��`N���f:�QC%g��Q��(]ڎ���j��k�]Q�Ew��-��P��k�;�a[�L�JM,D	ѱ�W�Ш�z�{�s���,�C��P����祐��0͢T"r�{i��J��}��ͥ�G�!����O"֜�c��I����v��m���Զ&qMEˊ���7�1�a����S��=̫R̷x��(_�h�~j�or
V�@���b ��? ���ڊ��bnM3���&+��"��HoKZ�9�[j����e�zt�ʹ�������l����&z��Ԫh4����&\|�8������LC�����e�px%v|����Gr���H�(�ZfY[��D��`!\7�G���d�����b�)2���n�7�
(zB	������)�>���7?�����y��p��|e���M��-g��͞�g6�g��@�B�-�B��[���o5�h'Q�A^YU\K^�=di�EV�cY�rh�3��5@��0�D�g|��א_K��nU�$��[�0-��ˡP��d��.�&>a��Q���ɽ���E)y�c�_x<�t�AP�3�6�U-��ԕ���(݉��@�O����#{��);�;��̳#&S
����>����#(oCtFŚ;�.=OJ��4ꢒXK0Yp�(
�c�g�x�&��w�b�|�b��d/�v�={PR�7V�>`�òf�-8��L-��\}����WG_ѣ%T�&��UN��r�B���g�4���Ж�-nCr:f&,`F�g:��N��6�D��Z������iU6e5>[X��؎^���V4%)�oР���o�X ���AJ,�5O�8%�d֖��.g���I:���I��b���q+㯊�Ũ}�sd�/�	��i�A�$�r7j<��*��t�+�:{Te��V0:��`Ԡ���31k=��"ފ��b��-���<1�ș�B�{���t�θ� _R���,��z%9#�j��8 ��#M�r>;�+,aO"3�o�&V\�:�b#���q�ڼ �;�,�!53��r���o\�!d��p�W3�+�,�j/]�)���qy�Vo���Kl�wX�����_��|��o�O�D�8T�2XM~�
�:K'��#T���d�ISDe��c.K�$'�t-_�:4"�/��Px�a +mI5b��K�U�P���	�8�h�{��D)�-"ۤi"�p���J�9pk�,�vv~|�
�� l՚ޜ�ܐ�#Qj��W��ʟK�\��EB����d?��+i��O���v�p�i������,�8*�Xg�t��s���!eZ�{,��lNA��<;/��;	��T%����687BJ�*������"����f�V#�^��v��*��B�F���f���(Dm�&)|ǂ<9J�fY�R�e��`��.�����\�v��P�W
�W�0H�.�TR���ޏx��xk͚^
�Q\&�T��82�}��}�y�TE����pf�ڈ�?�x2j�������Dӽ����G1@ޚ�u���h#)�� ��uƒ<�@.Z����"�yj�B��D���Mқ�����k�ɱ�=;�WXp����X�	Y͌���/�H'/�r�q��{�כ�U�SP;��S����/�Wjǩ0��/܀�9y&y��A��ŷ%�iG��v/ޒjN8o���'t8��%;�
9܆#����:/}�;zDT���Y���s�^�/�`Do+LX�F��K�%��(P��֬�ښ!�#f�����8e�4��h�j��6l~1���ZV-�?}s�W��LS©9�������Y����"-;��2�*ab����8&��2|ks�T!f�JO�� �=P�<�a���1<1�wB7�S�G��M��+��l�ߚX6j��y��qRL���Լ���l������E6��s%�ˆa�<��]q�VZ���1����t��p�[�jӨC�������n��n��������@ .��Ӯ_C��2�co[l-�(��h.+�u�`Jb�g!:�#�)f �*�s�� �
7X�S��!w�J��������`54�3JM�f��ƻ��"[��{�a�)�"|)jm�15ʻYP��sK�v'�I��($e8������=�U��VX̭���}7�d�o�<��̓A�jQ�9����n�C��(��R��%��6;��n��	�������O�S�P<z�i[�U�|�o������6�<�$_�<dX��O�q��k�WL�X�C��Ѱo�������IXMʑf�2m�Q������K$�s;"��C:�)����4�%l�O�J�^L�`x�l�c����;h�>�X�K�iCv�����K܇f���Ċ �_��%�C��M��0�qf��ֱf��`�p�e�~d�ѐp.:�4C�z�_�m��
���PRΫb�H�B�|�쭠/�����/�Z���d'�`�]�j �y��{�����ҏ��t:��H#�N�a�#d4ժ�kV�`G�~���sS>�b��T�9�F���q���t�^�b}����lD�C��o�w�Vt^��ig�x:��۫�?	�&����c���g>�,b`+F�E���%�����]���}Å��+�#N��7ۭ����\d�(�v��m�B�FV��h>;��>�0�����wvȯn>�����W�c��em�s������J�%,wӃ����hVŷ�n;t��0�Y-�&�A��I����}�����/�*���p|7����.���*YNo$��VN�@��Gu�n�e�9c�"��OG�P�	c�=�]&�?��0,���^g���7�\H�+PR7,�9������n���E(�)4�*&�]G`ͭ����<�h汔,;����:^)F#SE�(��8�K�3`T�+6�(0��ܷ
�a2/����{�mcB�����1����k�_m��/��Z�N�	��p�/�c�4!+��r���,���%=)4ҽ>d���WI���6|Ta��%���{ť��l�qع����Y�a֤�˕����ؑ���3���D@IU{�kȜZ`t(�D�6�[v˰��	ʏI�DD`��}��H�`;#v���̞�e)4�>( ��n���ͭ�`���w�7����<M�1X�,+�j������k��P";EL��w��ޛÙ��'6���\Ճ3�m�5Yì������������~�M�LlÝ��+f����g�2iB��L6�ώ P�%�xP��2�`�I�O�3`!a��k#���B�F
�4z�jcI�z/�?���/�O�N���2!yN0�e�B���WV4\��@�!���8B�L��E2����!DnH�w@R�7���i-P]
��Jb��A(����4]�C����.���h�|4�G��/v .�O�-���Zt}�Vi�qE�;��T�f�O�a��J'|�����z�KXy����N��������i_�N2�����ɢJ�Z��(�y�%#��0@���+�׮+����-��e֧���#K��}��[͚���iʎ�D�7_w����v������7T��w��ko��s�vO\�*�$.�r����|@��Wl�S9��B>��h�	 ,�}��y���S>�h�T�8Q���:��g���D	���Р��� �LL�����͠�g�T�[֘E�62 ��Wmk+� ��)dO�\�K-�f.�ɭ��ض7L�&69�]��Ҏ��#�5����$�:G8��jM3?޾~������^}�W��M�;q�Ov\er+�(W���3B�`���U,nY:/G�Q?Z��Z�j)*�h�M��{��J'��Ǔ���RY���a�h�?�n-�7q������,�
Xz�H�f��Z�`&q�D/N_�jԋ$Էs���I��fЕЃwa)�J��]���d�"A(p�֤4J�m}\�3����+0�[�=��h?��KŤ�#���mJnO?\a�,C1a�&KU�ndal�>Ĩ-��l�D�G��~��o\���q�kŠ4p��@8J��9���L�)jAU黆�naM���R�0@���ɑ���H��3)]�k�������(3$v�i�9uw���C�x�B�H.7[t���}Ɠ�.b$�Ѫ]��y�:+�����\���u�Tf@^L�o�Q ��d�IV��[hl��D��*37�O��7�5����
�@Q�=�Cv��Y��
��WT��7v 
��,4��&��s��j��P��35%�M��>r��u|���䒽��ڴF��᳘(�sн%�J��b|�m���`c�ذ��\=cK�!��%����]��Ӫ��Q��#FI���b �l5�����I�.��`�-�:h��	f�R�PH��1����]f��O[1k�y�H��\��n�pc�x��E�A!a�f���'���cX ��K~Ў�ڥGB��:A�͉{`"]��Yf���M㌙��V�U�����{��W����!:��P�-ɳ�rח�*K��'+��G�KL�X���ЊB ��7l�?""I���<WY��������*����E����V]ۦr�L���e����=mTj�Ĝ�<���ym�̓�9��tv%zC0f{6�9͑�d ��W���n��F��@m����A,C�<�S'�̶��B0 &3ܜ��]��й�j�ᄩͅ�v����G7i���#v�2y�(�z�}�K"��GV����������P�C�������|��m-۵�,A@�����{��(P�^A�^$۴L���,��"7rO[9ƥ��`�Wl�)x@'�[H-kG)CW �JW��#D��s�%�|�_2Ï�+z�h�>���O�Fӳ<��[1�ꢥ�*��!��B�G�&���RT��)V����*D�}]S�	���LUNd�"��)���.��w��r� ���&���_�,�����Mo0$�ĐVӃ /# �E,;um�/M�X�܌sAF,������ԡ��KH]�ͮєzTDrݖ�AQw����}��F:���/�_�#j/vDP)������-�MW �0Ƕ@e�擂Gc�)߼A�ǇC��!W*o������#&���Y��)�R�Md	O��{LP�!S�d�~ݎ!ϵ�6�l�C��Yq�d��?�U�5j��*(������'H��^xjm8ݡ,�<]*�pz��)M4Fr*�zJ{�A5c�EWFhYx �rvC���3%.T`7^a��������I��#Zg~[�=s�62��#�k�{73���.�ګ����3��N��ʑ?o�q�X�,ُ�P`ޛZ^%nL_��rP~EĈ�Y%�A@�~�VF���ʠ��H��	B��ޗ�$�^��d���l�}[˪ş�]Ɋ�^�58i� 2�D�/��7rh���_-3��-�]DqL})�� �|���OD6��B2�H~-V��hj&s���w���N��d��b�]G�ʊ���d9��C�*50��iB�N63_��(��@����H�=�Є �0�-ˊB�6�f����`����vV\���i��̐���nÔ�
�O�J mz�3
�K?�Rlz���w��a	��:���?VO߶�$�R�.9=@sr��ǣj9J��6��*;^MJ�!f�(������pR:q-e��'-����c5��Bp�Ô��5 bq?{9p��\J�����y����૰��!Y�dj)���Eie���vpS8����$G�*C���+�g��L���P6�������!8~A����2S)`��U���6�ǯE�o��>|�.�G�c1�(�?P�p-V�펣�x�n���3GeS��+�'���>��-�`&7(w�Рa�I��W����C/��֐4��ύfA���I��.�0$ڠ���mp�aɜ�2|��"�$��|t��J�t� ��͜�-��;�cTu]Q#�%iB�-��C[��(sY5͒�	��6�1U�s�_�xp�H���.�R���M�EIJ+F��yYe ��s�Js�\)��8�b�2��^egޞ���c&r��DU�&Ac�"�� l?eX�v��"`G=5M�dj�>�K��"]�֤�EH�Ό=~��2����`��u��3'�د�'!݀����gh�r�����| ������]T�<bT�g��ԅF�%��ق&�I�"
))��@JPO�^nIxg?V��Fw�p.v�do��>XP�f���qn�H�(W����D��ǋs-�P��*ۂkP��I���x3Z޲/�&6�(�\:��*{*� *Y�������,�J:��9p������
@����M��Ø�VcE�������������Ťp��M�	Ql�o� ����l�,AS)�%����:�J0��EJ��+)��%C�Ax�Y����#�S�[�:,e�?���.`�L�5���r��Q�],��	p��}�G~�`��@% �LT&�ە��8�:�)%��ADY�TO�Z$�e��p��w)���]`�*9�H;|s��|t�ZD�bI�մX1�VD���� Q��g)�LKj�<;�]���	O�9٧aÉb�@��� �w�s���I�i�x"S�
�B���VJ�>X� _p�.�3� ��"�T�T9L�z�D�0�񈐑N,B��`'�M�%�8y"�Mx��:|�N�Љ@�WJ
�4�f�D�U,P%?��C(�R%�+g-��u�s�D�k��dw���=P�TQ�O��^�P�Ph3M�a����:ϰ
lzK"畨�L�0F=#�����L�ݫ����X̶8�Qa/JZ��,����� �����1~�4�8W��lD�������ᇔ�~ȇ���xvm����^���u:�?Ofc�����;��O��R�#O�~���Hڷ�R�0��Ev�ST׳��c�!Ӳ,�B&g,�I]�݅�Ļ�EKp��E��K������}���8'�b�H�t�\H�#0��o�#K=�V�˙-v��[�����;9�������E�`���>3�g�H_���#˩ӁA�K�'P����5��7�4��k.�	�4V5�J5�pw{g�)jz��Kv��&;:�%W�v���d���;��ϕ�c,��ۯ���(k��p�Y�ᗃwC�Aʷ�?���N�t²O��6&�rQ�N>UU
��ۻ����p���O½Q���d�W"�i��C����>�����4�m$Ȕ�(6���X�sP`��x@pp�+mu8Lc�d(ޏ���f��*2�%>��|e썗�6V!M��"�9��~��O8�zܢ͛nTa�8Kѱ��/��k�.��o�x�WE�@�V�.�����{W�f�)�DSH���Q�з1�Ws~�R�8�	��23�x
������F>I���ϳ�n�kz�g��Tj;CV����᜙gS����[����S��;�V��Gj�����/|�Ӂ\��)�����LES8�]�x�n�L�e;�8�N��j=D���m{�3b�9K��p���Vb'�Ym�tZC�' ���O n�g�yc�f��ufu��dT5[��M���,m5/0�a!�B�L��ϳ�^wǧ�v�zYLvP���dj��j�Z%��eo��3h��$�����rB�=�O'
#{�Zde��B�gn�t��@0�xT�-���x�%��>�%��~�L@�Oa	�-"!n;@�:�w�2���P� ɩ/~�9�`�+�����O�47�-{�}�ڼ�g�>�Պ�yqyC/�SH��>Y�w��Z�o��k+/3�	^
 k���g�?}������6kak����ڍ��.�y5�(~�Qg��A:\��X�`}�p�y��f�,��w�l[ ��7�NLx���ڮj}�Le��d��}��JSZ�.u�WKAˋ7�s^XM0�������"p�1����|ޜS��+��n�=��%�+������q��H�底��B������	>	8X=R��xa�H�@b��ؒc#�f06Xa �SP֮hn"?+$i��%�O�U>���z��.�M꩏j#7 �Wcg���J�����?�t*p�To5(���C�R-����#]�	 P��C˵�:F��n	���@����")p��[ Q��̬�E엲;}K@)�����z�訫C�t�b>�_��0�i}�9Z��r7�'c�p���r�����7��EW���$��	��h/v��^���f� ��*�~<���Bd�#�|l�PJ[_�P��س�w��imozx�O!�6H��nm�slj�R�EUz�bL�uHE��MF�v��՚-n ����j��慹]���M���Q�����7����������-�|N}ed�U.t��	�g;H�{b���
e�����A�<H1A.uw|.����V�	��˙���EK�
�ܽ~�!�)pGQ�\��fk�]��7�p���B�
30��n����F;n��ĠCV�b-8_��z�x')�Z�<rHh������5-4���Iϟ���A�w��E��~z�E3�?�?�E�c �M+��a�$�����S�@�	���ݲ4��I�,���5���G���w ?�!\��8߮Dc̋�aND���T>̓��) ΥE}��ak ��H�&Jw��&�>g�������������HH.M�w}�ʇ�����N��a�e�L$y�v�}ɛ#B����<$�B�q�JD ���1�M�R�'��[����=��3W�Y����9E��m�zQ��t�3>0S/">j.%��-��V���w��o�q,��>;[�/! &��N��/�B�[Z�x����^�V�5����e2�0ӌi6tR~]�(��}�4V�'��.g���&n9�{��0f xn�\f�UI�.�` ����N�Y��@�����,ZA1t0 �*S��04=�b34#U�`������B��f��Ə�]��}�k�	P��_�#k��L�IR}�U��Е��Ȏ�@�*}�Z����|��'q�B�G�V�>>���+f1���1�?'U��ªMn�U��h�Ij[�<�n��}F� ��.��쮞Oi�Ֆ|r|>�<���=��jJ�f׻#g�(=:�s:��S6� RNZ��P<V֧i9�����/Iz*����?Ԕ�uz;�5"��},�l�p�[���ؤ�l�イ+����	~C���M��L��/��������������a
�����X��e�t�[u ݼ��^5�V�gď�,���Kj��3a�ˋ]ZI?��\��o�I�,�;q���Q�H}��H��e[��7�i�D����F�0��nE~��e&���>�/��?�э�9���:u�U�PǦ�	F��E�����������n}��O����o��m
x�=W&S�6���m�-`��-NZ���7D��f��3��P��B�{rX�=���ڴ�ߠz�e��ʆ�����&�덹�Ok�݈��`ô�v��e�	�+�$xO�M
=�:1X��o�u?r@�8ߘZcs��)>�OB��0��_�L�F��x�9G�G�>�gնF#N�rh�gc�7P�F	�%�����n��k͐�%1�ܑ)>,�]�gؾ�Lu��,*[$��v�+�I��G]^�%I�n%���+G�	~�~9�0�Q��}�	Q�y�0ƼJS��)� ���M��Oy�=��I����|s�\�n�lb`w��{�G{�EX��i8o-@Ջw��0J�vn����̫o�!*��ʷV�4����6�ՙC�@6�Lsa�6�<��ف���BeFBu���;�����O�H�@�QXG�e G�bIŠW�Vn�}��1�a������F|�,0��LtJ�"X����Ǫm^�q�T ��1	�{�?�{ O&mO(� K4L�d��/ W"`�0}�Qۤt`"r����֪�b��ݢ��l����N Q5�HW���ׯ�Яh�=ܸ��K�뿯�hH
?���L��
X���&|/C/�V�v?��|VIF��т�n��ٙ@@��"4BǬ��&,S9�T�nl��R6bK��`m�h�Y�e�M�5�aNj������&��ǵT_3{�J[��m	�J�ct0
JȰ1����͂�Fu�$����C�F	ٲ�hDg���P������n�R��8��F����]2j�5R.�� =�3���K���G�nX��L���	]�ad3�t2���l���=����������M7��syIpF�C.w ^��W�JCP1�݌&��9N<k��=n&2�X{�ˠDk����AI�Ȣ� ���Sc�$��� �c�m�_�Ĉ���f�t �
�97#l(cca����������/��i�	�.�:���P��� ��)/�JdS��Y���Ј�H����,�F���Ɲ�Ky+c���)� �,��U
.�օ����1��.��K�_x'a律�V��^��߳e:1��,��m_zŹ �Jx��ÙK6�N���J�]6��{�r�bTyz��!�t�2��XvV�j���v�߃,����e����G妴�o��#��N*��rk`ϐ�d}�+TA�������)c^3���"hҧ��i^���#Sx����YR@��zy�MTc���[��/����r<�;d�����~��*Yχ�uf�v��W�b����V����,��hԖ�7C�bG��Z�L�m���4�:�j�&Ke8� {��-�,7Ga��7V1��Z�(�3�Άg&��lj���Y2$^�!�p���gP�����E�5>��"r;�D$	=w���F�ȉ�m�����D�+&��x
��-hH�� ���� �1㱞�l��i�x</�"F��B����s�Wrz��y6��X���~ݥ�����o�O�֛F(���G��Π�E(R_aB��uz�.�8G]%�.����e�;*�O��>��ܺc�Q�r�`DZ՞����Eq��/�IzX�m�f�?��6�QUL��qW�pB��� �s������"G��vW^3�"���C ��&�j�F��ﾷ%��%Ɠ���%���wK��ؔ���~p �}2ZR�W���V�H1%~}�<-lP� 晨��~q�_��/.�<���'p�m�V�:�����y_�93+сǜ5"(�<�(g ��F�	��F�[/�'�חYwX�4�?�*�K 	��Y�y���;���4�0��=6����ԔH����D�bx�x�x��i!		��ʾR �x��]`����[��F���T�;ڡ�-Z���e�}��ϣN^ާ��+{l=�+=��8�hV�N����-.����Q��Id#:�Ì �����rJ�\0{�%��\�Ԡ�i;?"k�IlV=�Q�x��6�q��o"5#J)��{�`�H"�����{�g��<e�Ų(�>�,tp�﵍|[M����)�op���V�W���%"M:r�����anle'>�����^�	q���렛�N�їc"�kQ���p��Z�n�o��U1>�H%�b����i`?t�������Z�c��;���a���*�H��Z3A8�y:�<y��O��cR�4�_���UE��b°��1�[����m+��֩��`��`G<���>�m,~�������mH���C�Q�Y��r0��b�,:�e\m��;�P��M�9�h�G�v���*�O�p�~ ��re�=���	J�F����̆��ZBZ;O�:vխ���4��sA�r�X+S��]�`57��!����w�LT�nR�X�08��R��z�`4�b����2�f�)��]���+�F���*���V�|�+��0�GhY�C&�a�]��*�{��\P�;�E���՗��K�� �BUS܆Q��!��ٳ[b">���EĉE����:���	J�%$THE��陱�UFƶg��:��*�L?M9%D�eI�7��`�Ai<���lrޔ	�郎���ɂ��[e�U|=�o|?�7�y�9ʒ2e��ۑ��]��.�C���ѣ�z�n`�	p��l,���[��R�ٗE 웳��+s.���[��*���f)� #���e>	or�<�/^����`h�1�g>�[۰��<�V��9�L�\CU�s�޿
�ZLˊk6Z�O��@ 8,��z ��(�KN���{z3y�%_!b~��=L�`�2
8�n������/�.��J��L�/�B�8-��o�o�S���dP�4�:e�&�=�m���=�j�'�+��)KHS,��nl.]�!�G]�'�L�O��Sq�oU� ��:�=�h5M��d��\��J���xD?�'���7@W���7�ZݪξB�v����M��{K�eHPҲ	�u�5���E��C��^��U+����l_�c��n��+�M.���(�J��@9)��^��K,��V+k�&���L_+)K$�gkԢ�M3��W~�!&��NI�uW>,P���R0zbUU1���/d3�?P rۆ�Ε�DWE��ڲxrs�ޭ�v�r�~K�hd�8��;�6$"�=Ƹ�q���(ȷ�d[	�|�P������,��^��b|�?�P�03V��-����~@P};�1� 68���ۊ��P=���{�'jy�DMC����&o.�Xc�:F1s�EFʒ��Zl��0!>n���"9œ�F>z��n�J�t����<~�_�U����@���Q�x�U���]:��Y!W>�A^��5q�_��-�L��c慔�A���h�������Uv
䯥s\��t�Wx#�?O5�5�!�k��*Ype��S�	�f�O� }��e�I���j`�2����!�@�����g
��~�����;�^��{��l����������G�!�Q!��H���Uk�7?�P�Q�B�W�$�}y��S���118�-��fd3�z`��6�z�	��O{��\Y]�]�������<��8k�v3����־����C�lɳX��Äp�\�涀��<�g���k��_y����C���l"F�Ȟ� 6N�,Մ2���~�c������W�3��&/���������ߛ�3��W~�W����m�_��g�?7������p��U��W$���J�㵒�$�:K���3��l�o�����V�6�A
 vn^�4�I�Q]� n78x�>��{F��(�<y�|�DfW�J����%a��q���Ӹw���n�Q�OfsTJ`���:��s_ gs��c��?{&"#�d=P-�|u���Dصj~j6�1o`B?��[�<ͪ�*�u�WrL��F6���z���k��5���Y6�a�D��*ީ�:5�D_�6&���s�2�U���� DN����&�r�������������=# ѬlVB�`����F*�­����z��0�$� �E䧆ݕE1^�̊�c��9���=hlD�ή(�7�齠�����..<���X|���Su�Z�Oj�9��m�����$f��Z�cV��$��hh�v���D�x�r����Z��<8�7#���<�c�S�w��h��Ԩ��V�w'u8���[�3M���a��ٕ_Z�t���B�w��϶@�b���S{7�vETÌ��6q+�W ����B}�Lby��vM���&�M1���b_:p$��ZL�]Zd�� a��3�<��u���	����*��6�P��KJ�qiH< �'SA\Ѯ���!Qc�0гK̄��D��2�J,�}T�`D�?ׯqp�'�t/2�A�9�x�4�\֊�L���MA��?�����-���H�Q%�xr*��d���cY����z�Y��Ml�b��o-�\��=�HK"��q8F��d�@ v��� ���wE�Iں��U�u�+��.�B�����-m24C!㤄�M��ָ�wk(�k���#���Ɵ��P�r<��&=�LyT�$�{��@�u���_ ʔ��U�5�u']���(#���3S�K��Y�7FXrd��u����.�,_�%�E}���` �tޜ��}i�5��	<'J��*�꒨gxKN'� AT�r���c�\�#���I�.�mR���Һ#m���x8����=IU�t˄q�&�h�2b����~YP;�g�|Q�X��hcl�A���K�,_��o=P�Ψ�4�؇mz�q�7�3���n	'c�\���J7��^�zKE��K��ɺ���J�J� dj̯ο������F�I�ˮ�/�T��#�����
V̤���2Ijk2mt�j[I`����J����"�{:ޓ�%h�a�tru�*`����08Йtc�����o	;&���g�ފ�i�a��6=�߼u�J���>��O�|Щ��)$U��,���:�
�\���-�����8���~�-#���}y����Nx{Ie�r~P��^�H�2z�����?�5�/�����_��Q'f�\Z+D�w����&���,��T=M�;�^�y��}����,DPOs%[����M�CcU��z:Ff2fX"�b����f�zc��l��j��(7Dw��YHgİ�Չ���
4� PMx�EW�4-"'� 4�u5�)��0�S,�X�Mvl����� 6�*|C�l�EI�p�R �Nv���4hN����g��z6Q�;`8�W!�zB�ǖ���D)��NڤeO�������S���:�I�!S�a蹕��\(ǫ:쨧�^�H4~�F6B
Zoi��\-8�xb4j�0�P'O��|�����M*AC�HY �r�	X�\���3Rj{�gQ�8%nњ��|�l��ç��{��O6k�}�%d��O}�|�돬�#��2��'$t���&���Aq�%a���Nvv/��62�n��y�l�cl��Τ0�:dH!|>�K��u��\8�5��O,����r5S>��/�Vj��?�}�[��r�]6fۨª�Hg��h9��f�ѹ�>�Pk�y����@��)��[#���(�1x���&:�A�Ŭ[����l��Hc��=���Ƃs"��i1�X�C[��܀xfId�똪��vΡ}�R��&�?}ǔ���0krђ���x��A�Y�2s�S7�z tqغt�Z���a��|C�敋� ?��X��0�?�\P�@�;���}*�U�S�fڬ/��X��;�;�Rv�V-�-�蒱]�c����ҡlaw-{�~���2�d�&��S�)�#78d��6�{b*	G�,E������ns.ŌNP+['|18����J�"���z�E;�+�*��|��'����i�X���ϫɳ�OS�'-��@|�b-|T"f��f)b8Yꩁ�T��\-�i �^�%�|����96����A��d��Фq� _���R摒2+\4*��
:
-�c@�����N�t���Z<���_�oa#lp":PY��|���t�#�d�fNp�4�;�;[ �}\�QT2�_P?E@[+��(?���� _�@��T�>8"� �_��oJZ`N%aJ�%ò&N�%hT�/r�Gj~ld(�� ��
�@x���A�NO�PDV��>#�B���'��6�K�B��4o*��?jy�|����0Ye�@Ň�v��)��C0��#�>����	�ۑ�F��qՕF
'��T�lT7f
�ᔳ�-��_�6�A�3���B�M�����5Z�
#���{�|F�����C�r�A\wB��C����S���(�S��x��$Z67D�I�^Ɂ�N\݉�!��Z�eFO�A@�������f����և��a�����B}��t<�6���}�-���y��4�l�G����J�Y�qo���A(ïO��j:$�'I{	�wʍX�@��ԫ���
���|��4���w�{���ɾ�2pѕ��X5������ۊ���gx���
����$�;s���	L<��;�=��������W���2�ƌ����i{/8�̪���j��8�����&�=�Y���q�21�Wj ?n�ߗ��Qo��[ci���u��+$��k��Q�K7�C����'_y6y�{�������_�|���Nk_�s���%*�S�����^��j�~�:��feO{����N*�義q�yxb�`���(	!%�^/��}/�DԶM��Ku5��t �V�ͽQ���$��᛿�0�h�@�=�M��9����,�+�̷�S�]�C�e�YBh����<��6^Oy4Յ�Ǻ�����V�rqU�͖�T����$�<��fh���L<��%>�ڸ���$���Z\wΊw �W$��2����i747$_�_�V�F��ov��6�+�~����T�(] EW��Я�}�f,J= T�i��˙�N}=��Jm2��k �#:�|[�6����9^���l��QRI j����Hm�NҺ�ΝI�7h�6��JX����f�w�$r #L���n�W��آ1 �>/ˏ&���^�8$���^A���_��4�YѪ2+���(q�]��h~��� CL�=��.&k����k�P�gV�D���y��PW���vG��������%������A����Ǽ�nzW,�s���|I�yJ����?9o�D�\X'Z��)�N>��.�O>Ư�w���iV�GR���LN�C�|�js��2`��ޡ�K�E�[*|��n�}�NԵ�����'4��lX�B5#�O�Io"O~Au���o�>�wV�(R�u����'�(ʢ(��e�G�ov��n/�g�4^:�w�_P>_����)A�D��dB>����,�����H4M��îމ����"��!� }���j1N�L�L�֥p��H�4@���#�S�OvZ0�1���~f��'X��8Txy�tq��C~���LU���P���),�A��NVbWD�<I�å�є�Pm>��������s�֥ M�WSķ�Q�'��	� AX�'���(�m}��Z&9Jc��5nAl��@V�!!�Z!�;�Z�|���:�=�z�-�UAI�B���Z�a�h��_�\��^쾋�(CN6m+�	��v��j��!T�x�܃��4`16�����il���W)�Jy���#>��,��ug�@ƪ�;���2��i�>�}�1��kK��@���A��v�R>K��Q���QW�yN#�nT�����{9��� 7y���w�	��I@�t�Q��*��v;}m�A�N(���MLGi�hA0n�R7O^"I���8T��"):CH�b�5ζt������ܽ@e�Dii�Z�d�5^�V���N1FX���㌸�k�먆;�T'��*>���Nx::2��H�o#�����!����e�5� O��х"Ҳ����؏��	㻌��܅��pe������i=��p�ŬVi�����Z8A��i����fq;Z2,���X�����o��<qf`�?��G�|�#�t��28�y-Q�[2�h�%��ȵm�,%nބ�#�0�p��1���P��8���4��0�菸/�2��χ�I�Zf�V.�2O�n�0���E�=L�'���P���v�x(��m�mx`�s�����P ��SY�&�)D_�ڤjg����SSg����=D�d C^��Y˫���sc/e��Q��V:^����'���N`E��<� O��K�ʵ~����4��<������^�9�l���\�߼_�hFT��ά�N�ӟ�)�Ϸ�@��瑕�V.�*Dr[����k��~���1*�S�L�k��ZJ���ÿ�Y��)6�>��+��H�5�$���d�u������q�t��d�@UkU>�P�D�/9j��#F|��Zm���l��:P+P8��I�U�j����|]	����p
��>2��#���C��ƿj`{��\�09-fr��B������{�.D$����򛁎�]��~��͸�ձ0����Q�j�y�	��*����5G�Ql����:zB ��\b��Q�:���$�c�A�6�(/��hL���'i%d2���oW�햖�p'�tN���Q�ZƸ�m*O�e�� YLB�H҇���m�N��i��,��Ҽ8���]� ;��tZ�� H&C�-#��聱�~nc5�(�qv��^Pz&EJ�i� X��w���kJ��P��E_/�Uz����9�����		�������ĵ�J����6��ߺ�N�١�/�A�� &x�r�,�	Sou�`�'���������l�R��&hQ3���d=Λv	�w�)� �Qfj�l2�5;�CȊ�x���Dֶ}�E�>�� ���z�Q�'`|��Rv� ��K�S��9�̚�i�Ϫ�z��l�Z7'�Ev(��Vѽ��F�J��D�����
��V�5L6ofߵ���30��}�Af`��2��s	D��]ٲ�,;�����;�(���+�>���K��a��0���/�M�'q�d-��~��h�MG�s�t��S�q��18LW�ő� ���Z?6)5qp,�����P�wx��O3���D��@�i���"XF�#Q���模ڕF���<�T
$r/��R�(3�,�݅2qnwd -��*m�t��b�s��H�gH>��_c���I�Tiǯ7U���M<���IP�Y�!`����`���~��|g��~/A 5�6!V����I #[�(OJ��۹��GM��.
܇���'��ϭ �%�#�.6[���&�z8mS{�rI�Q�M�^˹D]
�M���>��Y������+V�C�{��6Mmp��VT�Җ;;ιrS�`�0
e�|�f4�E�#:mI�E����h<	�/+l�cP�����W�>���%Y%�sy���\������S�AkƮ��%tW����L(d���`�>a��i��Ĉej�E��&�b�'��q��-4���5��"B��T��%��/sq�e���0�]��Y����2�>��ugI
s����b,�n��L9Ȣ�{
�Y��_3FNx�$�sV��,�D3%�U�PP%sBrg� �p!��E��HK�j,�s�`��1u\��U�~L�l�� 4�F��y],8�*J2	�D!�ʵ�� �r���=��ν뻍�5U���i���EtNU��ҷ�tX��>K��sY�g��O���(9�.�7B����C]E���S����|d9>T&'���u`Q�����J=�� ?8��[��Rm���>��l�8{V���7�r���؁-��u�f��#Ƃ�d3G�Ac�s�=��p³�-{�7v���ח��)�!�^$L'Dp�h��q$�1��T	�W}<�����o��(I�ɇ<�c00�Uds�9;��w��X�+�K��<m%h<�8�=��d���wI�}��|p�	}$�����Y�W��f�/���Ȟ����)8pS��Κv6j�<�o(4�o������r��C� ���@k^/�GJ�i0����1�J��W^��ay@mL(n���.@E r�S|`u����hdc ��h".#
2���b>ٹہw,�KG�%s𰒪��0����wݏ�p3Z��݅�9��Vsk;K�'��g���-�E7*��o��q��ޓ�j�"���o�{��ު؟�ֿ��$�bJ+gmKH�5��$��Q��J"��Wβ>TS�~�g
��G^�l�:����E,����3jR�O�|�3}�U��LfYU0h� I�b��7E�x�=�7���]&�����h��L7�On���zo�K�L~�F��J{��%H�qD'�����fsT�w���I'�ǻ�MY=m��!��S���F
e(u	�|_d��U���a�n�F�vVTf*@��_�J$Љ��lu�����*������<����@YX�en$��wyn:꺯���OZFʮ����x��y�AL���&ZO� �Л"�`�0'��Z@ ���f���M
p�m'� A���u��^ٽ��ԘO����l������䯑�@<�߫�����*��>T	��Fb��]��Oq��+��x��1����)�@+�O�ÛU�8��!ݪu"5��,��2
ܛ�^��,�:#Є�=��e~��N�x}�Ҩa�l	%ʡ��<�;��K������^��v���rN
m���h�%��a�5I��U�zx�y7T�*�:r�,s�0��Œ��K)FHGG�$>C6��^��EK(�`�H|�ɭl*wuO�����*��/뻆��� ���+�F"��.y@F�NЂP��K	������¢�ve|2�[AdȖ{�=6;�Oz�_76���y�"Z>]�1�� ���2F=�MsR�����KE�6���1%��)q��M-g�B���9ҫ%��B/�A���dػ�.O�2+a���<�~�Q�7�[/�3��� 3�#�9Eg���6�)r�U�A$q@b�/}A�������*c�6ن/�"ޭ7g9&?��O�~��)Z�*SP� Kሢ��r�N6[M���
f욆	br�/<eO��k�y�[UA��Xq�Fe�?	O�{ȱ(Q�z�#�ᐌ�I��Ë��/�u�r�$���!�	'��ɱ���|�6zM�
�X��$�^k�K��"��O�������Т�_۱{Pnc^w�T�C����8-��Ç���'W�DPق봧�<���휡>7>%�2��Zaõ:"��h���Q�Z(�L3�<P+�Ί>�P�����>��n`��oYԟ��LY����_~q4�O<��Q���,7{�<��L�t^qhq��!h�֓�R�����l��I ��H��@�+Ƀ���8 �
����Y�aŘ��Rk�������J�Wp��U�X����#0�)�����t>î< ��~�,U�eF�|J��&�Y��l���ɦ�`�i�$냇6H�0.i>`����G�ys!�1e?h{0}ë��Ҷ��E��C�� ᷨ�����p ������f̥j�|#|�8�������,�v�� ��S4!8�8îq�K��.�a��-fx�Ó����m/jb�;� &i�d�y���65$�Q���c���X�#�i������h.7�oI#��鵁�����ޡ-�ص4>�7Y��D�jw�;�)��Z��*By�&��`�ܰU��-�����oY� ���5���0����?�9�$�Vڇ{4�V� w��2�w���,�KK�ܷ�l����V�����{�2���P���7�U��NUÐ؁�u�6��Q*�\f���Cii��R��Z8�14��\H������+�,_AJ"��̼��q����,�W�ߙ��������i���	-�A�/G+�+f�/�`!�� �~g�D~P�~�P��j~�?Tt���ܭ2�����I�x��{�꨼���Ώ_J5jƗ,����7	i�1�?#9]{�ji8��;��P�����B܊ �"���,�*�`<���T(��5GS�.{awD��pY5c��A�,Byp���a��� �Oor��� ����	�����|{��B z�"Y��JHR':���3��}�7�q�t��X����) Vh�,�v��М%p�7Q�lF�}ھ���d�Jd�s0Mm�L�1Yk�5*b��u����]'��a��c6( ��Xř�uy<3Mdq��x5Sw�C�al�o��1��Z. ��]J- 7h�^$��$�s�앎!��>��v�ܬ�	,٫��ʮ4K&���^\?�C�7s㍜��/���Р��kg�o\o�N��u��D�(�����2j^ ����!�{�/L��&� /L��R�_Nm8)"[i�TRr�=w��J7��a��C�"�ϓ��R�E�b�P�Dc�#�.js���m�S�<q
��V�(�m��f��)��G��ձ��!{4���=EF1H�; ��T���xi Y�(�Y�A�Q�#�#<�4V��Xhw�ݯ�~�Vǵ?��g��ʙ��;�������]�r���x�VR[@Oܣ��%Ӣ�JC���H��*ECpd�̸��I�Ԅ�����\��l�P�T��d^�Z�	D&�{@��+�7�\@��flp�)��$\�Q�kXD��z�dc"���⒕�R7V/u�T����k��JWdVu@1nj�Y���o����.H�:3M�y��	��d	���=~�"n�ǜ:=mY�^%����Ϻ^Q�*_�Eɠ�(��܄|��
�
�W)��U�SR�	��t_e-�;�;��'K���u<�_���Z�5�N��o��_��Q �Q�������x��|�N*�W��D��F}��;K_�/��"x��eHYV�˾4q�2.�JC�vK,d	Ž�Y�Q�ݨ�1~�}X}H=�'yi�|�f���>�b5HPޱ��������Z-��|UJ����V푿����p6�I(�:�5��M��<&7�5Er��8Z�)H��!�tG=���P�Y�U���m���m��jC�O�~d=x&rQ�ܖ| �ͬ9����tw���qh���YL�g�h���)�(�g<��I?���ʌ�!m��6-��ƫ���"G���pr~=�C S�m��5�g'oP��Oof�!�	��Aֺ&["!���_V��U�hw8��.c���j �[��2?D�Y� y:���y��s���|����&(LnZf�G���?�5��E��O����&s�1r}$z&�������Z)I͵%��ι���u�6��fAP�]��|B�T�5�vL�w����yJ��h�ً����IV�#
�s<��J�ϛ�*G�e�f^*qhEQo�<h��k	$�$u��<�0��������$#z�����[�5't���̭��@R�*�6^;D/� $�� �䬒����������Q5<��f����ֹ�ˮ��~-5���%H�U:���\�^��������k4D�Qfp}�v>o8C@��{B�rN�V�]w�pRa��{a�ݿD`�w]U���ʯC}�������4}��G-;�9A�6M]G�+>M��4�nK��t�w�'?��Ȃa�L�8�l ����;� ��!˖U�(5]v!�L�b�ŅS���읍�v�c��ߝ��n�kj���1��΀�]꿵1���}*9D���d/-{�&�l��3�m/���x-ޮ�|�>eoN���������F������=2zJl�~��8�;��a��,)>�I!�l�[NR\����=��pw��b�wy8 �>��ˉ�"���tZ�2C���A�k���؅̶0�9��� ��E�i̞;K�=2@9����H]�j�[������@�M`n�e⬌miǪ:�U&.x���c�Wm�Ls�V�l�=`ô�N��;ЛO]�Ȫ!@:TP���X�����=C[�� ���*�Xz����R��rt��V���)����FAy-���(		s�4���%C����v }������y�x�A/@;Zl�G��\�;D�M`%�	��B�P���5$�	�Xu����4�\�<[�`��Е�K�4�x�/#�����3{�״m��Dh�x�3����Wg`I���=f��� E�ߔ����Y�3-�Bu�B�/iE�V�l����n����];v�-wٚ_�a+�I�w%i� ��v��:arth)h S뙈���G�K.a�Ѩ�=��-��%1�4r4�mD��H�;h����D�#̘
TC�S�-�;�i�b��*3AYgw9�﷝Z�H�����!��zļ����M�rV�{-��5����I�X1"7v��o�pTb$���)k��~+��4Ni-
�&��&2݌G:/�r�&�e�����.�O�sF*8ۺhn��}���@SM�]�q�_BM�(��0�m���e���ӏ���X-�Uj	Cvi� \��_U��)ֹ��q��O'#�ϐnO���&��3�c�����r���V/=%�2{%�7����n��%���m�/�����ۨ˅��M �+ �KԴ	Y47��K�\	H%]�k�Dݘq�l�Hu֝msT�W��fu��������R[�vq�ЅX�4	Nl4��n�.�Ţt��I�
y��c:gI��kͻu5ߴ��re�MS�|]r��P����������ɟ�;�ֈG!	+bm6rɠ�C ,=�WѬ�,�� (5�TJX���V����y|�����t��׀��z|�bf)���̦�I�Jg��O~mUږV獮�����9Y *� d����bs^��B�)�遦����f#$tخ9���(��X�	���-�0B툯=`	��j��M��������3���f���_�>����ԕ5�	���X�т�>��f#P�Ϝ�~i�0�Xu2���_9���/���G�?��hH�9��H�	���ď�i�,�~��L�)��M����|1y�lh\'ӎ
n�n�a<n������{٪b�C� W�X*�hA]^�?S���K�t���e<�0e_2p�z��:�ڠ|t��x<bv�j�دc�M����~%�b|�&?G�MD��*���a/�彝WiG�.M�%��6ʜK��k�'���}���a�ԛ����s��sn�{u���~c����Y7`��P �9��C��5).Z��M�wX�X�K�94�)��@F��!�T�'w"�)�ܔ6���[{�s0x~�B.��5B<�8���CJ��uw^o��8�C�|��u��FM���؝s?���{���mN��h�H�~�Bd�	�{g5M2U¶^�!�j,��%��<>6)e�9��,~�ʷ eR{h�M��K��p��#T��8M��%���(�I1~�ˠƛ�=�?�_�U���w�y����m�X�[�m��B�A�`�YT���(�$����z.���o8�����S�F{�.{�M��`���3�z�*,�ag��`�����`�����ÂW��<{���	+f�e8��<��<.�����X��Jni���0MYwK��(B��%���#_L�8��$�Ţ*���,�́[ۍ|ִ1�\5��`��y� �c����ʂJkM�}���y�(��]��[�8�S�m�v/5�]n+����i-R���G��#�`JXC�T���{��I>NB�BXТ+�S{퍔��~�J�P�o�'x���J����o����[�+%�y9�7z�f4b9��*�P��I�V��y��2��YX��jn�bf�y b�h�%B��q)[�=� �ͰsPW0rgnB�H}��L��z)��G�m3ǃԻ��?̿���Z_��άLZ�\E����Pq����4�a�{��>]�b<�<�У�I���q��J��|)����U����:���zk�Hp����|������j�����s:� �Ŵ \�SD�%�hT�g~��V6�xFH����g�ƠyŧtP	{TC�M���1L��*�����مN9�7#��5lh"�	tEG��r����?F⨋�t,�y�/�\
��5�n�b#"���� *:����1�c'*�ǋ)9�!����R���5��Al�.���M)�S��2w�pg�oL$�����}����n}��
�T��#���!,�-��3I�_S���mSJ�Nz,��[�m�����=�)s'M��fюD�C,�6
�l����Pn5Cf�P�Z�Y&�[����g	�#��
/��m�P��޷�i�t��L۲[%y�w�3�FB�N�"� IB7(~2�ǧ��_v�� :�9�[(��%84l�֡��P��i��j�� �Ѣ��� I�e�y8��p�b�峋6��a7!��il#W��q�v�sL�Ma]�J�g73�Ѹ���B9��S��uY�n�+\���e���y�`��J
\�tQ��-���]����DE;puW+�'�&l]p� 	1lsN9����M�vWFʮ����cx��q�NЬj&�E�]�د���F�gE��)���
��&'ѡ?s�	�bw��o-C�A��H����]"��V�&2��&��	b��k�rs�����2��࡙��Q6g���qnJf����bC�?�yѶ(��/�[��2:e�����b���j�T��7�~t�$.]��_4%�u���$K��w�ݕ��g�V(���u��)'h;kx�9oFwyIa�����x���Jw���iU/F���������̡����� ����w���j�ю^I৫�~#��_�(���'�xƌҚ�!�!��;5�Ռ�7��1���̂W�OF��F��Tj�I%g��#��g�*��]���#m��Fv��cǮ��
1M���ƾ�[� k�A]=�����w�W�F_J糧Vt��!8�H��#�qJ�@�ͽ� VѢ�y~/U�1�M�ʟ)�Wv+�r[ ��]��.{���Px���������KmgV��R��{���2ڔ+z`����>�:/$Ѣ��F��[��yPy���/��Q�b�`�Ԟ.a�Qk�ۏ�r��c}L����wlVj:y�^%���|�+��-���2X����%�2?f�\��5f_8.k��iҼ2���&��	�V0���W&�t�̈�0 w��r+Y���������)&Z�=�;Υ3��Okl�6�C�S�	(�ș����7C��K��2�M��A�U�FS�YFG�������{\x^W�J�"<�i���0nZ���NȚ:6\�K^_���%�E�]���01���h�T����|t�šKe�s�LJ�asx�b��<��d�I1b����=XH�h��R`p�����x"K�gNY��ܓ��n=aʁM�G�nӎE	#�J~z���hP��QT�u���Q:1�����@T����Y�:}e��M~q�n�lR�b1&9�V�&5�~�X)ڤ�9M?�����n�wg"ȣX\�H���j]X�;������sp)5G��eSލE���u�J��L�nD*-����9p�9��ww���q�U2��T���wW�����ύw�x���K����ۦa��7�UqA�6����v�Q�����4�����&�ە�*^��&�b�7>��X���Ȏ�O\�+���&��C:Q��
�Y�o1Gz��������X
�o���6Ԕ�}��(K�����$\�����AL����ތmb�ɨO��zO���V7`d�ٷKf���N�|���%-���t���W���Ǻ�x(YP!3���A^�Q�΃;{�H��]1;�j�����v|�����S
�O�i�cGA� k�O�o~���B����<4��j�4���A��7��	�R�������f[�b,�0�ZzuB�&����y�|�|/wn���$��JY)�����qA�[ޣI�T�u���7�C�����mYzP���X�#&P4ԍAĀ�J$�{����Z1T���צ���A�E�Ӟ��T~��[RX�	���J@M-Њ�	{�+��z�n<�� Tv܈�7p~�k����l�<#�K�%��[��\aI����hK�v��-�|�*G����g��i��Ye�q�����"��~C���sS���(����ѩ��8�=oq;�y��֥��FRa���,0�"3������v�Uc��G��[���=*q�D~ �.�xr����z�b�楆ͱ���JJ�g��a�}G>+����eB,E�!�쳻tzh��&��&�rd��/ޱ�xΑ��7ч�7T0�������Dh_'q�����CRR�p�o�%Vx(�iG��ou�]&cWR��}�2��W�H�O�2�ry��dA�d=w���f;{�J/8�$6�La�>��0�q���H)�%�!I�b���%?�aa��k�A��}x�J+��T��> �%��Vt�v�m�8\�®WBh�\��c ]����)U_v�s�W��j������R���p�X��E�-c|Y�ʼ+?�&�@&�u]\��ׇ�.��Ӡ��d�*s(*�ѱ܉�b:i�v�/�}�!��-�~J��8���{��j���X��`$��F�� ��`��)2W�u�	��%����I23��8�8S�[��ǲ��	"ń�@`�� `%�;%��APV/J����b�2o$;��p��H����^�#�0�� ۨl'����{�r$kRE��اK��:�ḇ�֓d�p���
�J���5nmg���|$�k�a�8�#�Ywo���[��Ou*�U暠M8��[ݹì7�IM�-�8"������}D�P��QL9RHA�
�B�zO�G@�ly��ሥ�AJ+<z�y�vV��E�rL�w׊�Xc!�m�w@�>�e�8ΰ��u�$��Q���0���K�H���`�A�~ц��ˮ~���0�ta�S��p@��a2��:,b��E�:|��N`O��o3�$<.�#�Yۆ��n-֜�n;w�q�8;ҥ�A���2��&��5rQ�ȥ���Yh([rC`f�E�:����x��
8���� ɍ�(���Cs����t!��b�r2C@Q��#;%�,ò������� =��Q/ .��xknD	��Q��.0��K+q�`MQ��M�_.$��1��r�h��Bc����m]��s�}������o73�����¿_�&�dD�,Q�>�}�v7#g��g�̨�u|�~�(���@6=V�=A^&xX����'ԊW��5նC�'�&�p���L�ڽ��%�s���\:֚BZ��KՋ�Ѧ3�Y�1_�e]~)S..8�n�g����M�N�\�,�ӆ�%mz?"��2S� �}P��k/�
U;4hq9��1V�t����rF[��z���^$^� �.jW�lh&v�r$D#����B�	lf	��,��ϒ0)0���@��S2�,}�o�ʀ�v�ǎ�S�t�l,�٥�"���3��(�] ��}��Q�h���ե[{nx���I׫�AT�ߋ+�EL��ᡢi����Qb�l�a���n�D�����kC��{�t@�P<�h9�M榱m�R�b�1�&u��U�/拸�D��`y�6���4ϳu�Ôg�Y�8�������\�ɦo,�&l��Ʊ��V>�@hWY���]�Y��`e�:ʁ��$ҙ�o�GF
�������@P�$�UE�~l�+�n���?�Cp� �t��͓�I�/��G�ca	��4�㌗�u�מq$��B?l��U�h��I�1����0pbO�T����gDDt�}�|���#�!��dk���Q�J�#�[܎�Y�!{޷2+C���G��__׹���#XvVB���H�4�QS]O0��ԄOq s~�4GxA9�$���0Q��]y��8�Li�*/߉~[��B$���*G{8��U���"wѼ2߸ҷO_�<LK�@�X�+YNv2�	�H}����ـn|W#qyD)���n�`�u?X��o�wdu����{䌵�pPY�>�gO��F���$2%� pd���\dϓjs>�'K}�|��X���#A���;�LX?/bѱ�wc�?/r�Ǡ�\� ��B֪�˴ޛ�R���_c[擛O����y8$y���������λ�����ik!�;0�C�[��.�u�(���,��E�hQ�N��^���=�%o�nY�9z,����Nwvٷ�X��'RX6w��o�Y����8�OJڝ������I���	�">��B���:n�e4 z�d3���OC@��y0Tz���T��;C�`�y�7T�wnO�A�Zg`������c��m�z�A�1��B�d��w>��T'\�8���ƴ�Z�qx���f1�R~�I+�F�%3*X�z|������وh��x���`�<��6T�y��]q���NM7�,�
|�8,"�#7��v]4Wq�zk�,~���e]�`ϒ�{.��]kKx0@��t�o7��]G�h~�nS�.��gL��8�ީ6�S��3љ��+bE>w�7�;�AB��z�	�p�<�ƥ��z��ZSɺ��'�ɒ=~�"=<|?K�H��A4>� �IU����>Tѣ�}�U�q�I
�I�oՂ`��0F����|��i,�Oq���ŁB�I��y��MW�Gz����.��Hy�gϡ!f�젮��˒q4���=ė�ᤀ��6��p��x紖�Q%�5	��f)*l?п�H�E_�!�N�7(��:���g�fLK;���m��f�&��1��#gI��G���X�ɠ@���9z��#. ���_�s��v�EݟO����0pv ��G��	�N#~��S�˼�ֹ�:8�	�U��u�n|<�1���5�5�D����8螉Y�k����g��>M�&��&�2���K���A�>~m���\U�F��EnXc��큍S�}�v��@WK�w����H6D���Pw[��Ӎ&A���p6���RWi�^�ρ�VR�ގ�Ȧg��p�%�][~�������%xr7�{��x�� 7����ą���Gw<ZY���W��`'����o����;H:�dmX)\�#/$�M�u+���H��J�Z��dU��`�y��VRW����饰�e֟|]������z�f"�l1�y�E�x`����{�^����yP����� ��|�u"��2��G�}�T�O��&9��~j�����h$k|7x�SW#BQs���>)Z��a�P�m�|7`��fi���XUy�D�6�ސ ���j���k�i��}~�.C�B�����7��(=lit�v��='�����&s��(zq��oX���pM_�))٪�����P��.��z�:N��i�-/�'b���,2���q
>lr�ߺ���g������=�&@�'�o�k����A>z�G�/�y���ca�a�׷WKc���a�y͑Z#%�K�W��i8��#��&2`@�F�jw�.x��v_��W�������)f��ٹ��*@a@Y�j�&��ל�i�CO�,KDg���;����ҠtP��օ�' ���VˠP�=KM71e-N�����Û�#ʓ���������R�%ʣiqo�a+��u�1[��Z���V�VLoQ^h�+����̛��)ma�xC�)����b��y�"�@�԰�ޥ0S
(D7����t�T�JK�L�r)�?��,d3���D��Qhj<� �5��ĢC ��Td���wW��mǯѧ���|�+���4̴\�]j�%�6D#QW��>�8��H�I[Y���X���@*��'$�m��f~�u��l��AGV�i��k��W(����'c��{= l�'��J����q'�sYsh��*��2��&����u������E��ʍN����V�ÐЬ�0�x䴍7���:�@:�	�8����p더TZc(����f�cB'�ù8�%�:'��N.�$=HdJ�lVs���Mފ�M��9o|T�!�j��)�8��ֿk�q��j�řF
���0��ͽK�o�5���㥓��ս��`�9e'��Z���B/�\�D脯C���8qx�HIBqҗ�O^KO�Mx��(���.9Uz����4,�����a�]�Ń�(f�t�#��JP��,�A_��D��m��H(���-5Ѯ�kn�àYE��Xy�RY<��(��^�������B�y^�<1!�`�W�PA?�أY�x�-ERԚ/`-oe�M�3e-�Up~$�;OĴ�5BW���VK���N��yt�G�>� ��Yo8��0pc���@�s�Mx�M
n+�Q3�JӧE��̿��S�,�#]��r{\r�� )�[�3V`����`��j��)�ҤPј�x�1.kB�����6��]���[����!�e�
NRz�j��;gz�M�j�C�zF=1l��6	����ZJ~SJ2$��I�)d�hƨ����?�R��NX���m��CY���
�o�o4W�-�	� c��* �d�p�-���Vg���ꁕ�4.F9���y|f���6]N���-J�ׯl�(#l���{��c�DŻ����*.������B7�����Ͽg`E �ĶE��l!U"ٜ'�_��(���o��Mȷk���!���u�8ʽ.��D�H��Q�!��q�<�A��k5>O|�|����+wu.�I�.L�	x|@��=��e�{�5P�6M��OZ����j�b���V���U�U�㾤�����G�p �yW�<Ɋ���WTm�����a:���&k�:�G��a J�[�!�c���~Y����%�����%���0K �%�˅���Un�'�t.��V��;pY2�Ӌ����Mc�S�f�C�U�K�4�E�̏�<(ι��l�Z���
�V�aa�GJ3��aa�BN��^���S�F���T�?ޏ�ʌ5���(jR2�N��GP�褷J<٥�W����i8j�y=�<����&�)��S�aG�N��x�Dt�a�X�%�4mPo�F}t��A�
��2� A��_&ʷW��t(�8(�;�0DYlPuJ�.t�j/z߈ɡ(盋8���$�k�Í�#��Vl*dc/�X֣�a��8+�8X�J�e�.����TV���,�c���+}$�*����W�B l��D8JB5�A�yE�{*��Ee�e�U�1��������$�~̂�����]�\c5{,�;?���8c;��R����d�f]�e���)d�wQK��z�)�o�P���{0(Ώˈ���}0�MS�T�7!	��cy��a�-}�\�!o�C�L��<�!��8��7!��;��2��O��� @���gVأ]�e8:�xֶ���^g�~yF�YzKs}9'�ԝ�p	!Ը\�^B��ru�R�]�J�@v���.��9n�\��j��D���k#e��h�!�׸G�0P+$ZuÃ�M��PLHZ�h���ʬ�5��'=ŷܦ��Wr�k�3��U'3�⺓�2�t��)�e� ���>���O�E%?��f���pE�2�3�m-I��)]�Y��q�Jq�A@�v��������mj�Eq$��8^p���v� '��$-;��$�2/�y�Ur�궲�ap�ę+{\����U�T.��-�.��܀�v��^b@=���b�	%��}��|�ճ��M{�M!>��"Ն�u�HpG����E%]Xٜ�!�M���
^�L����������]�%O��@�6�k}LK.��C"�K�w*+ME{�Gӷ�0
�]-H�W��������$ �d'u�	f�\�|j��<��Ӵ�bi�R�w�ڒ���V��F��~V�b��������fJ����
Vz��EP3��{+av?Е�`�k��ý��T�J/���c�;���S@��+�$2<����B�8*�Ӎ����b�4`���t5}M�|}x��~qӥ����$�:�9YW�}�e"ێ���_1Sp�CW�mipkP\xl1�vN���[���e��Ze��:�+}o'E�@��d�1Le�")�hKK���ä�o�k�Σ(K�M����R'�J�7�y�k��G$�Q�(����-�+�IS�2L�tS� i�2�c�~2��$��<X�.v@���8G|�2B�i���ͅ���D>g�������m�t�l�C����1W���������_W�����=�iӟ|��&�g4���C Z��LY�X2��q��\�=�q�jӶ�h���\�E_u�I!
��Yw��U%+�[I�p����e06�^�$�W�M��a��/��V �T��PsK����,M ��`�m'tQ���0Zk��m0����T��o��B=���,�n���O��m!}\��H��}��UD�����Hy&����W��;L�&���d1O�,�U����� ��`F��*�s��{FF0���9/���# �P�����2�&��Gi�����v���� <Rܘ�q!x?h�3?�=��8&��w%.7��GjÀ%�(�~�hUfH���|��ɥD�~�Bz/�VnmH��:}	�f1���u\�?���P�H'��̱�0]��3�c5�= Rv�<"-�P�a��?�/�DX;b���pT �y���זG�9������L�*n�h�J�:O+��x�m��r�g�N�J;������&W�xd%�A
�}6�}S��u���:���Q�������>M�S
딺�j�����J���	ߒ����`�b���[.(��]��(P���4pt�Iԉ~��_�B6����� R|j��t�t&e��z�p�`�tc���R�s���V�&��~w���KB� ����8��h�@�|�ԪK��"�u.�C�u�Ƚ�%� ��2|rli�UOC��y74*���s\��jl0�56Xs�7�lWޖ7�q�e�+��߉��~Uz���(OmH���Yߔ4�ۭ���@ 4���=$~��n��`Ol)���E!�m$��T�K��^�ٸj6��Y[K��KF������rAh)Dָ��_���IR�y����Hb)'�Eŷj�c;J�bf�����c~���b�@WB�ԙ��1���-��������9��oyIg |2{�'LYG����U|/@o��z�">Ky&��Q2�I���0�K��k2���v9p�~V�� ����X������CHG�����
���8a��um�J,�H��5�\�d���:!����IՍ�I�f�K����>b8�H�ӧ�w��MThEt�JF�O��kFv؀ar����[��z�)8#��*U��������!ئ��E	$���:� +����1d��=�5��>�5�g��%�?�Iyܥ���=���|炲'�R�3�8ʧ�
�Z���O���pۍ�^_�@{���hc���/ �˂Z2�d���W��rt���/#��}cC'
T���(�1;� ��.W0���yz����ݞ�r��~=*���f*��_q��u�x��� XQ'��%IN��|���+�᣸D��aΙYN����c�-2}k)H�D_����r9q�T�!�H��;xo˽��%��������W�������D��{N�F\�	f,}�����ɺ���U�E���@�r��ɢǈ
�L�<�(�ۅ�V�Xc�d���j<E�����~ȁ%K�JU�ZĚ�t�dZ��5�&�P(�OҖ���R��u]�y�����*g[��-	AΕ��&��S��f2�� ӵ�W�T"*G��fQM�΢G���^�+�撾�Az�� '�����3�X����Y�r񅚁s�,�ɰqo�^�5�Z<� tS�q��
�S�?��ȗ��ii��]���xp�[��ܻ��P�GyI�����	���q 􏆤�;������,ɘ[��e�쓥
RÐSg5��%���¿$m�g�H�y��ѱ����@�pE�yo��}�����sK�����`-��� ��#g �k����	����'�} ]����KL������i�<$ŀ!	J�:���9�{�U|:��]Y�5��H�֙����P_aګ��J���˗o �`��m���l&`�	K�CI��W�\4BI������j�����/�
6+�*�2UA��J���p\�M*�'��1�,�G1�o�a�������A�{
��=/mdy����2�SWw���.�9�n� \�(-�nР��Ř[{qY��Bxs�l@�e���&�����\U�nӸ˃�x����zO�[���j��GT-�Q�����4
{Y)�%����*wUe��BK5t���M���h>���};�������~o���bǅ_�;�C</*�8������̒���fI�H�q7Q�~��#�6�b�e�e�l�m��WC�x��A�Y[�:�U�֎�^}ΘI%�6u��p�~�֒-��3�rl���� �8�-����W�·�g��n�vsz'A�ʣf��� �s�bL6���eʸqR�,����{�u�5���C����ACI~�lXʿ+*x���Ԍ�Sy�� �d.��N�_���R"y}v���V��[h���8N��q�tk�&!���x�d�)Ҫ���9�̸,ƹ h�C�0|�Ǯn��tg?uQ\���`x���2�Iw3�R�HL�T�o'��f-��rj��c��f�_�~ ��D�d��j���}�<���2H�0�T���p���X�UOoZEk��^=ޮ�iD�0�w�<��6d1�`�ҝ��Iia�����r�$�,�S������ڲ�O���<���ޣ .A)����O���7�LvF�&h��|G$F������7�{��yg��⬿�8�aY;"}�����~�9-�g7�P��i9���`��JX�#�~p�:������[��[h��S��ħ��h�]���3����s�|`=�t<�^�S�*�mZ�]�s,kn�?6)���YqJʿڙ��x}�~��\�	�X��ǂNtϨ����2!K�[u�;�����;��}�۳��ȡA�η�L��^>�7���%�s�k�rzn\�q�9{M�͌?sy��͡����%��5XRZlȝ*��}���Eu-f+�U�BX�FE!�뤨��8��C��1�vNWB^DWI��}���������m%�2`׃��4.��7�+���W�����~�6�,��oj�"�V;��ZHX��g�<gG��֪Zi�/;�l���T�kW�q���
s��*�SY�i�I�dAl��Ӄ;8N�'W,5�*U�� �t�vcx�6�nud�{�3��st�ރ���b�:D���|��k��$QHj��t0��TM wdC�i�Ђ^�w��E�t�T�AX�9P�^�fa��y����0��,�V�(����L?�+4�	��vC7�^���"�c�J�lك�#�s��H8�s�IЇV�F����>��! ���-��*�Hm��	�H��?o�ׅA�u::�N�X�R<EE����r�a�L�~�A�PƦ,�*��=��op&$��la����)��Ǯ@�P$��J.����'���8���A��܅Q��s��Q�Ak�8���;ɹ�q*����w{܇�K?����#oX�@L���������)&~+�x�{3Ԇ%����(�#�U=����ed�䓲�ND���#�����p�
y�R�{��UJ�D��秺���&���i�Ц߶�f4&�cʜ#���MB���5���z>�Z�@ׁN�4��Z{�>�ۮ>u�0���s��P�2�n�&�-�DKW#�O�ڕ_Ip����$��Sx�Gޘ|�b
8�A8Ѻ�*�*�Tm_���_����fc���.Ae��!��i)/�:vt�-3B���j�Ѡ�:��}W1}ي{�=�< �πq��oA�*�4���`Ɣ�f�8˥��܋�
��[%-�Krm
8[��N��U�b�ݧ}���"�o�������
���F$����𚀂����T�Q��G����3�)��_ԑ��J'�ɜ@SsR��];Ӱb�UY���'ah��jT�{��;������/��@d(Y�����÷k輋s��(������
pp�Z���	3�P�$#�==9���@�s49_]r3Ɋ��M����X{�����.lv��E�k�f;�#�sAa̧�.�P��,�v�M$������I%}��O���<��L4K��x&gW��`���Mi��M�c���z@���(�5� X��8Ңp3c4�Oު�${oD@�m�O;���!N�Y���Byi�yA���>ݮ���!��~�|���&6�=��iH:��x��E�1г7��Bv�efT��<�e����|�^�{�;��;ظ2���/���dS4�~�)�s�6����2g|���P��Dd\��8����|#;�rQ��]��וF��F�@��9�z�:_ Y6�]�8'v?�#�L���b�����B�6E�ը�(�����=�%�����ϵ�ϑm�f6<��BQZ+=�>�0Xx`���������(������ �<�VM�47CW �T?'eu���s�A�����z������>�o�#d��Ό�B��oo��W����<�����_�cm񲓾/i.))nD����3=S+R��_3������r`������C������X@��ޥY�VJ��v�C�[i���k���#j?��F3�і�x����D��7�`4~�x�kd.��c�U]�)���<�,����qŤ�9����nrZ�����g�1N�Dl��>e^���ɲ����Su�Z��00�L��K��c�dL��&̺B�
L����'��ʌ�qE�>*�
�'Yv�i؄n�8�I,ɐ7ZN'�a������T��9!:b'�_2���1�>�����r������K�VxK?��͍	A�hDM"�@���K5����G�w���y͌�Ś�a�Ņ�.��x��.�_I���7:�Z�y}�0b񟒳)S^��8�0�N��O��i$��jY'\<'����a{͖�\C�A���e�'՞@�g�H���[��!�M���|,#���r)42z����#���P���� �7�Z��-��y`�ke�N?_�Sl�e����JFj��s��������,T�/� r�34M����ǳ�7����;����ӡ��C��ʍ��š�\	��vm��l-��� ߨEh������0���������H�ؓ����y$�'��@���.~ܻ�EU��y�c_ǒ��~������	�g��1�K�ݯ�����̯��g��e�3���S� W���V��)�Ue����U��L%s�Y��Qw��Ov��<�1��N8/i]�e�&{����-G�ˀz$���^���)���j�F+]�K~�X�FM��m%V\m��el�	`-\�X2>ʺ����}�bG��G� �:,H߽'��	#$��
��}!���w ���[�a�N��/ׄ)�s)i6�1�
�J����ΰ��x�Y��
�Aw�:hAaPg;�a�����h�*��*׫��yS��/(���`�*;x���(���9��,�N&姚��RT��t�pO�p���U4S;��%M�}��0lZ�#�p��xqҤ��۪�Z�/��n�%c��U��q2U��XI0ҵ䬦��C#gr��u��cU���gn�o��i��ּ�#�0�ikM�;�����/� ^s�싎v@h6Q1���6�LX����b=6������l�KL���r}����cUj�6�o��46��K�B�KJ\��'�H����(>Rd��@�şK��n�3M�Up�����LI��C���7�ԋp���9jErJ��c��|�n�	����XE�K׹ؗ���p Ģ�W������nS\���8�yښ������S�a�}*!��/�<ysB&���. ޚ�����ę�D�{�)��G֎y$(�i��!��ѓֵ��2	��T�'��]zP�a���,2��$oZ��O�z�;��u�?�I���
��*n�4�O�OE�fa�J��g�������z>c0���ZE]n��<z|�|m4;sPp�<���2#���o��U���X���y��9��o�>7�ӡ\7������t�J۪S��0�I&�6p+LQyM=�$�[Jb�:��ô���+��E�N�C��q�4=���+`�� ^
�r~�5D&l$�벘DTX{�F��k�gBo$n~l�xb.Wlx	6������5tп���-7u��*_�}P ��;Z�!�Fc_��Ir�Wy#vҬ%Y0�/��_vE.��G���/pB��Z�p,���G�I�0(5'χ{�N��Vܚs�t��(J�T.J�F��ӱ+��v@��IN#1E�(Ӎ�+�J���œ��� ��p��R"��zBr�!�É��H��0 ��˔��[�rS��X�^,�E^Q]a)��a�h�v�ѐ��By"�Y�?��2�,R:��ͮD��|6����z���Zn��{�>ءuE3v ;��cչbN���y@�`ER'|����+�D��L�2�?��A�>�
�5J1�H=]d��C=V,���v�ɓ@C�ְNTm�f;��Z_Y�q)�'�{�tx"�Id�j>���͸%��O����3�O	EY�{V��_�FOy���iڗ�_>�cg-p����|&�|c�<�.����:x^j���*-�LwfH	3�3����+Wy'��$KUo<;T���*寎�8)��]�ާ;��m�#cZ�1.�e�טF���Wu6'�ׁ)��X,P1�.�ӳ���q�\/)��{�Km�X�)U�2� ���~usH��e����P]�:I�&��&�q��gۙq��&0�n 2��$�A ��#���l�rD��8=h/
��d�
��iv��b}k���k~S${c_&����FJ<b��`���7���(��g��ҽ �{�I{<C4�3�Ռ����,��;�����Ѝ�����΅.d��)�#�w��Xt��(�_m�X��)�A��ْA?t�X�؇�T.�u����(Gd�� �jxE=L��94�<��TԀ[%-z�yџ����7�b���ܣe	��vSح�����8���%�q�W5�M����i��*z���HX?����G�z�~2�g�P)��1�=����T'��w��ec��ptW���X���J�~a7��F/i�Q�R\B3�u���ܦE<��;����4�,Ql��y�i���a����?�Yo9��ϛ�z,�:���O�a���us}��_Z�I=xS&>�1�X��g!)�ld�&��|\��k�i�o�{˗?���'�`l��3q�NWڧ�'�/X#���ɏ>��潻(B���mo�w����%ͺ�a�h��SMDjXUM���8�'*��-��IA��d#/��SV��j)X��_v����2O�N1�-Ux�/j��-Q�V��b�>��,\Y�?�9fɺW�.�\����
�ʆgb[y�E��&	��Er.ߛ��U��I�nL�����ó��2��-�űz��#-N�L�Ԇ�(�(�����qU�u�9��x8�%đ$�n'gvU`m~���`�gk��v"��qy`B���mP��5��f�K����|Vsm��5���(���FB4X~ ���LLE����<��ׄ4�f�c��-�Z>n���;�o�V���u�ȷ]�� )/��"B|�P�{�^���8i�ʜk�{�o�@PD;�f}}�IggU�M��66�#�"qq������F�p�M�J/j�m��Ӊ�E�hm����`����
b��w�M��ph��V1l;t4�J���+���MpϤֽ�\9���O͠���T{��.ʿI5\J�λqD���3qæT朡J��j����O���f���Ej�%�F�C����I���R8q�+���Xj#���8��|I���v�A��n˒a0X$�(� |)Gm]Ð�O�����7e�����G+Y�kp#��L�ǋ��j/�[6k���)!�+�Wu֔�Su��dV�>�U+�D6ci7j;��n����&��b͐ҵ�9YL��C*�@�C�g�9�O�������EJ4�#��@��W{>G�TH���d���+�.U�$��/��Xj���ݵ�0/��@:p�� �
�h�0��xS�r����r{����5NT���u��O����B�X���h�����q��VG�43꣪j�;e���O�cI�d�A�-]�]��!�C�{����5���Lfс�� ���C�{!5)=�q���+1HƝ�N�r���T`�_�D;7����D��7��������pD�DS��e<I�U��d]O.��� �V.�ٷ���R��J��c��?(�'}�|�c��α��R��,r�H,��Lzªhn�mT�/�C�〟������;�_�O���W�2�W������Β���lN�y����!eb����X��`�����zeuE���K��A��R�%���5�r�xI�	���$e��_ؤT�m���{�Jh/{w�oAI���������	��`���T�I�V_?K&F�R��Q)���,1�x-%����Yk龱%G��#^1�P4T���S�S���_�Y{hA��$������@�İ��9�坂���?����a�i0+���� O��� 'ё��TCb�V���mU��� ��X*H��d9��Y�N�T�Q��F�d�X|0_��J���D�(���
�9c�N$�)��Ǻ]G���k_	��J�=s��P��a�3z�'�Z�6��� r�UP��M<b,%Mz��8|%P�)B��U@<�>Ԫ�������� ,�ؤW�g���XŬ�X]���z��K��dCE^3.]m��1����I����D�Qe��R����b�H�,�Gq�VJ������y�0V&ʝ�|��5�)�.p�,���I�2��� ����\�/�N��e;���ꮯrGddZ��<��� {���V�_^��R�>E�����%����t�p��i>@�5���k��ӽ5�>8�-e�<*w�%� N�s[4���
�0k�sBd|..T�P��#�c� 4}Ew�{�Xn,�q�7f{���:�E��>�ÒHi�;�0���(�'2��vCg�&.95�E��)/��^
m��RO���M��xq���g}8�x�5KU� ��Hxm�C]� ��q��|7?�םm�e�>]��[ı���^\R~H� ���hs9������
��g��?Ͼ*`"���嫑����]Jv�A��o'97 1����1j�֋f�d�O	��˺� ��N(���
��O:v��U��K��pKѦ�dG�6a��q���[(�������w��j���|�7��{6@ɛ�x�C��jd�fK:uc���e�B���B�i��\�e}�3X)���pz��*~/
�vl�-��ոVP>�G�7�ܯ��e���pJ,{�'vj�Z!�������[������C����Χ"\/ݢ��#^*���C���z0��ԟe�&�m'f�?ehx�����+,�����N�Z�]����:j��31\������`.��d5��{�6?3�7!��5Ƃ��Z����t��x�i_+��!�nR��w�]v�.�����Zy�L���_7��nÕ������@����֙B"u�6�=�m��L�V��K��kǻz����]���ۣ��f�$�Yp������9�����/�\�P{���@z�>��<m=�(�:J6�_�[H��9 ��L�}ݍ��4���R�;���6P#zꡋ�.$R�|8�rʡ���"L��'10��<�9�+�9cߒ��"���f�C��U|'K��V����{?-��}[c�-v�$K�����j�qw@�vb���(�𹺁g�,��Qx3�u9?��M�C��:��KC��p���ay����s��WD�A3Q٢JN�~p�!���"�r�Ǭ��(���Z�v��$4e����1V=6����X��16����?֤(�o��A+�.^����T��3����lD�� ��j�x�D)n�7��&-���7cnB����DlE"�tMF���hZ��^N���?�c22��S%�j�����>.\��>9_I����P�<�G�R�̯p�~�����*:p8z䙵L �٦T��&�YA�����Q6ǅ���b��]X����O'���h�0t�5�}�+yrJ��Z�ͣ��2>�`rW�t��y���-	>M�B���':��}a�;Vl�����	�]n�1�{w-B2���I��-���������S-�t��}j��T]�]�Q���9iћ��Ze�y/����_uQ:b��w�Z��\T	��l��?*2Z���y�p�ߟ���Q���1�,4Ҋ���"�k�Vs:���Y����J�6�-�����!s���C�5^?�&�1���
]��7�;\q}����o (�))�	CIN�������i�׿�m�rD��ȣ�w�
�����G��S��g��"�o2��vo��*�k�����g�W/�T�f�_;��7�V�~��|�=j=j�l�P>\��T(�{�HP�ki�3��1����2�{}ي0j�����y*��}��i/F�B��Fʳ�&��Tw��Ѿ��s��dvk��-5n�m�~z���� #����;��\�;��'���&Hn�YL
*��5���!��,u�M}�/��`����nt�ٞ���𨕫8����B���J�^I(���^�aI�k����hÉ��SBaV�Ї�Yz"�^Ƃ�C�tbv���yΧU���1#����Ty�/���HZ��-կ�s�p"��,%���&���b�K�VK�x���V�M-�o
�9Lk}�!���Zv?��R˳ɷ~���Hl/F��j7�HA};#zja;�5r�n+qk�򫽡���z�T 	+<�
���I�
�N	h:NY��r~�S� ����.��V.k���Y]�Q|��#4$lF+g�+66������jy�a+h�[
\g�|.���Y�i�.s�W��>;�9��^v)� ��P��/X��F��-�P�u	�^�Ճ�����=�!5"S�9nBM�@��vj,���E�r��\�MD�2ҩإM_��[�p�6�_�[{�E�@��B�G�%�ůvb���I9�	�߂ڦ�u��!��35N�X΢�э����Ï"��W�{�b]�����Ú�k�^|W���(t�o�/}��qb�!k�ꢍ�P���w��P��&�x�HP�.�zF��BXs�U8�����q~^�G�qi����9s������ $ٟ�e_  �<�	�b�CB��p��yz9zn�]>�C���\��W���ו�z�n�1_R��"%��
��M���>�&�qH�*ٿPǒ)��ۓ^�*s��A`c=�[�}4s�y���7�|S�0Af箝s�uI����@�AGB�P�^���ЩǞ��(tI�����4�����L�em��tY��yh|�w�5�R͌��<�v��� ��5v:3VLb~����	��}�J
�&١+��L1�OΨ�Y��)\,��Ĝ-�|KǌA�3>݂�r9�3���L���p��p���f���2%����uv�S�ʙ�B79��̜4����FdȉD���h2�m5�\�X���-���Ymi������DNR�Lu���83##^��䂻)�}lٍ��BC�����*A��9��L��<Z�K���C�F�|���樂Ȧon҄�(y^��������K���Y���
�Hd�4�Q:4
�)Q,zֲ�U/��|y�'�Z����o�
�Du��ޯ5K���X�LM��6�� �1G8 0�X��,��j�0��"c�`2�
����H��G�
����d�+E��$+D�c7[�q��'XJ"���z�,�F��k]lnդ�FM�X�[>àR�[�@H��
T�V���d�؋: [+W(l0�w6�C~��,��#�no�:WM�Kj���+�͞H�G�17q��L�9��?!��&�7G�ކ��&��𚨥q��G�-R� S�"Gn<+c�9,�fZ�� D��|�� zhR���%[A����S�[2)���B-���8�����7�1���6[�(��� �bvQ����5F�#�Y����;��{�N#6�����t\�/gŒDH�rR�s�"�� TY��*�0��I%&��V�sؔ\�D|Ք0�b�V�S���[��~Z"]a!��9�Ă������n�ð��l�&!u&����r��n�g,S�`Hu,]7=���M�u�K7�y�x�M$-��G@KFE��BM}�ɌP��U˻ű�IFz����K@�a��="����V�.���$n�h��c��}��ԕ����l�ҝ���ʑ�����3�R�k�kk�fL�{������8b���픮�m�.��@'b';+��֌ 6����·�ܫ�Ω�ȣP��`�WD��Uȸ�TD�y��#9�iϖX�Z�[�m�WX)������-�Q�S�%4�p"ᓚz�f^���_&�GA�S�*�]w��w)Te�c_{����ASZA�)��W��)�^���a.IH�w�����]�}֜��f��>G�v%�#�Ӥ�DŲƑ�K᣼D��]��B
XZ�C%�x%ڈ�� ח'ָ�C��m>ժ8l8�u�·�R�ng�K ?рī��n�L_��t�?�E���^g۾���������B��7�"/�1����!�]%��^�����QZ\5�^N���a����o�n�^�%��4,�je�����6��qN��Dp&�0,����{E�G��OBd���n�^0���T3�f����vzr�s�F�2LSV�?v���gk���@CR�� �Y���&"�
,C�L�1�(y���7n,+9��C�2��ݜ��Y4����U�T����bB:n���������v��GKO�H��r\���M�����7NCe��tg`j��s�(��r	�J���`�G� ����L�����;�
���TorOY�&�#wg��Z�'��p߬�w�e�S6<':���}�㇬"��yPU�4Kp:��\������ӌXNc�ͬ�D���-�^y�{�9��7�:�"�`� yR��k��)T�&���}����׮/�d��z���k��=��&�g�6�%=���G4�>u���)��G�:���L#UQi�l��
=G\X%0���v�mv��>�͜����ذ�$y�e?1����:	�	 �>�n����_9���M�9�'&=��/2����!ɬ�lp���,:^_�}��[�o*���]ʞ�aQ��߉^D�ovq�zI�WeT�߾Ȫ簤���
��|����ᆾ �TUٳ�'uM���;J0�2T���b���/c8�Bgx�7�����w�/�g���=�t�s :i����Cc���~s������g���b�8��ԕ,;���$7E�J��*�^x�����/`���Ŭ`�c�c�gЯT�a�v��T�|���d��vƅ�
�P���J�ĥ�޸4����NW�h���t}���i$X6���6��Q�_��ϥz�H��S^ijE�/�p�L�n�8�e��Eڌ�^�(�'4�5&C�J�6��y
�M��U��|�k���E�䨪�v�4�K-:;(�
p��vD�h�G���$Y?�S���#
@��%00<f�� �a�p�o�?�y��q�i.+޿�>�,��2�����i����c�~��!�T������5����X�e����>K����,��ؠ�	��\�5b�����f8��t́u�+G>/�9G_�  ���&�.�ٸ#KJ�uLYav�@��+&r�2|*��b̡M�▾�=�yt���۠M�V ��k�;=z��S[|%�G}�Nq�Ϩz=�0(:x��l/���*�U�h��ʷ���Q.���bW��1��M��6���n:��e*�����;9h%ФsI�Q��q�ɉ���̋����J��mR��,_�Z��P� #��>Z��A�I9�{���-<Z}��:5��S���O��%�\;��������ߧUk�c����������x�8�c���cߝ��5����
+�>fØ��<�Jۈ燍7���b�P��+��l�)Jz���E��+�-��4]�\��Æ��@Z�U�6(+��O����g�\�SY��ߚ�ԙ�e�����h3�,�<T@vS[�m��'.hm����ŀ1�t ��4�T�	J"���uo4��vɃ�9���B��$�ޤo����>�h�S��D	�#ڷ�|�+�C�s�M˰1��+�9A�a8a�r�c��\lo�?.6;���R��u_Ht��.�/�z�{��è�^ X���rǒ�N����2��P.5֟9��]yŠPkzQ���c`1��lVB��7V�7��Mm��_�e�
�шX8d���>��^�(ٱ~`�2�@פ@-�������[�Y���;wg,����U�� h�T:��ʹ��7�Z��N�n�TJ��;;?4��iu-��1s���@����FB�~�B@#�]A~?�-�K����H`W�5G�{�V$�&����l�{E��5��U��t_T������.*X�L��D�-��Q:��e0|])�����6L�	�dRl⥦n?�7>8�;m?A���V��ࡧ?: ��� "h���{�I���$FC�bN-K�����B�){�%24�j&�3L��V�-2�؟Hw�ht!l�Gb�Z8�1]����Ϛ��f@VxVR����ŭ����c��5�� PQ��	<�e��U�)",)ضһLO$ʍe��o�Cc�]��.�n�^��^�7±P�����X�+R� ��	u�Bc���Aq�?��Ȯ��~�b�H��%�4ӌ�� �l�����^��50(L�����ȫ+�3.Ic���n.�
]m�E���d)h-iN�X�&B�	բ{]=��-Z�{�
�sT�WzUr.יi$�z�S)�l�bc+S���W��Rh����'l����S�X0EsG�}�'��P�"����V�M?<}��ʑ8��H��H]����=�f�)��)�@�	^���}&�cy���9�+!��ή�7Bg��zN/��M�bU���6Eگ�����)�AK""۳ø�`d��
�|�G�zW�X �1I��^gn_�~���餋�����u�M����4���4\`��$v%"��R����s^���&N3�@�h����q�g|p����OMdHN}�T�ڍA�wv4��������Hw_�&��c�����]�)wd?���Z8HCXĦ�BVۂ�;�@����F�D�Ro2`�[�v)�XS��P�m��SA��&�]�+�[�/�>�`׊{^O;TV2<�ö�=�/K�S��k����������ʙ��ԏ�H'#�4����j�c��L��&� �R�>��H�Ba���|����߮E$�+�j��~m{m���	��B��	�($̜=�F�$�naKӆ�/6%"Giv��J��$1�D�DՠU4M��0xX��ѿ�
k*�������d�G�(�_���;� �wU1$߫/�����Ns�b,�e�zR���$��T��ir�A�����M$�5�����$��%~p��tW���:����Z}�zm\G�%M��?汽���C
c��a�Ы�7y��EW��*s��?�n��h��I+k�X�bP�K�~�xܢ77�V�옔�������k�Zg\�n�
_ۦSHӺh? k��u�KNsۚ.z>y��G������ͪ��쨼�H�[}Ǧ�
�s���O8��9�Wq5�!U�[&�`�A��X[j��'���<��^[Ug���B��H�.V�4��NB��]��+�F��QatP�g�	�͎M�~�d�#�k�y-��,'1��Y2��W��GEmP���A>>s�C�l���\*?�:.B����iA���uKPgൈ���q�@_v�}z�z|���������h���0�!��}0�|��HWt�]q�$�0��@�3!�N7,"Z0��F�3aK���4V�ӵ��_�˾~E���A^q��}s�L�U5�\fs���+�7Ն��e��XE~H�bߋe�-R*˶�[��"���r�߶*7@D��9	-����ώ��CT�2��i#��%�GW�Ռՙ@�`H� v����v&���B۔��ȇ����� ���n�;�_t���كK�u�� ��ܭ�oEEts��X�]�ʶ!�A�uQE���3�ri���5�^k�����Q W��4�j�X	���q�����6�1n����������"+�FF�̇�]sz��1�lv.J�:�.�Ys7��h�0��.�[-����M�$��:�1�- �HW�nw*D'w��^-<�z��u�% 9G��K�8�6"?��4��k.��ۥCD�]	�����f&!��cX��s��J�gW�،� .��#��Ǻ���F0��I�IL��BloI/|�a�#�?��ý�Z��|�]6B�)�_��-F482�!a)A��1�)����E�� 4@���a�@��.�@rq�B�����ͼ�g��y;��i��Sp�34D��}G�a�u�s��\�g��E�@�G��D���r	p�E/�hF���n=�	���Q]EIehF��(2-Yx[���!P
H�ڐ�	[��Yٝ|�a[�"����`�2�5���+�j9�g���9��{Ƨ�W�-��,���݀c�|�r����R�������޷#oZ���ɇ9�&��)&�\\��=��q�b�U����i�y�8�eG��YֶLUG�i��M6�Go�ƔQEV����
��X��K�N'�iRu��u�e��*�0j�F��f ,�.
?�jP�}O��.��'��E^2�8��PV��q�5�Rf���Mo��xo�Y����7C �#�L�YW�/v ��zo_�
OM�x0���P+���=��0M��:���~#�>�<g1����� ˛'ݭ���Ճ����1Bk�j>Dұ��z!��eCR���qN1����+N��*�<�e_��n� 6^�*ƶR�F	��Zr684� ���D����^9��(�	ˋ�2�e#���]��)dEQ�#�j�{�6�]�V����7|y��ǡ$#��|ə�-F�uq��w��>�6S]�E
���-W���b|vA�mBǗ�!<>2���ق���-+� ɺ�L>c
�wLNcH$�p���������v�v(:\@��Tƅqu� ��~��R�l��z2�m|��~���w�b�zR���!���X�9���9W		�ڷ3��
L���g��:�w)}q�g[��M��+_�t��즳�����r�;��A�]D���k�����|���:OقuR����u"v�9&C(<t����&zZ�:Wy1���Z��T|\%GhUf�"�Z���.����f^QǤ���*��H\�e������L\�<�b{�b9�%�Ltm���P�}r%�EbR��݄r/ϟ���j#�Q�F�Z7a_ku�S/t��:�/���QT�o��v�>٦?��f�S��l���ds�:��>�`��ok 8�ȂyU2�s2�Q��u#��D�<�ӁLz��k��`�vb)	qm���H���Y�s��o��?��螽�|�1���p��3��)h׮P ��U�Y�uk��ɠc�qT�6��Z��SP�,��v�9x�xF"*0e,����%�(��!�ϊ:���'��s,)�}ͱba�|rl��f�^�w��M�Qs���$ Ͼ�ɢ-yw�!y! {��칽�FG�X	6����I
��+�����Ώ��CO6}z�D}O�A'�a�A����a�)�� LE-�<�zV��,;"#h��񀀦�#7�����v��2�����������0�8���M�"���!����L������	S@V/�r8���EV�(���)��F�Hk����dWV���\��Pu�Vn���kB~&_��(297�s
��d��Vw���eF�X`�k;��s��l�s�8�a��9Qn�E*M}¿���g�#�`0G:�����9�F,��УcJ�t�3���xЀ�	$�"ż����}y��݃�:)D��<��#�>�W3�3:1����(Oqd���"�C^�� �W�|��z��<�����d��W"a�ڹG�����o|�S���/��~��⒢�
i�l�e�����8�t�n�n|׾0h=	}��wW�L���R
.�>o�
�˹�L���Ԫ�,#2�	�g���T�K-��;|#<'S�c�֬�.�s�,�l��C�l���o�G?<3	�0t��r��!3V4^EF]�	���m��yz�zgq�A�]�����c�C�7]��ݫ��8����7���"?n��Ο
��^�Z�������fFi5�%${����w�ⷾW:�����љɷ���V9�Y�5=P�]��@!У���������T�����ⶆ���C��=2fF��8DPxa��G��`/�/>d��f��H�� �ڬ���sr���3��KY��KpS_�/M�}��nJ�6�䈅��1�)�\H��%f�����k6��
+κ�<���*h�E�3罍�7��{��eȀNv�3���˹�|H^orӦ4Mc�����Μ6���n�a�����/������UѪ�g��C�[����;�oNMMa콳�(������$u��r���j@]�2�`��U8-+�{����*,	��o����܇�{F��	X��Ox�9���>D�;e�KO4�J�JQ���n9prZC��Z;
���yr�/�%l'ƚ�u4M �#NAv�:���*�G��`�s�!$�{��3%�����z������+��?��fG��6�6�=I��[e�L[9����G�Ab���6B��� v��'Y��R�P�_�,�R��_[JY�����$��	"��t�N.��N�ǒH��T瀦�m���b�^�jWJQj�^�o�	�,�Fs�PԶ%]}�58�iTX{gӀ�Mz�wHOc�(865���g�>�Z�6'���,j�S ��{�;�x��P]S-�v��o�D�ow�r���fY��qgPW��Z*��8��xY�f@� ���t��1�Vt��y\Oh�&��Y�8ܯ�?#���ٍ�;�+D�<��K&m5�0j����cX_�`��d�~�Qp�#���:4��_8����EJ_Åh�N(�Ӓ�a�օ�̈T�%Uz�Nş���V����X�@���֔M��&���N�ZWt?@w��S&sj��;��;vI�?�!�=����� ��s���~]�fh-�����\�{G��*��ʭR9C��ASz��W��4����8��*�pd8���ʥ+�DGh.��@��9�����.��w����H��;}S�]j]���
R�a�֔k��+,�?޽�(��1�d����W�^�b')�����.�\ZjMZh��c�L&�5V�~�D����d�T>�oJ�0�q*��BJ0��$%mۋe,vtj�����unDY�^��w�*B ݮ ���N�L��PJ�P�Z���(�O�j!��aR�IG{,)�Ħ�+�q.��H�,7ֽ](9��B`�Iv�p�*h�)5u�!LǀT�{I8��'
.�.���G!���4�3�*XN(n��>���0�᳋�s�	 ��U����6���Ų;�NjO��B��\{3��}V_��#�Ja�Q7g��AL��K����te�m�|��*Y����d�&��%:<�n��,h��I{�N>�$NA�$�(��[�&KF���r�/�s ��0"3�%N�bbogL�#M�w2~�}:�.Ȼ�&�* �?ӕ���-L��h2��̘�j��?�P��J��\G���t<�|�ox���O�K�J`ް�-i���b�hi���O����vG$�f����O���lB�AL��Di�E(B�$�OY ��L��Ty�gW�`�
�h[�����ީ��i6Q|����ĳR�0�l��7������l���Pa��\�m����g�!k,���r�d������ݰ��=^P������+H��7��������r� ¶6��AӌN҃ ����o�c�`Ȝ.���4���`!t���r�%��i��h�������3��#�ف��ODk�Ŷ��D�?$5y�T�c�yBc���c��&��*RA`i��y�m����%�ըj��rY;ɫWK�ԾB�0۪�r�n$�G�	��Is�hfLU��t�t[�F���e�����'��)�����uaF��lb�{
��r��]�^E0�=����G.�/�Sޱq��!Ee\Ոk��,gU-�\�b���;�X���ʭ=��Few�۫�$�%M(om+��t���/���#�ø�܄��6���A7���IO�w�	�$ �����>������ڐ��Doӑr��s�;��I��E�E/�#L@���yV�۳#����(n��{�d��9��������Q~���m����6}�P"�a#6	���g!��}���(Ʋ�P�Ć��0�6g��ޭL��Xշ��Z���B+�T_g���\I"��Gka��2Sey�Hr��㇠��|O���{H�D������֋��\u뫮5�#c�I����w����Sw�EL�6�۽:�ٝ��|YL$�%.�����-(s�m�|�ㆩá��1���g��!��r�����I�w���F��5��YZʏ�T�{%4�Ff�pyD���G;'#�����9Dr<O�c�r6	s������F<��W���Kh�e0�۪��^�?�(.U�$�U�� N�厝�J���Qy��J�}r4� ��\�������P���w��~[V^����[6���+���Fq���U%\}7<��\nc�k�R��M}3���B�&"h�>M�V#H� �L���B����)��:L0Ŋ!�"��'Y���C@ ��Q�OW� R2���갚��߱6�����Zu��ZC�0�,C�exin���p(���6�,��O`TDנw�� ��4N����Dz�����ܱU���$x�!N�e��[�o3�/�#̩X��$�>k�p��\n�|Q<!�::^�ZR�5�m�ƽ7�%�5@Q%N���H����.��J��t6vi?�BB�] �%~�O"_nۀ�f��}��[I�4T���8�!>�)B`0����ۖ�?�7J� ���O��~V����X3_޼'�'��r�ѕ敄��k<K2mu!���J�P��U"3�2��˱Nb�7U��!%A P~��
Z�%��~a���v������Q�J�B_냏d˯N$	wr;E[� ��_���Au��>���c�n�X��B�����T��7s��x�"��՘�e
ᐹ��?��� ���g�p����ǃ�˅!�"k�d#���"My���v���qq.(ea|� 0�뷱�[��1\^��A�$���n
�.:��I���%1%�{c��+��ף#}-xH\w���gb�=^ſ%���M6�ȏ_+_t���n�@�y�'q\�e!E���1����T�QA�
6i�4�q�� (��e��%*�L%�:7�z� ����廄�r<���1�.*����|٧%n����D��v�D�?���j�"�����HU⩍h���� +Swn�U7M��48���ʶ8�e�+X�{�L��p�|�MO�7e��� ��L�Άֺ�G�4���0\|�,"t�iN�x���_ <_�k&�_�O��<z��K�E���e
Q��\)I�y�x�}{����ǎ��Pgl#�Z���.���Ea��| /r�hm��o?�� HZ$����1vw�˻��O����4�!�@��}���t�Q��[(;p��F��@>���b,��f���>H��Wz̛$�Bz�'�5��M(�ty��bʯ���7s�Ŭ��K���ux�$�7��+ʠ1�Q��8�sb)c��竍��i�N�P�=C��������()��-���+���Z}^�b�h$�;3��cp@[h}4Ѽ
�\;NDȁ�k(+��w�X�VnQh�$�?h�@0\0�n��7�J׀f�v��Xc%_�SL법�\D�T)~���~��fk�[��	��Av���%I3�Ï��sD�O�cV��6�6�1���.�
��T��l7z���и�Es�`D�ir��ki��]u2�<KVS-�^ZI��4��L���c��a�/�}��R?��6H+!м���*��b�)K�0c�_�ͦ^��k�`�����` T���3I��r��Wu��w`��c	��%_]?�*���u=H��>�M����7f.�h�;��Xȵ9{藇�F��J䧕����T6-n�q��󃘸�G�v����o�&鯡~��P��#Ӽv�ΐ/���O��� .��f����9Ϝ��Z�x�A��U;��i6N0� �5�w���ެ� 4Fd�?L}Q���RC݆�f�X;w��߇�}��f��K��E�wSۢ�|h1Lo��z�^|���Q��~.�B`d�����#TgU�z)q����k1t���,�Ϻ�
:�.�3]��[K�)���.�#4��*>��x������=g�M��kߥ��E�Ty�O�`�X��=�UԮT��b� ��sek�9�P@i��&��Q��^�U�/+�D��g���OHw�G���	����=�*eC�؞�y�)(�r����e����*[��X����*(o��R���
��#BI���Ob���|��{�Ȥ���T2�(<�-׹���(�.vp[1��='jc$c��]1%�����V5\�� �*ܐ����.20	�*��.Kfp=���:����־��#���A��m{��I-Γ�	o�;���dF_�"~�q�P�I����MҪR�Rwr����yĂ�~�B�'t&0�%+������{�� ���(��[�'Ѷ�X�/�7(�z��&*�-XQ�y�������"lG2�t�(��LF�f]Ǝ�>��ܺj�s�u]���n�쇋8G�����*�;*�0"����C��	�P��Te�'>�]F�#� ��9�b-����e;Ч���v���� <q��zW�>hr	��ĭ�LJ]l�
��� ���x|�Q�)�i�U e�Vڔ�=d�����cǈλ#Р3\�ሑ"td؍�$gg|ըvy����t2U�g�ooY����ۂ��X[�m��hvr\[v>Ƃ���mMj��T/�;���w���$A�<4���Zr��
��yq6��zn��d��+�Ù-�<���n�*�w�A�`R�;�]�n$!���$�j��ݸM@�ʇ�t�W�7��>c���X����Y�H�K4���:J����|k���Ƃ[�>:�1-[|r"��o�uo��W�3�ߜ����j����,�N�����䦃S�|0C���x���$T���2n�\J�K��<����X�r�7��7�@�ޏA�bVG�Uy�6�Hj������~����6�iɞb4�yő�5
XҮ*0�p��E�y��+6M!��+P�6��&�u"7�-t��fT��eáGu�F/�0�?" EξE�

d�zDW� ��г
�'"��2�1O(�!_M��)�w�
bU��v�̲Z��0G��ow3�Ob�w���1q⇟��ʈ�xU-�_.�dk�8����R� �=Rp�UFZ/��\:j9�`�c�ꇱ��oG��j�ڡ�b�C1tQ��`��CY{�9��-a�w���r�]D����S�.�t�}�c���3#��Ey=A��Sy.N�ǽ�O�5���^�M��
˟�c��i��oT;qA�N�'���ͅ����6��q�sL�����y�	]b������ ���e� �W�7����j}���E+"�:�rs+��v^������P%NX�o�Eh~e���~!=���b	EAx�3P��m`x��s��K�
�,�F�.�2�efWM�������N�2�=v�`Lvеf/�롼¢�ͦc�2�t�E�aʝZ�ZG-@�����.��l���ݐ����׋�c���|m\���e��w��B�	�]����,۽\Y�?�\����� O�/��؆}�rK��|�H4���g刾k���+鰃64QكA�K?7���]z�H��\6Q�q|N�
�g�]��k듌T���gQ9�
{�^ �c]$`�iz�,�]F�^e4�9w�������MĜs��@�3�]D^�uOPڋ]��Fc��,NeY?E ���+3&({Qf`A��&m�Rvu)����o�M�c�K�jNR��J ��T*w9k�A)�ƛ}ʰ���v@ӮQ�� V�/0�H���y&�X4C�%g���-�A"[ڋa�M�_��NƲ�U\�G�yK
Zt\�̍~.�e$&�F���m��e.� 3����W��_������y9j1��#3���׷���GU�o�se[��BoJю�7ݮ��O;ϵ�1���s�E�����kh�'�����<�#ʗ���s��E�|t�?��A���QHׁc�����O�BfBwsz�oگl�6�@9)�u;�꺚}�I�,���i������������3���r2�@�^�5r1�oe����.�+Z�_m�, �L
�*&�&ٷ�O�/����O}����@�,��{p�1%V���nh:+WV�#��q)��/��W��0M8�|����}��m[�hFP����4�m�E���#v�N@��G.�G/�����q�{���X���|G5��=���_�_�հ��ʈ�q�_�_qDL���q�;&&�,l�"e-�	����{-�%��c�X�l�jjN(d���ԍj�2�g�ss^�����Ea������w�������^������=A�2M/7 ��I�j��Ix,,CK�O� ���3-I�I
�/�͎2[� ����,���d�����^��t�'�eE���tx:�\�S�l3|v�I}<�ɗ��8m4���Db|�>����R��U��jv���
�,3;�^�x���=nmKdJ�j�4{�Qt-���E���h��`C�B�j�?�*q*U����}��1��r�.w�sXJ2jD��ۑQ]���x�\�{Dl��F�p���x]��,���X4d��Ӄ$��v���4\�&162O�Za��ݝ�	�bR�/��D�3$R4���Q_�'	)Ȅ� #Ҥ;�t J蟸�]�I��K��j	 ��ZD�s��r up��u~�=d��{����R��GFGy`s�%�$&�[�Ǆa�J�x��琊l7��P���E���U?T�UNIl���נ��q\N��=�rb��i����͓BXЦ�H���2x4��F6�p���zìB������� ���YIH��w���Q����ǝ���4��B��H�i�`#9;���`d�y�Y��ul�VI�Xg��w#\&�=_���D5�,9}R�n��_vW��C���D����U<�!�A�j#U��?PNW����W�Ô�ar.�WP5:Y��^	ME���t$��2n���R�;d���V��Xh�1���(����m�o����T���1t_�����J��H4�\n�H6
_;��H \����_�e��`�����@��>�p�����Gc{����[�`^������%h���m\��C�}��Ie2�{}��D��s@\���v�	|����M:�`0l�U��>�h'#fѢ�#e�)@��{1Ș3��ͷS�m�#�T��t`�>��FQY�RH�t�HRE6-�H!S�	G
�W�������9�K[�<f�M��e��U�{5���6�jjp}���T\ &�5��r^>��9�P�bY��4�Q��B#ﳩIw(�=#}��'N��N��R�-(.����H{��!��r���
��㖅�M&���jЙ�	E9��h�Z��;�<�e�(�V��(�G�J4e�l<�\v���Ʊ�� _w$q��j�̒�Fˠ�����D�5#�zTy�M�*]�*��������2l�����l~��{{G�HO��Xp�U�gԓ����3RN\򐻠7�j���r�P���/qa<�}�] ��^�˥!m��j�DRG�+��瑿���=!����y��̐�-�X>�率�kQ��W�Kv�_Q��QdI"����_�U0��md��#=s*������w�ӈ���Y��w]���}#��c���6���m�_�F�C4��u�R���I��_��F�S�����h�Q��j0��_#� /�q����giٷ��  h�vS����!*��f��=Eh@��I����%/h��5�a�	3oM+"[�+�g>Ώ5���uh(-%���X�c?�4�U��ض+�[��f��.���k,g�����-͏��S���t�{"aI�������D�#�7Y��.3��xYI���w�}�f��c�x��y,��5+X$�����A.:iPf˕S�e]y�	_�ƶ)=�bf�2D{�Ș�k�,j�wc^�7ȢwS'H�I;Je6����]jo��N���NE����j����T��V��ܸ�l�\�@�1'�HDr�]l�i��,�,�t��t��&�Y�sMJ��ߢ�>8�fc��J�9�S��(�[�%�%(���A���l�{�o��|7`F2ٵd`u/P��wI��}]���u�|�Wd�-X� �t*���]�Z�T ��$F�g���E�fws� U��'.Jk�����UqU�2Ɂ$�	�}����0���:�ǹ�4�ش�z����u=��%�e�_��C���4��	�|��/�x
w,o�E"׋
*�ӷ���1��z1�UUi�"b5�����/L�����T������s��+H��p��V�1���f.ҁ�4#�5c@�"�B��ӞJ@^pkN�מ���G�˿�6��բ����G��Jv�*�a����Jԁ{W��M��c&�}���IML�>�9
�<e�v^�zWf��&�A[�
�d�+n3����J��FP�����KqfY'\ �ΐ�g���|�T�b�,ŭ��7ʵ�E4��YV���_��4=�԰��q7�d�'خO��&a�㾾�F:�*A�}��7gM]w���=/^�a{s�'E��$�F�?ɺ�
�h�޳8࢓���jY��2O�
�b'��ϳ 4ƛ��|�L0�/�y��Z|M����*0��
0�r�
�����A_�଎N�;k���n�ri
�:�z���`�t��,�N��Y%L��^={yWe��~����R��7�J3ٻl~]�i��w��a�}���cwצ!�	���!
yĦH~Se{~�*	���V�N���	��W�$�Sa5�) �V/�>�3$�g��% ����'�
�-w����d�	༏�&��.D 2oa~"ui���U+�� �Q'nQ�������3���H�	�.t���jَ�׾���2=���#����b�=i�˷�C��� ����e�է���-U}�
 ƻ���d�E��r?���LĐ=c�Fy����or0�RN��2�M�����:_e��A�_���VV,�F�5}5?{��9E]ˌov����q9��:�h��`R_��qP�'��P�h�P��z@Dܷ���AN�d������j9�<���Rn�z&�Qv������>�ŏ��e���ufM�.J�����A�c,����]�.�=�Z6e�s�#��=՘=`�����H�
�=��&ح��)ɿݞ�8M�,*��"g>�w}1!�c��hD�J�.pF{���f~c���y��p���'H��u,���BR?^3G�M)ix�jc��a�jiz�l�*�S�	-L��O�&���YӹyI���J�l�+z��Q�M3���!���8�J���^�<��殼rV�҃�&-��BT,#�SX�>
��:�ӗ�@^��l�Ʒn�*t	ǌ���\��I #�4����V��k��	
�?>fS�ʑ,�{ T4�*�{P
��Bc�����a��YJ�s&j�3���"���l��$H�<VV�-n`�r͐N%V��#Y��znc���w��̡x=&�|r[%��J)hiqR�ӑ �	\K��+�/���������1F�GX��Ģ�*DZb��bmL>��;��cDrG�ZMqw���3������*�]�ZF��;�4�#�f��:�:���r)��:�'�y���S�v�h���kk`͔B��5]g!�����_����v�k�dV � "�Xܗ��ѡ���9ᆱ��������@���53�=<s�oK��?��5��keZrf���S���M!�?�umg��o�v�d¸`�� �4��[�G~ѲL3i�}�#u����}��VH�(ί���-n����]�!3��RL���m�K���r��n��ׄ���'��s/}�ƒ���3����I�|�C9�5#�[�z��!F�u�3�^��P��b����k!�Ú?�J#�^�}n5���**��S���0����z�$�c�j�[0 ׂ5��>���T
qH �n�Y}ѝ:���k�H�C@Fc��`n�P�����g�e�v���8��7�yGQ����:�e�/��oKʯ�ۈO�ɱXװ��֣�y�ly8�z�m�H��3'[kBL�0�H䤡,!�ێӛH>$P�Z�: ����7�����y�Ԅ�Н�v����\Ik����x�l�(�&b���4!	�P7����_)}r��@��������J���V�Q��٤��c����6>�#��tSYf�/�����k2�k=�]�u�q����2�!K���������tp�rz�%�8AD])�b�G
ӭZ�Y�����K�=ڏU��Mi��N�+�B��L�s�����%�I-<.Tn�|��L�.����vT�
����3���.��E
әP�^:�^6��3w7�|2�ѶD�6�nԉQI�D��1��֘P8�:\�O��ߪr����f\nJ*��X\
F'��'Α� �
b��r� �\�K-�g�N�v)l��n�(-۰>����mē�%�.S��������d�U��B,�
�5O�^�ev{���PY��=Q�?�0_�rwi�Q e~@�r�T?Ԧ�I�ɴi�dWǯ����>����4�_\,l\�������"�&�@r������BFXU�dL}^ <u��\g����Ifo�z��qJd�ˎq_;��A�2&R�/���C��/��7Ȥ��^VvL��1ޭ��5����b��&*m�D6�_�|�C����M�S��uB�|�:��`�����qy��C8���[{j�P9a��GX���=���c"�Y�!�T�..S��/�2z+�ح��v�"��쇨�$�VI`>��_<|�����zD����<��PV_6���^0��D�/�����(�H5��}����n1�-V �n�t�^t��R��Y� PZ�=�81Y�	a���a�L�$�k_�l�PF��秦]K���8����+O�����xۏ�~�$l��'/n�DEÂ�q�w�Ŗ�;\�؟��؞�H��;�P_H��8�@�3/���4�Z�X`ȴ���J��B�앻�I�(�ZDB��07��m7������������LMJJ�
q�����la�ݟ,t�y�㟻iE����lreNc���o s���Z~�۸g�w[L�b4��Ƃ�w�y%��@HJ(�/N��b���2Y�Y�Y�|���FY�P�:A0�e��蔲} �v�`��{��׸X\�p�����X�s�N�@����y�x��?�b�O?tAf��>�VY͐�;#7�6���!��dI2�~�kŘ�y���O���ZJ���2ak�B���x"��-.�_q�t�Q���$���J�t|A��m�8��J��e�mW��ާg�83���)��E��/?c��z}\����=S�,B@N �?�b�῞4x�+�sռP�M�p}ӁH"$��J�����}- F����U�X]�n��/,����9�=H0@Nc�&�'϶0W;p���0�����G�ޮV����$��Ǘx��Y��Ώ�S�l:�c��O�b>��3���C~��G��LT���W*!{,��b����҇�"&c�t+��/�?*���*|#��FR��|w���cA���e+Zٶ��i?H 0�i�VX�#�����I����G=���C'=�Gw�b}<��
"��A0��Uc`�҉Ca�ga�u��S<��I��C���\1���PG��JV=Wҹ,�^zh��3��slɓ�5"����#\o�c:�pv5���deb~YRNTC6��\�4�0oi^;;��ư����Y[~���P�ZQ��`A��Ȕ/\[+�``֌�en%y�;���rx.�A�f��nJK�_��u�=m�f�����r�l�1��D�8�%�
񗊊���`��W��m�4A�|�R&ּ^/[��7�C[�+��@�\Y(���2۩ĂQ9u2%�ы)Y.y��9p6Yi��ؓ�U_m���Wj;��hI2帍�I���ѦK�&�R3I�Bŗ	H�&���q��dL�N�.1�����0��3�?�����ۑt}��"��HN�;K�1\

�J�`��Ż��v�>
�"=s�txK������{ZC?9�;�S�@���R�_��6�8π��`5d�@ݼTH������4f��i���ڜm͇���㻲���9th�c�yΠ3/� 3<����pV�|�s��3���O�.�鎣�!���,HM����Y�!�m�"C8�ȾMjm~���0�&�#<��n�A���W�� C���}tsp]P�&��8&YVw�p�ؙ_��=_�{���`�Y��~ ǲ: rEw�Y�������I}�{�h��gf��X�ˇ_�H��U���;�N�w1b�����B��"�$�����7�-R�b��ʫ��#��9Mn�w�{z�U �n=!�3�4�,�u�~�8a*��h��}�Gଭ�}�Z	}U�F�^rOTY�]щj�{��i\�k�'J��on+����xKwD|ܰ�j�UyN�͇3eÍ��x��Cv�1[�%�h�.�	�2]b���`�vԝјQ��� S��k9F�bf��V*i�����5�׍F1�Ԇ�����SQ�y���2��ĳ]��-��/��Ǔɤ�`�U�l|}�ä!�T��x�כM~�9e���K3��J?a����1���%p= ����]w������b]����p y�9+G]�&}lH���ph=qT_�����Jj�<+?g��X�y�>��}�&�@W�[c����]N�Fa�;�ZsA�9W�v���͎S�n3�O�}�Rݺi�� �q�;�?����
�sh�X���L|���g��*��o�.&�rx��U
k4�͞N?|Rk��
`C�6�f
;�F4E������g"�$��$À�����z� |l�cEl�/�,��{�t�.��q*ZvYe:~�d.���Mf4-ϸI��w,l���5O�̃w��?x%B�r��p����<U��W���OA�]S���"���;��)������%���'mRa�簥<�su�W>�y��oC�K�i�?�U���q9�=R����A�=��k��\�H��=�eø�����&�&�t0Q�\�_vs@�^����dt+����m�ð���S�Pf^-���������	�<6��&�Aԡ���]غj��e-����m�Q�#侟z�����}R��א �g���1�U�9��L��B�鶗iӇJ�=��O�gF=e�N/�զ$�ir18Nq� P���y�m��f��Ո����ԃ�G���B
������/.ӕ�Pޗ��Ws�ލ�ǫ�@q�{�y����y�܌������A����:aD�k1+��9</�A0�\�t�ΥU��՚r �`���

(w�B���!�"��"�Ț�s�g?5�M��; �l�.����%����s�o,2��R3��[�f�j�^��"b�L�N�q�v�@E�&�MG>���fm�.��:�����u�$%�x4�y�x*�gܘ`�#b+VeR�J0=Od�S���_s�6nuw=��uC;H�ɮ�,ɄP퇡S�'�>S�S�J�Z�g�˕���Y&�,�
��5ݛyU��0��#���\sf/B�,̠��:���)ҖW	�}�>��vg�ͯ�ky?L�?���O�ڹg�2��F5z�8�}�U��$���;�qZ�)؂`��˚�����;K��>z��s�_�[7�2�o�R1uZ4F)`?�&<��(�Z�B� o;)O��P���)h�\>���C~oה�۴��~R�΍xv)t�^~Q�{�ԥw#J���X&�ج"�㼷�+&b*�?E�oΧ"��)%����"�#�*�jR����TR'\��%�)�ػ�P,�0@��fNY}(v�rߙ��i�֗�S~v0[W3��5W3���"��L�ß^X�Q��v8F˖�s/�=�M�Cl�Yն�g֍�I� چ!����/ U~�	8�_N������E>>�ѥy*hd��&O���@�M��ĉ�T���>��]daIM�G��`q����;$]��s�3��7���w�A�Z�)Nz_LK�d)'�.�2�R�
���E�x�c�4Y&#���@���YOj1Jp>Ev����.߱9�]�
b�tk�&�,T����W<�%�CO�:�U�T� l1�LhZ�[l`��ڮ���W���:�4���Z߻u�:a'��ڒ��̲��m?��;���љ�>�AJM�p��UL�@p�ޯ��B��XU�\_2^���ĝ5�AS�*���F��<�F/�c׳��U<���g�g��[��Z}<��H
*���+�����������TEu4x�i~�� �O��j��d��ම�8O��d,�<Wõı��[�[��l�C��uJ���T���h��e[0�VY���������7Ƃ�PP�:�R��<���D�Nv�:�+��8��;�Kc��\��r�hkh�*ܫ��A�x�G��n@�w��$O�P5��XׇY9y^�o=�3�gʤ�c�b�!�ea\�2G�o�w$݉8z��T;٨��D��-�뭮���\��y�CZ`WT�����i�F�V���"T�Xb̯�D����ɋY^{!����殙Y���=�rj��_�r�ܻ�p�����P��4���gX��&�������rq'����z��i�n��V���v�z��G�9�@h�
}�� �(�|Q��8�g^�+����9PSG'��`�[M����P�N�D ']��i�1[���y`��1?�7�^L��ۧN.���:��5�PP�J��U���Y.�V��
Pg切C%+=ntU�wc�mB�Ȧ��e��mi3��m�x����<��<����ȉ�D т���}�`�'�n�4�o�9��m�V��M�:_�uO(V��["U�J�����ѝ*B��gN(���\Tr�	��W�&��
geFQ���hʃy��E���?
��I�io��/Cs��������Jj������Pc����x8�XG���$��W����uX�R�l���H}�[�/+�aZ���T�N��H�ʕ��� p_Z����cn�r؆!�$�����1&��C��r~����F-��"�сYw�̅f@-V���"�'�@�yY/N����Iz׎�w/�d��+"+����j��=7�{�V"���GunNyLϕ� Z��W]�?>�58/"�����;��&��Q��/����s:��u��5R�b�`z�,�7b���ص�{%g��b?I5�2�aH�D�;�1�H��?O����I."=|�Y�LE2Ӌ�?D�u��������9�(t�ݾ�jJ�2V��]����_E��Y3��-��:עwp���Rnt�K�pqTnI<@�`Ƭ����ɚ״��(�f��v �'"<� 3�S���I`�������s[1��2YյΨAw����^��ٴ�xኚ��	��k~����+�<�����v݅�1���� O����}�ר̗zr��ؠ�в�,�����c6�t��ŏpV��UdV�3���w<3�k�Y��f��&����'��x�W��r�[N^=��s���Y�L�;$c��강$Q�S���Q�������`�K�X�Ih�6�k�ɛBۋ;2�;]ܒ�;�j�C���d6(�A�l���}��;"VBr	�Ļ����@�)�d�t�`Q��kys.u�z���n;�nv�!�Sw�Z��bQ����I`��g(��LC�04�d3w���k�e�0����c����XםH����+㌒Z+kZmq�����zZ4���L�ș��,`��"�,u;�0{4d���,�vŅ���k�r�V�* m(���yH����,v�~*a
mV@����)�����dNy��v{�pbj���5]���61g	Q�:פ�nS��M0��T��Ψ����P�h�k)
��]�֞i��~���/�1C v�&�v�/Qζ�񁲆��E�~�(L�%�pp9�)�'��U�Ӧ;��7�H�G�\w��J����|��f�`�+Gf��'����k5��Fg��8KɼL&�F+H-N�:o�`)�S��)�p zw��iy�ٻ�ܛ(����>�ti���s �i�T:��(�˴��p�FZлm��Fʊ�#�`�l�A����L��Ve�\���F�OkD����>}a|#�����*�_�N�-�Ќ������\	��*!��	lf�k��b�(K��ܢ�q�(���̌���L��m��uJ�)���� W�P��*�lS1��NkK��w!�1G��I�)����Or�.�0sy�&χP�L������zo�%ԇ#?�b�:�<!�����C�Mڇ�=�dC��p�^��X�D��Ox�ߨ��I�̄����	1?�d���C^��S�A���#������;�~��N����3+��V	�Bb�%ׯ����\��a��2��h�2Pb7e� cC� ��̞"\`.\,d���Y����BQ�n@�n�=ڈK�T��bG��6��bVG'ȴbU��oM�Wۘ�dh�R�M����O��j�
���e�-S����"�~F�·n�D�7�eH�j]�%�u��A_z�K�(B��7�KuvH��#Oz̷l�~�9�M��<��A�K�s�ˠ���ao]���\\�Ϥ
��L�٨�!YFTNy��zp���g�'��W��OZ:�ȸ[%���ΛǜN���N�?LJ�M TCaSt��Ga��|�d�J��l��Ǯf��w�TM�̒A��=<m_�H�1�G���3ڟAxE��f�6\e�P[��_$�W���g��͡�����wp�gm�x6-U	����fK���1j�W�	묡�@�L�?�>=��&��y�ۖ��<ŞO�)���Ի��s�_&����n�>EΊ=.��U�Fh���@�F���zU��Orniq�8^T�yp�Op�[��rth�����J����!#�"M��3m[`��u�@�+���a�o�(/�w��x|za�T*@){e�/��1w�8�k��uB�;���7�c!���Pd&*m�BP"e�a?��'=��5�m�չ|�:nKmm��W�v�]�8�����B\1���s0���89�hg�[�=a.�u�<���A[� ��uM񃈣��)��eN��	�O|!d3��FǠ��i�L|ߝ��㤟�F.�E}�0ӿ|�E��z�)ڄ9m�8�0�O�6��������:�T��n����a7 ��l���M���Ď���ϵ�e���gb�-�ͶCѩq��q���D(��3�*`�zTk��Cq�*vuq�Q�P���Vx�=I�)&��U��=5�vj��p7/y�}��Q�z���z�6M�D�l/� ����-s��zt�vyQ��_�v&+ɇފ�g��c�W��1�\�x<��ܵ)6��Ck8c�ن\&ØA��+ʿ�9t=q�Ye��s7פł�^��vd_�����l�dgC9�\��]t���ӣ�� ��j[��Q�pCPb�e�j\ޚך���]����0��z�)��r��!�Aq�Tʻ>A���L��oN̟�ڊ2���u3�ו�p
��AS���A|�+��&�����l���f�k���E?f(o�{��~�ao�錃kÅ�!$�^:��<T��h���6��P�:�P^U�$���ޝ`1�Fa�) �-=>9��>`�%��4�LS@��#��|QF&T����v	\�{C�}ngV43ܟzK���t���&a/A(�]1�|�6���uCh�S��7�ZCBE!�}`I��B�������QdWaڈ,�ڿ��1�F�o��EA���jo�~��8���*���y[e���h���l��0[�xE�~Gq�YKȆ
 ��U�)�Z��@b���;�_4�=�R�W'l���ZbK�X�jP'�m�J�7C/��Cgɥk#xo�T]Br7���3���*��PN@��K�a�1c+��/��W��v�J�h�ԤQ��d
d���_��\�/��j��X���rüd��ʐ�"	I����L\Y8)s�,h�dk"ؿ������Y�),��Wqg��v�9�,K����~�O��5h����o}چ�R-�(����x��{Gk�ץ�'�7#��.f��5�A}�V��E�r���=3����=NXT:]���4
�oп;,Bӷ���k��/�ǥC��.���u���qeN�_G����$WP��͛t5#�
t��#�%f��X���p��U�tp+�i1%$F�9TM����# ���hsbP�g��~g��j!�z�t���� ��]#����PL4�EP8�1-Ӵ�5l(�A��6Kk�;!x�_��㬏���̠ZL�1R�P���3�������E��o=�<�0\��M�@K0i�L�6թǀI.�j*��C�@��.������������j�����N���Ά�:X�Z���&Da+�,�!ܛ0M~�>���'��"r�Y���G�ݧ�U��>����]�{݄-�NSÅ�G��mv�Fȼ�ǌl��7�>}l퀟��;c�o6�/�%2&�L�hl����㸺��R�T�dG�Tb�p	!0���5N��3���v�P22pXw%r��5�tN�f?׌�T䙞�����D|8�=J,��4�l���'д?�j������m�\ش���뙮�LRöyk3lb�M��DI=i�%��
��^̬[�|��.u:�v�-Hf�p�ICߗ����p����1yJ�e.O�ICw�=�6�r��сy:T�k��h�m�c5����Mݜ9%(x�z�)��X�=��v02�V;îc$�g1�Y���NO�$l%�0�#�[S��7;�@�́��3������T�OV\�ħF��i���
����C�vQhm\l�{��Oj�^�ޝ�B%q*�vKX�E��֚䂸Lsģ�Iei���ͥ�n�[��0�^�X��a��V{�"7�.�D��]
�hU<)B� �8]��
ʌ-ʞa��=��Zg�to��&�Q�u���#��ޘY匌�l{D3�Ԋ`�Mp�~h�K����d5@��5j%��Q&�$�2�x��;h���O�=�\gۅ�*Dۤa�	V��ƐM߃V�4,
.w��Ǵ{]�`��q�!�Q�3ov��������*}�w��ׄ�^m&�Ybo���W�Y֯J����,��. RO�9x�.$���F>K{�+����w<�4�Y=�C������;+���E 5d+ׂD�T��&^#幞��k����n# :ް'ߚo��q�Ȫ齚����_���ղ��{�*�E/�|l6C����đ,���2�Ao�I�AJͻ�%�N�)|�^��H�.!�{l�tg���Wu��pi�<���:��ea�T�������A�?�pX��Rk�џ��f��KvT��.���y?�H}����<��J4X�U�4������7��a��4���x�\߉ttl�u�0n�Q�G�����X�S�)�������+t��:�NH��=���rW~������M��߆��6%!bI�X�]&'_����"�*S���R�FA%
�{��[�iyɨn�s�eq�X�������ݽ��A�y[
l��)��8�0=�2k�v����y/}�-Ѵ��	E2l��p��G�G��1lp�:v/�Zw�Gő�%���#?�%n�1)��Y�@ֶ�����ż�󵇩��tG_�q�>>I����NP��h���H#��bp�(���M#������I~p�S�`χ^�!��h �s�pN� �ϓ@����V�q \';��>_�9����Ǒ<N6�AY���6�E��2/�p��7�QNN������@^�)di�W�1tU���B�Yޠ����9�+�v�s\Ը��5��a}WO�'v���{ˡd�M|��m�����P����n�d���I�V��u	(�M!���@���)�2N9������hȡq�)x�?6j����0+h8X�'HE��cB�)�sE�q;�q'�Lg���O��ԟ�Op3.	�ϕ��|Bvk�*��*�~菰I���v+MĀ��o� ����m[�C��5s���6�%����)���;c�/��Kך�%��4�L�,3B�N���@�0�ivN�$�m��t��AR�V#��죢SGM�?��U�Q��&D'&ڒ��s����J�_�['�
2M��SN�~�?���OHɤ�Wyf��2��.���oW�����E��t���oؙ�pܲ��������|#�8e���� �U`J��h�����Z!�N��XP͒^U��� a U�HT^�g ��I �>G�9R�mU�=��|���d�Q�`�
�U��oV@0Xڲ��y�M7�Y"������Q����3'4����cM�Y�~%[�H�(˰��ʗ��>g�F�Bh�
�9�$�gA��Z1*e����xB���;��y)}W��<���-��RL�
�A�rd���)�qy�\
Q(Q*}��e��l�I��ig%�>B�93������}n_������I0��V�7�4=���/Z[<�zrxgF60��NԼ�r߉��G���_U��#��x��3%�v�|�������V 6�t��U>Pn�� ��M�k�?�i�l>�fGet֦_�&V�;U#�ȿ�IM���T͜o9v�q�3����Jt��-��cM�*��*w	��$g�ŭb�-���O��/ά �%C�c�g�83���3������6�0T��y�=.ï�9�Ni��1Ԯ2&a���@L�0g��ߧ��ߐ��>���'n�*?������3�s�/�X:4�ڝ9�O�k�4�Dx�|�{)�4 �=�e�>b�I�kO2u���]���&�n�r_�f@_�3���r4��D�&W���?��s�ſ��V~�c[LǼ�|G1�A��D��5�����ο��\󏷂�Tӑ:6b�$䱆�Y.�7���ݬ[�07T�W`�@~Co�JnER��Bo��V�'X��-��]S��RQ��9�Δ�VF��w��"5؁�Dd��Cʜ3�#�����YLxn����UE��P�����'�ْ�� O����r���"���\.58YXpe��������°'��9xl�)=��D�l�y�({ө���`{9v;Ƅe;�h�"����T��	�mS70.�zW�E�e�a}ķ�D���H���{4�J �-�D�\c�������#�+�({GD�
�=�1�&��(���[ �x�g�)9���z�mؘf��ø�唈j6.��N���nq5 O�`�n ��q�R'�Rv"a6_���^�b��۽~�lF9��SL���w��lޕ1i��)��q���)�� ����k�
�����(±�Dj�����`'BV[%�%#�۳���k��_7G�`�)��ő��}'w<�O����6����(�^�F<ɿ1�$�U�}���S�~u>d�կ�H1*�wc��y�=qx���j.������g��X�ev���+�R�,&��Q��x���KQ�[�-�;0t�R�/D��b�6g�U��^��͚�iM�dy��oz�m�Od�W�y�i�����u+0�?�Mu����H?�d0��K��9����y��"1TǞʂy�yτZ`Z��wR]��wu�!-�Kפ�	S����L!��u���<��;�{ʗ�>mZ<b���fQ\�]0U��z���i6�mڲ��q�W�����������!m+eHr6�=��h����P�h�o:v�A�'�5��|��"m�[���[tp�J%}(�u*(q	�s\|��bK��v���l�C$1�/�qq1F������ɓ�����hů�$>�d�[�P4�r��T2O{@�g")�C��e�J&�I�K_�J�����6Ia�)32XC��q)�O5.s�t:���
 ��&�a�bm��>��<��&�w6�8�K�/�-a�j�/5*�Upf���ܬ��Ǔ
e�a����pc]��PPz��</��`e��Y=86��-bmk�j��ot���ET�Ѡzt}0o����
2=�x3�o�����+�(�i�`�X�#�If��7�?�tbQ�-��a�� ќ:5�'Ͳ����FyF#���l��vɦ���K����P�$�W^�1���e�J�m�VK������-��[)����>��js}�Jȭ�t5����F�� I�4�+���_\�X�d�`�!/��u��q�__g[uBr(���ӿ��q�Ί����4ʀ .q�Sz��ݯ[3�����C�w<�*}n�*��;1��q���qџ%�u�J��eVT��z	m����{����EI{���!�wx�>���C|;��-�,S�F��9J���;�8�V˗��0��'����/4Z��	����b��&�?KFp�����ӎ���KE�Hk_j=���B:�דn��(q2�F�t��
3~[�f(�9��/A�i<iJS�R�f�u9�^��w,��������=�S�8�>�5��ɶ���ʚ��we��	���w��>� 
/	�cջ:"�#��5��WZ S��� ��v]WBf�Ȁ���80�ǔ�R��*�E�C��R���b�~ɵP����Үws(�\��q �d�N&Vj��V�{S;P���|%A��Q�=�@�� 7��F� �o2wI!�
NV��)��/���D��`D$����.� F�<�w
�sc�иs�9q�%|:��D�̤��P��,U�%����0Va�@v"������r��2C;��:ni]5u�8!n�VM9\�l�K(f�?	�q��&dw+��S�a���N�)�� �O^�{��F5�[H��;��RX}��iζ����� Ĳ�%=f��Q�Dq������ԫ˒_�m�So+s#g�S*xe��!��l)7��:'a��ۍ��M�t�����'o���&"F�*q*'�頨:��q�Ӝ��G�ANq�1v����]�T�1��8י�n4��a���[Sط�P�ߘ�˒3&.A|Gu��2�]Wa�Ñ_$8�716:=w�3#�ƀ>K+�ʮ����VN�p;"�N ���J�Jme���2[�K��0R�{v�w�'�I����0���ش����*��>��b:9a���Ҽ�qN�(8����2�f��|ub��o�R����� ���Z�DYFm}�d@�}���4�A��X�O}w���b� �_A66l�1�1"�����);�������k�9V�䃫K��F�PA/�Y~�n�FK�H-�Lh6�%�
I����w�'rG����6!�d[�F^������?� �U��_r��[9�B��x^�R��N�@l��h��O��.[�)�F'��.���;����a/D>AJ����a��ϴ�] �{��H,��*)Jf���/;Z]]��y��:oJ-�xݜ.q�Vt�k[������¹��2��C���0d�����<�m	�4Gi��c:��oN[��%k���ب����NE��,n�@v5����o��X,�j/�A���F(s5��57��{\b	�<2t�e
ɵfO���¶�������pD��ц���Y"�q�¬,jħ�Ϟ�{�1��g���n�(��v;!܏:iٮ�.	E�n����Ob,j�R=����y����q��K|���@W��Ʊ����t�����&��H�X�(d��������u�łnm�W��K�+��4�	4,THV����}%�U��$y0��X/�)��T/ _
1���dq�)K�f�K� �qm�g�H9Rb�n��(C��C\t�X"��!���a�~��������i�d��jrM{�51����kӿ�p:��5!���}�>;Ք���R�:Yx����m�Ԟ�&�a(D���j�N�u�{�x��%�qni��bL�GU~��.=N7�A�'����V�Ğ�.7�0�2,���z�3�� 3�I��3w�S[��A�ݱM�λJg�ŲR�,-�*�d����35x;s�1���J�/ڵh8*����'�"��4�5�Ex���%Z;�����?lT��g���Լ�:�#�J�������p>lz<�aa�D|�E����r~�֭����أ�>%�P?�,�M�~W��8�J��m�T}aQg��]_$�� jXc
�`��L� W0����H�k�dL��Z�C��q�1�K�d+өS�c�g+"a������`O4F�D�,6�~���wf�E%Ov��+��$�Fx_��d8����nxe&3�![��%њ"����%��eft��<���v#��^�F܆�볛��"����QS���m���B���EMe>�2%8�	�C��E���m��ݞ�aeb�z�KFRڞNfI[�lt�~��ڟ�p�I�7P`m�$�~FY&�z�N�h$��2/i1`�w���n��x)A`�(9�Xa��_�s��}5����zQ*��$�݉u��.
J�n��4�S�%�͋O��Ҍ���A˖`�U.z�O���qi͏���èB��A�N�26�k�
�z&�TFO�s�-�5k�_g�[�ȸ��u/�jЬ�3�>{@f?�"p�J�d��S����H��!�%��j��:0���UD�k�����}+���}���0��,7C�/ZuӃ ���a�k �#�����.�~���w�f�Ds4W��2C���l���E �9�нnQ���50}ϟ��b(ފ�Ν}OĎa��wrm�h슖�dq�Ecюb�xS�ĜS������(�Xu{K3��}�pf �b�묔��f�;k*@&�����<�9%��(ٙ��rϝ���_�+�eڙ�AX����<eۋi�D]���薾RT2�3Z�(|������LI�X�gi����]>��$p�U���2f��Օ���gۭ��y�TǄH6z�5�FP<��C��[.�j7G8н?*Kh�`����I�&.y[��T��*9�Cϵ�����E/�!�V|V`l�1۫o���#�C�����AC���P����["^�q�AҔ�a��m)8t���~���L�e\z}ƲN�0t���������P��j�e�黷:IY���4�~�oSM�������Mma��C�R���W���;��9��~;���r��Lw4';ߢ*�R4Hky������q
�.?��i�1��p�ף�f1t���$�$���%��dV�.����/��D�9�?�����:�u���5�(;�$��`|����~v������mC���40�NU��/5��V�"n�8��\����wa��@N!�
@�j�m;�.�&��B�ph�g������K�7�y�0�m��bN"����z�@*=M#����'?��^^��ȱ�>5��(�+�.���&�@չ���1����hv9��nw+�@b�r5�R���r�<:��AT�()Yv5T� ��@��!����9�ΛFf̑n�%ƴu������f������_�Z[�3�ױU`)rz{�gi#B���F+�Mģf�E15[����E�~.���ګ�e���h�G���i,z#�7-z`(1���~�\�)�B6������V����"՜Av��RZ������-w��	��y�xx�P��{櫮��g���ax��^������ˮ\/�йw5���{{4O��G��{!x:�cI��XpP�˃�?sׇJI�Hf7;�e&�L�q��ߺ��{M� ��
��~��@�y7��e��O׷��w��|NC7��l�#�O�<Yr	��s�������9�d�E��ځ����ݠr���p��}S�H~���UkXF�E3�/[a��6��EB ��qCn�N���9��D�[�q�������!�j]]�7�Ѹ#eS�Xd˩��w�q��%;W�F�(�2���	���SP�������5C�<�{�������+W9��^+�G��!׉��Ibp� �7�{T���\#��g�.�z�w>�(��(5�;M�����#�D@�1��[�,�B�.�`�|<�!�If>=���.I�OBu ��� �Am��?��a�?B�<���:4���ZjVr\��B2�lIr�.�Ҍp����D���E��j��������a1*$�l ����W��D�U|b��/�V�[[2���սGFݤ�c�bPs�Z�씢PR�{3>���Ԍ�xSl�k��%f���W�gU��,�,5j`��]�	G��0N�?[�r'(��DZ��*�<	�핌�����-�\����cx��鶑ƥbA��I��E$N�duYX�a>�Ms���x��4���`x�2�̵,l�\�L�F���oNv)5���jb�h]K��T7w6���`'Ȋ�]�!�5dA=����AWNy�ʜV��;�cQ�eU�&�GO�3�}&{�J���eMD/ػK�Tg��f�����c���Ƹ�����������=x���D��D��x$�8!T��{g� ��.GA�kc�����W�Ir��Q�$��)��I<�kD���s�.�>�����J�������m��w�l��?��Sl��l������kg�$�BF5Ԛ��==6�B"U�ȃ�7K�ͻhqt><Q��D�j�_�엖�I}����C�,p-����6>Z��� �[ˈ%		��s/6�7��;�������~z���<����[���ڙ��p�Ȱ����^j�u5J4��.O�J��̍��%B]m��Qdz����{sh�͉!�	�裞�H0Mz �K5}�x�J5,Ǘ���s�K���ڄu_��%t�SK�ϒ�id��=�:l"(���2J��hU�.��-����
m�//���{��]#<��~�y$ȅ	zE��f;��>�vb_��˿�ۼ뎙�!ɷ-���)�!dŗudW������z�-���c"$��S3�8�������+ҩ��*S�E��P$�MGA�N�r���(�ab��E`�����a3����&���f�G:B`x�5h'@�m���]���6u���Y6�iǚ�E�[Uy=�&*�>��k����]�"p�r�M�G�͟����"�,�]_Zɋ��uC�0���ܙŎ(t3��В��{�9��?[����N��Ƙ�/P�f�_"��J&T�x?�Ҳ�~٪��5L��Ә���"�Bm�}�� �6�������=u�v�N/"��6_G����FV.̱W=�-X"B��LD���ݺx�<,l�x0�:�=?ݽnKU*ٲ�̱ ;ߝ��e�ke;�-`�@ʱg�q`��6��K��7��5�CZPTѾ�F�A���]����H�[������5�����W��"aOz3� �c���!b�,�^��:a5��J���}EJQ/JPH29_8F�d2���]�ݟ���&8D���0�'���[w���=��B��=����n�N"�Ҳ���Oe��1�˾nh��œoxI\��;���L���V�t��䅩=�+ą��ml	�U�=��B̛TX���;_E�Q����q6{�E6���xG������{��cb�H��ޏ�Gd�&���*�_=u�WAr��#E�B%�������I}`�u��P�|؎�b�(l�=��]}GmF@�E6_r�I�*�(�kc��C�y�X��{{��2����<��4�(W[���B0">.aH�F���wL��l�埔�V_�C��8�k�OA�4����'6 N��ͅ�OJ�-"1�SN(�r�I
]-̔�K��62f����{A4q��y<�b�����B1P$êŞI��z�,��)\��tc��	�}j��N��򂆯���>�D� ������I�_�\/T_E�Cx�#�^���O��)lRmf� �,蛱k��>4��d���w�ϋ��A�a�\KmNJ��f7�xaȼ���?G���Am���W�ԉ5 �W6t������K�;i���>9響���9x�:���	p��B�G)gm=�o�h F� =��6`REPK$��[��C/og�����P�����*�򐎕�Y�恊c��Lo� \�V�)x�����L,�Y)�~(���كh'��-��k!�������R�IC��fg6��4$��_�+fᜪe�?�/k��ϭ�1�+AR��섲�Hæ����:0%�����al���[+ ��s��9���C.�tgW<7*�,��r'?F���Q�bR]'���ΐ�KJF�g9J�,毣̅Q:�uB��q]D��_C��٬cĻc����ꝕ8��H^�����4�Ի�O-Z"w�d��v���f4�� b��8�H�0�{g��z����!�W�tP�?=�.��e�ҟ:�J��S��yw�C>���_@���B�T��_�C�]����|G(���C�-��L������s_P�[S9&��M�R k[�)���g~��*	B��x�[��ģ�,5|��z+�#SSI��F5��G�Ҷ�V�gʢ�kA���<���Y;ٮ���F�P��r������y��R	�z���>�i�AX�\�����f��6���b���3��vHP?\h��S����zo=uGUK�<P�h:N�7�p�^�g�O�gS�<�l,�#5�\:�U���ll��"A>:n����Ϟ��#����`@s�t	�'Z�N���?ƃ��=P���1q:�:�:(,�N�λ�����6�(;>V{e2d�l��V�^�${�ݜp�5}��.aêCy��F�Gx����ֲ���9V\O	�Z�Kl�
M ��~K����]�qQR�|G�r�f׳���-
Q?ڧn��N�U�4�k\�Y|�+G���U,���p}A�xL]yûs_�Y&x&TL4jd����M0HX|�I�~=�]�I��}�#��&�H�U��W~�'�;H~r������3f�\�ּ���5�3����	�����6�']��d�.�_����^z����A���Nj~44ŉ���Ehm�`����:�����&T"�F'7������R3�`
|U��� �����u�ڪ�c�D0mPQ�+M��L#~��L�^�.6t4����2v��ėف!�*E��b�[c}��۝��8�|�P5�M�J`Xf��W�a֏9{@r��iK���S*N���S����V{{�Ŭh�c�T�k�]�����|H����N(�TG&�����M����h�S�H�v��IpJ$K�M�%Ǭ@S�ԺTy��d�r�&����J��Aʀbda���
rP��)Ҫt�*�XӪ��_:���K	��k��(���O刦]����گ���8��)��6��K��Ҽ�9���#R59c�F�@W�ڢ��W:�A��Tޟj����B�٬�xN��eD5|:W�vc�v�E���a�\GRS�]o����F�51��pPy,`�s}h��X(X����G�ڿ@*��^ }=�ž�]	���b�k�z~�'�}eܬK�s��������IF�Fc�~K�g{���EH
�W��*5BF=����z����u�;>@ �{;��I*�
,��fZ���T�0f[v��H�L�(���c�~�V���K�O�'�N�D��Ué���2k
�LG�ة�e�����v�5���E�TE?	6>Ȱ��;t�|����8f�_��t�[
�Fxa�|!�w{_�6( �p(�P�� �si���9
�;''s���E�`f��u'�5�äȵ���N%�qણ�\_�zIOVP��CS�{�O���JJ�u�JL-�p����(W��Х�bb:��F�[�)C���s��� s��zĖ����g,�kX.
�G�!A ��G|��7u�*Q���#H�'�q^�:̈�-���ڵ �s���n}�Ql͆r�R�x��#�4:���c����V]U=!f5��x��}������~����ӽFW:�{R�.�ۮ�S �LC��5��)"4�@�*��n���l
�4نi`�7��x�n*�98=GNfL�����O���IT�/��4%t�~�Yl�9���3�P����@�#!���,-���@��k�@O|7���F)�F���h��p
����nF�Y�M�]�hf�lO��
[2R�Z~��F~�X�����5R��;��9�1BR���ri��;�ˊ���*���������)�	^�z����:��(?i!$�#b�]s�}bf���5mt�a;�מA�]w,�zږd[�{�uA8S�1��4�A�NZV��%�:���#�u��C�X�R���$?o�:B��
 �%�th<M��	���~��0�!��w�����,����|FX��E�~k5���;�-H�FL��@W���1��`M�5����m�������{�G ��ߣ[0��S5�xGJ��`�]�.�V��R~d�k7R�(���W��z�ʶ�A�A���l�T�ܳ�5�/�>6������ӛ�Bj?X�6Ȥ}.�
_f	W����>�xd���=��b��s�>PW��뙛��s�1��"ٺ�17 �*$y�D*���ʰq*�pj$t��k]Z}*��T�*U?������J�����]�K�0q����)�����s#�I�!X`v�5����Q9�ǜx�)Q�]{7�U\��wT㡤F���y��2?�Ͷ�i�^��g��v�*�\�1a|�&v���o��WV���x�E>'��� ����a�5��!@�����9!ZU��E�JT�J_�[�"-~S����#�*<����Am>����<#�է��Q}�=`����{��'T%���~�������R���2�G�Nk��G��eºx݆}/�s|�Q���Tp[G~���џJˍmN�M�ҕ�Rg�����_r�v�(�v���bN��9=;�.�:�_��
pT&J��`��E����  �	>�q]�p}/�t��;u��i�4J9����mQ�Q����ն���?���R�b<n��:N�?D�i���k�:hLS���n0��5��÷.BG����љNc�o�;v6�\[� �ߺ0<�=d �KG15,.Wg��;��]�gs��8�T����;>z2{�Ԋ�`�7@�6�����AU��!����s�{��rW��Tk'j��C�*V�3	���(Bs�W�[-��g'��kžn5���!�TP�A����N����t�\��
���{hз��{���&���?&�㿋�<��G�6��)��6�����������7�:��"�Zq#_9c���	+�pxLhQ�|7ݣ1[X����p��Q�j�1P^{1�{�5�&�3��ن�rx�(��m�M�d�ǑnX}���o���߳��ú0���A�����(!�I������qI�l�:rT����ٝ'�m92f��~}[�w��>qMY���M�Z�MP�Fn�p��f�O��a��~��p�L?V�����&��?b�zf7�A<�xM�����v���	��L�vg��v����S��n�t�K�<&r.��Oy?���*�A2ߤe��5�HY� e��'�ǵ��z������媱��hE���o�پ����#��m���@�j�����R�(��^� g�7�R�#������`WՆ����Bt�0B̌�5����ͬ��C�s����Y~j�DK�% J��ڴ'/�!�}�Foj4��o�R��i��#C�&��L\g�ێ�ƾT�>�E��r�MQ�_A�>SA- `�3�_�zy!48?_v'�")6�,k� �@	-N<xucd�!y_-r/,ԃ%�2L�9�UѨd����Wg�6҈W�͛��;�_,��'�߹s$Dwo%����2+�DF��N8"�t�n�t*!�Bc�N	:u(���|��S���M�����V1F��D�����5��s70��"�C�;B�	�3P2�R��[���|�+H�'����2K3��}�	�19K�Ӎ�U�^�5�i7�P��2�G �!͌2һ���w�b/DC������!w�sJ�Y(���X���51�[������|�f`5���p�� C{�O���R�SX;�)+X(~��(-�&}�Q�'1�X�ϓ��֙�"��\n�]���F����҉}�#�[����	����
a�.��s���L�y��|��Z��դ��J�������1�LT.�: �����Vx���(p�*{���aq&�]��o��*U���db�&���#�U���v��_��6Ҥ[v��4�	O����1i,󡕸k�8���bH)x~}Ņ� Xp9� 45�nN�݇��6U���W� �Q�����T?y�����J��'>���{�r?7zfY��E6Gä����E��G��ez��[��V��d&ϐp�UY�F����ޤ4��u,�w����w1�t�{��u7�oLVŉW��N.3��fw��/9�&����H2/���[����g0ڝ��]�������<�R��Ӕ*�<���b�@4���AR��w��0Z[J^�w��D��P�s��O2Pnƨk�6o���G`�Q����w=�#0�<��D	�������p�c$�T`Ҥq��=�ρꟕ��
��b� �@��-04PP���V˙f�z쵬���H2�@�jX'�H0s"�j|�d�)-�hwG*{�^Pkcr2�)���1H�.1W6|j�ϙ�����D��rE�"��>&�x}��z��5P�����p���U�"������4P�3�?T}���G�O�(�����V=�xq@3�OD�5� ^M��e��7�����A����X�>J���X^7>��5f��I"��[PW�h�[%��%�r�.��]�޷y>�0n�exq 6O�D?b��*�.��g�#� ��������������3"��C���=�gSr�v+�i�����˗�� �#8^�ۨ}����]`����7ԶP��[M��c�12���3@�eh�q�B��rv�.zOs�,cD�C�'v�o;���K�/�lK����c�G{��zP�m�<�a�b�I^0��΍�PM��r�So �����G����d�+4:�Bi�I�|,\qF����M�a��{��ˠ
�]&��]�R�R'	(Ky�c�M�mL������Z��U�$���wvM�zz���eiLDmyg���T!k8�n�;�[�^�"y��N��$�]�]���\y���$�,Zf�+��oxB���n-(=N�����C�0����qzbx��jkB/+7c]����Fxr+��W������h���xq���C�ӳP��N{3[-U�ً����P��� t+�b�Q�M)鋳b��t��	�=�J���Q������e�{-��8��>��Y��K�����"v��ԍ'�+��C�\?�<=�@�Ʈi���e��jYTbl)��E�GǓ�v�����2�P��}��1� [�5G���b9�t�&;#.���W�˓xv�y�̿5����l̔�1C(Z#k}0`%��w�MW!�4?s�EK������,��x���^�?T&t,k֗��7R�~t���]�� r�7s���fg�ǰ�<}�!b���ft?���;^�c�fԬ4�v��b���Bf�Лl+q��id ~��D՞f�?{d��Y�&���C�m�&h�e#j���1�g���No�����x�`I'M[��6����L&�i%�T8FU}�8���67Q��$m"�v����̦��h�V����_�Uͼfs���w`��īTKOӘ,�#�N�J��ӎ,W,,�H_��s��a#ռ�wBh�9�j�Ă%��@�%�VJ���b́"���I����� ��rH���������d������H7\de�O��e���=��qk.��j/DŎ����y��CSO��!/�#~4�@:��lЯ(00� d�n�8�X��F/aP��*��sm�%vE�k���z�p�'�E�<�8Jjw�p�:���i|3�A��J�Q�]mMZzʯ�E�;n"<�;"#�n�<#�p�iY��9����"����ͣ����n,B���u����@^A�H��xM�I$����J���2|��ЌjzT�����@���&�T�U=�����VՃ�p��F(�zP�M*�-���cT��ߍ��@�p���ξ���ԋ%��	�e�\�VDJ�\�+J�:��0�(2귔�?����	��T�xB�U\�g�	������v�p�؏��ňP�2�@��ke��>��[�҅�I��T@4Ն �S%ʦ��(�{�w���o(ݬ��+��Y҉wn��X�J��{54`�.�;�,K�r�|�T#�H��}�2�Z�p�gO�5ػ����h��;�U�/y�th��ZiO�ż6��3�	�D(������_j�W"L{�6�;e��i+�A�u+��{��1c�iV�&mL�K�^��Ӳoc�ں��:���p,�C㸺��{,�����x�F$k�ö���6��s��Qv�9梑fs!�ӄ�W� %e��Ɲ�&�<����'X�X�s�j&��y&�%C^��3H�S7".Z�q($�?�D7l�i2Fw��8�0�&����ݷ����(�,F�T^�1ɀ0��;E�����ڙ�AKo��\��Ǽ|��y"���I���b��lwmg�(�@?�ϙb��"c��{�CJm�qO����R�]�(�Xt��z��S��lW��?j	���K�N�D��Џ9EV���6�\�)R-�?{�޺��t��O�-D��ȵG"U=��N�s��WB �s0i^Ф��M�q+�=/�n�C�]a=I�q�3W7��:E��?���y*�Ҡ�w�Yy2D��V�3�w��o��1�s���hp����4>�b�f��G��IZ&�%t��.t*b��!�8f\@����U��yǈgv6c�0@~ȶ��0�*͝W���ؖ��)����ֶT��� S��k�_�A���;߼ ���p�9
��jD�pTdg�Ԧ�]��'�[�_�ݿZ#��p��(�2J���!J�Y|r���݄���-�{��'m�g���|f��?�I���E��k�F�	I�a���I�ɲ0،t$8��U:��<��e,�ˢ)�x*.��ϙ��5Ѧ4l�?�,���q�P�+dOW�K)Y��>�|}Dj@�^8�_@b�|�ot@��c2�;g��B"]�&o�����-�ۀ�W��Xr�
�e�[ׄP�c�6T�E~Y��'���U׵��q�i�%�p�R<�49~ayO�X �0��6W���]�T2ZG�� M�t9G!gjY����0Woح�X���
����G	��U5��t���|�� �nb�8�Y
���ÅN�B����%�+���aVlĩ�_��\R&뉚���M6PK�<�R$��X'�YR�����9Ǒ&X���C'�b���@��q>���> �x�k|(����Sk@��e��P��<��_�{�B*ky��5L�s���i�ag�k���o@~��q�i#�#}�}�H��_�y��jD�#L�\^���F:3#��4)��ի1���5���Rl���X.��Te>w��C���^�H���F��lQ�X�����߅�w��e�򉠚�+Sx��#�z�/w��D'�7�A�쮞n�m$� _$YSqC�<ʖj�6��qN9c�Z��v3j����O���M�W��-=�6�R���7��L�;�%�	 2����6M�v�C�8xU�#�:��E�ǝ3	�[8.x�i�����R3���+�f�����M���؝�*�r�`+��d	A�2��-�s|�ӞKn3@�,�c幤1wY�oE�و�&P�?�9�'�ze�,z{y�@���37���NRG�4F��d�|'���T�+�--j�W؀�ui��������ڙ�^J=��r���u;`6NkCG���(m��U-�6l|������v�s4J(Nlk�)o�=5P����:���F���,�d�"�n<c_NG���(��`a|o��D�wH� �l$Nzaz��@����[�ڤ7(�i:��]2m��<�AkO��,�B_L���+<����Ӿǁ��@6�{2=�K0��N�w��N� 7�o��oy9�-p��߲z�� @��I��W��.W� $%47�e��E"nS�V�?�Ǉ��|����JqR��4U%��?��B� ����&Px���T��T\�6�Ϲ
Tϔ�&:����H/a�
MyA��+��2��{a�~��2�0�Ѩ������1�����̠*C�4��l̒,�����p���Ѯ�ֳ<۸�����i�8B+�����S�!YϠ����* ���I����B#���%`o�q�����-#���:2?�'+.�:�'55�6�A�T���+��4��x���ĦS�L'�W��͐�Տ���H�0�+�����"�_�Ȇ�T9(%%)�x2y�j������N��G�!#-�bP���=�R����:4��>W]w˧ �b�Vb�����t�����d������ɹ�U��	PS�L���P�2�k �j!���a�J�`��4��_fmڦ�s˙�!/������_I(�=����)"q�5�'�l4��V� ��o��}P���\�I�`.�
P)�娎�R�G~ݺ������?逿-��z��,t7u���.��Ed�v����2����O�����굑�-�Dgb����H�w��Ƶ����'���ԔZI��v0td�<PZV��n	�������Q�Y����2q�+�������xI��6�SX����W�u�����s�pi���:�Eh�]�y�X����T�ۓ��\?�eQ��S�O���yW�3E�K�U�,�� �}�u�!ZЃ�3 Ē|�O�l�}�`���.��\�]�*ͨ���-#��v�%�c�A�~��7�GZ�7_~9���{��rP��Ӟ����Âs�uT�o�)~⑸��<�����P�h�ڬ�J����<֓80<X��m�@�y-�������#�qƌ'�1�b�>���ݨY(�@
6�~��|��P�j�df@�JRW��\�ڐWJ>.��:B�۳/���sډ:�_Q�o�R�Y�_���z\�C���S7BT=}�(BEcD�6���J�����=�v��w-�|Q�*DL�P�>Y�R��Th��҄��D�D�/�sT�[1���1#F�_�_�2�S��-V�1 �_�3�J���m*�O��RE���Mc躢[�<iu[*c0��)+�̹��^h��
9�D��Iz������M���4BL�#���Il�?y4�l�"�p��J��)u�F������'�8IC&(w^�ڽ���*3f���o㼴[&�3�p��wV���u�W�qYd����h�]d��f�m5���쨧���m�1��աy�f���g�	{f{�� :���Y��"@�Ҟ`���3&$��ʞZb��.$��hι����a����+�7c[������2'���sdM�j�;��	�@m��PGP�:�H����.#W������H���?�êؔ�E��Z{6 �/|�S��
������PE���3�}s��d9��-5Ec��S[�7a�!8���d���M�,�kT󨲿�N	�$�/��C��ܹ��Qn�����|*�(he��SF�}�1��rI�T�>�p�k,ܾ�Z�gZ�^y�r�u��<������ǚ�m�fv�;�����р�
b�,�J�ԧ��e���}�#�)W�x\j�AO4f���j���/M�P��l��ֽ�Ϙ�5�����#�k�rִ��MOe�O�[/,'�W���.����sCG�P!�u�����$�Ed߯Y\�[;j��0Qam�F��Ő�k�8�!3�e��;+6���Z��ފ�A������T��S����֝;.Jm@�,rI<i�Y�Z"#�tv�)�/���f��ꖫ���^1�<4������$��6v�k�ɻ�DD��'[lIi�}�4�	�������ZG үY�\M��ᏹ�D�����ퟸʱOX0Dr��:Zu*=�V���*Wₒ��Z�@��{�����ӧ�A*'��_HR c��*R�6B(P(g�pe���� �Ǚ�t�h`��&�>/"5p�b���UI��/��c,�e=�v���ϲ��/�\�hl\ތR�����sSrrܲ�j]@:��K��9�%�O��<m4 �ίm��(�ZcK��Vd�7�쇮�H���G�7�$~f}�.3��3�
��l9~�Zp4h���l ��b�/WPE���2J�+W	�8� 
М�KG�ޝr'�K�WkCO��ڄ�,լm�@����D��g\�Ϫ���&��0IJ**|ع��bOr/����sr�	���C8M+X�i�c� �*g�(����T򾮥��΁+ߩՒt~��~�TK�0�tے'#�����D�v������X�" �p���PO��R��>a.�U%mdrU͌�{C��I(�0��D���D�%��NR�#��}5����B�WŸ����G�U�dT��G�K9a���G��/��� ux����}K�=s��q:~�؃�EnX��fkd�u�DU#v�V{S��k�6ĽR��ZJ����w�������m���~�]E0nb�7�!fr�1� �Ow���wC�ᩣ6�$���j���f�,��;�Gd������Y�!��g�=t)�E
"��*�>��Y�j�|Q���J�uG+?3��^� �g1���6�Z�-m.$�������Y�D��� �Iz�G�I->���Jۤ\M~^�.�ߠjX����]H���s�Nx��, {6���8r���3�ip���YǓ5�?���D��5tD����o��F��������zM(ՁAd-
�%�P�Nж*�P}��U�>�f)��558��*�	x���-85�8LSD(�^�X�~��Z�1�g��)���GE��y�j�ziL܍����%�v��Н]�`m�6�w�֣�v+��vD�
�Z#�Y�T�:�z�
�Η�</Ǎ��N,�y�ziV7���*�Vn�0kb����̚`�����Y��^#����m�x��#�,\�3��)~�*m���}����S��HR��ԣ��0r��86,@p��_��Ƅ��f�9�q�L���ׯ�b?nfC%@��w��Mv-x?<ﳖ+Xc��C�6�%�,���OCc��G����ߦn&}~
����q�/3,:���C��U����!8�!�.D�D��$�p21�Sg��aN�m;"D�E~h��m���1�
) �y�݀�0�����n��-��ٹ]���{��!9�6�T�Ԙ�@��ӄ�.Y����ż� �I�m��t.绠���F�|�բ҉ �����8��ꃮ���X@quҍ8`A�X)a=��0��
�%��|5�!k+���4v%��	��[1x�=�Ani����7��"L�t�&zdFAf��������~իS�S��;I�����w�2j��� V���S)%�ܨq����Y���	�*��4��MaS�W捵��q΃�L"��v��wl�����A;�w��=p��uJ7�6s|=b�P�XZ����v���V����Z�ތ`\�E��D�a����/������퀮]�\��.Ǿ��W���U�j���z8���s���z�;�@w<{ז���Z��9���Z�ak*Z�S�D��R����R�d�ɟ��D����i ��������:�5�~���y�{3�	��{��zq�BI�(sXa��V�X�7�ϴ���1N��~>%������4>2��hK�$ۂ�5ۖ�^����k�1ɯC֕X��Q{���K��y���
Ӻ��:�S4�v�VZ=�D͹�j��}�E�Ӓ6��,�.ȅ���p��po�r�hh�½%�bt�����{A���RH�#)LJw����o$Z������n�Y�v".W9�)i
�S~Lz^]���ɨl𖜄�^������*'�����y��g��<K�a�ԧ������Ŗ̉R��o]ȸ!��=�m�|�]OI\�-�U��K'�����f~ �uByE����?_�2�d�D�ƣ��6��rqrvƃ���$�$W@�-De6!lW�3�a ��#s��z-�s�s�ļY��'�Zb!��b�al2i���>Cx���@�#� �I ��XV�0�f�im�" /{sk]��"[��x��]D�c��$���o���VL�{r�7��{�Sʰ��c#젫a-��_��]��?��=�	�e���4=|�n2=j�쳚82i+���H�쵽�=�x���5�0(����cg������G�}�j�[���$�0D��9Goú��q
)q�Xj ���y���c�.�/�61d��y�3�;ʬB�)��Kb�w��,�0�cE�>�<��{T{�8f.�/�̪�5�K`�A�1G٧[Xi\t�����@)aUy�dE��Z�!��%fF?�J�)�Q��S��9:��� �\�in�!V�i�6������(7d#W�*ۛ�9��r���A��u���[������Y�.���Z-*�t[!%��>C|�0��O7�ٹD��z�c����(7����=�� 
6'��T��>%tF+��C.;IVgN5H��_���O'��rhg
��v�����E_|���9�ol���Ꙥa�l��[��|JxƠ�,52�E����-Ѥr�#�Y�ۂ��/m��x�H�1`6�-��ƋOIO����/���Q)�/�s�9�/�X�D~�\㉉h�JN��0���qmo_�94F�Q'�ր�w>;��N�[�P����������)_���dK�,�f]�N�^D�2��h��Υ�Ro~����1�ː�P����ݳ�f�-���r�\K`*;�}��j��]��o��+�~ T���%���ݞ�q�s�3��.u�$�'���9�����q-H����m��Gy3���ԋ�I�|9pӏ�G�2YЌu������zU��R�7�-��e,�#>D����7��X��,��sg1�����~�9yRn~���?l�.�&������a��u�,�60U６`5	�K�AI[�&-��D�� �ѱ�{L�R)��*	����'��J3��:�A㛢��9d9+w���NH<j-,NȮ�� 7GŞ9���X��g�`��6f��D��C��l�3j*X\�,� ���xn*ju�N�o����R7���tY_�&���oV7��&�\7������N��6 
�qk(vAk�k�]�Ka/���T��Z��|���ܶʜ��*����0�>`b�
V�6㼢��N�k/���ڻ�ʮ��j��In����	ͬ부]Ș�KB#��'�y�/C!V:X�[/��V�������͢CTY��Ͱ�	`�nV$_�`j�e��G�a�;E��9}B!Ԑ��z�ww�]+Td���|�Ͱ5�:���ᔰe�*B�!��	EJT�;8Zo�C�iV{������d�IV��:ѱ��	L8�ߊ�)�R`�A��İ��\֮�Gu7�$#��I�AMh&�y |ME��m��·1c��,�c|Lt�����_<=�yj|[�c�|C����;(�kP
dI�|1Le�p:K:��H���r�{�y�Nسͯ� s��ҩ[ߏ�yMAY�P�*�F���<����������K�(��q$�Esy*X�I�Vf�C���+��#�K���4��h�2��f��5��E�?�:l��d~���.�"<Q�4�ZV@sc�q�$�s��ijjie���ɲ2�m���hEnI���$�4��6X)%Q�A��wp��Hk� p߽��ɿ\2�*������� ~��z1�\�k=Rd@�0u����Ѷ��4��.�(�-�1�!?�Zӵv̙��K���2�뉅��ZS#c�)���G�����1�!�k�5g �F�%���u�{���_^\�:�F�o=�/Y�L1R����������$
ڗ�T�HtCoffB)/y��ݣ��>�V,�*�''U N�i��Ž��%�X5��
��ye����C>�s_�p|z��@IRRV[2gd�r�Ҍ���CM�R�%�{��M�z�:�����9�5��9�(�X�I����c���CS���Q�KOe6�cp�t�0Ǭ��yB2��_Z`j!y8�М�
k�ꙻ��:P��z�� �-�I���"E����o��pT�sȱ��<lR�A�$�ˠ�v���r�>�y� �c�V���x��5�������:�hp��������G�5�-�Bv)��Ώ���n���E�@��52��ƨ�)Jy&Cc`EkD�miMK]�1��`^�?g:��'�����y���8���ڤ���^)�#�2��D��>��.2�V/��u(����S�3�TD*Y���y/�}� èμz�k������o�Ȍ��R9Q�b7�z�E���%��.�=��"��;������sm�0�b�O��lه��>����~g~�Uq�..�ئ��)^M��7��R�i�,���BS��*]���͉�A���������Iɛ[Y�W/�߉�(S��}��3W�:^euZ?���
���u��y(�Q­ �4|��6�W F����s��� ����	����p��\M�l?��H��qT_UMz`��WϘ'�\ߐ����1�<��,���|���]��<W>Xǽ���?9v�-�;�9o�S����B��uj��v Uu����Np�!t><DQ�eo�DWMދ�VX�i��;���5�� V��M�ԉ�3�ǎ5��M�O���6�wNLk�Oo�7� $��X�]a[	���W��ƿ:�q�9����⅃C���В �qjv�q�j�ٵ]W[*cc�����Z*j�%�3���3K�}~���ڈ
��?v�d�k@�! �+P�����}�VyNAxZK�H5�8H�9�f]�T�-?�3+�5ӵi՝�oܣ�Ϯ�.�ն��B���q_ �Y���t�r���!��غ��G����܄C͓��(���o��_��-Q[��f�BHh��o>�]?i[��(F#Կ�7�?�t|�+�`�����z)(�	��HQ�-�
�w��nP�&��0r��x1�raI�Li��k�`i�:W�Q�r�yC���~"�^: Q�
C�?�`W2�[��,�+�~W�ͣ�]�Z�윛�g�����	�-��m#|ugWT[�P�aI�3��g��v�s%sE��X�d&P���V"�rvC<��6-�	 Z۲g�f+8���z:�Ω��*9����)2q�>�6s�1ǥB��9�wu�7�3<A٘J���Y�r�0k�&��n����a�c���~�t���\�v��н�Y��{�
$Xփ��=�s��&��쩮��Zs��o)��|��FZ��TĀPt�~���p�Y��C���n�z�]pb,����QgLۓ�ɟuk;u�Ĥ�FH��D�t�UuH׆\H�I�~�xQm
\b)3���r快��c��WY��Ou��h�G�j]����tE>⦲�jf��P�և]XV{�������Q�qջ��s��q��}w�v���Վ�z"�\��Hl�M���߈7'�x����� MI8.�UL-��ق~�PJ��c��o��'Һn z�Z"��R�<�n�BNR|�S���@SSH���9=���7DLu�5t���L%�\'���q��L8!��_z���?v`�;`,���wk��h��n[���Ź��ޡ'p��0M���	M��.Q9jm��h��T���VE7H�Q��u9�ީN����܍(�E� ��?�&μ[�0E��M|Ks�S6J�4�d�/4�[���Ua�`?p��پXP���w��_Z�p�����
���z~PΰzH C[l�'|օ�;pM�_���5����I�z��9���!%�Cը���,�Ir?��K�43?��Ը��!�4�b�3x��٦�X���$����B��l]�D��|�ȰѪ�)����YMʇ(��W{���zC*��lQtkH�rǆ�V�$��8��5'2�+��<7ڼ��?���f��R��k��Ixd�$�	�PZ�+фi��/u�:0:���'��Y>�E=�f8�M%[a ����1���L�n��چ��$�יO�#��wzM�"�#
����;�w@��Ke��
�K���@!�}��O����͑�au�K�o�6�4*�>���E$����
r���Lޏ:T1��#@zH5;�D�j�����7�h���po�s�	V_�؛����N�F#,8&��;˰���c�������kd�iH��1n��Z��� ҋ]��H��0�bVb;G���IHj_ʱ;T�w�R���O���,#�����mRSK�%C�� \~:zr�5��2rq���,Tϒ�)/�#���\�f��B�9��[�L��,c�%iG��]!���\Z�>d�h�}N�kQ�h�c��OsM�W��+Ж.י��?�Jō��>��f�1�b��R����;�DWu1\�o8���S�;��&\_��j�]@�Y�!	��-��K��!�)����輸��o�S�Oxa\��<ξ�q���%����
p����P��}�Ƒ;�Ы�V_��_��hPiѬu���T���v4���[pY������f}���K��f���y���\�LT=��Ql`ѻw:}�����W_Ƣ}�$�����)�Ӎ��7b�:��j��D�!13��X���b�Y�I��I6����(�5ՅB�[����k�����ZW�٪f�ob;�C<��R�-��7D�k$�㓐��-��1D6�ج���:��O��ZJ,Y��c��w@Bw�A�����]��(�ս*=%����v%��"g(Kiv�?����Z����.ř)�8}�y��au����� �k�[f�/�zէ.�/�3��X�:|�9M��x��nėz�w⼑�,l��k�<6{{x�x>fFO�;�o�Md�;�"��$ ;��0�;���I���h��QD����L'�S��"�t=g���"8�y�Ĵ�n8�Vu�V�K�l�
H/ڟ�]U RR#�F��r�\|�*���@���\�s��3�9�3�v%32�)S�'ǰ��
�`�%�����OW�@@Z?A��a��G�串��7x��V�Slg68��@ż7ޝ���Y(�=pA!���ɛG�oO��d�� �!b�.�)��S��������6�$�'y����r�D��۰CD1���п�ǫ/��������Q/�ш�E�\�2���D��}�7+R3M�Y0�/;� �E c>կgA=ӕ�sw��������R�RX��q�ul{=��Js�>Q,��/�����C��ee��c�zu�p�����>�)��0SI
�:�X����Ω�ݧ���G/'s�}��	��f�&2���'r�r��k��+~j=��G�No"=��w5-�g�Q*���+�Y51� �%��
I����$o�v��0�o�KZ�P�w�0 ���3m��[����@�<�9>��a�q��ob�F��X̋"Q�&s��I�oɚ\�"-n�d�+t�|�~� m�u\�I�^aW�xDyo�i�5!�S�d�(���Z�ѣ��ٗc݀�}�8���S8�;AW嫰�S�Go�@dQ�h�#����|�#�[x��Ȕw�V�� �1�nJ���|e����F�ɼ���͖���W�Wa���j��0��6�v�|M�WG=��پ�IC^�,��1���:�`L���cb��WZ«�Zs[O!�g�/EV�2�Y|?,ҟ`�%�C JIdm�f�E�#S�P)`"�?���� w�3��ޓ<����"��"C�@��߉r�o���� J�:9�^1��NG�Y>Ց9!��e���T|��ۑg���q�?Nt\+��g7^5����n)�[/�F{��;oA��I�Wc�fO�O�.-�R�a�/�mc�R�o�q͔��@� �?���0}h!Z��.�kŶ�W��G�s����d/[a�1r�F�
k,�ߨ,,�_��#7�� g?�]��������Mx�$�H;msn,J�̿}�q1�Ypa��ЍH^��	C	Hi�r���R�r�g�sV��+��(.oÕ��F�Оt�#���T�w��K���ԍu܎z����[���T�3� �ER8�� ��W��
��79�qx`4�7im�g*�.�m9����Ǣ��h����v͋2���k��g�z�CL�2�U�1�{��PvRyB��F��2�Ĺ�xz%.E�]$��Y���~v3E��ف�^w-i�n�e���B��|��gJ0��}�N�
=sdq-����/�&XK������S�+��zy���J(�Xſ��e��ųu�f����m��m�ը�����$�Ӯ����b��H��H���Q�Fn�{}R?��w*��e��5,��ҟ���ɩS�\S�ĉ��%����&�go�q ��� Z�>.�6����J�#� �k��!,w���П�rwCfjp.����%���i��mu\�Y˜�_�
c]��E��wn��"�5�g8a��]��z����5��=R��L�A�=�`tϲ�N��M؊?�d1�Y�x�5}c�I-)��1�[4�u�RAN�P�յ ژ+.y�$6y���O.��!/<'AHL�j8+!��jZn�zͧ�1~�t���XR.�˝dE�N)�j�wb{鑍{_��Jٸd��
8�L��Ǻ�p�4���`��s�e���6.��X��{��٢S�5~�iD�7���}�e���J�i�!70�:KT���7eK�ף�o�d(6O�l���3�i�c$��eu�?ʌ+}����T��-�)��ޜ�A�� �������3�i�����9JTBӟ�dV��C\s�\��eOg��G)�u���p�e��(��:�r�!g%� X� �%۔X������ل�:�!?.j�C=�f��R6��%��t�`��&�ͱoݮ�����.]���-�̓&Ski��~N���y��"������8++A�*j]+a��[lg�O�l�>�Ϛ&3$�T�8u�V�uU"�O��Z�;�M/m�����dr�}�������f�bʐL��{Ξ��_�>Rӥ	"?eM����V]̝�4r�ȕ0��\<Y|����j��j��҇F�Y���_<�^�������ts_���h,��#t�������=���3�F��ڽ��@���!�o��V������0(۰e�z݊�X}�"�&���]��DF@�zI;9hQ�߁�e�B��:�7AK�;��V���ǧq�p������<]A�`�[p�L6���S~��'�-��%+�(�#�-L�w�V(���� !�{KC�ՅZ�qsq���υ;?x�����|�m�a���aF)kk���(��z�M�-ڲ![��"ȇ~�����6{��/�b/j�V����;:���Z���g�?���B�&ȾDc!G�l4��i$ ���� Ξ v8�z��$.���}ڞGP�ӊ�6ܭ���ԟ�������79�=�%coAk]o��0�h�X�������^�Jo"qJ#�$m�GK�Q�dB�Z@f��36�{2��47�R���Q�r�]�耆e���ƚ	S/�a��3�!a%($����6Q���4�}�I�Y�	D8xE5lS*̐F�v�?�PI~l	{^�s�v�XL�-˿�n���|�R�d�EU.�5l��0x$:,­��PBo�O�Mj�0� :�E��=��R�Ny*����Ԙ�/K�F�{Ư�����!������Ɔ�՛���ٕ�5���=~�4�-e���,�!3��n��l����������<�o�䲄n��=_>�vŹ�8SQ���=��f%�拭B��$3��Ŏ[��{hC
@�%U~��OpX!W6�-?x�
��oR�O�Ԑ�"ỳ�o��Q���*�.g��c������S��9|�c���\���vh�b8���z�������^�4�Y������f�Nk9I�ɟc�Τ���	hz��bY�{���"U���ؼ�n$'�X���"\�z�<�8�Yg�|�_�`I8qq�큒���W�$��`1�JON!��74tca�����pS�!dJQ3�5�R*Z"L���R�oYMI�h4���N�)��:�k����O��*��x1���GMj��H7jc�Pg��t��^�n���hsة��r�~�ɓ󄽂�M����90���4���D����������>#:���2]]�4�S��r,��w��*"%��j�a��E'	*�#@K������E�]�J�e�j�X`J�����UN��i��t������!i��K��U_�L <�[\�`=�{n�����]�Zz��N�{3��Gr,^�љ��BU�u)_Dq�^0W&Lf`�X�[��R�N�%�ݹ��O6�~e���
��?C�����؃O_��"� wmC�C��ͳ6�=���Z���N�p'� Z�'~]k3&11֔ ���u�8V��B]��2>��m�qGb��SeO��S��~�6D'E]x����p�d_���%B+�5��>0���r5��)�x�?C�I�	��d�eA��:H�,��$�1[â�(o�/F��;�
���y��K���m<���.�]<C�����5ս��������6��U��?]>:J�f�(v�����PӤޔ`��XX�������FO3
"�Ip�<�z�"���!��gv ��x�ߺ8JzP}��@H@�k�\'���YT�t`�b�fϖ�gU=ӧx�����ӝ�D;h[���A~s8I�m�� ��:���)����@+x�oknH��)�UV�N��8а�;�hV����t�L�Ɛ�t;>���xyq#�o�M��y#}-�D×BJ�$����/=�UU��,d9a$X���eB�'"� b�i���� ƌ
�4�h4MBv�k�7��b����	xȫm�p��*��ف�y]�*`"��$<	��1TXL�*i���eP{�� ��]�j��d+���<uy�U�M����1y�څ ���-dG+��D5�Gj��W�!Ҍe7�A�~�w��Q�q�/be���rᨇж��s{�NU�n��?��_`9�M�aDY��y�R����/'~��(���������䑛����x��(ƀ�r������T��b=�e�#ZiC�ז<[��H��B��՗�V?��F�9����xB�҉GnC�.GE�B��@<�%sV�G�T\�K'�|�%��kH�&/Q�2�.���>¹(s�Ε�`G�6���r>7~�!}����}E%�氕e���>�Zg�h$m*�쾹@��m�e��D`�\֜� \��d3�����g�D��ޭ�N
s �#:�4QV��&���'�S�:Z�-��5=P}3�/����d98�T஥e(�^�}|k����	&�`U^��Č��:�3ͨ�h��"׊������l��.^���9�ʤ�	��P@v:ֿ/@.w�ء&�7!�>�E�C���+/�N�B)(Y��2�������M��QV���8.�뇶_���E��H�]^t����W�����Xxv���;�Xp,!���s��8��������.�wt�}x�n{v�ԕ��H�%�={�#W��"�k�|��kat������J�ٰW(W8�d�A0G�$�#	z+�NC�� C��������,C}��[�D�,��ю��*Ϭ	��K����Npm���V���ԅ,��FJ-�K!�fRp���k0.-���%��0P�P����5֓��� ��y�0Fw�ИM.0�KdI �?��nG�WX��ף��9a���i�:y�KŘ3��2*�����ց_'� J	ިN���W��B��v�ͳ[	6.��H�v�;B}�ճ#�������L�1�V����C�v���tP�����v�U�d^l�*����*���2�o���4�X�1���ĝ�T��k^3?;�Dv���y{�T��w鋨��vx�k�����琬_�U� Í�ɚ\�gv�}��7~Lks��z:��!��-���>���T��E([R �.�|�bG�a��'_�D4��j1L� �9�
Ԯל!t>�����n����3� �wͬ���K˳>fs��&8����#�]S1���۠H˘g��at���d?&0L_BszJD3h"���V�P�)�4O�o�.:;�l�n�`�W(*t�}����c���D\]tC/�7��9*�����Z&9$#�����c���Щ��G��|4/�h5{���Q�����w
�!6x;Mm�Z��t�;q]���Y����1�%±��!.��
�?txxJ֑�H�L�Q@�o6l��3Y�����D�2�|�y�s���r�u_V6n�Z<F��#�g��c�yzg�������n����z��X����.P��_��FkP�m��ք���������D0��isE�S:K�A��&�0%Jp���p�"/�0�O�#�)����w\cp�~Ix'����eC�<�-�����봣��}t���L���[3�\���a�%|���&Q(ѐ$U(�{/#����>w?/�d�
�hiMR�悱1��&y.F� ��=8ѿp��`��l�9.sPr3�t���⒅���'�;m��}Փy*�:Yӧ�9�D ep��`"��y����S�׏ژN�rv���;���85��:L	}v�q�+#�j�C�o��o�]��YB�ǳ���Z4�n=�a0�&7�|Zz& ����Z���A����pOr�B����j�E��Bl��8�,��6���������қ2ʫ��oj*)�ut�rJxcXu�@γ�8��F?��ZJ�����v:0Ʃ�N��Ԫ�/i0]? B��q�|�9T�P�w���8��+;6�R"�)(�|����:�$\�6�ϖP�|�{�&�_�7N��+GSi��^vH���:�}���`�-ᄳlD`��jDw���;ΠN*u��%葃@��YI�0Cx�� ��	�x�2���L�!Qn9	���1���|�OL�扛��S��_�|�}��	˷�S��q��-yu��BMl���]���k�x0F��."K�.ߴҮL��
R¯-ZW"U�+���p-.z�U�4ժHML�>J�n�Ϙ��*<If̮o[�h�n��>�'U��K�k���0^�k�I��`x��'��"��	W�_e,5�(XIc�ſJ7��\X�����6��(���+�H�3�jg2k�8��D�	T�p񯸮��Y�Fb����7�'/S�A�{�T���v<�>]m�1
�D�Mg��25�k�O��ʔ��=��-|t<bk�_W8[��X�wzl7��ZKT/sw6	{Qo�}K)�:����v�Vl�V�4�gtlP8�)x�7Ns��uPYJ�4�����D�F���V,�)�?gk��͕R ^�l�~�ٮ��|M��ˮ��kq0�0���TFt$V��z�p������d*�d(9��:HИFD:�7,����(��C�tچ�؀Ν�I�zm�� ����2���N�QYߐ�:1�R��.		`;���Q�m���V�Fm8C���̀$�[Ԗ~�w�i�Ǵyi���+���Ƀ� ���-�u(�`C��񋬞�b����?co��B��:�)�[.�Ճ��y��^��afbm��Ǒ��E&�3O��P�MT����4��|�Q�GA��x�4�s��o�3t�Hm����:� ��A9!d�X���,��3�Z�E�}����=���s[�(_�Q1$�*,U�������co���D�
�E�Cj�L�i��X�P0)F��{D�ģ�av�2Ek�(�p�dR��J�}���Z	M�V�4��6B�I6���<vy����Ë�GL3�w�u�@���:���Ӥ`����d�u��ku	�de�L�nȆ8�W���M�c�~gx׬]C��)2�pW��<)�W�R��+T�׳�Grf^��xjJze�w���j�QS ��I�>9����)�����驑�!�ї������1d�2�b�"?B�����.%'�g�a)�eh_?����h���`|
FS�!ۢ>����;2�_�*���Q��ۋc���}L�v�z����sB�S��z�*�c����n3j�',�<�D�8�GIF�8Sڒ�<{�كE�-LZt�D�c��]1��U�z�=�_V}�Y� ����:j�f����Y-�.�bv�žj~�>��()�C�b�'�L�j����Z͚ܼ�A�^����/:˒�RaAPtd]v�J��o#+U"�":MLgD�����-���c���s���[nh�.�2��>��l������%Z�b�f���H���!k4
\�k�#�}V�7��4!��o%́+�괘�\�1�&���^E��N�]�L����.+��i�a��Ή=>�3f�հ�jz3�ʞOт�4npZ��K�Sx�o6),�A�u�0�9��bG{#��ᯣ	����̎nR��#X�'%c�Z���{vt2��kȋ}���� 4o:HR���+x.�%4�)˸�Q���nZ~22)���Nk��w�h�iH�x���u �2q:����?C/10����j�R�e�۾)/ U�k�Qa�cq38P�+Ȝ}���� -@R̍+x,�L�>2��`o��]��+#�W���'^^mt�����\x��ɞ������lеy�U�W���G���鯙	Enɑ5�I甞H�zOE�$_ߵ@Ȏ����y����_��52fE?�E]!ps�d����%��*~�v1�Qb��s����al��W�.0�=���ʜ"�A�zɭ>���%>��v�6#�q���#/��14t �4s5g�'Z�Oq����H>K\�t���x0vp�<)4.<��ۆ��:�>�7*�<ExU
Ü��Ыi��C��f����f�_XA�����C q*߇c�w������~�*=>�����M O3#D�����V&Tא�R;�!��U��0i��$��a� �K��v,V��E>z-!w<d�����e�E�#��ĸ��.S� �㦳�޷��\[&II�?wfW� Wyգw������a�&���&�$��p\�b�f=�j�OF`�&ȕ}99�U��.cyP$���S�Q\y���/7�_��v����i���Q�B����T��[l���	����i��ΏA3���m4�<�w�|��+���R[u�sڦ�1�"��^Q�TZq˯��i����q�ƺ��,.b�[SR��jg@*&�R�!5��8��C�M�¯��h�"�ce�كoW���V#ˊh��[����wnQ>���]�@��U���L�%��"$��-��qJa4��PkW�����X�	ZQe��*�wxf;Ogf�9LJ?~��1բ�-�էH�)�E��!�~�1�s�ț������qX���>��ʧ�ʆ4��4�ȵ��	��+=f�?oD��$�*VY�Uս��{�^�L��닯�}���+̠	�������Р��(��;6�g�n��*�l_C��ѫ�lN�;��K4�ĔE{�S�^�����I��*�D-���w�ScU�j��D�:��6\:�Txl�=��=�g�Ք�!c3�$��4��`���K����,.�d�G����i���/s�e\Vt�]�zH�!�4�������6%��Cr'V�b�<\%��9����|!�����L�9��*��o����������7VDI�D�q�U�}�}�W���"�����IR��%s���%��@���E�m��?��B�	� ��Ɠ�Y�KLx��8اp�g�hjA�t�h��j�p�S��&���s�U���mX4y Y�i;b�,���<���L��"o]��� E57#�+�b�v���q߱�:O8�����R��o�tO����W]I%�6qT:����>V�[B�`Ð͏N)Q?5����2��$Zb�`�:S���vD�]����T)qh������&I��͇ש�� اũU���b�����'��"{�;\ʣr|Y� K`�<t�{̚y�!{_1���ck����5Ÿ�|�S�D<P�3����#i\�Y9���B�L�U;SK���h/$eL���9#w�@��A�}aR�c���h��O�L��W��O��j��E�i��)U�=�9iif���,4^jM�`��F�M�U���Ӛ�&twC�[�I5:*�)./TM
��UU�B�����P��"�(���r̷8P�xJ���ɰ�o J']�wk�xK[�y�٠~~��	�U����i<f��V�zLSP'L�.a�t��(�R�߬ޕ�}�5,���6:�yzP�׌��F�Q�i�[pD�Z� �B����w7�"�V> ZR;:](�'�}:��ѕN�	�aJaC�R���L���/D���A0�}��������#G��M���p�	vDu4X|���نk�b�ӐHE��ng��gDhaR��� x�)4��m,|��ǈ���p���M��a�]��I�3�g�3�`-���:(��"���k�Ǒ�9�
�h"ⴜX�r"`�����
e���L<���(��!�L���v?y�Y��M*e�r�M���S1b�G|�ٸ6q'p�T���C�rA�7X�&��)٣�ď~�������6>q�䧹+��fxXÐ�-�k�+?��F��B�����rZ��P�ˋ���a�-s���lF�{�\�J�f����Lb�d��|�J��e�~�-�J���'S�g>���E����:`;BW���%Yu��a��d{^�g+��peR���N�|���"�I��%*�Ac����{�?�8���G�����v�a{}T9�U�ѨF͗�h?"�b,�Jٶ"+L��w�d<k��2�+p�񻶑_͝�V��	�er[�!|+ݰ�!�]�E�"����g��ϛf�S���Ѵd��c�V�SǷH=0�U ^�7�.��B�0�(��@���������o��s�R�Q�u�*�p��q`Z&���M�<�,�߅�����7�[�qD���%|"C�/���ׁVƁ�@�`%M a?�������;�Ϝ����9�������@�;h�R(B��#�� ��$�\�e�\��4T��n_��ĳ�:R����7#�[ܘ�'7�(����C�1���"򑀽��p��� �㝇��xV7O�z`n���T��|ХRUCE��
tY��� ����e�%Wg�Ԓ���G�����'r�%�]�*r�� �z*Z��|J	�U-��k�R�|�^κc�%VUa"��@��c#���{�>&��2��Do`p>d7��Ä[�M�Y3΃�/#`~��l��0j�8K�pD[N�`׮ȬK���ŷa|jMY�[������瀱�o@�HE��Si���D��	¢�f�8�P��l/N�A@�k1jA��G'K�~\n�,��&�i��8��4�$)j���k{i"�*���?.٩'�Ӝ���/M���@�+�4�s[��A]`{����fsW�&톴i����{�*��m��=���1*�i�>H�.)��l��<K�<֝EťA��Pҥi`B��,�LE_F�W�X���Mթ� t�Ldi
�Pm(��H��Y�&gq�S�V�Z(���Y�P�� ��ႴҦ	��4��Ӗ�x�o,��׍��h2*x.Tl�$��-tZ8^�<UV�����g���1�����{a��t�%q����N���rt�� ��U�>:�EEs^(ꏃ$��/x.���a�ī���5�!A�"1v6�9[���i�"��_K	9Xu?������c8��$qF
qS�g�&��]��=��0H���x	g%����Ub��T͜�)�5e�?�%��^�J����&̰r�z�):6�q�w���: !�����0bHȰ���'�uDG��*�nıT��鎽X���[
<��l�H#T�7��:��#�����xk�LFu�$�y�6�$j��l���K+J@�U�O�K��h�p<���?���1����p+�j��%���{#0�.r�ȷE���O���jߏ�2T�Z��5K�I��Ƿ�N��^�~����-��	�3SkX��;`y73+�l�v6��ͱַU��m�S�N@+#;�k2p"`��5��v�,Z���}Yl�-�	����V�'�=� IMRO������� �O�>:�j�V�:��ȓ�!.Q��U�kHL��j�p��V���ةs�I�:���+/�J�7@'Uc/!.���q��7T���$����P�a�B0�#miN*C��m�����z/+l��܉�P#�T��0y�<T=�^z�^`J {��M�{ `�Q6r�3�A��7}�q��*s�ok�I��M��� �W�s���{���� .n���b���:��]�璮�������XF�WI\{ц���}�\�b�$̲�����w��9G�ke���4�Ť���ۉ���$C����cH��!v1*� ��L��z}^��$��0���Բr~L�e�x�.0"Y�t�+z'y\rķu�*�
��x���31Ԁ���KA��jY/�^�dm�4��fu*<ΰ�{������`F��n.n>���<�5��B��������`ڶv����v$�xR�*kRP0�7e����l�A%�_�]b+��[������
�L"Gۙ5:����&�ꖿ]����h�.��k��jZ�����mҠ�%4���x���e�C7L$��W��a7a�BI��{�p+Ȝ*�V�;Z�|���wv�x��z����`>�`���XZ��h�d��a{�t�Q��~-�`
�K�\Q?��	����9��i�VU��o��\���wW�H�����P�U�W;6�����8*1A&��%��p��MT��r X�8�@ݵե�/r9c���t��3~��@��S���\�{H3q+�D���%j4��q�TO��^,�B���&E�0S�MH?��r� {N�%�
����B'*�$O�\�|��,���~�b�G��{2��y.�.|cwV����A�W�O�e�6H�%~�䝓2V�:^����D�qL�ʆb��Wly&6���O;����r+R�5�N��$�Ag/I��
�!�5NÚ����-!y_��o�H<d���T�pcW���1����S^�uo��Vq���D�p���{�"ML��=>�D�ڀ)�g.~�2ܨ���t$����'ʐ���x�~�ɰ�рOj�[ l8µ��C]�Q��s�(X۾2���l���r�$1����=�5�����tS���rN�qe�H�r%�K���ȓ1M''�֐+m�BP����~��i������?n7�	�w�Ἂ��C���dEEZK���bbq�]�i&�!DO#�S�:;@�]s��_�H4Q�����?��Jp�2W�@B�/t�K:̥@Kh
�i,���[�J5�.��5��tJ�����?�Vs�����K�!]���ӡ�T�Ѯ��&�:�T�^�όd�.��ʏ|��v��#ց��.�T[�oą�{��{K|ԡ��=�rx%�W4����5O��"�Tp#��ί��z�mFA�c����/4D��Lnu̖=\s�?T�6"��".Q�Ҭ5E�I����5y�ϸ��[O����Z)���Ǯ�n.�p=�i0����p�����1��JC&�5�1hd�U<��V<T����?�]�t�u[�#�)$�1��1��lN?uϺ}Z8^ӱ��M����k�E�y,���(���x�}g���,
}A�iTP+~A��o���4�j��v�B΁B�K�(��s��z�^F_'2�tv��e�R��]ћ��)xwF��Bk�>��8	���M,�m#}I5E7��_ĸ�;�U��6gi����ȆF5��4.�8ML�����<�E�����Ǫ� ��a���m���#�/l�{�T��5�i�~���� ��ǘ�b�unA�i� ���}c�5Ŏؤ���GPs1Ć� &�Y�O�qppdz��9�r��S\.u�Rl��J�0���ۆ����mI�a�z}>��@^�橕��	�I�� h�Ҝ�����I��"�Q��1����F?Z򆃊K�پ����jcQ��dԩ���M��e��鵘�]�[�qW�6M���Ƹղ�1�}��Ű���"�'�ŷ�N�Ǳ��~�_hOxn��arB�d��-aTU�����j�Ж�5�Rح���E�}����8վ �ois���d&L��d��]���{��x�Q�ӱ�_�B��"}���k54a��}�l�m(�吁���犗1mKk�}b�d�]��׊������?[����ލ�@H���$M��(�T��������hz&O�D7��
�)>@�G�
#�	�2�� .��.Q�(+��4���;�������0�ZPA"�)A�$���>���Nn1B�W�04��������t�ل0����vX��YI�:��#I`jh�G�\˓���h�2~�>��/����%A
=�c'�'��ć��`#�Q�����x��"` �i7>-J<=���g�

�Ǳ�\�k�j���j1un��s.�����anǒc?@}�t��>k��������p~�e�/�#���4d�S��=Syu�Ql�?�#�*D��!��Ć�*�Nr�
,���F���ʘ�^��Ԍ����7W�&�w'�s�q��1$�H�WF�=_�o+z��\6k�jM��	�ɶ�iV�䭵:�u�����hفd!�M ��1G�l8	.c'^k���{��.��v��0��ܟȇ�w�x�K���e���
���6�@Can�q<�p���c者|[.E��>���~��=�����r'� ��W��r^s�j�+ib̽|��ݰDf��QY�_X|����\}Ĥ��nY�^���Q�?XC.f=�'X�E�d*��T�\�@E�(���^$]��R���D&b����d���t�0ѓ��V�L�j�@E���t�Nh�0P�6���Rd�N�4+#A������!�����-�@�MC�s�=ߩ1b���ө�O��~ݪ��Ƥ'��׉ �t��+SFJ���N�BlgRsl�?�_S㧥�xj����O���#�O����,?�����:zZ�<3����fV��#gZU?b³�B�]{&��_���B3����N���瞂Ҳ-F5�m-K�����mA��)=mP�3�Y�9�}��K��$�"�+�z��4��H�WŔ��y-��� \�����;T�ȐZZ2�σoŧ>��
��'ԯe��0!0J��?���a����%�X1rz��7gq�)ʷD����� GKI37D8La״_ʐP�:h��x
g�VO��3�>�s��L��7`�k':Y�9�_�,�Bԡe�_�����E� `CibP_���Ƨ؞�Fc�j���>I'�����\���c�-���k@@]�縌�b:"�S��ϼRg�m4����o������lwas���
B
-��`�}�iV#+e&�g�P�dN���'CA8Ц�K�
�~��b�d�Bi�dYb��`�I5��x����m��s����PhH5d7�&+vm�d�J�cb`�>�<�[���_��	�7�>��ۊ�,79���S���տ�ʹ����%P�?w�^� ��:eO�b(m�Eek�ʽ롺V��p�'���5��k�'x�DJ�9�C�D��\W;�`��pM�s9�PҩVUzlUH�������0����_9<r��9͘mi��{\1�Q��Lv��'�d)�g�AR��*hy����|�\@Vo)���O؁�y�flc�]8�p\�)i�m9kn[�2z�g����؍w���cs��J�,.ph�}},ð�>������I�D�!DRe��K�˵Rh��A�{�M֬��8��5^�S�uՄ�������utU�V�5T-��I�\v!�5��0VMlM|�'�����	]8]H���Ϭr\ B��7P����yX$���2&�Q���)�9#-�3$�xI�	s��N<(UϖGb�x�'�� B��MZD��,)�m%���o E�8��
"2~g	A�.�:K{M]�K���<��*���(wOy�-xx��/��ϊ9����(�X��E�7���e��Nd4��p����S��=��ST�����������Է�e,�X46� �dXe_���I�H�R!ݪ<6w3�0w��)�|ӋhбK�|A�Qmd�� H�*3c*/9^/ˠ�$cM���]?����b2�3t8QmR���H�Ѓ�	����Q�ʣe�q������� ��6W�cD�0;Rx[�Da�F~�,���l�\��vN�(r�mb�W�{-v�o�"�� 7���yc��&5�G���ΪE�&�hיFgp1[��6^O[��nŉ���ܟ\�<5MH�"� }�R�<��I��D��4�N)`�Hr�ϓ؏���(M�{L�Z�H+�@� b��v>(��t�+T���N}�ZA�ѢI���34�H1��ɐ��,��E��I�㵞�R�'_1 �E!��2m1VW�G��d�LO��,��V�Kx�_~\��� ��6�{����_��sg:��a��*����L?)K	@��PMlLB�$E�j�5���3��R��M0�Y���N��B���� +@��mi��,�9OfT���LEo�Tg�\j	b�A�)������v��^k�r��P�E�[��{#��|���R�b�<du����.4��/��$\�a���\��v��v����J��G
<�D�ǎ[N�eI���W�4pb<�����_�]�z�+��4M$�u�)<�-�o�xV��m����a��oh�!f��,B�A��3��f=���nD����Ɯ���	fA��n�"!I
�o;n��'�/}#�[f[w�=w�r�h�OyV��g���������x)[�\�&���c�3�����X����+�Q�W�U�d��;��y�����o�e���&�%�7�o�I'ҡ\�k2
 ?��acg�_��[Lh�|	�g���!ŜQMX9��IG�+2���xw`����4Qzvgs��y��lմ*2R*�g���!{�e1���#�\�t��	H9�9�14\ ����j�5yu�Ku*	8"=���zJ�;h��(o�l2���0e�	^�B� �`5z����3�V7��P���ȸhD�'�yI���I^�sC��I3Q�p��16�ә�zS���eQH�J&uFQ��)�3WL�E�Ȃ��}�$I<���%���l���vaqW�2>+��+F�Nj%i�`e-fN��'�������R�㶋w=�`�W�i6k��<#�g���E�EH�����M�'������;�#'�?B���"��N��T��
Ǭ���Z�ƒ]JE�k�z~�3�L��I���ϩ��>j��]�A�$�����X3s�Kx%v��RR��2���Ӫ0�z�!ۤ�'�MC�\�	 ��M5��:@Fs�h���6�b���(�ɘ��)���1�D�	�
��5b$��]b��m�����>�b�4oȹ#ǔr����H�з���-AЭ�� �u�ǀ���6����mV��i�Q�r�LQ��ݲ]"�����T���yT�$ʑ��3'G>�Y颖�ǵ�K��y#Z�y���0�#U��X�W0t�o��3@v4�i�hw��y��њ��/�s��sbŻ�(�͜O7>J�&�W8U\b��#�tw�F���wqF�M�B�����(&f�A'O�I}�����"�y��Gd��j�:��qj���h%z}��4��ugUrT��[��GKk�K�za̪\a��ts���b��4�Qח���w���" �j0X�u�1p1$vE��dg�?�=��fS	���Qכȭ?�'i]���f�t��e.MDE|�{'5�u�P����KJ@p��t�Z��C�,>ˎ@ೣaZ�N��id�<����]�	�j��/W�׎r��_F����<v9d��'y�'��;��\���&��)���'_T6��|�eb�%M甴�vZ���ɝN�zc��#:��%8L#bU5Y�D�����vη2Ђz��:���7���� ��� ��L��!��/o=/(�d,i|9�5���33��c �x�`s;k�\ ���/$U��,tc�oÜ��W��@�C���b����i8o�yp�|�
S#'��/2��:�Fi�m�`��Ks�d$ÿT��\z�8�/ܳwA�����ˎ���38_�r"���Ъ0�vf ��l�~�i����\4��ڏ������uU�����L]# �=���3�tvI�=r�3C�W|VM�pPB�܅6�]���j�a�����P�Q������:���ܪޜ���pc�0��}6�Q"�^�����D�i[n���� ��=F)�U[Rk����V��u�v��z�CW8�}��͸{RB,y�<x�3�4���;lW-s�|U��ݐ	T� gE�"J.4���4��5-뇐rV��(ت������8�M"�1��d��2�P�\ �@�!=g�����9ʸ�v�n�SM|M��vK�=?��\��#+��ӂ���9�
&{m�"�g"����%�#R����Z	��,<��1�c�T�՘$������}�Fw�Y2���ʡP0��P���0/@����(�\�4�ǄaP5T�n��c�LW�Y�c$#�G1t͟������v&f�y9������j���w�E[8����q{p��j��4:�YtƦI�ue���'P��q7�(ϙ�6�A+R%ș�������H���I�$-� ��s�����$ݒ��>I�Z��ek������S9�K.&Af�G�S����ò��A�z=��Yw�Gӹ1�+���7�ES38�4�ww���E�GR^��:�)?�x@D:�h�q�E3��xC� h�հ���Z�/DZ���I ��A9!�`
I����EY�ta�Te��%cA�!oSu닥r7�����
'�*��ڑ��nm)��.��?�
�9H{�.f�������1�񱦡������m9��*�]�����%��iB�Z�)]ځJ�`8W������m�4A�Zk�yD����E�C��x`{��҈����!57��o�Zvv��ص�yW�d�p�^$�j�u��k���0.4�Ö3��
V{�ȌM\��k5������ɬc"i4sl�
��-P��_l]���R�t�ť����/���c!K��?����ED�OUJ�{�x2�Ğ��Tj^<����d���.&%K�{2e�?�^���%|�>�JC�*i؂S�����.a�j�p>\# �X�{��\�0��xY����j�2�FS7��-W_��x��ifյf���ō���G>J�M��U�h�q\R����������V[���ć2~f�R�2*���a<^�#;�=�l���C[�e5���:�����!],MBp�L��:q[�0�� ����`-&!������;[R���9�v�
�$���sV�s�`���I���:�9�É�����T�'v���^�I_�D̐|ETA�o7��55�4��d��+
�E�����mP�A xĘ)��<x��_īhM�^����NB=����;��R��gЉ���Fz���:�PWR�C��}��y��+�\U�`��O��|��U����tA�dj�pV靼�\�̠���=k�5r�VI
��>�hC��QTVD{�?���FcB(���(7��k o���t���[}j���ج�(rjc[����p��C�� �K"?vh���h�ě��z�f���G#�5�86$�C}9(��i}"��;���sʕ��-�9�Ք�{bH��N���A	�5�5�0��ܺ���-P� K�qؤ���\�d@b`����i��z� =���\�t�+Ʈ'6N3J�\�'����v���8��(���UQ�Hlo�̈N�����ױ��=�����0�@+4D]w�g2���-��b�d6Q�9�D6)��t�4����d[_	���0�?�!3F��-�B��!���`�G!	�B�(J�U:��)�~a����vA�N�G��A��{�_�;���g3G�`(�����2���M�o��̚�/�܋��=���C���^� �JN��;靌����J������թ��m!��$�L5���~3L�E��>S��G���Bs�a"�WW��,�Dp��r9�ٔ<@`E+/9�m������X�?[Q�&�%��쾾�!b�S�{!Әv?6���I�nffχ�O����I\ݱn��S���*^�2�<!���%���d?� �U�W�n7�T0��8�R�����1�d�S[�,�{���~���sG�ɢ�7'���1�.D�+[���	��m> ��S�5�8�O!Fv��{0;%s�x]��?۝/T9���w0}8�Q��s=ɠ�(�; �:�ڳ�ާ/�;�3l�V'�9 ���d]K�=�uL����Ŕ��8���&���
^���wR9�[a���8� !8~�օOýŶ��+�he�q����`������3\JLs��Wa�;=&5���q��yXZ5�V�O��\s�T����o
eJ9��_�E޷x�N�N=�w���$i������SkE��r�Y,���ͱ3|kՓZ1AZU�2�_��C{%:�Z���E�Q�4q�?�S\O��N!�pFY�x���y�D�)_Z�ٯ-+T�T��W>I_��^���>adi{%�&(�<E��o�(���$��%)����`\W�;�$�h/��!pI���1��9��ݨ`�%��*.1�l���ڄ�D�����U
�]X�*���~w�����|���%,�|x�G�E��G��%���<i`qg�N*�&�m���X���}����q>i�K��� &f� �q�!_��*h�@�/	a��-�d]2�ȶP���@.8pc�Ç�>���% h�����C>M��S �V�(��3j!g^�$���6�^�h(AY��pn�$HgWCk�&���p���Ĵ����%p7.��9���3|q8U4�y�Qt�<i��y"��(�\�䋁>��{L��I�ʢ�8:�W"B+��J��U�83���:�vܭҢ�� Y��U��J8_Gk�ݍ���ļ*8�����e�G�����G�}���!����(�����
\RO1���.3�������rA�@Jϡ��ÎRP7�6���:���:��cb�?z���9�TƏ�-jǕ�]�E��=�����6	_�Y�[SmvDU�ul�Vc%��MQSy>���*p��Y�'	�(��N�������]����XZ�jc���p�c>SM9��<�-f�׿ݤk9�I�؝ʂ�Y�4fe?�3�M��hW��P�ř̦!�B��RnVr����l��'�M	���ys.ä��47S
��#�!Z��3���F%ǰķZ�C�"�����ꗩɀ�.�Z*�-�����lM�(�Hų8�i��n9���]'��#-�[�CC��P�.��\z�HW����4��C%o�Ӈ�T~a��{5+�D�%��`�2&0+zO��ķ	���):��X��j�z�8�{�]��������A����g�<�-P���Os�#�-���V�ƣ-�r���]1�T���h)�A��@t5�Ds�@�|������T�萍fcď�Y�[*��Q�lx<��P�%{�&�%߼&�V�U#ON���ǡ�����Ì/n��u�A$�y0s����4�+��<�3[g3��\1���c�s�;ǟ��?B���G�0�z�x�Z�bGZ#��� ����� cPqV���~�SLڗ/\JZ�P&3�cUU�H��h���r�w˕;�,�a��2&��؎���Ko���aE@��g���-*<)W��XB'�=�i"<W� -���Ku�b8��P�P�ۦK�@�)�������K(��봐�,�.��_જeoA_�r�}SC�x�l�ߏ�����[�� �5&r�@��Զ�����C��-~e�Ȋ�Ɠ�oD#���ʚ�l;ZfP-���sq��{��b��p-8�>Rm"E�D�����rB��i��͑J�n~i2����,����Fcn�4�/�M��R��\+/e����D�4�/�2m?��ADt���yR�W���F�3�yd]o?��F0cɞ�gZg�0hVi������؍��z��͟�����K~^\����E!���j�׫f�"�h��.������M���m>���痸�{�hu�M�����GX�w�&G[n�n���?�S[����A�JK'OfOS`"y�Ѣ(�AHS2[S���x���[��Zjf����/E�����V�<}	1C���2��9K��M܏��0��������]�j��8?Hk�#Ԣ�̘�L�-��_0�{����$ʂM�ҕ�b����J'�x�tR��t�!��Ф��ޓdl�9��Z$N
*/x�Y�4�ǣ+��#rCqi0~��R���JOl&�Q"��IxBܲ}�^	��]T̓�.���;]6`��-Ad(�t�����a1XЪ����Jq��ɽ/��(�u���#��<�=���|�9m��Z��fHnTKKl�w@j߷��S�X����vG��C��>���I�\��o,����<������0�v�@FF^��Y���2�yq��C��
�zu[6��b����\#~�
n���¬̼b�L$�p�!˧�a]>�H+�Q�@�6�����|�M[_G_=��}�mmNW*mzV77��Y��t�A��r���%V�~ ��Zs�C��(�1�q�y������4�/U�|�w�>z�v��G3U�">Bf�{7J� ?̐�:�@2@�1H���ii�>SCФF8� aڐ#�ٻw<�NЂ��"Г��uH EVZ�MS]�����~�s��^�I�o.�fi�/�;�"�8���o�"�5� �B�Dʫ�~7'�ڃ�$mq���+p0L^8�����Y�D�%fd)f��^k63��0�����N�g3U���d�`Ob5��@�}C��fI��u���X2F�;8/9lݫ5N�T����1��ݚu�ى��π�,�i���k��vj�K�H�C����[
U'��ì܅f�~q��k�v�E�ߕ���h�Y®dtU'�oZ,�g���hq�����p�pCi��x�M��&#&%��f~�c�IČ6OHh��Q�u����&��?ѫ����Wtڻ�Y�x��l��t�E�1�>:!6�-)�^{T�6t�w�~��N$��"����;r�
����n�;1�v�=�1����W�b��Y
��.p_%��i7@�1���c�mex�����55'"��X�������$�X�]�-٬i�����J��|��q�2�u�Ԡ:�" �j�ɷ���Y�A�*>6 �����@�T�Ā�
��p��^?g��O��MQ���W]�SW���������quj��I�X(�]��af���O�m���
��b��A9��2�TϪ�bom��T���;��X�Jcj�Kuqn;�׷f֊�3��:�"�����TT�5�rh ����'EuYm@7Mb��xx?,�P���|�����R�"����#�R�/��4��p�����Ӻ���[��UP�]�C��v��c����ru�Y����y]N0�b� ���4u����x��y��ʲ�`�^��#&1��X��֬v`uht�w�>��d>S7���>fa�6�u�N�Ꭴb�ed���)�:���8���v�:bWu�#�s�����R� ?�+�B�
y1g�1ɀ1��9)� ��O�<��3S��: 'R��;ok���M���Bu$U@���~u~��l?��U#���`�&7� ����Ě䓐����0�O��<��R�7�q�03� Z\$�Pc�B��ҍB}b�(]
�npf�]ŪV$§�ر[��v����8��)fp*n]w���_�5��#�{(G9ܺ�������m9�&�Ht��)�g���L�����9\��d�{5%#��f��.q�D� ���T�U� 6n����]N�qc]Ϯ$T���F�)�W�u�1�_�������.��ӏPl<��||����ݢ��In�$-���6�{�5����#gd{��?X
���X�a��D|�)�rYX�6��1��$�l`��PL9d&]�e�	��,�{�O�e�N���� u
�Q�V,ܱ�j���@��bV+ơ�q���2��"o�!�в;�xJZN�lh��(� R�����xUӅb��k)�৞�2�Z�=��PɮI�"����n��]p���{(a.(/Jn8a��ϣ׻����,�W�������|o��P�b�<�������*W���^%�v�U"E����zF��5��0�b�f���1��X�:@�u���^K�����kz�|��ɓA(����q�q��EJ;����j�h:4��
��pz&��N��^N<�)7���_�j�~�7�jT-�Enu(M{��a����t��o&ޱW �X(�Ӕ�;$�@�+#���-�y5=(]`p�<�ݽ�(�D�9��=�eB���K��Fk�����Z/��¸��Sc(���4�5L�g�^��m�:�y"��#��i:�\=�x<�@t�7y�_�4}����c6.G�N^��VyC(�wK�o:��\���0��6r&��)���M�9 �"��&���KuSI9���{���9ol���O&�9g�����]��gG���W��2)����r���R�O��6W��0$�E>�:9��h��?<�@\S��x,��]�(�ȎKl@`G�BvæZ3ѷ����Y������m�ua�_ȶQ�'�@�Z��b?����Cy����&f��6gJ,4�)i�=���wĚ�i�^���n���0��<���6�I���8!����]7�#���T�@�{�P��Fӳ���g\�x�8�Ŀ�Vi5����|ܥ�_ �j(����P��aUE���Lc�B� w�<��|T��ʖU�"�*V��Q^V=�0H+%�sc�b�KǏ���R���<��=�����Q�B���S�vA�̺~�=� Di�ϗ��Z=(�Eeݭ�9.�]����RF?����@nQo����4���[}�<�Ua�$��_��	u���!�ǫa��:)�����\z;�	��?|��C՛���P�0p!�z ��!
=\�Z7���k�6���F$�T�b�O��7KwULЯ.��7��m	dేa6�h^�@��4`�Ԉ��Yl�������a�|I	���b�h��
�pFz����#<�H��U.ĿU:�lh���bY3�����onT�
������@u{��`3�Q}2J�T�Fư����󖑚sL\6�w�K�,�G>��kp�D<��� ������Fv]������ǎ�W�>`2͇?u�l�RPo��l���K�����S)��ꁎUm����s��j�ۂ[� �\,f�0ܐ%fL�9\E<���~��L�,�� ��O��]@�t٤h��1ǥ����e�g�ٔ�ᾄ��?|~�_��*�J L׼l�&��"U�]�Js%ԚX�������b��"Y���L��c���o���$�G���oν��Eƹ�WU3q-F����߃���<��bgHA.������aE2����?�Y?6�����+ס�D櫳�oѩ�>�h���A�O:��ޏ݁��A���gB�Ĩt6ʻL㰱z�����A�+:`�u]�p�D\��Z�|�I��ڕ%��o^F�0sz�1��ђ�v�xj=��P�nm��j�]�E�E�?�tu�js��V��u�nbsk�Q������pc���#�L�2E�а�� 6c�������tE����|{�������� +�G�U�Z@��M�[>�T�ݯt��q��Q�s>��T�f���2�	�^���Ovd���c��٫������/h�h���w���H%�1ʱ�<���?Ѓ=�XzF��r����	@3��B0�a-�[��������3�3�U�<�F�fvY9��Sj������.�I�۵x#="t��N�&�Q6%hf��<!�Zq��-���ƌ���Im�X���?yFg�@d�J�8{��jg1X�Cy�h����s�وh���
;����0�ѓ:4ϗ?�%w��AZF��'by����t?�~���L��mIZ�i��[�I�bc�j���g.����b��d5�J�S��v����N�{�T>9�
�:j���HF^��֑٢!7֑�<�_�f���*�GOW���/RR�V�o/(�`����,��T��I�����ü�՟�0	M�̲h�-�^2���vHӪ�ɢ��a��X��.h�rw�I�O�K(������|�*�H��ƣ͓�7��l{k�Q,��x��R^�8R�Z{���?��A�V�,ҥ�k��8VD������4��w9�U^�`����Y���뇔pu�P(���&���N����W�.���O��֖ģՃ�;4��f�$��K�������CX"ɶ�U��lA4�Td���\���@�&!*�Dŵ���e��!�o��?�2������d�S�����>�V���]6�t�GAE!9T����=����N�3o���8�ƾZ�c1\7�ճ*�UvB: � �F��v�P8�{����p&����P0<	@�y�9��S�R��	��od�#�)+���ʔIH�q$�#Xd(�����k7� x$�d����Ľ� I�#�RЮP�:�IT
Q��"�P�1���702E����r��2%��	/E�e��nG��{��<��F�N9�K������2�%��۪ٚA��,���yD�Ƒ����<��)Q�<����+U����86D�%p-���@w�oW��9{ҬՋ�cr����30n�B��ʽdy��N�!���m��k�~��,��%����
E~m}&|�h2 �e��E��v�[/�X�r%İ�`n?�[�$,�U���,Ә��R���$a�f6}؜훌����,�֯�R�r_c�C�0�(-q%�tU�`�&�Y����\���v�8!pJ���Q�p�@�'�H h�>R��kq�wN���A8`���I*�a��R ��e'����z�L{���%w�yJ �����u��M���Qכם�<��X���ѣP4�B��0xg�8AG�r8#�=B�caξ�|�G0��N3-�s�7n�D�8���N[8k��k,�N���?< ;ay7���α�5h0�h}�`_�m��$Km������>�Ò��
tZU�n���XH�"O������3!uêZj9����H8P >���m ��]��
�`d�U��4�KW_/Ⱦ����GtDܜN}@[����x��ǵ��g8��f?e!̏� ���]}fZX�ȗ�X����(@�x_��dzCT��A�����Z�������R�`AaF��>�*#t���)���Z�S�,�ܻ
�5)
4�s�� [����Ϸ��w��ɥZ����Tg;�:����sb�و����B8����N�3�Q�^8�5�4�/iُ�s̢�X���ެ�t8�����D�/[z"r��l��@2��ԯ�)9��qhR���:O�l|3�,��NK���Y�L������z��Hk?��[���8��B�kz�K!��V�������2�T���;O��X��<�+�����.H@
��Δ9�`Y���ً�Di����u���W�3�,�LbR�K��ۡk����Q���f`�ɚ�h��f���")����ᄧ�4)��oWQ�.%xW���M����.�Ŏ �dW?�d��X�.�s�$}jb8�-:�D���{��V)5�64����M�T�7(H�	'
���<���x��}��'�Y����^u OQ�w�R�N���CM^�EߺI���a�LO���Y�ŬL�w���|��UeVQ4��tH�?��*�UR����RJ�\{����B�/�@����r�%�>HY@�'��ݐ��|�Q퓗(��.��Z���E.���G��a���=@Ը���5�,�N߉��<5z'���Ђ:����8j��@I��k��,�������%��~&��Q��8M�.�:چd�=��-���
S�|��N��L2�(��&�b*}u��<��7݅��E^Q_���J_b�>�/�zP;���Ȕ��7�s�BG��1�]~-��[�����,�	��?��!.���	0j��{� a"��ȸ0w��-�,��N�-\F)��Ź��@^���1���N2�E��A����[ϼZ�ʊ�]�^�'�Xą� *�Ɍ�?&xO�ܥ Ќ,T�Rи}�<����W��<lk�%X��a�AoQَmx���aI��<(辕��h�y���Fա��R2�<�(���k��J)y��R��6Os]�@ �I.�f��5 ��Gd�����]Bw��[k;[��S�eb��TV�mH��SU� D0�Dt�P[��a,�5�d��pq[�o�����)A�$����Vw9�\m�3
�M���d����b�#j{Br�ǏygJ����"qK7i�Pp����-_��:�y�	GՎa�`t����Im�J=��ԵߩE�6�,�.�@aqn�5H�W,�?Ҧ(���W�:�X��+�o�4Iw�y��֠����wVs��y��=���Q�'?Uai���!��>e+'�� 8;3�&�x�V[Bu�����v\!A"1]�n��0���V��\�A�N�:Y�m��V��
(:�W�w>Y����Sڤ�	���Ae+R��X��O����v��Z^�i��AgM���5nj�uʯ�AWd`W$>t�<��Z}��o�Kn�|h�R�;��Lt��':��܅g>��l(�P�oX
1)��)�Ҁj�i�������*�\�lQe��c��[˩�M�9�����1�U��6;���l=j3���ۥ�+GZBS�Ҟ%Kc�7��륦�/=��/�V��s�5�|i��]ХB��ٻ�y�\��2�j��jE-�!��Vϸ�/;-�f�� � p/�b�B���R6@_%�A�k!�t{N��O7md|� ���1��A��7���oN�4�g��6O��%}e"�~%��ȵ�Q̛SH9��O���[%Y�ա�B��������)��ф��(E����9[�p��q����N�*��o0��X�oѕ�n�+P
����O����×���з�9�\���,9�G"?HoTzg��rtm�o�bZ2����w�20�9m��9�sT[������%!�F(�,`�����r:�����z0]B_�E�BTZ�]� ������X#���H[^�s���܃_���� Y�=��)�^����{@\�//��N��Ȳ#�ȱ6���\�I�V�Jd�*V~��QzK�(y��$�$kG-�aH�����T��<^��޾��;�@�І� }��Ȥ<�jm(E��le	�YM�p��ָ�?���>tp�f	v�T��9v*h����n��-��;vh�0�棇�ur��|Q5��
��Jc�x��x��e��Z���(��i�i�ڈ��r��)#ݜ����Xo\��^o��4r8ϛFh������R��E �� �EXwx�*��`����x��6�D*_�_��8��:��g'K�_��r���1�Ȩ�݊Gp��3YލG�(<e��g��!S�B�?)�]qX�ʋ��L�i���G��ӈ�u�0 0V��#��{>}G���Q�����Ze�������(.P�����~K����EK�c�7���K�hl��&�}B�X�I���V`~����-Yk0[V5�?�/�Q�r�,�l�,RNP;�^d�Fy���	a ��a#���5ja�x�̳�X�k�-˫�+�C�Q��
T.}�����Vb,�R�l)
���12�=�tEp����g^�4d��(f��C���u�Ij�u%�$%��y�ih�\�|}?O��l����k���ux�}kc,�$7f�$)ŻU~��3p�Ȳ����`p�/��<!dd)�p8Xo3��pm,����]������$���ü#��c� �(h�N�s�D#yS�顿Dc%��id�� ��nP#bη���?�>V��(r��`������+r=�t�������ř\*��u��>;��nۈ���'H��Y=j��9��I����]Ԇ�vw��/��M�U��)Tt�z(�\ m��UC*�.�h���;ϯS��$��ٞř��%M�C)ؠ1���3�����j5��ԛ��5QF��E������\
��=�o#z�(TƊ����F\�����k8��]��-6lR��Gh�*�,�����J{/g��l���a<�sa��彩Gm�,�̌����r���}�.n��8,dնHt���9��F�G�J��(�7�a>��^C�J:�qg�܀z��6�j43��28���%�gM�wwe�uz"~ =m~6m��x���ݓ���Ç�'f�E����ԩҿJ����5� �T��-� ��Z�t5�SO5�w��2�Ndc��5)d?�/�_XM�9�]�%�E�((��,��(jd6�u��q��[���z=b�I��o"4T���AP2��2$�w6�� 7�qţ���7w�ص\�(��а�P^�;D�ّ��%A:>R�^}F����i��W(n6y��oW������^��)�Bp�q�[U��r׸�����-<��0f�K��%�>��Yd+v^�
��$XӲ����_]�˲r��t��=����-��@#3�F<L�d��vi&�ë:�F��f(ʞs�Ϛ�?�%7zU�j�S���A$9ו�[x��Z����/r����E� ����(�5���)��~ ��im"�:��H.�	x��F���Y�N�l���&�X���;��2m`4���,.c�-Ӑ�+�x��"�Tn��a���0��J�U�o�#z@���ݐ�� -��G(��Y��>�:�B.��[�v����I��R ��INfl(�C��3>�x����g?.rh�X9]3#I��}T1�pM��{R7�)���0�����r�Cn��x^�<��2�؏��O�S��&�Ȕ���f;6Kx��)���(8�qh������u��
y�oج�o���\a�ʗR0>����o,ؤV���ȷ�֖"��#���p���
�m
��T�Ae���ܛL��GY�Y��4&5K?� ��4h�p�,�>��X��M��UX�g��s"gs�
���:C'�y ��lK�Y��ܲ",e\"�~��Is0"��W�R-��m�(`Y�5*a�_ͬZE��x(SڊT����<���0T�/]�>]��K-�k�-֭�$Z �OLh��ł7�I���@^UF{�(�۸���L�ֿ����M�<�sVf�g�Xhjf�Նܸ^� A�n9�V����cCX_�i;t���Bq��l�.��,�|r_B�B	��XXDRL<1xɳ���sU8e�%0�� L�'X�e��T�_ɞvZ�L�V1z����� @$�}�9in�Z��R�{��i�+?���?KG��E�n(�R���k�w�X�Q�+���{��Oa�@a��ѓ�72 ���|���UEKL�g1;�m�z�wQ�f$ʁ8��ʢ���s�r%�6`~/�֪c/�N�k]ө��G7=�?�\�#X�`ҳe�7�7��UF^���I ����1��ǯź�)�"->w���I��[��0F����K��M��gQZof���ٴ�+z��I8X�;7��J�pZN{��xB� %=������a�،�ȴ7w�6�R�\������s�NK�Fk�NtǍY�OP٤�:U��h������3,$@��(M���5Mߦ�e�'�
r��n�7NL�IYu]���6���0H�����(BN������b�\A�\�Gd�PN)pȓ��ZD�S�G�Z�)��r%Ԝ�o�^T��.�r&Vs����dD���;������O�t�����;�`~;T+RQq��p�i��^??��e�Ñ%]Z��9�۳1	+��M<��k׳�u\��R,�q4JzlX	�id2��F�rm��q��4S���(�j�b��_�ڠsc!���6Ζ�$8?
�N���z�TңeQF~��j�7e'��c� ������(k61��8_�P=I",I�྄}BN��Ø����c�E����U]����_[hm%�r�
��f��%%�3ڪ<`�0@R�)h�R%g{���՚H-9��k��"�!��w2N͖ޔ�����\�%�!��}��2�uJ�3'�!e��IE�o��s��s����Մ 0ʒ�4H;�FLX�]Ke�]_*��W�Fn?���:����{ҕ��;�*�Tx� �uI� ���k'Z��Ѫ�W=Cf��ɷ�R�o9	x,��~��A,p���	] ѩ~�����+n������9���h���>������g�v��:L�΀��!n�/a$�+��ө�O�*e��ֻ	@j�s��&�5K`+��w=M��	���(�>��?��/`�iT%�i��a���>aP0�<�P�W��~���^��� D�˫��[���L���e�$εa�� �����n���%/"�@��}��]q���'Du�T�IY�p73����	�\�С�E���J�}�Ӈ��F@�祽#�o�+1�M	2���p���zӾ�-��[܂��$�<�g�f)q�:,lz���D!��d�����XLWI�d!��=����h�5m#9|T�����2Иm�ZR�n`��M�z$���V_�*7Ȯ�Y�D���%����l-9��>D4�r_�t�Ma�Ԃ)iXCp������X�J��'�^g*�O�V�0�A.J�A�_���(�{l�����9Lu�T��Tz&z��&H�������@���z]�Z�7`zٲB>�CÍZ̏���T	���a��&^�sO�N�� ��Mv����-���̦���S�زi�`5d)�	d:Ԕ=�聡�G[L�!��o�^�v����t��	jH�ǽ�����	��
�o����E_x:\-�j���}��d�Ԭ'p���%C�t��!n
;mé�!��"j#��'�w��5�ѿ ?�3"bWU�{;����H��=x� � �1�%�l���n�+cEN�b��Ş����T�{>�.�m��Q���Kw0(y�a��谚�IZ�J�>$�D�S珞T�y�I~61�a���G]��lƵ�ek9���F:���F|X��ȣ<�ĀF<�?W�3U�^嚉�0�v��*끀�n�Ʊ���3c��I�,#t_��ڇ�jb�co�nn�"���O���= q/$L
�CW-���r(�Fn�����;
��\���/e�{aPD�(��Պ����S�_���ZE�::�u�ք!1=�n��u,'��d����R��g�����Lle�s5ʍ�UNSCs	g|�Hߵ��%XÀ�/��C1��X����_���þa7lU�p�d�z��1�2��8߂8'���.�|�\	���M�$'.��֩~{D<�j1=��kO�cK$i�p��2�3a�1�����3�d�ӯ�����+��4SV��ݘ;e h��L��p{��#�(l��� T�@���m�O��Ak9��Čq�.bW�؃d�	�����	^��{̽�O7E.�GS�:���I/�Gf��P>�wR�K�����j�0�Z%���ߘӪ��������#�c�#�.�-������#����V,!e�gl��\�|�1��*�V1[wo]�	=ҝ�6DB����O�.�͍-�tr������~2p�laAc'�u��c����]�l+��8�=�[ ���� �8��%�4���A,
2�0��t���O#�������ȥbH��}�1m��ױ�4��Mj����pm`@����X�6�u���R��c=RL�F���̋�<	I
���$w�����O,�&2�FJX	)����B]�y�z\ɗwd#�8��]g3"����7Α�ՂW��1Gf@4�FXI��&����@Y��_��[��=@]�����3�6�}�W�(c������T�c��!��9ռ|5W�5�����04P��k���0�Zº%����i�I�{,HJSR�+0�Ο��[�u�����ط��z�wѺ_.S�Iȱdpm�N6��uT�F��{���+��jS�NN_�ү�fvk0�nВ\�T��c]$^&+���V�s#|^��D�i�F�`�������Ls�V&z·�	���&�q�	�	2��:XH���jo	Fx4r�!��ޙEW��Օ��'Z�k�K���fVG��8�2����x�=O���)?��H�jN�q�z��	 �����\�!�ͦ��$ɱ�a��s^Q�ߘ�{�p�'N����,t�o���'���?��W'��Ԣꢚ��E-��5�����z�D��?%R�P P7z�X~�����Љ����m|��F��s/#i,���z\:�=�.i��)��Q��\$�х<�vq�̩� ���7?E�:�@�ǡ\�\1��[_�����h�4Y��Z�nlf�������dt��ڭ篲�%�SC[�����;��[`��*�)*p	�T? �1�&�0lQAx���"��-j�`�%2��JO�=�x��3p2��r쎸
W[;����e���J|0����7��}/�>ѐ�s���>����/��p�0�I��Č1i�V�Z�8���#�%�X=����MH�m��p:-���C���/�'��e,qQxą�n���k_?����nP	�T��]'��#�=k�ĎhȂ�k�ß:��L_�㺇v�"��7k
T��_f��|��9�3�dѮ���o
����
����YT�]>�6�x�����PT�m�^�.�O�.�M+���~�4�gc&��^���,������x�S���i�3�f�X,WY$�.�6��. ��Id��9�bxQñ���e�zo����X���oh���Y!^=?&��I�yl�����N���cߝ�SZ �)�z�r�dt6�z$9�����Հ
�Tۙ��iD��sO!A��R ~6�@�����n^a �Q�U�;�N�&�D�6����'G:���[�ԝ�wiN0�O~�;gǮ��d�M��j��PrQ֊u��iw4ȅ ���B�;��P��ڬVG��pD6�֥�Paty�z���Pn��I��T[�����$��{�U7�Ow �FCWNd�]���0�(�����)}
�	]C� \k�x���Ȝ�\��b���]�y;�O��v��
�^��C.W�����m���/=�5,��
����{_Z�>�QGS��?_�	o��-�)5�� _���w]x��J�t}b��Uu����$�MZ�_[��Fji���e(]ئ���ˡd�;�1���mV<�S!�#��܀;5 ' Anfe^�XW`i�Eޘ���S�ǒ=��>���z�:|���C-?��)��މ3�~v��|05�Wu���\��NR�.��g[�2&aM���V��ORC���=��n��vdߥ}B�w�w;��V�8�,����� )���C��ot9�cY��<�Y^�x߶�k�E��������Eq<��*�O��赇K�*��V��צӋE�.S�/����L��Kk��J$�s$��8��T�]��1��OHM�I��E�h#�ȠD�afI�����6�S���ㅸ����Q�i�@���t��v��:|U������<��C�>�Kڧ��I�YkN#��� ��V�4OKҢ���v��� U@1u�Y]���!�\�,T%(�n��;>���m�'Vbá��D�V����9f�,��J�hy�!li~��5� ������r�#*����u�|��_�M���A�^�\��ϢG�⩋=q�dj_G��^�Q!�z�<�`�`Ǌ֑+���s����s�
��Z���d�}^��#s/�܍�@���[��Oͻj5U�2n\�)(��QDq,�+�Ǡ�����]��g<�j4kG1Xà�Lr�v��.�.{�q�@5e2&�v���'�������Q��E���5g�Z�w�4��I ѕ����%�t'^�x��~pٟ���p�6 )5���P�^���yǊ'��ʣ9}�y+d�I��k��-l������B���Č"5B��}a�S����S����4��O�uJEF�Lo����_�6Lq��U�;�h��#��g�u	&n������a�����|'#�D2gtO�����b���?7D|}Kp=hu����;�8Yhm��;;����Ve]��VpE�!q�r掟��mj���L��Mg�Q�z�iD/^���'pw�j� �޹� *��,:Q��^=����t�����a�;�����wIޭ���O�B�����q� �J����b؂����E:L����4�O,_�r�S{]�6��#�;�w��|�
�N�^�ȴ��?
gJh#�6����&{A�{�@����0q�a�������"�i��؎4f�π���}#�no� ������7�ܗ�=�t]�+�;s8��ٷ�-��Yv���[h5>X
T�zz�Ǡӭ�C��Rkc�p���D�I_7�e�v�Tl�CC�f��6�`|���HAf�ɒs���g5w�� �q=�`ŋr0Um����w��4�Ο�lJ�ϵ�(O}I��+M�K\?=F⦵a���������|,����.~�;mir��+�����2TR�V�vzTr�Mv�X��hUUi���`�$ɶEYb�E�� �K��(6�Z������/��yO�h���r�N���.�~t҆?��MH<P]PH�8}�m��b�[��#}�Z!�����#.|	�A��q��C��mma�L�xJ�Y)`���c� ��r	.��s�ˀ��]��;�$* ��M��l|,�
�a���4� z�(D���(E��q#h��e����c�����d)��IBC�zz���JBdŊ��β��p���}��舧���k��w��%���CW�Ǯ%OG��Q�}�g����r+�V��]�Ӡ\����'}�'�3�j�<�ײP��X� ja9�&g�J+va>�+u�����밠��؊nmub6����, �������̄Ek����BA�d��~�'�k}�#��Z�d��R��G!ps����w����|0�N8��n�z�a
����A�a�����#˯"L����y��h�E�c���_̒�p.sK&�*L�E��'��1� ��XDx�J9�B���%'�r�u�3���~*s�)�����0�%^3F@l�F��L���a��e�bY�B�۷@;���ݝ�]�"�[ek\��W��w���]0��tW��,��G�#�t�w�mT�i:Y�ɽF4v��:;Xd��7��PYd�b*�	������K�o��t�����~M�����9Pt���A�C3�����N��(A��G	*���K�g�qK%�Ʋ�hr6*�V��ۄ���H�Ó+ȩwJ��Oztw�H(Ь����v�d�~��$��I��E���Ү���Z�X`����{����ꮳ�=��@�$�U�L�E���#B��Q�hNm�/j�@ՈS�C����t����}��ӛ������Ȓ���<�lH
���R��B����'�eq���M 	�,���ɢ���{�����l��W9@��1y��n�,�$i�6�u���0E��Z
�B��@��:�k�?#ԑ$�x�}Q#g�B>l{̠�O'Q���>h�f%�d4���9��u���AOT�������!&�SS:�6��'�����$T�PZv��+�ܪ���v�˨���x@9�ơ5��)�$��]w��ǔ,��\l�F�En��u�R�rM�}L4̐��� 칫���Օ봮=��zB��;a!�����%�\�]�)��< �C��"1$�U�������$a���##l�]sV!���H�u��Aj�}v8�r@��3>X��b��Ӎ#��QQ/
��%���͸�r���&�ea�~4�쇐����2Ӫ_�y��j^z��(����u	:�$���YK���0O�r��I>�_����[d��cD�p�a����?�oΫ ��s�ێ3;�m�[���[;�O�Փ ̓C��.���e[Ď���22�p���%�m���o�gJV-Mb?���^!�e]X~���SR������k��t��#�����_%{�b�"N�I�����D�">V��EB�ܗ��MߌL?�$���w�a�Փ��E]�N�iD��i�PG
]g���p�<�X7�-V`�'�	��^�G�۽�_�����9�V��/�*���B4�ˑ9�G�6�{�y�OID ڻ�W��k996` �&C���
Ј�iu��H*)j-���@uB�y�7��h'ZFK�B��5��vD h��ݩ���wT�G(�s�RVÂ*#0��A�X��Z�k��o�����`��0[ŽRY;��Z۵�r>��i�N�`�/��D�RB���@�߶
�h�i���E�٪�r�l���|��>r����㒱�JÿE��F*Hv~�����u�������
����������\�j�	��	2�^�U<��|��3(N�M�'$n��ؖ&�>;{}İwsļ���@�-�W�>��\L���������8�b��=؅85���[!�$�t��(A���MS��|�Ws�֦[�m	V��U��R���g4��&Q�D8�}XMj@�Q�ѵ�1
2�k?4�݌�O�7K�&��'��'���JhVWϸN���s5NU�D����Γܕc�Р5Ԟ��Uc�4��<qwZ*|��
~-֝��D�aH��WƬ�M�((�Ue���>��2� "�%�ʺ�"�`ZM>!�~�Y1�t��O���ٹ@��Z�Tޅwo�t���S�a�3d���J�x��0�8U�+6�&Rc�Ì�8V}�)����Q����r��$(��VJe�,���0��K��+�X�e��b'`��!|�@�g6h���J7-M�E}M�~�w��I��$�3��F�R�r�H(�D%|�P��~�+�b�k(�+��h�D�����54���W��A�83�v���\�H�8���9�s��-Q޾#�mt	�ycҋ
1ʐ`u�Z���3?����2����s�Tbf<���C��\�l+q�ʋ}�����1��0đ�$}RM�m%�%#�>o�Ӗ��p�dF�@A ����ݓ�\�"��=s[�v��@;# `
�J�a9Н,^�)];G���9�\k�%��'XQ�|��r�����/qU��ѧ�$-%>e��Y{]��})�
TY�F,�����H�����+#qp��͘�HFKl	%����|���Ue�����2ڕ��C��Gr��v�qS��R�|�W~�m��?��,�΃��<�4ab�w	}9TÜ$m)� �&;�[����w�Hn\Ǧ�g�K
A@#jz��+H�(�J�$���P���C�6O��9�}���n��y'_��H����μ��OYCo}�1��!�mC6[�`�]�����c���*�0:q�w�ϠA���B���܎��ګ?_��!�d�%�ٮ�(������c���<i��"[��2�+�Z?6���U���f^ZN��9�U�o~�i����������^�z��j���PR��~��X`�x���݈^ӣ#M�W��ޮhu���B>>v�� ���ڃM���i(t&ɄS9c�Ew�cr��r3	��Ѡbj�$b�
T8����F��H�4�1罍�۪B��yW�CE�x�`�@?�1��'�]�1[�9�Sw�5+qC���Ç�Ȟ�J�Δ=�#�����p�de����7��ё.cv��L��b���5����#K���f8K��f�����~"�� ��?�T�F4���-���$����s��r�"�jS6�"�
0�R��\4{A�&��XE����8S?�����~&�&w��P��T�$�����fA�Az�����OW��5:K8s�y_�����'-b59��(/7��\��� �FJR����~k�B{2��b�4"L��@7��3���i��ݿX;j�����o�=�����*@x�u=i�H��0���z
U���hQ�������Amv"rք�ͻd��#�Ɔ�{מc����~g�q�F�H/�.t����ex����b��E�9@�n�v�D*��E����ٷ����!Q���׈��@��=U��kG8!��Gɂ.]ʶN-��	udZ[+����C!z�[��n)�s�W����+�������م��«қ��}��r�#`�V��o1ؾYa�C�>x�:B�DYѥ�Qj��yyh1+7�5)vU1e��N�>��c�(�M+�U5|]>c��������ˡp���""�O+��c��u��N�B���S���!�{�Ɯh�I"�9$c?����s�37A��UR^�Y���>����,�q�<���W��0!�y& ~U�������L�;T���=��ˀ>�Ӽ0=�_��]ڨ��Y��h��F�m��=�Tp��@42v��\�����b4+�8��X��a2/:"���Iqb�����!���>�S��������g`��RdjJ*@2������'�9j�W)\k��g�H�A���	���)�%	;#|�=!nl�w��@$�3z��͆> �]̜�Br���5�-O ˼��颯�
k<�����(=.�4'Mr�H����{U_��b��ln()N��AۭK�׾8�|��V��|�NeǾ�Sũ��K�1��y)��K�����*'���H�45�`2��]�%�3cȬ:S�����t^�@��C3���]�N;���a!͠OnF5 ]iMO��5kQ
4����5���L�����GFS�I��y.�bU��*8mc��x� ���O�U_�7��հo
F��o��n�YI�O��W�B؁E�a(�.�����A��r�ON��Ӕ�lբ?�N	B�϶/"����h	�d��1�}�B�L�3U��c���U��'X}���)�JV?���#eǝWۂm��E(�^2�9r8'h�l)	o��XBAiec?�Z����_���ڮW����˳A���#$U����쾨џN�<�P]�`�����s$r���	g#�iY-糘�7����R�0~z%�PN��F�9����'u�c%�lvg���W�E�
�yB?POY _���0{�et;-/����r5��F�����(T���tq��97�^�U�`�9����o�y�rf��ډ�6$��e�B�R��k�\v؆��9���y���/�7W%�h&2@!ģ��KhăJ �q�$ߐJ�L0n;0��{p���\�ً�mXa�+p^k�O����/e�$F�%xA�?0�P�PH�B�������*�n��69ܥ�l~�����B&zRV���}���9QH�E�-�Oq�6؅A֢��p�ZϜ��*i8��!k�����8d����Q�Q�s��OC<ma�u"��qn�q�u�L��vVE���m��[ E24���lMVc #�ԃ�fB���ʵ |�yƻ�����X���*���
�(��8�q�2�&?���NKjqCc�?�3np���]Ր�.D�6����-�}�_��k]��|8�<E���LkB��+��ą���Yk���b���Z36�2�&�l��럢:��"n�,�"t���L��3ˊ �]R�lM^D�z>mt�[��O�V=����(�Id�"����+]��uJ��K�N�7��XD��ƺ{ �\j�%����� (�O���l+�U�}�n#���2^�=l�4��ɻ��\���6�>#65�����Q��|=���X���;imSí�<�j��+���A��+䞍�r+�<$`h/Y����Ul�A�����
���R}�ڂzr�YTp��n8�i~��Z��<02, ��YA6�##�����m\4��2�W�h�m]�|�l�&C�q��'�Jlo����qmZ��msyeP�}���<^#�,��c��
��QFA�o �R��klnBKP��y�6�*=3h�S��ͷ��@`cīDpt(��`R�,���V4;���A�%Ϧ�F����4_F�厄�*s�ځp���Kat̽9��	�v^���1�HP�wi.��*HS��/�L�?R�mD�\�ǳ�-d6Bb&V�^������I�i��TrJ�l6�9�z��5��������	y���V�����f�h�$=v�cv�f��rt�R?$N��Ms^�f�63�n`l�Ҧꢩ��7BA[~ەg�9�fj=_G����a���*,�#D���D�%h���^�@#�����z�$Hf2k��F��S��>��\v~(�ך>k6/�=�µ�+�G����Π��w�ԩ%���+ ��2��!t�&@s��Ň�dX1(�N��G�]i�����~��SA����xoY�e��	ҥbX�!#+o�G�eb
���ٓhϮ�����j�.���m͢
_�'���N��]�(:��4���a�9��&��+�~F��gg!����솦�j-�������͚���ڗW9f$^`�kL	m&TB�^�HH�{S6d$m1���+ڧR3xKZ�����\8FgQR�'��E@��߾io /���>S��mW&���B��0s����u������|?%$ 7I�Gn9�PYs���4*6�X���ٹ����U/�`�g�n^��$��S�؁O{�o.[��c\?(����CWz��&3\��=���]�#�D¼n-�Md�`r�"̎2�m[b�'O�j���&T�=�9�wlSq־?i�Z�.A�׊����T6F
\�
|-�e'�!4��#w��ۄ|�]S�N63B����~Z9���A�Lj�A�=%��l�`2�p��=�����FG��ݺ�r�ͷ�'NcOzR�6#S:�����U�8l�V���׬�5i�˖ӊ��?2_<X1A5qq���-� 7�u���S|��r����}�W+-J��K�c'p,�d_$��G�]�eVM���p���(�2�c�sC�#�.S��%��Ӊ� �l�)^x��� Q	�>�9P9v�����M��Nb�Z;�bS[
��菐�^*��W��Mb>B�vw�q���r��4��x߳��6���o�V!����ՍF�Ъ/-=y�p��ޭ�&k%�F��UO����)m��qG:�;g��g���d��)e�Y���z�"E5e��n�/$���<�QSTO6�h���ۤ������W���H�d!S��:�*�⧏�c#�B�U��?�u���v������9�hM����G ��UvB�t+��V�~fk�ԫ�N <��q�'��,.Ot�k%ٲ*C"���>y% �7�6)���؃'�ʑ+���(�ܲ��T�둒w5���	�K�����s���\��t��5����cm@ծ����FG�v��d�m�3̶�]���E3W�S1��	��e�7�	����:��n 4�)�^#f�O�N���u�͓�6b}z|��h%�-*�͆㉈���wU�E%�t;4��*�^5U&!�tLL�d=�b�ji���){ B�|�.��0]�Z���/�9���:]��T*ҵ�E��_�+�
6�!9݂���7�X�b�}�RcN�ѻ6}�I)��,�(zM{����^��ۉml�������>Y��Ρ��T��R VN� ߰{bf�/����u!L�}��Y��{lWP�,d �P���%מ(<@$J@UE8\�c��G�NU��e��q��[/�TY�cy�=*�w&l+.�
�m���ܻ�ڷ"��*p\��6���u�H���P�5Si�{"k#_&�ς�ufQ:���'�/�f��i'1�(������D�ܪ�>�]p���Ki ������+B��D����
�[������uߟ
�5�I�����O<=�8�7�3�ɰ
:�����E����8+��9V�^�_L��;�lKg�̜~�]~̡�/�I��\�B��M�B��J�u%P�U� �3Lle񓾭����x��K+�R��W^4��s��9�G��,�W4��lI��U?S$�p��c
e� :Ǻ�W�3����-����ɾ��u�fsH��Tћ��,(&и̯�0~f��6|渗0�SNQ}��؋M����	����r�ku�K�f��q�ç��� ���.V��LBz�F�01M�3+����ޙ�u[�\� ξ0D�ʢq�#h�4�H���l��4�� O��'�s��:��$�ӆS�A�vｗbb�Ķ�ꒅvb��A֖#e�C�$�� �=������²!�Ѳ|�A8w�V�?��Dx�+X�I��o���R;��y���R*�Q�Nߚy�64W6��_S�oř��W�AAc�q�^�MW�ݱ$" ���:G��~��Wj����W�b�N�w��5YZH�-�5t��a�f��n�R����ZS�N�[����dqB*P����G�M��C����ϟ�W������;��mc��X�������F:O���)��a�5��=�|������Au���]��"�ݚ^hҢ>���DR{{�Hb�
�\0�DF{�`�]>VJ���80���D|��Q�e�t�T5�z�,V��i��^�"-��xGQϤ��R��F66�-�B�@�U�|J����^�X���a���Q j{��SVy3�\���1�$�HR�ɡ5v�6ظkuv�N;����&��a�	1l���ӥ��/T�=�L�\gQ�:~e��NY�߫���Es8�M�.�JHƹ�X���$����$�8����:'oz�����*L��j_V�l���ז�|�ŝh��`�)����w
��2�L�[/|n��g�CNxluB�	T��a� �R�s;��Ӿ�����}<�d�'�1X��	�]�y�k�(g& �����	��IG��s�*��m��$�l�d��[���.K#5g9Ln={�{�+�����ר?������d8��#m��qge��ϐ�U	ԩE�8[���or�����:o��!ß*Z6�$�dNN��w�Z���s̅?�Vx3M��}v�����oX��VU��,�U2�ј��~M�=��	+�[w�������k�M�t[�R�a��f4@x�d��\��08B�K@����&�o�2W��'���uJ�� b؝&�p�C�F@��i��i����*�(y��>�BQn?���
70����g@>�����Ȝ!ŢվQ8�i�!$ �i�!i�����HX����`�(��^�O-F�ʟ�.��w�T���!���:��E�X�Yְ��d���
)�B������e+��ye�|��Bo}.��.��_��ːOrwZ��z�$|�D{���G��x�Ki;�v'�\���ݿ���1�TqO�������d�ێ����A� Ib�S� ���ͥ=��Zۘ��C �:�y�!сDZL�w�1��j�Ý�iwO�&3���Hׂ�4�}h�z ���(���,�AG��^�u��F�y��>Z���7��ˉ����e��F�g�`.n�"�ѤaCz����v�e�C�`j�N��KT�0#��{�rOݨ�KZ6&�H��Κ~�.<p�7���;�4ٽ'�p��Q�".���u�� 62x99(E��j�<��,{��Ѓw��h�(=�
m�`�2V�6L�~�!�/�*�m�x�|pc�������>���i�u��hH^�r��zho�H��Tw`cU�A.�v=�5��_%J����`����B���L�Q�kQV&��YܭaB����~p�G�FY��o�k�/hV�rͮ	�E�*>YHAj� V��23�$�AS#\ y�#�Ld��,�k5��-��.�~�c:.P>G���/�^8�f>o���L��q���hkd��{�a���(K�Z�m�g�=�k�K>�4�pN��O:!T߲�:ګ��<S���io��JT��M
͸�ܹ����W�<���Kj*VꚐ�mK	�,�F���Q��`a4�[*z�Ŷ��\��ex,���+�8`�1���y)���"��Ŏ�mPѐ�K6�n!�S�|����R�`?�܄C5��|[G3
hd��g*}6���2��R��菾�h�`��lL��6���U�&���6Layh��Z{�Q�W�p+�i�$�����4{9������X�!���u�D1�iED
<��ּ1����L�1�KN���$y���8T/ԯ�!J]����iu�=�xzx��N6�LY=���<�bv��|-~d.V�M{��.4�r�L����̪��j"�wȽ)���y���v�._��]���9;�1�#~W_fӖ���q����s`ذ��V�Jd�1��'��
%��5���z�Wd>s���id��y$8 P�Ҵ�[ȎS��2TK�r����3��,�}J:����AV�,��}���Ժ��s�h#�_{5��C����˷]�4j�mB�J�hz��,�DE1��L�|�}��Ֆ��H�C�3�Ӆ����S�瞵�z=���J����q�M���p�l�G}x钘ӖN �uL��\�<��0ر��G�^3V(�s?;I��]���b2P�,�8��Y�1\9ώ�9��*�����<�H�m���D[.��Q� "̕��S�4��2I�@Uoz>�\.�ɠ�9g9��_�(:^O�6^D�/��a�ɩ}���b',x���Y��q̺�k�͗i�D$g�[g,R�6��o��[�?���0vT���F���^�>1����,���V�R��i�0�x��u/�֍��e+�E��Dl��C�jD��
:�)]j9��	�a^�t��<�D/+b��V�������[:�Rʷ��=���T�w��c��jń���s�v��2�<�VMMO�����B������Q��x�#(h�_���*=�PK�TG K��>sl ������]�-i�R�n�6r����e)��Vv%1d�BѦW�G�ݍ㊹Z�KJ�=�MDؔ������`]���nj�I!4�J�	���f�����a�Ý�<�M�#ѕ�v(o#0H�g/R`e��T�e��(88�_=�R��b��`�]<�qi�A�-�����l�Q������k��݊w3->��9��׺�����[E�W�sƐb{gf���D/��65}T��2��%�-t�P��c���H���D��QD&���
>J�L��km�Uǚ������W"��������:�	�Ƞu:���|0��$�RT*C�-5NRy�&A�5�@	�"gH�4(^cg����2���^{M��4�
��7^e�C��>}׀�ҫ0x�Nb#`*ݬlC�S��,"�I��h��$I���V��������ޜy�$
���n7Cz��Jh�?K�3�
i{@;�^]�� a������r���+n>+_:���6��m(��n�\DT1�rR�APX/J�fZWm�Lg��BOڱ�}+�R5s�r@��3��^y��U�24����\����-�Y��0�~ч����$.3
�� $�߃#e�����(�h;��GF�meӿ���6��p��Ȇ���[ȹ�$�%)$g�R:A>�s b�b>ד\%n2���h���R�vL���^���c�l���2ΖƄ�������	Xj.�p	�v4��5���N��%Q�~ H���߷�ەm-�T�dI+�yb?c���v^|�+�"4����t`��iq����v!s��S����}�����\�?W]��(;'��ѹ��m~��)��q��ee:<�P�Ę\�f�r���mI����R�+rsDFT�C:�4����ϒ�\�^���R�k����\P�%j�����Y'�+�ޜ�$���݂B��!A$�����Ǿ?*�-��(8����?��F��s�VD��K�)����?2��+[NY�:�s��P�d���9�y�wͦ�G�<'_�L �����TOJ,Z.��ZBڂG�$T��&�M���Zqb�:U��ME8�S(@��`?c���$��*5����eA���7 �_1��v���Ҩc3ɫ�P�*��OK� X�l����s MO0�F!W��߱I�	U���K�V�UjY_��Q����\ce��3	Հ�D��qb++�t�4�|(NS1^c�?-���aTn=h���M!m�Ŧ�ƻ�/e�j%��z�c�fH��t2��Ga.�n��ajI.���<�Vd<e��hߌ�A��	{h$����#���_��]�qxMڮbPM�� �r���[d��9��i!�o=�N�KE�S��XuPP�_겜?	 K�|H»�0��!8���p��#��nW�5���s�������(ӕ<��z��y�9̵����ٸs/�0��:�~M�R���.�c�у*	��S��J����^%w�4��@���� n��jy�_;D��k�L��"]�$���(��B��[T���:sD����(�]�ɉx������i�(�n�o9�H*����� �{�"aPp���j�jN��jE��Y���U�
�YG����+�'�T/�D��B�=t�z�zFR�g��Ci,q�X��)�\�����y�h�h~u�����	֘�8���ι.�Hk�#��ȣ+%R	]� ݸ,�����-��r��xձ�:۟�κ/0�R�ɟ|2���O�г�9�^C�Ɋ}�s,�;��{�D��μ��4tr�(�4��8kΙ:%����ŧOw�����$��N
�͏ov��aM��>OiCBF���U����L�㣬#5��̫����\(�	*�:'u֢���^mB
b��F��l��j^����$��SPO�
�C7�Geb����X��;i�� �-0��w٣��5b�E2��c�4���YI��t�,�h�P��_U\(ԑ
�� ��y	d��k�H�o�I�gn�.��|�0�I�Z�H���R�g6�� Z�p�2=
�� 0���ފ]|´�_��I�gvȫ���c����;囦,�Q��R�pS>���I��X%�y��D��0'̒�e�i�ɢ��Sfs�i �ҩ�������������n���|	�71y�D��ʗ_ ��B�y$��:Y���]$��q��Ye;����hL�eA��g~�|uŁ��b9K�E�F�Q����L~5�����HX�2��7n�t�h����8s��5�H7ڻ5��|���m�|s(�h���5IQ<��S�s����JoL|.
��W2o�Z�l��Ȃ���m���LO,����d4ό�6x�S>����le,�JK|�k��k�1���/�C��^����]�v�5~Ns�l���G
A~-'��}���C'p�D�6�����[`�'�����Ĳ�j�z��)��B���O�/��_��D	ߚ�1�4�R��X�����X+S��,_�t㚅ØS1($ax��OD��`�kEJO�*#zB��\D��2�7�EU��u���D$����;3�6X���7���q��	�<����N����w�^�mh�Z�*�ߒ���My�uCSV�9�ms�{�pu|�
���6jCt��a�	�7o�G��TĮ�K��� ���{�V,�Mܒo큈��m�<$4�����3Cf���\�1��|i-N?i�����m�?͔�2��O���]��@:vP7��+K᪊P�G���
j��Ŭ��5���;q>DI�����Bm�ol �.��Rׅ,�Gr	��?��G81�%ճ��\����C��P��j�.f7LN��S�N�_;x߮w�������0��3�2�e�f�w��+�,�!|���vGv'�	�\�b��Ձ��QC��N�8hG�sac�����DC5��Raz8��oQ���	�w�����۪
�(�vӝ����H�"�D���-��Z�5`��X�=l՜�?{{�L������v�ѯ6ڍ��z�Ff �C�FF��(�W��W(�Ӆ���\�h(�7�K��Y!bDa��(�̇��ux���p?��SP�jN����QN��L��r��;w���|�缝3�w�UJ5��]��-Gc�C3��	^p(ѐ�J�<�����H�Ӗ�]M	>��D�yZa��X{pp��?yn��W�L����-j<y(�����iv�z��`��(@��y���e)��v� /y�a} Ӆe���!���Xӆ���!�T���9 >�Z���;��=��(���~~��b T�|ס�����:�"���Яf�՞;R�I��Fv���+��+q͖��3:����c�d2t���%6���#�h^��G�d�����0,�}7�3xdE������+1ΏM[�ED]AEx5#���q��x�S���z�����!Ƙ�����n�z��>�ZQ���+�	��_�s��.ݑ�-B�c���e�����Թ�A����q.��������L��>�9z��`k��f���JT���k��vԿ]F�=c�n!^� �ż�z`}=�|%�L�f7����]ڣ`����I�{�+�k�-�wE�_���:�~��(G����K�������>z�O�:��O��3�lՓ!8��%�f_-����eeF�Y��.7�4�H�l�TJ�+�U?{ �Q�Q�.��O���й���d[�5��m9�[���8T{�Eb�-lЁ��¤�����A��t'x�)KMA��R��u!���
�(��%���p�����!�����u��u�@0? �'�Im%����vJ��HlN�ʰ�*�k�����Q�� `��{ET��*i����� a����F�i �c���fV����c	S�̭t�	�hM�\�r���P�15L�e�`�C�s������!%*���{�����NP�S�z����u3��Mz�-B��"���̲)�	�#\fi�������ð*n]��dUS�F PD�����pM�j:�9�[�������%��qX��[@�r�!0bra�'ޢvc�az�It(����Ɠ�:c(���X]>zp�A�Hu��Tj,�J��|U�,�q�*��+�Z_z�y�#�^_IlTM��
aj�M�,�������4kE]N�(SQӎj=U�["2��o�:)ɾ���Z#U>����C��*������	�E�=�\�E���>��c���7n�ki�[�� ����M5����ǅB�ؒб+�Hn	���əwI�~En��0D5i���@F��A�:�;�����e��h>uK���{E��9��Z�q-��/���D#Z��F�)k�4"3���<uSJ\��N�p4U������o���l��j6._�0)�܍p��8uE�f�4dFv �*�RTՍ��@���_j#�� �Hɣ�������1FZ^TKM�.�9��l�z�E�Q`�Q¤�L�Q����FH�	�U��a��B��G��;hmA,�#��}Ґ���P(��ӽ��(=�ԉ����]��U����rQ�nY�%����Z�"���_��D��կJK�	v�x��Y������K��2���!�$�������dx=�ӴX�d��t���Զ��Gj�t}�/����RY1�GE�*�na��F:9�A�8�RQ���$+1�ց���2�9����svh�[h9�O4�͆� �H�hF�e,q�-�g7$"9
�T�8f�fep\3�(�q2/՛�4;�edV�IGTs�N�5�M�>�EWB����|;�����V����zM]lä�����n�O�DQ ��:��';�;p�?�4�cs,�Q�^�ޒ���} P��&I�}����pn�n>�����}�KȚ�|��m�:7R�Bp��Y�|-�炠��Ee?�U�|�!�L,���^k�șB�X�|Y�|E�B�V�����6Fp`�ʠ�R{����1�]� )��١{�������D��kbG�P�Q������f�n5��H2&  ��Eyw1��\t����X �/�,m�ŕ��*>�畁*̐;^P����@y��<�+}���j��"�n�w�0rX	
�N��&���Q㌊G;�]�Ĉ��oU��D㈛.v~�C�����K'��Fk2Hx�ؑ�lh� ����E�4c%`�#@&��2�v�<{o�ޅ���ͷ@�3��Yp*�׷aI�M�Iι����8���?[b��:�!nB"�|O�/E!��w����MI�:[*���n�QIf;�z�wyUۼs���B�[���q|�䡵��B��_�_��*(o�;���M��n8��^W��<�C�	�<�))�^?&R�Ш�3��b��W�U�$Bi�S�E�H�F�ջ��S�G!&h�~�>&Ա��@�t��}T����Q�]�C�nֳd�c�j2~�WE5��;�Lr�H �g��3ٹ����zD@�A��M[);�X����Oq���n��w��>Z��7� ��Io�bGh���%0'P�v���z@�.�f�0w2m��b��8�����K1t�C̫�+`��$/w'�`s��ՅF�K��?0XčWW~!7�Tk�^�@j�n����-N�c��	/�Hk��z��K��0���
�!)��C���#�9�XLE�9w���c�����w(���v�� BG�)}=�e��]H��P��H��ه����I�"�8"��#���N�7Z��࿙�o��P/��)��h�����}]���c���O�������(.~��r���~a�G$�%�����\+W��!�tq��{P�J�q��wM��՗Z�t쯟��A$�W웦��]���X��>�("��u�K1W�1Y���$$���Sq���y��r����X���Y3���I�"3K�!��dMan��}Ё�S�ND^����״��c�C|�ݺ��՜~�U���|���;�E[N���R\���Um��_?ߴH�/��qIz���[��G~Ϝ�}t^�1���|�a��j��c�E�#)h�W�:CNF`v{*�잀a�����?�<���$��w��^f�L`Q &����1���i"�w[mT��$�ɤؙw�F���<�v�*Q���e��#&=�X����ڛh}�� :���\�?���R뀢���Ee�8�]�ܛ�M;D;.���Z��ָ�}G�S��Ch諊˓�ܘ
�?��K��(@Q���\�d�Lo�O�ͫM/�>-0�&��1���o��L)⃿]�{����>W%GW����5,	&k�2�2N�D�_�ʅ������/���-	��(���eT��0��M�B΢5��eN$-D�)Bu����:�;�l�{	�$Mi%qH��?���?h��a�i �;��\�`Mtͦ��H�2ɮ�3|���2�G}����6��.:C��ѤTR�v�<����7V&�z*���f�/�� �5Y(��7z?vc�*�8��=-���ep>՘B�.IE�Q9CP�����E*�M;� ���%^r�����k����H{>���3��bG�+����DH�`{P�X�C�>,���5˛���Z�q#�FlsW
���Q>����L���1��~�+�S�,ͭo��Օ	�Ղ�����!J��Ο�J2�(3�`��ב�6�&N���k��{f�!�'�FMV�,�'t��	��lv��mس�6����Gx�eV�/�*G�D'q�J�B[�^n �9�|����c㹱<�H����&��R�d"7W["�i�{g�x�:��R+tz�]��RO�ȣ�n� x#G��۲ix�t�)l&�72�l���98�2�!0��6��������Q!U��~s�G��;L:�Q���/4�����\	����eL�0�|��T�S��+D�Ɉ��A74T�Ջ�jٝ7I�"�2"����w��{��;p�Kj}�(�P���Q"XNٙu��MGw"r�l�����&�/��"�wC����|@�4��s{���ȟ��OX�UG��&I��I�-����x�ո;�~�Q��9D�d��?�J����X3�G�4�ܼ���#w�Y��:�B}2
ɔ��5����С�/(�^�C
c�Q�4��ۆ�c|�W�Ǎ�M�G׏d���e��H��2��$����[#������.�Vr����G2����R��	cG�2�Vb���SW���sq"�q<���r;
7(��.fVO+1?�J?��١S7� �>�ھ>�Ӭ�Q�ؗ��$�m����E�Ok��0�Ȱ'� L��Òl����^@t�$n��Ie��+���}�M|�!J��I�1��G�}�Ғ�գ�jW�T��j )��	z�Ύ��W	�Qnp�3�ڛv��~:{d#����݇B�[c�7��`+|�����e��O�j�) ��3� �B�R����߬���j~�a��?\�s��[9_A����`Qa3`�|�U�Nq��L��Ч L	��1�W����A8LT�o/�Vb&�Jo��&�%�J\7ؤJj�<3�R��o�< 8����d����^���W4��O�Ŷ0J$6& -f���+�ݣ�G���UPS���v��z[{���rPd�����t7���(��ޓ�*�z�TL��=��>9.pF�į���=f�U���V�1M��y�m�w>��d+>��w��{�:�L�u/c�|�m��|~^�Z�i�b�s�z�8{j7<N	"�&������P�b'���#�S	�bj7����w�_ߋ-ޯ�a�Θr7�ӗ�K�A�;a����U�Σ���n҇�E�}�=�1��b)�6e3Ua�z SO��b�0%E����ߞ��
��C�k]��@'�פ�[�Qm���_�p���z"��#-�Y �f�-e�� �z4�z�}/z�lv�Q���� #
[8���G-N�Ww���3��j?tS�U��
}e�
��j�(��$X/��Ҋ���F� �P��[��#|��6��'t���1�3�j#�$oǩՄ\B�Ä�v��`A�Ʌ��� @�5�Ҟ�A���~q���!c���i��}�C�4s%k�븗�%2~��'��L�p�����=#�pM�4��\Vk��#�k���g�w�����1��J�������@�HS>I�Z�	3G �b��- i��"�����e�)r�b!����3,��mҀJ�U2?�\�þ.�ݻ�K��v���e��W�5t:�T���B��_�39|���4����tb��\ʩu�=�G�c���Fb�1�5�(;EN���ZN����ق�Q�Ԇ�M�l_#��~��'�̼3�|r�^ⱓ��:O�<��X~����}�z��UJ�T��ó�qr1��n�; �S@��)�l
�\I�x�K��n�c��D50�Ǥ`)_�-}g\�T�N�E��;̠M�]���o��!��Z�3�R��mE�����L�&R��;�[�o��m�U�dNbcn���I�������?Q�2OCOd*������Η���f�����I�Ĵ���T(�;��l��.�n���ې�1K�|�8Moi���6Z��4Nu�K�\KLS��GC�$3S�8E��%uf$7 ?��RG�eƊ�|���6T��]Z�.Ҟ�����ɔ&	�2�@@&�+�'�A?�u}=��V� �ո��m �a���&��'�Q��#�̆��28x�U�;b�3�����YO貁X��S7r�k6TH
-y����̫v��`�����%>P�6lvw����!g��4,���n�`58���@6��ż��M���~�\>}�GG�89� ��b)O\��&*���/�G�t1���tf���p�o
/S��Bc��L�'�J	��~�8C�h���|�_���&�C�:f�������G�g��hSKUJ�LpF)؃0���86fV��G�K�{^�~�*CW�~�T�m2��+d���d�W)���u}����D�� {R5�J�=�*��y�wь�F?��)T�:��e|��[��:t(��a�	�^�r�Dj�ca/��H�M\7"F��7�E�:S�ȷ=�����#�AT�.��)������ƶ�_niI��1�%��H�,���Y�r���3H�v�
J����R���g,�[�`�-�Mp�4�[J���֜]��yTP��:�Ϣq���},�'�k1�!��j,v���g�ބ���χ4A�����B$'���V���b�-��ۇ(~	"X��c�q��=�m�و���;�6��hnҏ� H�5�9B�b>�/����b/��� �<-� �ha�V���2�+J�[�uS�����{���j�]aF�oĒ�H��vzi�i�!:��)�6�{��~J�am�@T�%��=���;d�B�a�P�r�,Ï_0|�]n�+t���b��=5��ow�_�Zx�_
-�Ao�P�p�Gm�&�p�=OOjۊ^�k���_i��kK�6��� iܩ��N-���5�_%�/̋+r�����h�\�\A7�E?)�y��g��?[����-/\/��F�u|���d�n��?�����6B\��g��8sZ-ɹ�9y�G^��.o?&D�b�Ʈ���z�E�]��q�����(�t�,��������h?~��@�y��G߆�[�ӽ��x��]yh��_L��9�0���؎�ٺZ5F�j-Nko�Z��q�I��a�4�v�@
�lu�w\���������|X��/x!s�����ٓ9��c
���՟� �&�,n�l�D�������K��<u1�R�r���X���䆕�-Rh�8�k#�q��b{�y�W�Ĳ,���C�����鋨C�}_��9-���}PL�ty����Gyj��<�rC�K.,��d;eM]{�S�rYCJ�J���/:���G��9[�MVWq-�St�M)P�{�<���3E��H����i]�j�mU���_R�����M�ܰ
:2�b1��I�u����*��8)Iی�0_�J�[N������ ��i
.�UC.j�2�@��b�w���T���
C8@]x`e��Z� 	�gb�dt�P7YB=�Qƒбy������6�=��l�,����.Br��Éh�����SB�D��2c��w9��m�H/%��MF�k0�E'�,0�B�
y�x�/98
Sw�	�9S�����>�ʏ�`�B
�J��"Os]=.t9�9�d�U�Њ���	��W�[�,*UA<v�xe��6F_\YW���g.҃)���KD��$z�F��ܿ}�^�'��p�Aֶĥf Çz\Q̈́l�&�&������E�vu]�jH2+ԓƏ�����Aj;$��O�%�\�w���\>q��J�Q3��\]I�M0�#n�3�rXZ.�$��Tor&�&],�T��������̷:�m��������%/��b�����s�t,���ԏ�S|��h�雓]�ȥ����t�7�_�}k8�ӆ�tz}4}{����TYUd �T���n77�1�1�ꐵ�,+��;-��N�4nk�0�|v=�;U���:LAta��m?��	��4��X����9m-�>w!����v*����T>�E�t��I[����r+/�E���� _	�'�u����WюP��η��9�y�M�F���<��V��E�|.��q���#�lUy����H�����p�B�:�����-;߂gs5�����k"��j�g�#Gﴒ cŻ��F=>6P�ȝI�T�pF�W��kVCh���QrœLV5-~!C�kC4{�wJ��st�3�BS8�c2����ƏV3a�G�)�CK ]�M>��wm�Q.*{ �.7���R�3��up=K�/���� v�6�˫�i�ߑ��`9�p�{��Ą��"�4�5�d�����8����o��Px�1NU^jpn?�Q,�� ����P��P���	��@���Ƣ|�7�Q�G��Nِ��0N���}l!���h��t��<�6�@7�����"w�yN�$��T�nx!�G̋4M>aC'�<�_W�n_S�������fL�U���B0��*�GH��#M�s8�_�&9�g5��J
ٔb�7m�R���PE-ɢ��5�&^s^���N��7�� "�)���gg�����ҽXL���=���bg.>O�� U�%= 	Z����5<�L�?P֓�Iη�w :٢>��9���������+�zxW2�1�%r;B�:����U2����冒�.�u��r����8&Y=���#�k;��o��M:aSH���gЧ�iY��v��VѢNJ�	�&'�An�1�2�`Y��d�6gR�޵�9���9Η��7e<	eӓ8(~�mi'�9Gؑ���,#<Z#���q�� �?V"4إ&йQ2O���m{�m��R���̯`��S;���i�Ad���Ay� xշ��6� E*'�p�#~]-��*:ǝ���z\�BU>��u]�W 酭�9$е��)U��<ṉm�a��@4k��LF��m)�m�P_U%	
�F���⻅'|;L&k�'[������i�ET������:j����� G`�K�YXw�ì���3�Y�4H����׮��[���= ���
�]���Ck	.�����"r�3$D\��"	%r��z��5����h+4�{+6�߰���Hfd�Üqr{mmѳF�����W����]]�#i��/LOs�dR���e��Ke�逎�>��悹Œ�6��^<�p�xЁ����_}�S\Z0��O����~y|_��0���ƹ��Eq�hK~���P]H�0dh�Lv���ΖUئ��0�J�����ϴ|��_F���8�چ��
��D���)���Ya�:��̼�Q*-<�;��K��{�w_poB<�*h�)�"N>Qe�-H�k�;A(��9<��ædj�Cz썰�h���"}�0Ԙ�&R�lx���V�E�0@"S@;Q��Ϻ�.�eT�Ԛ�f��̓�5v��8�ǅ�$��Y'��V�[��G��k��L�A��;S4;��E�o�In14�v�m������^��u�^`�x�ʛ���g�
W���)�F�	����OmhV����͙�%(1�t�vS/o���@�wQ�ql4x\z�����<��E���73󎳣+,~&��+S{^'r�i2�y���o`�Ȅ��&Jy��̽��	����my�[rA�w��`���*�-s��&��uR~ǌgf��Ҳ����;�U��J��i^,���禼i#j	������v�?1]�I��~���,#�Ǳ\RBn�o3$O��Nrc[�VZlCPsnA�ߨ������\���4�V�"}+����XP���#!�%o�Mth��S)�b�VS�P�_%�);!t�����7nO ��B��� �����S�s�v��t��"�р�E���~y4wg	
4[�hX�E��#�%6�me�rߪr�C��#l�%�?g��CY���
��X�����t��!}.��6��j���W��8!*BM�tԦ�E%q��]EˆG�]	x�2�ʚLɡ��b�x�����
�>���������.�wȲ/�D=B�w��4��w�0���z��Tܧ3��6�����L��z�#S�������R��zmS��f���H8(��"��x6Q�H��[ӽnۓa.z����m��NW^�K��2%�� V�6{��O��4�@�o`�)����[)�O=��M�� ��.L�� �D;Y� ;hs��-�X�/�t�z+�����;/~1�wmS�@kk+����mZσ�;r���'��Sa,��-�#{����L�k�?��3wy�9i��\�)}r�j�6����c
'9��}.i�QF�X��{&Βl�>��  ���p+��L|��(����q���a�˙I�}���Pyց��	��Pw�
Y�[�hɴf�ι�I�A�,��$6��+� 8��V������p�$��3ɖ�S�	���\v�x��z����h.+�'��Y�k׭��؏����X�IP�#=t���WT}ǋ���Bai�3����^�A��0<Tq�36���Y�!�w�b��q��Q<I���=$]%��4'���D1�����3g��v�kJf=F�Ai,�^	�z��:u%�4�Mf�Y��2vd����+!U{Uc�M"�$F��D��qYB�姶��E��,��r�E�+����[x�U�$6<��T�G���RH N�����,���s3� T(O�Ǘ���?�٨��ޒ��n.���� �ϗ�̀T\SG���M�s�`��~f����x��J@�_��BP�m_m�^]-Z���}<�J��֣�K�g~��g�0.���`P��X����P�885q���g�RyE��m��x�kz�5f�38sߦH�!5�AY����Bs���D���Pќ��K�y�Oh5�OP����� O�H�aw�ۥF���Qd�uæ�oG��L�;sO*��z0{�������Z�J�cȄ���C�W�h���F��2|G��u��v���ƹU"��~�σ�&��81���lnO��!:�-*��KnҎY��c�j!U��� �]��N�?t���lfs�x?��jx3��!�Q���M�J�����)����<�\٭�W��z�z���B�H�pO��P�+_��oG���-��#1�JP��VUe��{A �R��A���Y��ศt�G4�� ��1����0sJ��x�mcVR�����������ƛ0���Dq�g���v��g��۞3�帟j����}
���7.�K#Q�J�<+_�����u|Ԓ[n��a��LC$�R2�� �-�'��R��u�\j�w	��������i���5���!��$l�9*<Ō���g��h�'�f�ғ�t���@�5e*U'W�U��l;���B�3s��r������5��&�ᒵ���/�kR�b����;�L �M��O�U��l�e~�W*0!��<�Jj���ϫ8}�
5��ð�Ъ(��OX�1%WL��S׉_om�/�r�b�^CgA̩%�a����Y=/Ʌ�������>�q��p���9�-fAm��x���xe=�F�Rk@����4�kti�3��>�O_	LH�s!-�'g��8_���a��â�������mJ�W$�^��S��W��=cv�E�J���q�1�UA%D���[;���P?d?��kQ��F��}�O�����t�#���V\p���;O?����Q�"]~I�l+��f(;���<�_'��y,e>�Y�����f�.c�^䯄1��]�������u2>�efT(�3�acv�����'���f��f����p�Y�?�;��T�i�9�����W���t!_@�-%����9c����F�m�x�%��G�-�~8�m��<xy�/�&@�Yg=Ā�1��|g���ZX���l�{J�q(�
���)��x��FC5���L�F��o x�땎�}�:�k!��R��qKs���]'��!)�t�ڄ��6fC�����}�������O����V�������^��k��� �B�Y�V���T��*Q�G��E}��V�rj�&5�^��NJGH���v%#c���ބ�oS!�CZ98P�X�n.�i8���5ܛ*j����/��FE�E�Y��ʊzg0G˽�$�![��`%7�6������:~~�#���/�����*`�T�� k�����eq��A\ ��B�}��gy(��Q�/S�G�é�<��_�h��RP��Ӽ�����'8�l�� x�>�w��O-\.7ʯ�����ӗm�{��W)�[*�9���V�AIBv|q���`��W�6�`O3�$���>3����Ƣ���M�
0�����+�b``3,x�VX��z>Ñj�r;��ݪ𞛅�u�s�[r򈿴Q�!���.�`U6\8�2�q�0�Dب|�f��dO�%B|x�,�	�Q\B�eŦ���'��ec-ϑpII����\�+����V\+A4���(̦���'�4�jgrc��\�o���S�
b���{+��]Q�Im�����`�;��]���B�p�Y��4�WSc���l��$9Y�z�>�u�YsKT!�9{�1U���L(��� ���5ʯ��Yc"�xA��jevN�*0��^�$� ��R�W�5U*"98ٞZR�0��_�Ls����9�
-���<�j�"Q\3��k�x#X�}���U/��ĝ�jix&���צW�{ѠM*;Rp�1R�P�����E�0�R�Ε�XΨ�)�N�5��{A	%��>�(��RZغK�m���֣³K&GE*L��[��J��~}��3�$:փ�qP�*|r\Y�V���@�n�t��@�J@�"}R��¶�S� �o	%�IJs����-�q��③7g����[��>?�e�˄�j��T�Ҷ����\���Yy����gm(��������@�Xq&^����{���NÈ�z�������HLXt�?������N�����߼(�d�����
��V*����ZC��!	�k�8ڰ$<��� buyw�h[��~.��Y<�+ZtZ�IP4�
�))QO�P�~TeG�H9QD����Q���2@�D���7����b���C���G�F�9b�%(�/����=_݃er� z�GA%��zJ '�9X�*r��-� R}E�� �tfS��6�_��b^�!���+�>f[lpL����$�sq��`�v�o�VS�ߓ���ԩ���v4�/����|��y!��ɹkW~� 0�_��҆��u�l�ǋ��*!`F0w@VpOxwU�Z�>��[�/x�W:j�;�р��vWw���E��P���. �������o��H��홬v�=�l�������0��<���_�d�je�8C#�.6���#�O�t��"B���8U�#Fݯ�d�`�h�J���|�NÇ����i�{�d��Y@������;�1$������-��M3��d�c:)&��UD9P�?�`;1+�"�I���ޝ���;�㏮�{��X ��D�Z��T��1�ɁQ���Jb)5�o���(V��I����i��x׶g���M���e�i�U��X{qҠ�=�r��+ГG�t1�w������f�X�J���.y;�u�(2�<Y�v�_i�l�E�n'5)yć��j�Km]��7*9�q� �����(ߦ�����~39cu��=?]9N�GJ��KS��o����y.tw*�rG�;s�N.V~��ީc�������t�U�uy��w��Ǖ�L�1�<ȟ ٝ��Wx ՍU���s*ʹ�š�p�͸�X��U.g�f���<���7[-3�~�Nd�r�Eƕ`9h�H.�u��P3�jQ�A���o��"B�S2�?�i�����y}����m��)�����}��<��N�"���g?L쯠j�Z,� !��<r�4R�V��Di�0؍
���5e���z�:�қB�w�/�����O �#i��g��E!�ٴ�4hh=�!7 ����^�����rI�$���#d�����1�__ )�vP|�@�F(@��<�Pl5�<T�J�d{�*RC�p��#ay����0��YNn}j~S
�"�F���JNx3�ؼ��|����P��������_Y���߷RR�	����xFg�*U�����ׇ��^ i=�r���>~^>��yS9g�6 �ɲ��Q�����U�0�6P��ǈc��/���1�	r=��3��� 
��$)<��^K��o�X#��k���w�����б�~R��
`ݳia^,܈��,�;��.�k��e���}7�		��$zVP*倗�Rr5��9s_�{������jȉK�!�YոOTi&{��k2���,���b�C�g6y0�e����h�lz��������R��	U��x�ޝ�0 �ۧ�0�~,%s�'�1�2� �d���Ԫ�+�9,��4�`����؋��������>Y�ʵgLiSl�hܑ���/b#�%?T�A�`��a.l�F�m�r�	�筮v�Hv��:����V�'G����
��G0>L�a�/�8�v�w& 6V���@>��Dd^	8�os���/��d
�$��YI�0�X=����¹����|�u󵅂b��cr�X��,t0�Qƞ,v����}�|4'Yu�쑪����'Y�^/�mA�Z���w��]����+�p^�%�& R�)"E��2�=�E���~r&s� 5���������<F�s�� vF�Њ[(yjn6y_1�.�3C�ңa@!y�N�`5#79���ڂ1<���p�7��v���T���7,�Hkv�p�l���=�гHD���DD�Ħ��G��#y^��<�}�~R;ŻCnh��7�7+������B�iwC�5�F|���S0�U4ĝOt�2j��	@@Z�{������"ɴ��N��WE��<I2)2¢R����9�}[x� ��J!�����jĿN�Lp�x0������M�l}L�šB:����t?��Yı�ɽÊ�$uc)��$��^��o�(Y�a���"�e���VH����|xj�>D��!��Y���#,.t
ު��د���7�]MϜ�G����pG��̢%q��xD�M�$�W�0Z�7��-n꫌fI��*�R!IDB���ν��v�w��I�1ə�[Gtg!��>B�9��p�w]���Q�`��n�Qt�]g�* ���(=_��DY��Pќ��8�����ҡ'��	��m����2"���,9Jư���ŵ�^`������3-D2v�ّb��mr� �]6�^��.�U;��՟���h���j�r$��9W��Z����[nN�o"2�cPv�%���ԛ#ٌʗ��4c�0�>ɂ={N\��/��W�<���C����C��2��xlJ�h ����c�#��`�C��/�p�@7���Qe�B�%����)�Y(��3E�g�����E�<P���M�`��2��$;h�����鋎���T�N����	�e{�c�w<znQ�	�Tݚ��`/PT�J�|�:r_E��0	
�"�6�K��pN%6���ܧ�:7�ș������[+�kd&en~Cd�4+H�-%" @Δ�4&��kϵw�&�#�ѰVq���d+�.	$���3��8v҂�(��q1�y��V���u|�n����DŎ�' 	+�j�v	��7$�-�[m��rO���^�n���QߩN�ooY���U]N����.��\,��w#����0
}�7��6)B[���.�$тZ��d��w��s�t��T��R�y��6�}���h%$z�Aj"u2����O�~b�BA���-�_T�f�BnD�D�&�����(��g�A�lv�����.��O�=��l���w�ѵ�+��I��Bԟ6�)�(�w&�f�[�(y�L��!T��P�[e-���* ��k���7�@�ﰨ�p2V�ֹ)&/�e�O%��t�K�@�"��¯ClU���K-�S�^��;���1����U ��7�B,8��_D:c��ч<-CMɹ�k�%���b���`oy�s�C�K;�3�=zF�L��*�h:����ͪMz���
�n����hB�Ð���F XhZ��^���M(wA�:�}R%��`���O��`�H:����/9�v�5@8^�Jqs�0�.Q�$���40�S.��@���w�n�=�g%�-�H��Z���ҳ�T���I�v�5u<X�۳6X2t�>p�,HO��·��V5Hf�JE�=9�
f��Q9�E(<"])(=90�}7��X��� ̫��~eW⋸5�/H�p�9m�<�ό_�F����\��l�ϝ�<�eA�����j�qiα���*#��`o�<�7{�B� v6���	E�Aͷ�e;X0��X��Y�ܨ[���8�T����{r�2Q�c�/ք0����W�����S��h4�~HAk��i�M쥘�Y{�[�����*��=���}��5 c7hq�0pl�{��A�@� �YC�s�ś�b��!�cla�����9H~��^PJ�B�G�@�w���aZv��u�s3�^\���RŒ��*X��-_Vy>R�AX�AL��_�}���~�m�\C����P�%����Exr{�3p@tf˰�W��Ev���ѡ-$�ZN������g�Aq��� �.#������׻�YD�e�E���C�'^h�U.��(ͣ�rԒ�bSJ���sLI��,c�	U���M]��'G�)��θ%���RP�=�	h�V*^���I]@Δp(����߃W�w0Hر�4�K.0<[���C�����j�r=8�%8ZuΜ�6�9{�se]�f�*2^o>��
�}��ѻB+Σ��g�2B(��k4����l!���"Z��vCt7�,���YfM����l0��^��e�;�}>J�Ւ��W�ʨ����Oq��`Ս
H1����)Qf]#��n�˧	v��m���6����,�*��N��K��K���w#9�r���[
,��%�k��w5�3�J��E�7�R����AJ�]z3� ������/p��e��c:�S�T�Rv�� ul����P4L����;!:Ҫ#�o�:0_�Lũ�({!�-�<�	�^I��� H�*�t�	i�y�],���u���~�{m玜3����ID�Hz��8Е����Q�C���*�>�,�Lǥ�?��$�S]�=�;���5R"b��n�-RP�Ķ��K�!�yV�du8��*9#p�ck�&mk�#K͸>����� x��M��2o�E�ܺ�#��^�]
��G��U]ױ�e�?s�Tw�-a�/3[ǈ������6VC�R�<?�8�PO��-Ƽ�G�8?x~LXԯF�6M�ح�����������E
�B���5�G�	6�P�"��2�p���bT�o�{E���b��S>��@x?h��}AE�Ҹ-�:�ٍZb���TZ�p�q�d;�Cш�n���(�l��c$�0���d&#�9.��n�n�e�vkə�7v]U����FZ-r݋�=�*��d F�_XB��bt$�:$]�EE�j�x���g��ʝ��P~X$o�<�+�рq�j�>���Ȗ�n+�� ��&� `�?g�c<-�Pu��.�@����nN� �<�c&K��	��L��
����_=�6���u�#��&n���\d�x�����/$5`�z�E,ކ�3��?.0�W$��نM�XU]��g@c���~��[j2�3�sy(�Q w^�Vk�`j;a�ԑ�N�H�cb�� gn�B����>��rs����v�Z@���0���t�%@��Ea��s�Il>��|�6
$�����X�%+}��5�X5�۲��c�J#��":�>`�*xo�������U��}��wP�J�ވ���=7��g~��I�L�GM^|u���b6�ќ4��Ї�|��1����8�����d$�3fr����\�#��(�}{4PfB"Mc�����*	b)���/Y���<c�tɯa��C���J�;��a�V�'�3�C��-K��?omĸV�dtq�4��F����j*��lN�u�-9팓�}p�a+� =��з�]�"��Q��9��)����	g��N3���ذoՊ��Ue\�8�p�{��-�c'��I�Z'a�a�`�e��\��)�(KN����6��w�f�;+$o�YѬ��a�uo�{L㐗�
79O�g@<����3B��ڠ��aY���Wd@..�����qz�>�d��1b��'�戦M+�z���"'iu���JǵZS0�>�ɛ��&���D*�X�;��kO���;��C����Q���S��VX4B	�?^��@��_��9���f�1 ��x1�N9k��ŭ��y����4P��r��d����� bAacb�&����
Ai�����X�s�d���y�V��4��Y�g1D��S��qyC�ݾ?a|:쳀���z�� �{�K^+S%�k�VS�Ԃ�w}��_�iV��X)i���T����0�
	
`��pA��d;G���T��&4ԯ���P����rcFB{�:���F��}u�}쪰�W��F�i�!�e0����r"��o�&����G�w�^@�v/R�3�"N8�ޜ$t���{?�3�g�Z����ȧ��f�����[���Ê �y!Ö�Z��C^�����<Ϋ�h;˷���-�z�E��vJ�mئ议�+=��=��e�x�s#���W�=&���(<�������=�D���sHp?�����C�1��dߞ��p�V'��g;+�*�F����l��gfM�GS_��i5���!G��!���S8�5<����8eZZf�ȫR�zW��P�$�����&�{,p��3�[�E#�#�cHD�ڲu���[h����f,ZIKZ��Z$N1Wu�O��E�r{ˑ�K#��1��v�±�8/����������u�������V�=��?��V��'͸<u*&��Ff�a�O����U��>n���af"0�#B��w$ӆ�
0����u���(�`g�H]WO���4�UK`_�eӵ�Kpr��:!� �[g���~�e{�������o���X�-Cw�6�v�������5��!t�4�G{�#�oչ;����`��m���9#b���$u�{����G' + 8d�&Yg���2������9�����(H
���N�)(d�O �S�)ʝm{I��4� �D�]�Ƙ�P�7K�ر�ѢǼ��P��pH�MZN��^�C�HM��v���~��3"L=.Ke�~D�z�|+����f��&�������j٬�N�H�vY�M��<��<]9���B��8�(���B�ۍ!޵eG?��"��[1H4��j+�3F�D�~׉���NΡ�}�ݙ�P���#�(!�2�($���x�`��Y�ҹ�I�f��n;<�l(�/�Ihxo��	�{��:?�r��$Nk�S�f���+���ikZ�c����
�E�y�4������
:i9����ýl�be#�l�i�f�q���R����n|OJ���[�+O1�3���(��&����D�*w?/�ǆ�vK�7  �-j"����?|�$���{�TRs�ʝ펳�N������>Uo�N�^�e4��bY:�KŘ�e:��Y
�)�(�%t��k�KB��oxB�Ԛ�5�B�5�%�Щr���t�j��0����A}���Xv[5I�Ճ�'6s�q�b3�'O`�n��~Hw4<:�>R�ۺnςn����R]�'O�n�w�!A$�F��ﴹ�MZ3�?���)3��72���3��Iu��~������,0PxV�6D�<l?po��
bD|�	�^����u����U��ޚ�.yt?C��U�WI��5� R�5z|�
�:����tgd�Ia�1!����3�g�M����E�O��� W��S�܁I�.�����C�ڪg�Д]�2��:7;�c2Y�1�6T�;���]9�`�>��-��ϩ�Ľ&�G���<��+O�^��,_�mj�ϡ?�=�P��u�j N�%-TZ�ǧ��sKe�j��8�>�%bh2y���#����jȋE��_��_j�~�L%�O������,���1��5�sW�t�YO���b�ٺ��e�)=�,��Aи�,�'�fk���z`��7*���R�So����<A��O�3/c;03_�?��h|���O���s�^0y�z��R"�cTA\�T��8)e9Wu�@� L�'yl��q����	��+Go2?[ń���b���ϥ�9y[�0��Ǵ����m�=O�."�<�$���]�_V��I;���Y��_5�ĔS1�
��P�-��2� �nȐ�2���{��&r����J�o gqD�PE���=<��CϹ_�$��+�ez�S�Z�T0�Eg86�W+�lҋ���?��a$��1���`� �j1�ڹ�4�{�8��~�wh�0�3$�UI>ܕ`��M#�:���1��E_������7~~)K��eu�&�x���=tn���u�v%4W�3N�^�����N:k��'�����=r�����I�].^�.��N�8�k�H�����."}�=��T+��I�X[	Sj�����l��h�}Ywu�qzR��ƺ<Gʑb�><�s	Юhzb�����n!�;�V�/r[y*;��g��q��7e�;��cˋ⊢ǯf�S\���{���tj�=������诱����#\
�!^�b�s�x���d�`��ï��_�k��O����ZգKW��h&��v2P�X�D�ޒr�_����|����fQ��d	�",,g�$A�2��0u���F�-��зUx�&��l�����w�\:e)���}�[A�tLR�A�7b���e��P��'����\��ŎY�E�f��p��1z�T�@2`�!$���9l�-�K2]��m�����7�i�����5À�u�0���s�	�Fu�߯�����1aא����v��N��`���b��� ��*�9,��U��ֆf�����#��o��poI
�d��fy��O*����Ӥ�M�o��GN�B�j�	�CJ�(�*>��Q}g��-��K:���w�R�@�,�ܹ�L�������3�1�,,S8�2�/��TfL��#�^g�"�7���qq;���V��@~a/>�5/��wC��KkB�v8�G��UǠM?��<�,�0ͯ��.1j:**rJ�c�-�^.y6�k�6)�;�]�*����m�
%!��9�~Mo0�M���I8(���$���0�,'�1��xe�mi��Q���sU<�(���τ٪�@�`$� �q?�k0��J�H����S$�f�K�X���ޜC�#7�h�茳#00˛��^�������E�HC(U��g��ZI�(�t�j�.��9�����jwX��e�n"�>c^������.�t��3�x�4eZ�x-��(��;@��7]
|�'�X
��N���S������g�/vW�����Y>š��0O������x;T���Y�Z$N���C�R{��~Y�E�uV��\	e�NkAe�]kP�]�O�7d3�4v�.T��:ц9n3kwF��c��yM^]~:� ��&L&�b�+L�4-�p�s��|������
k�`"��-���6 e��z7�G7��av.�6a`���[��*�̵+��>3�  �N@�(/�d�KŬ��*��Y����xY�����7���Ow���T�~�|-����l��Qr�T����y�0�٦7	l>�P�.mJ)���ͳ�B��1���ɛ��sl�m�y�/�SHՔ9kY\k�/�%Z%.�[aQ��?"?[5�������J�V�l,,�D�V=6����Т�[J,��D	>*���{0����Tp�pLB��5����,���Y�}��d(��)�z�2��j�y��@D;n�K�&!L�����y�f�P<N���pX�N
�)e�	s�@zY�@Rs�[�C���y✳��}�ų��eUb4��$��m����lU�}�^^@���)C������⃹(,�?)b֕l ˥j�:�>Ə�M�� 4�'�i*��=��[4朾�Bj��.1�[����X��OV������/�����z�tvfiM��U�S`/�"��2)�@�L��F��	�AlT�I�L<k˱�c�Ӛ�"�5�ڽk��޻�8������ZzE�8Z�����@ݕ��Aߛ�#�?+~s.����ۑ�)�f��Y�:c��h�*d�Wp�����Q��)��r��Gn�pU(&R��7@i7X%�i�1N;AZ`Z���H3�f�m�A2�L�x�!O��;߹���y���$̗�&�Z7l��R�d'È�JS`�&��\��f�*�s"	vհ�u,���Bt�,z$�]H�`��Z���/�ݑz���� ft��� C(�`�R�`��SN��2s\�a�*���.���t�k	��ש�M������9l�V��7l��*"[@�x���硃sWL�͙߾5�_#��I�lT������o}�KM7	U9�C�������lcr�pt$��Q�dkM�ϏØU�^�ǫR5�x:����Fws$��<��y���PHE8~���1;y`{p�����i�r<�+�0�~J�� �|"�u��R,� ��0����-�p�녣_����3�=e_�t��k��5x�v>&�t[^��TӉ'#����9��0&�l;D���j�p.a��f`��98NW}r��.���Z�����R��#J<��rC��ɸ�ec�s�KJ§��R�Q�s�w+��8'Cg��%ID Sh�↳�J5OX���*q��q�s�	Q�U����ihJZ�dpZ%m������9 ��y4jOc�^ͅ�N� +Zjf����i͸2��mٮ~�J��]�,�	8f��Ǌ�7�Ɵ��气qv{uԷ4�{>�gZ����������Gs����G�?���j�N���zDP���y��F�dUoS�`O�>��-70����Z�����'�v��v�fXKZ�C)�Et!��T��w����m�Hqޚ�����%m���L XL�@4�Xۦ�����	��������S����ȥ�F�qalqB�9����︛2�}o�4��C3�z/=��-�
��JRMD���Sf���J(�
8�OU�z=bۨ����
��R�e�:O}����T�>���s+��s�(�Θ�$�qa~n��>��hh�'q���\ۛ�1�'߈���L�mT�Ǹ��b�T����H��T�RpEQg���1ooO]v�"P�YZ�;�L������A >�vN�u��Wb�N�R�1/����_"�_��;n7>�'����d,:�k�ݵN`+n����cn�"8j��k�W\�S�#��#w��Aʯ���[c���]T���b����S��L�XK���~�����]���� �;�$�A�VQ��p�oܢGa��ؖ��@�����x{	�&��'�ߢƫѽ1�<�7X��{x<���S\1������nu��TD�kg�}�8!Uuf�ÿ�FP��8��꺢��$!Խj'�����N��,E�S��P��5���޺a4��w}<��^��>.}�� �R ��`"������O�I�ׂx�ڻ4�����!���@�ϕ`���i95���h��<N5g��R�sz�c�@���] ���Ks��زF_�<�`b���r,�b)Ǽ<t�[Q�i�nj�UL�)�=ޏ�FQ�?x�'��Bo���E-Sِ!�+�_Gk�$ݝȖ'�Y+�E�eܼ�V%��1��bq����h��Њ|{��������h���aU}�uvu_U�s�Fu��@�h�Ȅ���9q�h5��v�a�el~`dc\�E�G��-9��A�08��]�֬Ò@�Oc�1�a����`�1��~��U��1 }�f��w�ct	����=/����sҼ�@F8�|������)�/t0�Jls��cN�p�$r%+1̥�A2�x��H�9���w���%|���dk��hb��R�c��sX>�ї�q�!1�hk��u���x���x���wS_PV^��g����lĒ�WZ����#��)B��>���` $�[H^�Ϸ+Ï�s�Ȼ*}�L���3Z�u|������?����_H0�4e�|����3��P]�+�wd�����}�����^6�g7By���#B�rq%=f*��^���혬���T����B%e�_�q���o��`�s4}
��>���ڮ��|����q���斁���]���G���`%I��$���
�%^_��s����/�2h��_�́\�P8A�W�'=��q������B�{�@%�̦F�3�RO����>A2:x{�=�9�Z�ؿ�+����j�2�L�n̻�w��w��m��Z�q�\j�w�,�^+8dK��J9$K�w�FC%?�T�Q���23�B�f�؍(B��s���aJ��Ծ�D�z�Y�������*軷�=���N�ڶ�u��ک=-T"o���W�#ʳL��h �Y슊>T����U�`�D"�G���˔�fG�7��>^��Gd��> Wy�W�Q,�6/n�[�Dܠ��?���r���m�n��^D�:���8P��uO�߬E�U�Į�nTR�}�Q���Ǿbg�9d��:Y#���p�]WT8�c:#F�K4��o��h^�yOЧ���J�N֓�~�"�,{��T��!RY�U~�/�s���v�K-u�bӴd}z>�8���s�����(n�E˧�N;L,��G]�6khQ�I��A�Q_jXZ���ֽ���R!�?.��A�r�_�Mat�f@	Y��-&����>�]Ae�M�gJ��4?B�������bl��nU�<� ��B2w̓Ӹ�1]���:yb��X��;�©�������(�-1)�؟�N 3�H���$I�,���UO �V�1�X[�j��k�.�uz?����
���R0/Β��mNW6L$o˸���w;I�4��K�4~��rc�"��$A-�ܳ	R���	Nh`�	nb�y�'� ���{ ݿfP��\N`p�R�}g���Z��̘�:<P��W^���4�3;�}��)�˛k���J?~�B祈�	-� �)8����w��P��"���pÕ̹ĂdQd'�_�f��#1�������]�
[<CJ�;N&�Q�S���y�k�rU^�6�/�_nF�v���V=��V^�s�Z�goA< La	�B*a�8�K�� 3E�N3U�Y+�Q�̀�Ϫa��)��c�T$[H0� 3>�S�!Z�4D6>����b]���3���XS������a�G�>�,b�0�b�>�ۘ��aG�^���J�ܾ�"�(��4mz��L}=u��R���[�!z�_~)�d��:�#h�w�o�BiOh�E�â}[M��CB�)���u��� yy��IX;kY�H�},�9o
Fwu}N�o�10�� }DS�9>����P�	�	9;/,�-=���h��1�6>g?���������0B��"��ʥ�4a�k���se	g�W���o��b�G�(��`]�Ʊ�j�z�����g�d=/Y"7)h�.(���+�#ަK�`��_oeb�1����V�/	mu�I1yp���,"��1+�9ǯ<Ul��ip�����+��B����!c4gX8����c��?x0+������X�v}[ω=`�V�jA��#����GN1Iq�R��b�z����6D�5�=���mC!&��z�θǦ!���P�\U������(��0�V���=X����}έ���~��_ΐ�̲�#Fc��၊��$��󕱷����6-���D��� I�����Ƭ�WN��6kɧ��tY�����yXW���d���\e�M��T��7� �~�4-�U� D	���� 4��S�K�ү�!00�����U�e/xf֒3a����v.O�{,��<�5�y���G@*B1���s��,Aa��t~=fȦKda��n��-�є�xI�wD������ {I�.��^��o�d�~��S���5����R���K.z���P{A;24-E�o2�"A������ؗ�I=��H��w�υ�� ��FwhtӉ)Dz�`j������ٵ��2CD\R:�d-��x���Տ�~d�xR��|�<����c�=�!�y_3�<�R��"�>1�n^�I�֍�c�����*3�Β�R=�A���[��Ϛ7?C��3��a!)��S��Oz}z%�J&���F�����#���w���*,��K4���¿bK���ЩPݔ��b`�u� ��gH�lB��!~���t2m���?w��-C:~d����������t�-�b@g˽�i�Y��9hx<+97(F���J����r���h��ic-�Nዮ��Y㳎g����j��@��i]�EH�#,�t�,��F�\�Rv]]ϑ8�|���( �=�]��]�g@���t֩��X(�����_r =��T����$^T#�@" ���pD�Q��("�Hٞ�{�9I���ݥBX(WUCm	@�r�0�B}ZJ�� �~]�k�Un����l���E���
�|���*�P�4\�n��lܾ��`J�$��+�WY��"�L�HCd����Z�ba4��h�%`uT�]?������[�"#ljЀ�BK��-�p[sW������Z���mЊU�Kb�{U�K���a��tTuf��@D�p*��|��@e�@��%0y��a�49����+I��pAg�N���;{I�������6���\�K�	��t�]�pˑ�"'a�\J�4Qq��
M����H0R�HT���j�<�&$	,&�mW�lf�y!������-{�:F�-І�� �jMX�5�+Y!RC���ⶖp��0Um�AQ���(	��Ma�Y�5����|0��q�a	"���i���Wig�>�? ����`<��F���?]y��X?A� ��\/�@*aDV��:(��%�s��ǡ�*�����P���D��7�/�Ȱpc��ɧ[A��"Z�{Þ�b҉O޹P��Wx!���4le,��0�6r�Swgp��A�b��l,b;[!o�KX۽��"�qZU ��@���qSb[$���u9ޱ�0� pS佛��'��k�BO�W9N�0z��c%B�����<JU~2�֕xU���`j�bw�E�P�9�
�[{�>���i;V/� ��\Oo�h��V���!j�TDF��t)on[�i�zT���e� *���aG۫ P���B-*�-C[�$�</<���s�Bf�#]Y	Km qi.,b�ɭ�87��%"����i��4�_�^��1��%��$=�OdKǐfdNa@Z>i�Ls��($C�:�o�0<��I���-tQO�������do�8�B��d<A��W�+�ݑ��.�{F�V]�bd����Ij�d�����0N��,�����Z߃=��ƫ�9���\1&��v-�5,��T�)"#S�����9Њ�X&l� x���8�����o������3� �w���̈́��Ǟ���b�ZW8';���ws�ٮN翱�)�a���S���Ր���L�4&^X�3���{�^�S��L�,<%_�!%i��=�޾)�|Y�U��n-�|�@yiP�ڵ�Wz7���5?I��[��F����]R��1I�V�X�#� 8�a�ɯ�"�<�p���,<m"�|v��ƴٕ��ȉ�^�ï�\i�_3�	)a�|��j�z���q̒�޷*����!H Q��M���.e ��`�BP�5?,v�B��DK���+x�y���~a7��poȯkv���'%�Q�9z[v�V�Wڗ�ݕ��"�Ew�zl��Cq$Mk�yE���64�S��':Ձ�tnp��=MZP�be
���z�����r�4oLp�	�6XX��gˤ�H�^_.k��=V�Z=To5Y�ٹ�����:?j+v0zh�����=��{�d:<r��#m_[O c��jq�Xr���	��&����\�p��X�(�f9ee�bE{s�P
�avZ>����p��h%	,� d�5q� *��v{뚂Hݣ��_6�#1ytmesNl<���]����CF�%�fK �,л.��j����L،|��a~�qk۞�WNwys���tj:��ڿ#�	/���_vIw�.[`���䉐�?�8���͝��S�͊��I��%iǖd/��$�L\i*S��b�£�FM���g�<5f�I���#"s���WM�7`I.�"։�##;��@��uP�����;a��3A-Kbz�A6	�H��A�����%PʌUܝ�$�������2�V��T���0[?1�!�����9@�lS��gy,��Z:Ux5���p�\��qb�BU!���N������r�x���&�M���'���˖�|�7
j�%��7w���b7�}�~���dP��p��܅�c5 �;Y��7g��T�_��@a~�2��D���3� �iU�iH��q�b��DTR�1����H۹��O�8�yi�8�[WY�mZ�uB�x�%5�����6tr���	ڙ�*��GѼ��,�6Ϟ�~m�D��s�
�h;��b��)}����&UU��žIB�ݚ�Ģ��*���ʐo6J���Th,�{��%8�9��<���P�~~���Tt�x�R�[��w^1u�xX����B�`���Zr�8~04���U�U;�_]j�g�!<���{�0o[�Жbv ���܀���[�E�S���W�l5�!g�;up�!���S�n2��&��P	
���n��g����i�dj�+e�r�r���?�`n{��D˧��B���ovj}�T�i9������R͓aL�$7RʣDd ���smz?�g���X���Ν����k������e�|{u� ���1�ކz܏�y|�J�8��^Gv�:ߏ��^��<��̝�q�%c��1��z��^3����e�}�ۄz.�U�@5�"��f��)9g!Z1�XS�l�p���tb��ѣ}T�^8��؀Y��`����Ŵq�8� ��Sv��R"C�1�������������ۮa��\����$�ݨ�����"Ԅ�_��0ꬢ�FY;%�Φr�e W5���#ʉQP>�-�1	�iЧ���G�?��6>j�DT;�3yZ\�h�j�`��/����d:NB���sf�gw�);�t�w�H��v�� g���0�#ѵ�f�J�8�۱v��6'��Ou������O�&����m	���7#��tA7i0���kW�W��/�)7)�Yy��dor�	H�:�ߴ"+1vӁpET����������A�5T��%�O7�{;BL!މ
]�ʰ7�5��/��!�aſf��9R1j�!�`r�����P��T˶w8�{��Z q�>��� y�����NȚ��عd/yMA��,v�N���f��D4brFȱ;y��g%2������Aq\I��	�T+��_��o'(�8����?;{���]�os�UzL��3��x���0���K���Q����{E1
���p��m���a��\��3��˟oo���E# W�����
ux�A��������[���s�����ĠMf_�5��M>�K��J����Ala���˒�d��H�q1A3ݥ�;����3�d3�
�	�"@v-5c� |~�
�ț���اC�gvL�&U$��Y�F�m=����@�����h�B��=�B}V*J����A����.֮w��ԏ���Hs�C����<�Y��*���Z( &��3W�*�/e._qC<ԋGOw��CԹ�K�t}J��T`�r�����#�XM	�qc�V�;���=M�u|�Y���Ꮱ�@L��Tz��]��%��(۞jHf �TPs�3�|p���Wǂ�Q�����C�ÜA]Tb>ʖ��|3�&�ײ���E*g�=^0a3a#��u�?�	θ�[B�_S2��pO:��سx�[?T�ʞ����=Xj�V��zR/;�z+jD�K����S�� z@$��3&�ȭ�G���9ZoR{��
7&Q����-��u|��o�2��3��x۟~�k�G�6J�@�,����=O�ᨤ��Y/��",�k�EG�ΉSg�u ��y�eߏa��U�j�#F&�����u��<L��~�T�4�a�i��!�;W�ߛ��K$�そ&@3�w��u�~
F�޳+�`�h��A/�vI6Q�i��e�˹�R���^u��s����ia�l<��F;E��h�u�i�W|� �ۯ� ��Hsc��ĩ�#>�����y_cb�k:��3�ڳ�w�i
yY���ԇ]��v����� ���k4ZJ!8j��nR�����*�6�tѠ}Jo�>tٽp���b�N׋@Flc�����:%�Z�Mt/�����Fڝ* �f����a.�h���<��B�s!�g����q��Lbg�}��Ы���:�IU_�,�\,3��q�ьH�%�¡��_���t^��h&�+cu��e�q�w�y�K�x�u6*9.�\M�t�"	��Ө�Wm��e��<���i@[��;���D�$`�l�2�׻\�n�P�U�\t��kJ^S���D[v�xA�����莶�՛HAmx 0�xv�+f��<*�Y����6yT�n>6[R񴑌z�(�%�l�nn5�U�g ��!����u)z��2lg�4��9*Ѹ�N�$�c����V�}�V�ة1	TX%m-@��8��fa6��e�Ł�<���pNJ���{5��tGa��H�~�����=��Z�	�.��i�:ۂ�	7���fkS-�f��go��v�9y�;�����|߿����L?=�|�s'.��eeYPOD�UK�*o�P���b�[ZB�P���&���P�IϞ�
�H�#gk���v���%���K�
T��T<��bH���A*��n�	�$������ �0��W����4$ ��J7T��K�y�Ee��h�3xgn��^��$��A��H���W�3�u��8��W[�M���*f��QE���C��s-kҖݸ���a7�dc:��e�}���Jy�94֨�\��Z@���_��eF;b�-��oH�0�u3v����/�f�rϣ?��_Ȁ�#ð\~&��F|�����`��:�@��, �E��h9]h��ׅ:(�e6�Eg\ڷ�`Q����P�z�"`�fZ2^�r��0ɦӞ��5ܱ����jk5�R&f\Pfsg�c�>����y��bȵ<m�T�B ���e��j��>Aۖ!�t�v�R+��IFhe�n��Z��9ӳiv��������N1�FH�5a9͟�5�r~�N?&,���=����^Vˈ� \[+��kW���/�u`]��Dt[�̇���nF;���a��?����S'��i��4����F�2@a�8��P;^�LI{�bGE+ ьHc��#R��	�@����Ce��ߎY������4�N[Wԃ��mj�q����7�*@�}nA�N
�v}�E��y���N0H�L�!V?M,y�����2a��r��p}��P�����V�X=�$� ��]�1��E��Yf��f���
���1N5l��}��'��@�482�)�A���Y�j��>.�mBD�c���`ك�w��,�@�ѢHD<�#��T���fU��'�뿔��s?�4x.LO/о�ON�7 ��6���2m�ݬz!JĜy������F�+r��.�QD$z�ʎݫ;d`��%z��-�n[��M�_S�oiⱭIQ��1|����H)��ir%U�c�k�q�K�JtZ�a�[�U[u��5��,I��0��D�
�ߞ���.p���y������H�)#H��9����F7VCOn7I/�h� ���k~B��ے2hm�y� �ŭSm���<�ܭ bH��P�����,�(G�A�X�!J�-A0]GGN���C����/B<8���&�;fa^>�4�Ϙe)�7
�Y�W5�S1��
Ⲕ�e� �`l�=��*`$��W�<a��ȃ
�g���@�h7lx{�'��#ȣ��χ��題�P�+�
��$�K�y��&3� ݺ� ?_|�w+�.yV��m�2c_�\�Uy��
�>Ɛ-���UxO)B�c��`$��pT��l3�W�����佳C$�iy�[^� P�$���z>q�©58�
'����H�����;>�d��
�60�j�T7pbL!Π��z^�#�|�(�{��|6��7��a�%M�}2���jC����k�kEkp���2��qA��d?��I�	��v��������*�a���^�]5 �G-���m��$.~�K��F��L��4�hQA�E��:U�p��|�_�u�� ��=�3)��P�R���g�dT?��CG�1�E�t��4�唋"	�jr�HJ�3���B��`���}�Q�j���Z�^\dU�"�~�2ڡL���_���FN��+q��^÷[��q��n�ՙT<��w��
�&����6<j#���>�B�ʷy>\���P�2�I�2e*ʹ}]a��)�ME���4QgHzK��Q����/bW8���
�uU;���
0��h����S�CI�pZ�h��ya�b*��B	v�@�'jI[EX�Z��α����Q�됪pá^�L9Y�G��ΠO�)I?�D`.���}�w�'r�\n��/�k��~���a{�(���bt���R�p��Q���rb���fݚn5����.��i7c1:���+!��+>�d+���FM6*K���N]��!g����Y�|<��6|��Ȗj?	{���ly9����#ګc~�scv0йk�wU�٪�{���D�*�6篧�G�~xp2��������X�&9�)�¹�F���(i��e��,nP�7N�~���)0�u�8���[$+�Ya�N������L�:��J%���S�k�U� uyw<x7� ���b�\b2�V\_����/��Z�m�,j�!Ԝq���2�ONgU��A�$�a��$�
���b��qQ�Z�H��)�`uIm��,��aN�V����O;y͊��m5��=VNV#-��4�s���^nb��͋�1�R�!���`��)#�;%J8�^��T��b+=l��g�:�?��1��P�q馻 #]0f	�ȇ����2���y��ܺ+pc�)��U g�����E��S.�6<�h�"�F��"���a�LE�d�+�aJ]��a`�����N-*T�M��W��oG�z���q2EB@�d���R��gi�����J9Տ���z�{�n'�M_%�b��\�E�2c��Є�P���%�<�V�'��ǧ�.]�r��X�A[�R;��]�
qI3]T�6���~���y�7�Tt�|Ѭ��A����N���Aw�T�5z<��ŧ,�Z�J�l��J�O��B#z!�+���x��þ�hȃ��Emp2:dcV�azSͧ.�f*_���R��V��,؍�f��L��F���H����wQ������_�{l��tgg��e�蚴��w�y���1��Tal��9�B{S �9�;�
����Py�
�f�-�G�F��4S��:<�]s�qS���#��`��ؑ+s����~B���A��G�i��s��(�E��m�إ��F���XD�4�Q�m�g�8��p�ܡ���?]p$w�GZ��{%̂U)�C�;�Y��_l/�Ǉ�\%�.K*�:;���%tS�)���l�+�j�4��}��J�
�?E	PNoj�Uϙ2�[���p��'֚����r�m2�uڌڍ:�j�J-W_1w�s_>��Ц#o��x�r�<S�-�S�K\�L�u9�^&���� ���S7����5#P�����.	J6�t���Z4��7���(.��%�"��o�XZ;�PP��9s��[k�R�r,�	���޼�������G���<�-m��,r�VW�{F�{�@�M�$C��֝5k ��2߉��`�����$�r�o�	�}o�g����D˓��������b���D��׳�u|N �����;�����l��]�k�=Rk��o'�j����_�)�I��SUc8j'�˵��~�;1��Za�p��8�G���H0�Aг�iK�.�� ���\wށ��-v)�FV�<c?f��j8��T7w�>��=^���5�j�T0�v��e��;����м��`�X��8���@�43��/ 8Io�M��$�Gf��9ʼȮO��͝	q]�DF�9�'{wJzf��b��amP�24}��u���|L���ɉl��c�k�t*~�D-���r�����<󀹷���^{�˴���mK��edf&���ԕ,�P4}+�ռ,��b+.����<�-Y���L���cy��a/>X0��HH���R����i^�S|�uC�o����C�YSc��yr~&�"�w�SH�w��L7�p�$�Y��D��Qt�Z��������s��'���0��Ԓ��*��c��C�z�a/�E��+=NO�y �r��oTI��D�sZ���vi�p��^Y��ah�� ��z��k;N�<�/��,��?��`��d�[[�k� �͹B��ɳ�B�4�43K5��(��Ec���D�J�N�yTX����d{0D�:�<�H��*�<����OZu������&�k#Qld�����^��������{�L�7�'-���9�;�P8P�\�6b j2:�}������`*�,���͝�*tE�]$s�D8a�z�q�����;�I'Ը�JaY��l�=�;���'�lQ��*���P��e*�x��.��ɕW;�[�����1����O�M!�	Oϣ�
�.��}B�!�?@Y��}WM|�u���J�p��/*�N[|�R���X-49S�jrz�Nm�Ȅ��d��9¿�zF���ȈUg?�{d)�1�h/I}������� �_��|�〫BlB��@��W�4�A���^[]O&�b3�V�h��^��sh����m�D���֠�"(a�D�6!��tȧ�=�؆*�(���� 
m���zx ;Ɍ,���[W�3@�zHUHv�#�<�;GV�?c`k+{{�-�QH��>t�0�:6���[�2O}M���]BʋP��~߰ n�3�k�h{��
I�����;ּ�*@���N��Y�8���D|�b�Bx`|p<{�u���F5�ٷ�8��/Uh�h_��c	�{�k��\M�>Y�.���N_Q��*�$��l�&�p2	������h2(N^�E�,�%>`|t�-���q<T+�Sgvz�߯�.[!NCb�א�U3���A��U�3Tʆv��y�S�R����S:�o��;�`���[� 8.h�h�h6d��iV�W���r	��w�蜗�TF�����6@Uw�H�������'��߯-�}\�j����"��G��O�׼�A�*;Q�d�߽���&��U�$�/YxV ��{mz�W�m]���m?�����Y�J؀�s��C0�$���#��s��C\�Q��<�r���Wb�V���	|m�����Ȋ�(�y�s�r�&8�M~I��)p�Uf�v�
/ɻ�0?��C��8�X��e{Zx��!����7~Z�/�E¬%eގ{}����:#/��|l`��G��>���
.^�����*D���h��/���w�W�kb�NO���z�z����3%J�:��ՊA��E�8�ԗ9#?��;Y�툡%["�I��v�[���y�%��_�Ϟ	�Sl�7�)��Ë���Dc��`¬,a���[.����\$�������I�tߟ��I*����T3��}�V��/$�u�5�RY҉$܂l]n]𣹀�n����h�OMM�R�����Z{����Y�h�?�E!���L��2�Ԕ��h@#�ٽ4�͸�S��C����Y�E2:W �s���hw���w��.8D��9JΖ;�zT,��Ķ2�Q`�����V���G �#()l�ˮAI=8��	�iaK��-����gXpfJ�F��N��bNR�mw�U"��8�kY8U��d��?��h�P����������9�4�
�~�ٙ����.��_5�4����?�!D'^z�����9t'�dz|�Qk�%\%��Z��G�Y-���ղ�W��«��	�	������n���E���<�G�����?&��4���J��J%�N�crdܭZ�t_3��T�d��K���Q�61�<�,��7U��?t�H�kVk��\X���G���ی^�HW���wo��_����л��8���w L�&?쏔��(�?S�uY����_�gR�ӛio�����<��fb��2[S�g+�w�#���⿍��j��𬎌�I�N}1���3wZ0�F�T�����B��2�6Q7':��IvF�k'�wʋ	9����[a
-�ّ����IcA��^��$b�����4��zWc�g]Z��Ջ��J1������G��k-X��i��d�hi���O4�7�+�*�p9<� %]�Ne�{\�dب�ˇ�~�_}�A�%�U붚*��YS���%YV�%� ��k��cr�"c��z�%��,��HS
�T<��`�o8Ԝ�<���.�}�=����-6O<��S�i�S�r�@�>��{M���D����M����bY��L=��cчj0�ʿ�*E.���,�K����Y�&~����ռj	�6ndB�@_)�����q��?�ǟ*��{+�fz���N�(Iu��m/�����ԾA�|�����'E�V7+���s.<q�����H�-�}�|Y\���v��S���=��e��Ո��;K[m��i髢F���M�%���O���*�Zα7�E�����t�jr�2D��!__���Eɐ��"�W�c��=��Q� ��:nP8��G.b[�#/�ʬ��;q��C��}����B'v�S�fH�ܹbB�/�I��x%Z�Q�gPq/�ܵ��_}�K�T�o" �m;¾�&�[���(ҏ O "cd��}a�.����	3�s</,9�ќ'!��)�Tg:�esT,����l
�F/!��_O�P�9��+6����kW�ǋ�%��s
 ,�Y	TX�H�]��V����
Z��N�t������r�/����T_b3�MΘ�ʠ���Q)F�&��H�e������P0�H�OMXw�p�q��4��TvqO�����p��Na��B*��뜄3��#2d!��f�b�_���Q�7����1.��`i
��h?<���cn�\�F��C�t�/�42���"�3��U
����z�R�b~�j�էHW�j���b�Z�+�O�q�t4j���>��4OR�Al�dr�fz��{Aq��r?�_���u��,+��|4۽L����T?<�,�i�٦{����$K�2��2�4�.�y_1��/�<�ݎ��;d�k ��O�&(�P�P�;4�O2��hjL��:�ʳ��|��""�g���7���-,�����,�p�-SV�  �����~U��ѱ��}��Q����c�Q`����i�>@sqo��~,� at�s2A���-�P�
A���<r�+z�8�U����R����C�z]W��A4@��)�+���ￊ���}�zX��ktnr�/f����һp�# �x��`Bqq_�&s�Ԣ�
��@�7 ��9R��e(�T�/�X����R��[���5����g©���Z�j���-M�qSu�������7�ϥ�����1��EÑ�� Ԯ���p�Hف����o�����ڷ6M-��O@�xB`U���"��Ά�~k��
�B	�#�S�8�����q��EH�� C;����="��"<�O;Q��J"j8��/�&�"W`G-[�QdZ���,��0z5ur��wH�6������	�<ml�Y,?�B>��\�E�M��&�Ќ7)�ɬ�L.N��&�S��f:���-20�qbĲ����l���M��X��m&�š꟒U 6 �c�&/���ujs�'2���%ȾCs�����	���Htj��p�k|J ���0�^L[�"��d%�<����ʴ0DAɤ�"�nH��Aqi�iva;�W��m��Jw����puz��ey	�@[A²է�#�)Ckdx�_3��N�`��t6=���7������/^�?G`bA�-."�����6(c iT�^J��eqK�\f���FaʄwRD��So�5fC��/�ޔ�eX��.c%��%�x�v	V3g$�ɭ�� Ͼ6��e�c(s�u�'"˷ 5]Vd�_b�46⢮:��D���-k [�|2��#H"5HOl�(���DaL��X��/ώ϶T�	L�7��Do�s�!��Ք{�M8�vNhE�L�{��}2�M�i��l��oVB��o�!V���ϕ>]K�o�Ej��Sv����AI���p.�~���(���毿A�;�޲-~yk\��2�����FP]g�Ђ�h�[�OOy_�첔G��x9j�M� A�M�b��ѬȀK��:��/sfdg�)��J��,BAnڍǥc[��=p��粏y��@v*m���N���W�]��'T��xs����jbp��6ˈH�|�lzfP�=��j��w�DB�9��S���H��R7�C�4���y�&����N�Bt7C-F+���%�eę�Eu|�2���GgQ�1�Ŕ�Q�y!��q�ϺN��f0�c����ʳI�P[��\�|����2"��z��R�]A6���B]�����6���\���c�/��Y4��s���t�\ҷ]"�n�d@����� ���\�ɉ+��H:Y���9��H�<�؇�� Z��[�S����G]����H�V�T#�OzV�ֆ:��L��.S�/��G�(�;�\6�	���
M���	��=]bҴ�BEi�'�@Z�3���spt\����9<�'	�U����p8Q
N�~�4u��/(��I%{1��|�F.j�GU����?��Z�j��"W�9!��7,���+vQe�m�>���^OF5:'s��������Y��W�����e�J��mc�N	�+x�6���r��?��Pu^�j$y�^yQ�A��h7�7�h�jTAt�+� �Y�b��GM���Mb��"��,����.�e�/R���%@��q���L���nq=���(������R�����"eP�����?4���/K��ar^5�wMjy6��0I���u5寯ք2�c�VhGyЊx�%S����ӯU�s � �\*�}�����#AsW�����4��@�E7�Q�1����s��,�0���h]J��x�����ء@������3D[�g���ȥ����'Bτ���q�V���3ީ�.:f��Ae�	U��QW�UZ'����GR* c�����3�4;B�|���oZ��΅�l8������E��+`��0������-U9}���[�l��A�y�-ϴ��5���D�i��o;�Dl˯)�-�n�<�ot��W�DMI�Xg��7�<vMCR�)?;������;�����H�*"��7PsI������"���k̻���s[��;���}�y��wB�q�M]�C^YӸ��HY;��U�`�e�ׄcZ��/A=̚46�iW�n�Du�[I��ڏ���5�Y��[4
��=yGD�/odD׺�i���,�3XG��A��7�q f�����%;����9���
ixeB����� R��êQ��z�&V��
�k�����@�M��v�ǘ�����'�&���_��^�hn�h*h�&�m���ˊYm��\>��7�}Mv�[�c�g�o��ò}c���\���*����ИQ����b8�4Bv�>6+~آ��3JH}$�ܛF���;�F"� ��r�q�-(@�7t)ׁ��@5�&_L�
��3tA�(�p�d�ɂKWP5H�M4C&����b��'���3z�|�$�A5�u��Q-K��&@!�E=�G[Ƭr�j48/�b�6�.E��#�,\��fd9���~�{���.�x���iHj%-��㐙�H��% ����+�5�3��C� ����0��h���I���SP��O�# �z�ݩ�/��E<�OD���ɮo�ޣ9�Wx�`�3K��ز�iE�Ӭ�۔%:��rʒ�/��F��\v:��d��Ǚ����!\y�.󀌘��ɔd�؄fM�6j
PeR�b��Z9�v�lxr��+w	M�z��xH!��|��U�4PפJr'�E"fem�[���jh��iY�i%ͣ]�w�$����&*��m�d�q�^��[�F����w{�����*;o�!`c"ŋ��+�^oNs�&9T�ZEpg�S��8圏,���v��L��6�)nX���ޢ�hth����8�x-��q\s�E��G>���RIn�h3J$	��=��[/E��^U!�/�<e���E�-xT�K����I��Vc	����1;�S�'T�S*��C���D�t
���O�!��O[i�^N���8�������1��S�[f���K4��Y�K�`f.jL6Vz���`���o�6�,��7�-���5�����"c��o�x�X�nSJ�*�Lb�r�䉉�}���{���9՘<$`X��*U��Q���6mmˎ/�dB���*���dj�3���'�F��߸�ew��s��|ř(��j�=��e�%/�ޤ4��)O9�x����#v���
/�^3ޔ�_4x���Q�˒�;�Zn�	>"��)\k���#�S�!Ie�J{�yOA�<ӫ�M\͞g�4������L'}��o5���,�D/�o��VyE+Ei��;S�z��+��1}��8�P��������Qȫ��ō^������U�a t	Q��,D�h�5�S%@�Gq�h购a����m̈́܁�B�>|
���B���ٛќhءX��,��J-�K�4CY��6"Z�X�:\g&�%	w.f�n��A�h��^�P�0���$�$�r?Yz</���z �`��+���ٜ:"D�2Njo��9(<6���}�" >�?��R�e0W% �8�m�!V��ؙЁ׆���]�;Ϣ����:S1���+z�m��V�#�e?����a�&���X���\� [O8H�a��&�St<fz�Y�	Ĉ�`�2����1����Z>��W����c�k+eF��a��´_�Rδ��t��N�/F��N")u�[?"c9��ϼQ��y�)��pL@�c�jbUm���#2����޼��g�m.賛�1[�{k�b�Z_�ͪ�[J�H�/���Z�h�J@��p�X��,�8ų���	# ��}�F�'����)uJD��d�SbB��~>���ռ��^F�M�&E%���s�*�9u�{��^�)>U˶5�i�Tȩ�i'��h�N��慄*K������ ��iˇ�h{)��a��dCTX��QwjF�������^�,�l��(9�c�:��Ի(�|QL?#H�ou�ᾓrQ��Nj�P"WSk�>'��v��%lsN��������R��㋁��j���x��id�wV�S�S?S��3|�v�����No#�v�~TK!�VEaVM}��Y�R5�I�aЃ�������(n��H�ۼ����R=��w`h _�t�	�j1� ��9�o��W�{��i�`���K�(E*���T���f7�p~�#�*���d>wKI{B���8�k�!& ��(K�<���QO���H�6�W����h���ּ��q�ɘ��]x{̌@ojHmT׬��N1�}7��?��Y�t?L���GW!��;̒�X��ѫ l)�zw:��׾צ�M�+����1�`u�L��o�OD>�F��?CC�n���Oƣ2� )$�z�Z<��+��v�~2w@�fB�lg�S���ME�H�gC@>�uC���B~�$H�Xv�ٽ�ӹ	U�7c�s�O"��X��ڤ����^����.����=���E�Ǝ)�M>�е�=3_)� zGjw����g�L�ܜ٭�[��۪�gʑo�w5@v�򥚋KU@�*RK�04YH��D !���@i�����	h	�
t��i2�\V=�G�^V8{����z	�Ӎ��?���o4p����X��L+9�o�3\mx�{���3/�`E"y Un�p$/������=�����6`�#����r��A]׸��
#5Μ���A�w����Z�C☸� �m!�y���}����)�Nr�2w9+�T_��y�!�R�ئ����	��C�r|��?�NT�U@(Q3;8q8�y�SY�Q��?���ap�u���o/��{��B/�%8r��/?֩��������~�b�_���U�}PSqS���į(Q9,��C�:����e��~|aH���4�f�L�|쐣�n��l��ۖ�G`��C��d�L��97m-1a�Z�\k31�+��E;,H��$olL:��uӃ �u)�S�y)�]�]�y�CD���K�L]O}+�7�laVRc8�kCBgب�.}�m;�E����x��I���P�TW��X�sb�8�k�k](%��:���*v�Ź���l�vc�bt�v;��s�B]9��T|��<@(�}�U�<�A�մ�4.�?KD�muN�*K� ä�\�ŭ�G�VB�|�r�
:]��#a�,�ݥ��6DH����'��V�Z
�O�����F�ىl��6�S�-F�}���\�+��,��0�Nҫ1��\��i���9�DC_�C�����X���<��'r��[Q3�X����CU��l���Wi�4Bf�rs��`"�E�Q�6ω"S]>��Q�J��&Ľ�uj�
�
0gQQ�`DN���A����_x�[���6N��2���~qV�v.�
���tӞ4�6��rM��r����a���dO��\X��C췙��H��uk�����e��]CMv���&s�����Cn��U�4�b4j�w����/QgK���j���K��G�3�-V�`��u_N����w�>�����`��@{������m���FnW(NV�oȚ�K�l6��&1a��,�Zp;��o����vZ��vX�ܞHJ��Ʒ����g��T�S�=�Q�>������3)��tSɄ?��V�矐�֢�������O&����ꎎ���/1��Z{��0���h�p�5��'�5k�-0܄�����Ot=�r�0�G���,:��?�y�����o�-B�9t֝��]��xM*�X�rH����C���i��� �i�N�'5 �6�N��ҙ��dJF���H0#�d�@>��t���uۆ+eo��Oλct���\#���E�G�a�|Aǲ�x�l�#h=sF�h Dn��@5v`f�{�����G-Ώ3������1�qdf�%���'ar�g��7��`$���rӰ��=��#�)-8�/ȴ�����l�$yA/���6@U ;�9�ɧ7��P@�QNKZY*��&���$y<!ԕAwT��BioU�#��L>��	�:)��cpnF�� _IB.��ے(̸�ً$	�ğ��+Cw��-��*TF��v8o���P�3���8M��܃���Vy��Y�h9��.JE�RM��m���#����S֩+N�O�٥q�iwY-����O_k�9��FW��������uda�?���sꥶ�U2�f�^5�~�D]ӝ R}|��R�Y�Kq��&����Is|�Kj*
G��������e<Ռ��?f�yڋ1�x���IϘ���s�����3��u*e�^--^`Rh�RE�m*h���"�\��YB�S�+�M�{ͧ�?�4g�N���y�z‭�H�y�\���5H1��J6����wE�ȳ_���\�R�E7 �"䈢Χ��pEH�|�8H���S��(]+�^�
#�dG����2(Y���qG�WO�D�CZ���3��0�W�+��X���eR�x+���;ˀ�T]�W@�?BX��*�c�=C�A�n֞~�q8�����Kw�}h����Ό��mgɰ��8�jWB9�׈��4|"&b����ʀ)���]8�#?���6�b�ͽd*�����6���9H��H�P旎�K�t
ؒ�b�����s���|��å1i��aN$�,j�������W�K3�w� ]���d)���z��\�P����v;
XBg�}JN*E�vt�QG�y��v�?�š��8&A3d*65�R��l^����ޗ]�r���q��.���|��%1�b�j�<(���C��0��o������wD>
�>�s�����o�w��&��ʁ=(M]�'l�;�a�Z�>R�7P�d��&�;��#�G�Jp��(~�Oön�g���5�$���'7F��@��t�"?��Ϊ>9|�6?;��\#���'�[S��_3#ә�Uta�d��B��?ƿm�>Ty����Cջk��oTW���e>&g�vő�18��?>��D��o�;�t	>f �֠Ml���� ��A[85-歅�W���>��{��SX�B�iٶ*�;�c���@1����������m}�ClT�ܺ0/�æ?2�"��:��7D�����������)�ąV��-��Ī��^�� ��:���Y&}�j��˂=�����N�3D�E��
�-`�/4X�c;X޸�N���(�~�� M�àM��3J�Q��"��	����u^R܊ʏ�X��׾�� G>! <#',"�����{Kj�,�H`�ᔴt�'-}<�x�g��D����/��ac���U��s��C\��Ex���4g�-Q��v�)�F�!�r���8��~1B�[��!E���Zq�jtAH=<�nm������V#�S7Ϗye��@ J@(�%^U�| -�?Lk|;H <<�[�w�  � �o?+��l�!bųRL��)-4G,�$���3���!F�N��������n�s8�i�6�&1e�dX��E^Յ�s�I�q{�'�f������SEe�8X��>�x��1��4��ٷ� 	���Hz��/��H眸���Y�lRu���Ƅ�O�5��,z]���ywx!�M�[�1'(�K�r$g��8��&�N���)��G�j���}�D��$� ?�E-�i�\��N) �٠uF�!���h5�f��w'�8ܼr$g�FEk��	�(���|��3X�ށز�7Ⱦ�_�1q�ۛƸ���7���+���;�����	,} ]-#n�	W���!��q� @�P�:͍i�N���a�Oz: LQ�21�b|�p�"����e��d!4����*K�:fl�t�~��̻㈹쮆l��P�G/��L_����oyn���K���^��D���t�64�˝�D]�?c5����V��N�;�-�W_�j�&���B�!ZU[�]��9ŁZ/ك�:a���a �{�$:�A[F�;�0>����,�Þ+��EE�v�m�'��N^���÷"S�?n�*!͗;-�j��Y:��zӁ]���v��x�/
ԁ�pB;m̠A�ml �ʲ-��Z����-�"WF��N�3jgq�ـ���;C���|E��A�o�{��3�����c�������*M�s&�-� �7ݭ{�=qK ��xۥ����N�Q>�DdH��<v���(Hա�D[.h	&V�D�i]���&;1,ޗ�]=��� 	S�X�d��F�9Y�����ʟs�~:���?�Ƌ���H���(�`,����U��&�TJ��Y@��ݕ!����q?9�ܤ dR�k"i; /���<��`'Gz�����h�[H�����i:-�9}>X��\�Ҫ��<.y���w([�7��BG��=Z������a_�v.(�bI��F �%�`#�n,�ͽ}tV�M�׎v����3Jʫ��!���q`�%E��u�sj��3�0Lm�<#�����08�r5��͒�-������h�|}�E�%�mp�(S ��ӹ�������#� ?�� =
x �l*  *��>�jW�J��Jͫ3��Gke���&>�Ҽ��5�hɣW�8l�2C��jEp��!�T`$�1!��N�W����Ä���"ċ~���
�N�:ө�Q��2��2h�y���;�_���q򨌢0��k�ɖ���#6'�3;�.�-Z�I�,f��ð�Ơ����S�D��	������-܇�6ӟ�ן:�����	5�����?�k.o�TT/�{���������ڞA�B�`%әzЫ���!
���<�xg��+�8� _Bel�c�������d���1r��20N���t���7e@�����_ߟ?��j�9T�e���е)���d�('��Y�����w�x�_�CC�x�'���w���I�⬄V����(G����k�����C�D������	�Y�P\*��9���OD%�ߚ_�^Y��ӧ��zt���R��
:���tEtc�Pi���֎���ѮM�v��^8���U8��ZQ�1�=�Я�p>:�E�7o/������qnIc�˜���T�me���9�:�� ü��Es��f�t`�5w!�K*��s��k"Z�6��By�\�7�^WW/X����XrV����{Ȁ����c�7,Pрs`����dD ��]�J��hLImq�cHz2��Ҋ�ҚX��]�P��_�I!�9�8�x2�_ý�9�Sp�{����F�%r���!"+�$tُQ�~�G��_��RF ��@M�z?�֎S��MJ����U|�b�u�^�UVf=�{�ڴ"���ON߼�GX�Y1���l�p�s|C;N�F<����L��#]ןAl$�8�/��>��P��@����z�D+�bޏf�{S]oڭ�9��GN���p�"g2&䗅��������RQ*gK���bܸj���!�1@G�?e��s�9Y!� �n�<��E�E2�@��㱁OFB�@�uW�T8Hu�wm�4"'��t���������{M�u8���ǻyP����2@,�;w��7�^�"l�S���p����gy�]4ۥ����NE�D�*W��ɛ��8���I�q 3�A�h8��v6H?��%Y��E�#���.q5c�:C��G���@���&4��Z��l���"��؃��/�K����,���Cih�e25��5���3����@ai��P��E�\���U�Gch��ձ��p����BOQ�0�� 7�������@@�\��ʱp`�d���so���7��RBv̑g�k�O�����bi�J���'���'��!c��k�%�'h��BgI7S>Х�m�J�sB����\�!T>|~�"{����".�G�ׅ~R�%>������*��8�E������6~�+BK'k?J�:g)Ϋ���.��Q�����L���0�x�
yu�I�郯�2����>S4��*�����6��N_(P�ǒP�9���.a|Ɨ�D���E����P>y�� j��n#x��3��ؽLC�Y��Q:N��~��p����"|h����F2*��t\��ۍ��_�����pH�� e Z�(d�T������p�|N�
/G8\�|��i7݆�EJ�#�D{��1H��խ�"�b́��#�	Ŕ`Y`?��g�VÌ��V�0F�N��`�^���6	�6$��^���0�P��K9�U*�hד	"�,ᕛlS���j^Z$����Ќ�C����>4}2d��R��@����J��3�)�\�AY���T�u	��x�MoH� ȹ�S�f��7���T,t���ە��1]��3 �5��S��U��C#L9*�p�9��Fw嶹Գ��9�;S������W�I��v��.t��d�oer��J|��0�����'�w�W�'���a{����A8t|���>|"�����C⟱��^1#>��r�ʀ��-@����$�H�1����y�o��R�a�+,�fȜ@��=�_���5�i�6�����o@j�_S��i��mڶ�q�SNyWF��>���ۺf y*s�cf��웍�ec��>[1Z������*�=R�y�.!���Ë!�����;jm�[QJ�
���^��n\���(�p��*?��j����Aֽ;��Q����K�����:����L:]NJ���$� U|�ḡ�*Y�dNω)4��b�g��0��q���aƊ���Gh8�#*3���׼�T��1/υi�Jj�$�p���@�����������Z����Ym;w��ϩ1.4�;���9��a�V��Vn��?L:�d}f��I:=b������"=�Ό6S
zd�c<A����&��$9^P���:L��Sg$���8Zc1�7��`q�"�f������j՝Ċ���a�%ds{���R�A�w��wG	��)l�����t�
�t[w�5D�l����}>�@.�G9��T����z6������4[L����2L�g��}���ZW+����"�
�K�z��1�y�pvesr?|�h�֫5������͵Dw������G/?!E;A�Zh�;�ap������P�@5!�a��'�1�*=�U�4N�S�%ltO��ڙ?��R�tΡ��)���G`�
��Sx΄<mCk�# �ʺ0GA����R��ts�3���]���Y�����2�n�1DcD2�'b�nm_�,k�bU��ߦ����yE�Q���wm��^�P�-3�A�J���sG����N����>{֪L�K��� �+��l��+�sG��3�4�x���ҘWl>*L��^Ku�!�,j�v�����#���._�N�8s��r�8h	���k����"�d�ss�r����N9����,�@O�8�EY��TR��Y�Kt���֥Gp쥬����k`�3g��������u["{R>q2�쵼��Ot�	�dܓd�6x��C�_Y�kV���w��=�Q�4S	��e<$��7��7���x���:���ԉ�hgX��[Y�^R�N���*������@�����`Q�y�=H�������o�l:̧R��?��oJ'�Vl3y�"�찿'f���Ss��i�;	��p�!j/^֚�_���������_ױ2ho�͓q"�L���}7���9��-��BR8�
��s����P�������6���%b�)� ��7v�ģn,��j3Գ84�uWc�
�����E�������CW
^e#ӈL�*嶧9h���<��_��F�������u�	�P�[���v��+DW˒U�O����@��x���j>U���x١�(t��F�"��[~�[����� Z$���}����Ƚ������+f�eZ�'ùo��Zp�I��*i��ruf���r�A&�׏�4��
2����M��,�
���r��\$#D����7�.�i����L�]`_����X��g����N�J�H�̨&�`7�<<����_�� �IM|	D�"���w�M%U�����Yzpx�g׼��֠k2�OU�ޘ��}	b�L�1i>��_����ҹ)�RЕ�X�a��*�A�Ǥyt����w� ����.��H\#�R�������z.Wm2�C�)z�Eժ���H�59���v���Yc"t�b��g:Y�ϛ얖�}�����Z�g{S>�1e-���M3���Ĳ��ŭ�x��Tvy��A�1������y��S�����/���c���U���z�m�z�u2����1ڹ��� 2��&q`|���	��ޟ�my;��f)!T8�j��@�+Ԕ�9�HlMX`�Md�e7`;��	��#���Î!�%��eԮ��n̫���"o_s��~�i���-X�=��V���u=`���_��}΁���N����= ��T�҆�B�� �X�u�Vf�}��	f�d ���M�@�K�I�z����_����'��gˏ�e���[,~�7k���D �|M�A툅�59ʩ�Å�� ����#gɻj_�2["��6�<���	#̱5�rw�I�k�&�l)~�ќ��������D�*]z�i�sjZ`�4�63���Tt��u8���R��/�:��H/k*T�ML�B�����^H*��������<^�y~ �Z�uxC~z3�dДnM�"j�=���d%"��ȑ�0�[\�4���^��ȍ��|]#����g%��V�a��WC���!bű�/k�Π���<�y 2x��jŕ9 �%�0�x�xۭ+�
k���&Eɾ�,�q�.g�������BC��E�)�1[p��1='{�\�yW�^,ԯ�*d9"/Z��@ه�>�x��*/��;�)5���]x+�QY��V�=�AU=�)+C�7;�i�ݠ�6����O!���Hh5I��D/ N���n��Uu{��8��GWe�)�he�İ�q��	�� ���N� Hԏg}꿱E���>��N.S��T8�+��j��R+<��V���zi�4�S����>�߿��s.b����s(%�0a�ǳ��U��p � r/Q*�:`��ƳH���RֶBƳ�6ŏ����ۘ������2=���z�����Cr��5��#�\�����@��$d-4����Jm�-8E�`#0�Y�h%B[����ֲ��+.�0�{��Ej\,K��F����<՛J�>�s�0b'��n�*��獾uļ�C���j|@��=����6��A�ڠ�t_ʓ��㫚'�:�(�3�3I�O+F�n�L���ئ�� �V�ީ���o\,�ӫ#��	D����t�Ht�)W<�t$�gxkA$X����"p�Ͳ$ypޚ����#�}T#�T5�?�	I� �(�.�xϠ)�V��;���_=
]��u�g�	|�7JX=v[����Hc��j{w��g.ܢ\rJ�z���P	+�8�ٽ����]S~>Q���&Մ�sS��\S�%.u~`>�۹"�b�E!a��&r�؝S"�f?	9�4NCsy�u ѐ����(�9��Ы4�������a37�u�����%��d~mf�%�a-�$M�n����L0��F<�T,Z��m�����9Fc��a���eSم[4am�<cԁ.-��r`��Z�ҷ��
�V��E��U�Գ������m���WCƿL�����4Œ�_�N;�R������4H�?<'BF�=�r#�'��9��3�7*h�7Z(;��-/���(k�^��,�I���Q}x%�N�)���5��2��e�&o�r�DŔ�]�l�:����]	P@�����{� ­����%�F5�{A�� ��7�ϬU�u��M/|���O�Z�*x�����`��p�k��#�եp�v��M�wh8˔�|�{�6)C�4��{�A�s�W4z����g���T�~K�ʤ�ġKg��|i�h(`��<�OLb�w>�Wu5vn�c��Y�k@D	�/��/PX��2�$����L��/D���L
�K��|�>���$->��S�^<��=�|�<�v����0��s���y��+��b,bfQ��sԸK��*o�S��oR�EM�+��?��p�T�	��E8� t艭	,��k����^9�i)-?��D��PU�C+�+��ȑ�2�mc��yXj촏rk?\z��<{1;gs�hd���[*id�.����7�"�̼݊���7vW�W���A�ߖ��S����?�s,�n��~sI�YVn8��K�E�P�?�DA);'C��0����K�\=Hjk�Bx橈�}%�֝�����&3ҿ�O���V&W������k�N��2b����"��)%����dT,,���Eo-d���D��Ƕ��i'�©�*�h`�����:�K$�Q����,��X�mٽ���S"I���h;a�Q&���+(�S�?���S��O���o%`�nu��t�z�G~H�@@�Eϐ�Y��(�ee�B#Z5+�x S�疹0E�}���������j�"	{K��v��85|��#�Q1��"�>P����]��b>�
��(�|��(#���L�@K�jm��h�W w�I'�:^Dǡ
_��]761=�Ɉ�3��ʴ�"���WM�M�A0t�iϺ��5�g�����ɍ+PqF[��铓c�`h+U��N���M��ځڇl�kӗ���	U���@��=.Q���"�]���5��*.� ��ڵ���Zd5λ��!"����W�6���=8C�f����(�$�!@s�%�6h��F�TWŸ���[�c�[Ю�;�rw�!��X4�!���������X>�w�]f�!Q>Z�����.��w��[8k�z?`�˻7�%1l��z�]/�&#:�ga4A�dwf�_�8�@�V_��?kB����'�^���6@z,g�@,H���}h�߾�ķ���Ҏ���gc�f��e���d��5��bG��I��k��7�^���	����RQ�   E���a�l� z�n��d�����D|$������R���T�T���^��L��%P���E�N�e7��B�<\�t]�ާG_�iD� �!u������|�xY�Pd��%��4�����1ÀL,;;���0Or�yL�����t��ϗ�j���\��ҿ���ٳ!f�ia�@X.�A��a�-zȕ��t���x���f�U��N78^$�-�wr�N�u���bN�8�hU��%���3ĭO*���@�����k���
�C�>��Gwp��y�s/�ڡV�i:�1/�?Kˡ�*��_�� <E�Yy�M�?Y��r�h"�5S3���%�_)�D���H��O�R��*
H(a�����!����h׳�U�T3M�P��(��E�eec?T�4�µ K,IXhj�+���8�#G�f)�(z2e��Ga�%�U�3���K�?��pK���;{	�����K���I�0�M'Ⱥ��ְ�Y6����<�{Y�W`�z@��{f�. jT���R��2��c�1!�@8o�M��)C��2�jTUɒ]+s��3����JB!�����x���!B�+V7���?�!�X�5M8��ͱ]���|R�������%�w���^��54�̯��2��"�+W��)&���Y�Nv{j��?@#lW��W"�����l���U�<�}���/,P �˞<�:�&0��}��+j���g��m����D�~�%w��T��).$:.9&dwyV��j�yDw�i6��_ދo�F@_�ۏ.uά�*�L�`�����ڠP��������x�?�幤��#U]I�7%�>��<�U����ҕ��n���LD�4���T���8��V/������D����e��*(p�_=�MmF��:�4p<����H'Yd���9ͤ2(�����`����������ma�M���� g	z�����<T��+���e�	F��Py�DW�����6XV�].�nS)Bс��^�Tɞ�c�_�.�Sq�'Мmj��y��3w����q��OP%$\+��_greZ�=Op��ov@d����r�yd���9-�Q��Ţ]Ɍt�0 ��Uh9C�p���N��V6�!�b��t��??H��em��˽�D���lVt^7����ID�[MOPڮП5��������<�GO��dä+­YR%l���M݀��v����#\�yS�h<�B��^T5c�K���y#�&5s��[1��e�c�� �`I�Y���'o�#0�l7�7�&�t����a&y����6{4�����p�p�fJ5�F�$sNF\[
��]OmA���u��^_��Y�[�_�N�|��̣�	Y��<fW)�O�^��&X�춤
���W���!="�ACk�yD*�:.��5ԶC}����;Sa�E�dO���:���d�[���S�z��KR���L���݆����p
K�D'�Z������d
,<�p������32٣ z���� 	ps0�I�S����)lX� ���:��L���[nC�b�ӛ�bd��LV5��A[���v���{$��͕O������Jw�I��݅Ց�r1����d���r�3�xnO�~��1���'�����TOM���G>�U�f�[�g?؎b]�ѫ�_o��NJ�eXJ��P�.�{>���y�-�*YkE|�YM]���/�X�������C��Y�_��6�t0�0�W�J4�G%��������NX�ĴYIt�`~����H����$��eeK��o_Vw�L��s�����Q���[�����[��v�s�N��{΁)ކIZ�ora�6E\�,nl�9����fFA�"�WJ��FրS�|���m �#Qb+�rq�M:y[�I�1x
<]�d;�h�h���c+-�A�i����0�e������)��^��Y�6�!d �0<��	�xm�ן�K�F:g(�:�'p(�)�(�F]�N�Y�>���?O-�I�!{��`j��Q�����;\�"���.?!RV���ű�56�� ��Eu��'3;'y]7��� �Rs\_
U{��]�Y�ebL�l�Qwm ���^����br'HXN��6�$��v)�V�&
O��Z̸)9��kPM����5b�L�V��_�i�~Ƣǡ����K��8�	��D]�~�	<�礜i!��{XEKe~�D-!�Z84C`\���2�0�"	����	G� ��2�J�63��H��f�#V�8l5j�X���vi���<���C�c�����徰���`��mlGb��^� ���ݲe�t�A��Y��H�,��m&�*��B�ݱ̺���P�?#������Y�팲BC¿�Bƽ^i��9vY�Ɔ��F�W��O���Ub;Tfҩ���<c�_uK��M)�d�5����[?!{��L<�ڭ��6��ر773�1�������j{�T4sQ�I��gk��Y��闭�P�.18t���>�A6?�RBI��ܤ�<ݕH�bTH>���/Z[Kjx�=�ǌM��W�u��	\iW!c��N�7�!� �	���;���*��Vg�rA�����R.K9|���L���ͼƯ��@�΄t�au�S}� �pg��J����L`��5�
	N!�#3ޱ�!���`�;:Y]���3�r�&�N���=���ƒ
���e����]����G�6~\>6��w\�,4��b[ڡ�.	���Q�D�V��h�+*��9�q����U����)���7K|�j���|YM�-8����b�}m��9i�Z��%9��Z�}��H��&ʡ��L;��![A=Hna�db�fMC��_�t\\!��o�)��z:f�x���a��+�Yh:+�l|.r+�}'��o�QW%>�~�[�ɗ}�Psj)��oڰ�0�S%��^_ í�;�'�^��V�W�Ǹi*�/B@�j�����M�6@Q����>�&L�PI�W[u�5��WA���z_����?�"���o5�z�1ͬk�GMXm��)�.����Y���ޤ�1gz������'9��~�#�ہja���*p�V:������ꈫ��%�v�����r�8(Ąa��7���j-�Y�m��_}A>����f�� �̕�>��8h����u�t�;+
ͭ�P���4�ZrXz(A�U��\��Y�/��s���<���O����� �}TcGV���ev�Q�1��WQ���s6��uZ{�cV�vo���r3�gҦ/��EE�.7�ӹ�ux8;}PD���"d+5�I�����':c�k��Y��CO��b��f��w�\K?R6����&֢��P�������4��}]����½��7p�e:�Lw��Iz�D\@�c��8P�&��"f�+0K/b'#@��bt������@��L��:��^'���!;0(Y^v�&Z�5G����>|�Q������0�75v�A�����ኅzh��>u���P�q̳��e�}����xb�!}b�<���3\B�h�u�b��#_i�I�fh4�n�CKmw�E��b�������\�]��[tY0u7��w����p�y9˖AЁd����>���:��ĻW��/�k��N�o@�/��c2��o{�s�� �LivE!@߭�9�֬Խ�h��$r!��jb[��~=��T[J)ӆ�� 6��4�S@L ��^�~�Nߗ9���Z;��qU�cvP��9ʂ]�y��u����S��Bǯ\�8� ��32�}��C��"����ę�������}���F� \��Tn$�r�i2����5s�z��,a`m��o��K���|����[��Ф��$uyU2��jD���������C�ゟO5O_�Xel�5���䎉��� �����!�wR����+�L���M���� ��e=�R:S�����!O�U��-e�� p� �)"�f5��,��y��ۿ%-K �V�@����m!QO�%i��l��8��/�~�<���,� ��}���E�����+��m��l�\)���t��7�8	l�(�3�2^�ei�CcҒ�il'�x�jw��g���{�Id�#5a�7��A�	4�y2n�]�ŠLی)��͂��;J��?����ֱ����A���y�,�Ja�~��9:E4�i'������I��Vt���Kր,Qw ��3��w����(���Ǳ��~������Qo]��&�4c��Quz�(�,�N��6�Qh����A�8zH:�߃C	��I�"�4ٌ����s�v�"�pӾ�=��h�&�kA��R�wm:��x�j��^x�haV�I*t\RWl3�G�W�L��_��%��� �-���z��-�"�~5o���F�g�[૨�9k�#-�9	�Ţ�9j?�bUr)�=�7͂���ၲ� "��n�O\$P��s�_��m|�LvV $+�L��Յ㍒�Ȳ�Ȉ6x�	�El�pe�ܴ�S�,����-�45i��5���~M.��\ڲ�ڭ�1X�S�Xrw��2\�A���<�����G[W�L\7 �v�&dp���۴�Z��o�;~N��0,��/Ю ��O�M`�@����c���6<��L�XI�>U��f��:E���Q�o�N��v��`t�%�V���QJc�.|،�x#��y��� >�f ��X�0���=�0�bW�05z�w�[����_��ް��k���va��p��â-�9���J"�k�v�u�#[���KlV�"�u=�;@S�N�E�gE�]�9'�&h/ڸ��(�k�p��	7���Ϯ��r��֙�0�uN�{�%r�UD:nni�@'�>y�8G"�Rr�Wo�q�Y����H|����$/��?�[�<���\�1 ʫ�S��(&r�l��1z�q���#�8^�j�bKxѠکV�A��F�R���h��0��ub|K �L��w�V;���)UHnk����?�!�ւ��Z��D+��4iо: ���g�5Ѿ�Cl|����k{�&�nܽ2b��`�B��X�
s��N~ϊ}
�F/�+]�TT���b�V�ؚ���_9�(LD��±c2�+��p
�u�w�*�l �5���^(^�n�CG�ׁ�Y���&U �o��'�� Xr�\��d:r㽭C:��a�^���PK�[dО����mA���t~��Y��ɔO!~HY��(�����@@�2��kh^{�k��gr���Sj����Z��R�7W���R�eRt8��B�L�}�� �̠�O���0	$ ���O��F�u�7�n��R3�	��N��Q��5����:�j��ȥ�q��;O�����8�A��#{K����Չ<?�X13�Gq�Go¿��ĬF58�dj[�:C�����3[�����m�ޭ�[&p����֒
�7�i8�nb
���Ճ*�?�I�2��75�%L ��b���)�)�d�6A��S�|6���������V�,5�AXR�����j��ʗ Ku��� BJ��Sx���){�ޏ>��_��!�t�w�e7� ��.�+�����P�fǽ�=����Q��a�^����84�p�������6K��OC2Y*�?'F�׬�]=��6c0U��	��[��6=o��T�Ȗ�w�,���%�����͡��}4����hý+Q��$e�2>�H�c0|+��=��y$�o%,�DxR/ ���`��Ie΃tygn�Y�@�R@�=�m�������j��ޙQ;�eC��!�YV�;�$Z7���"�2���ӊl��a3'�1�%�+,gU*l��S,�(�v����ʵ�Pv_Dq���cH�Gh���5/T<Ke�[�׬W@_K�5
VB��k��	4~a��9S���a��ޥZ��l�������O��M?*_��%���0'�->�*v&��}��?�&4�rUA}rV-�"�&���L��g��D��V��15��=��C�o�������r��P�CB;���-q˹о�Gr�q��Ν���̸�)�d<�wOˎp��P٫1�c�{E/m^�S��#�1E�Z�.�v9[q{�^�0b���Yd!�^��F>��Z�FI
�<`%��4LÑ��*ǔ@���]�ڧ&�I��j���$8):,��Z�|��ke2V���9����/y��,fd�������B-A@�����`	6Fs��_/zi��vnN�Dg�~<�[��U�z4����[�&��8liKLDc��f�\V���s�{��v�0I� ��,s#��ZZ)�*�H�}-[���;�C������]o��U ����u����`H%�uY~x�D�^}����|W֝dN��cVU|���DP���O�8�o\�L ./���4���*��ʕ�Į��Z(��$*XG��o�o2tvg#FN�ڃ�!'T]��W�V�>��{j�ti��4�\6��c'���V��Lk����\�]l8�K�$Ԣ����3L�P�h7��S��t��5*��2��X����Q_Ġ�
.$������]�c�,F�d,��rH��h���w���>^����r 65�v5/��@ g}�!��ܘy�����0,�M�-c�BK�B��IR�nn�,��fL����̼�
b���<@��ɧ1�)P7�4)�Cxjۭ,�H㉥Z���2��-��焜��A�S����ҲN�k�m'��}�ñuB��Abi������Jld�~�n��eB�?#�	o�m�^��	`�U�fSr�8�f�ր�����������1&�sJ	��}��4h��c$h������~�,��h�Ҙ�����t���%�S��3����ھ{c�@	�iPn1q��#ݴähg�ۈШ�lU
�p����h�g�	-��)!T�����OD���s��,���}T�h.�ih~;ev��Y���ǖX�$����Ub��;E�ޒ5�1CP&q�� L^]`�>�xI��J��Um�}\9zx���@�q��:��o��s ��$�(i���gK����S���Gפ%H���lܐ8���q��<���3ؿ�{�����LG_�<q����נ�I0z����f�$3��H���iE�1  ���^�k�@�)��#�Fah�$��2D���6�@Cϙ������"B���c+��7�hG��v@�
_��#G�P�����w\�8tm\yH#45yv2)��V�&�����e�&0P.�m�񥘨|�q�򏅯�p�b��{*�2��S{�K��C�� 0��ɱ��P9i�3� 蝱�^#b�g75�@�9��I��BѤ[	`���M�O�Գ=LR]	0��v��9o��~l�~� R�� �,9�>��2�CC�~��Rl��9\�����-!V�%J�_2���n���6��@�V��]k��"��h��1t"8�R��ԚP��Dz7�["EJ�_]��=��	y7*�YMW<���ݖ�Bg�@ZA��Ӹ�$ܒ�!��Cqfz���.���did��\����F�X��,> ֦����H?�W�ej����8�< �6�����v�v�'ӄ\�.����G=�j�j�}G�3&|C�	0�!���qՂcS�z[X;Aq�|$Cm�M��Z�N v3e� W	��e�\bOL� P�ǟg�V�c�Lb������2��اv6E�n�)�.u=����hDU[��$؎�/�Ud$xH�6��A~�U��4�3��Z��bF.%���4~�}UM�K����V bg�y�R��W ��@ݜ]rgJ��_u^��>�	G��
�7����a���V���;k`-���rH��R-�O��fD|���<B����&+ZE�*�i+9��/����M��$p�9�<�F��oh �%/M]��������,P=��G�BF�0���H��5���ŷ[����ڐn��$�`��3��K|u�׫`���U���s��%و@#\& j�~S%�� zπWE}wkw��J	\�Ğ�����:2*m�wH`>&`rw{3apEt*��H�(�'��XYr�W������3J�δڅ�(�D���-�xƧg����]W�"�����?em�c�X) ��� .-�_@�!����`~K�k�@��{L������>�(>�u�z�ry����o�W������ _a�vt�����푘i(D>7�\8�id.9Yj8�|_�b^t��9������v>X��F����ϹPѼ�s'�jP'�&8�B"f���W��sA�ᰔR|c:ǌ��y	����
�x�C��xσH^��PW;����w�;��9jܒ�^j��/���6��%g�T��p�y�5�-�������P9zO��9��Z����'|2݄8�ו$�E�	�"�m}���|+�j��0'q"�1������I��"c�FF�g�S���0M�Q�����!"�CTشD=r)�ú9W��=��V����#v7���M�	���w��m_@< H�cv�=�YO��%���(�����R
�k^٧�<�K����Z+	ߍ�4�ʖ��;�9q���}���s��	�S�8E��q;p��0mJx�sl�ڱ{��N.��U
�S���;!��0��4B��VĞ�N(~j���Lť�<Yoa{E��;_��n�&��i�l�*Q셼��h��@�y��p~��5�r�BI��,IcHc��cF.�Р/�6������E*���j#b��8?��-�È�{4� ������{����������$����	g �����Ѻ��~ ���J�O�!�ㅤ�,��� ���H��>�����yM	���Q��l�7 sv���t^���xU��~"P�/>(D.��SLn����޴��Ӓ�׼Aw?v3�[}稏�Đ�˔�B~3��5(S��9�i����1��C,	���	{<bD9U_(j���n��߶��b�u�9��xj�� ү9��(�]MlTȘ�lQ��F��?�e�u;hP
�ʪ����H~lO'�D�]��/�����#�{��E� �t�MC�5 P�`5� Sϛ&N>��

nmz0���,�>�{VF�N7;�y�K6:}	e8Q_bʬ��\�i/�;���:��F�t����i"�󧓘@�hڟ��'[�FZ1�FZ�%6���A����m��Υ�toE��籾w0 E�]g��%]jl�j��s�\��� ��ӎ#Vm�^�U4����������F�;��^Ѻ�"z�����茠����R��E���ꯆ7��P��ms�a�����(fط��=O(!�g� �y��������������|+'f�݊[�9h���I�{ ��(���I�4�̶;^r��G5Q�)d��\$�x��ebI�K�Z�i��P�.e�}������hK���N��]���2R�	�ҡW�F����G>��B�,�$��˽�:�e ��IgX�A+�U��y1��9�uX%��#y%�����
����B�@�'e#4l:V(�����)��`q&z�p$�:�g}1bKyh~��(�H�N�d`V�,f�s�>�g넝aa����*��0C�5Zs��Ȑ�+'�1�����*ă'�~b�*�?D�44meB�/7Sa��U�5�ߦ�a�.���};v��)XF���81�������%�ui��&��D�k��?|;o��YwC��K�� �0f_�	�#w��c;��{�*�ۮc�ٷ�M	j�2Y	��T�)������jw�h���ӆu���`�π>�+$d�E��u(��#;�:�hqa?e�������ʑ0A5��uC��n�F>x޼!!�zm��������hbu�A��1��|�����䛏yc�)�U�E��k�}��"_���5�nă���$E~�;�'�_E�*���������2|�K�r���Ly[�� ��N �����=����fd����W�'���2;ѤFN�ݖoS2ƛ���[]@/����1�h9r���Nz����c��U�L���>K+�9�	v��Y��F���BK1�*�g���$V��o'�	s%����1j�^��Rw�:G4�X�q�R�d�yc�\g���:-�'h��tO�U�Na��d&o�-���}�Na���xpp5��:���ZR��������c|
3Ŗl�S�kDŘ�*\��2���d�*���ݢ�"�Mj͛oj�?rNl�5(8���?a�z]��W���K*��H�C���Ê�v�܃�������>��/i*�L��7���i�Z ���%[F*���y�NR�|�Zx����Tm�}�4������=gu0Td߂�����+�̗�h���VFw�����vJh}z�ݿLC��FNE��I˜`����qK�%�x�� ���r��>k�[�b/����H�=�g��`|�X`�3f�������_C�%|5�������ކ���o<�̨L�d�s�W���N����%��p��aձ�,���H��R`3`�k|� \�N�6�m8P^�+		��8�ڏE[��GRB�Ԗn8u[�8!������eɈ`��(��%��n���=��/�4W7�}��Sgx��4��c�ڼ��8)��\DoR�FY��V&ޣaZ�1Z��:Օ���4vb��#�j_�
�p)覆�A�ifz��B�M$���-όn��Y�^��3�Qb��Bb����.�5C:<^�/�]�6�&J{�����eE��9b����v���ժ{�i��*��|
|sI[���6X:�~:@�9>G|��㧒�
�E�e�p�����A+�I����J��W��8n�T�0�e�+%����/S΅z��Q$a��_��"��hgO[5_���n�ս���}x$�#��+V��S�$�@��#{�뮁W6I�L"�e]�b<�����B��ΎNg��̪��s^\��1E������(�<��kugF�y4��m������8p=y��O|�Km龸o���-�&/n3�Ϛ��Hm���A5���Z*�mȴ�ω"L���>�V���O�m�A@�J����Bp���ӰV��FJR���$`��'���M����sBN���b����&6��A�z5t�����V��,�xju��S��;��dK\���398O����ߞJ�qN��Et�"�ܳ�JB6�H�d�ϬQ��i�潢N��b���7k��Z$��OPVb~��i{^���K9R.�)�^Wvf�۹�I~M�NK�ډ�kf�sc��B����S�2��Fo'�(t� ћm���� ��'y��g����m���z#0���e;��W�;���e�k5��Ȇ��R���L~�`��/��?�� ������������0�
�b爏~&�*%d�Dp,�T$�Y������u.�H�x-���<��}{��{��̷�u���6�B铄����ST�p�&��\�n2�N�����C`�?��r�a�,�h+�+�4@���,cM�$?D�����<�/�'�
�J\n;�3��c���]�=�fM}P����dY���{� �1�S�C��Z��P�"@�b¶x��.R&����ߝK� ��+2�
W���XP�M\k�����L���̎�2{pb�wg׵�[n jJ!6�{&.^a���D�+�mf�1����YZؤk�}}5�
1�?*����.��Q��t���}�ҁf|�n���i��S�Ո�痍;q��{Oj*���m+��ōp&8l�����T��k��h�&�KCƼ�;胚��$j�������l�ߺ�P�G���h=�ûb/�S�t��bb�TvH��sKu���֒v]+'g):�7Ҍ
Q�x�}|Ș�Wh���"%�����cV� f2��������>?�	Z�s�&�ZZ�6�0rm��i��i��W����~�G��>�9┊t�O�Ԕ�z��>^s� p)٠Dj�n��I5Ne�O��'d�ˢ|Xs~�g$Y�7v�K�������￩P�լ},5�����y�'rݰ�Η!x�!�~ U�,뮸�J�抈���?}h�.f?���)ׇ����ed�j�؃�L�#s#�W�|8�{��I���M��¦'���Љ�?q��)��dSW��ˆ4Y!N�� F�w��������9L����8�W:�{B����cZ��5J��ɂ86*��K�b��k�.Bg�wL����U�$A���ڊQ�/��"L=��n�'�h唸���77xq������6?w��yC����i1w���W��s_+laNz���\M��ΐ�1=c��7�w���1�͞��3)�<���I���n�*pS�԰����"�S��p?����;��²�7�j�vނNRA2�RF���A�з����A8�^�d�+r������hK�37�������N-��Qp��\Me&��;dE��Rͺɯ`�����K�_�N'�Iy?9H�.� �_�n߲{�t%s8�qS/����>?��t�	��.]Ic�'�����0�����T�@A����/K5�s6e˃s�;J|�IK~�:��b��׬�(�i1;�D��þ���8fK%S	��%�J7#���ֈ�m2e���q��o�Ջ���֒�Ϋ�[΄���n<B>����\�Ӽ�~�#H��~a�����������f|�8�M�����L)�|�>�xK�u���U�L��{�jIe3��K�JBCSQJ���[����?�^K#&�,��&Lj��+=����`���%n�ߐt���̨��P��65eW1�-�GQ{P��޲�>s'�%��~��o,Hs�a���T�PM{���P���%��7!�D�Cq�"���H"E �+l���ݜ�̓�{���瘏��5@0�����S$\ �ϡ�{Q��s.i@�t=@�����t��E�9ql>D�'�{�ݛP''�^�t���}tI���o�_� :��|4#�����N�f\E�2KqD�b]��aF�
J�ϩ6����g`�SM�BVcRbv�5����� Uߓgn�/`��/�T��K�<v���*ߔ�T�s�p��*���M4j�j���`���6-��RpZ�q^�Wt�����b�0�v�)��ư�l�c��G?�\�&�	�ߐ1w\�Pj�i�Θy�Px�k���j�ɂ�r`S�B�Ǳ�Gʬ�O��Dxp��8dp��VYuZ8� �����0��kG�:j���H[��{n�Jٴ�����|�P ��T}m9�(p�}�K�����07��"�q /!P!:ʹ�����dss��a�p� ���p�=&��pM�&V��͆[�[9���h�e�{#����j)��I�8�yAkTW��N��Qm	�z�������p6����n>��1�`0�2��s�L�ӿ���92���J5*W?1�O3҉��#к�;�����{3�
��N��T)m��&"8��ӤbdAlQ	�APw����[�>]���m�wE�A��%$���az1�dW��N�T��a��Ҁo������C�T�8�5� �I�S!]�YUF��ɇk��H�����.��͠o� U{�S�ϙ{-4Ap��!�������c�yI��S-�?u�s O���?����=�����Ij=��dP.�@�$����ZL�D����NG5��1��'�.$��q`�=<�D"x`t�p�� vn�^$�\L�����AP/Q��[�`e7�7�����۶q�x2�
.�4n��<�Ɋ���w�4#B��W�¿OZ|��sw�
/�%o��)�+оɺ3�L` 8>}���)���鏨�Mz -A���yϏ$K,�&@�_]a<|�t�b=�RN�!-P�0 ���$�n�>����H)�єnԸ���$��G��C�f($X��AG3��`��*��Y/�i�����-��MFlo���~������7��u�83a=|�/�/�^��$U��u0E�*0b��Gq�?�(ʺ�	�Pюnܖ{ȴE���cُ0�;�� �����l;�	��"�]SLoM�����Ɖ繨��X$F���p��nS&�f�
/LM�Bx�W��Pl�������+ ����%��^Խ#-�,�E^��jUW�v��	y4�L���gŋqI[�"��	8�Х�o3�%)�H����5���7�<H�	ji�6����j���nl���{E��~�ĩ*���ot����5��� ����p����K���'m~��cjx��!��&�G�H��.�,�������U��u�O�V��dB�["���4(��?�>�����i;����D�ۢF5#��x.Sp*g@�<pK�K��TY���;rn%� |�j3��]X>ʅ���a��~�;��u{��+���i�A���X�n���׍����_X}��n�� �V��zMD�y����A�!��T�$"q� ��C����i�����Ma�Z���IVi���p���l*[�g_��<�<B�����,:�k\�?���_�`��~��7`@�L��.����$n��U�2���G��s��^X�A]�U��T�k9�^�P���sH��lm��t\Q�3�k\���L�>�G���]~�T;ϖ��D�hJEw�G|��g��Qᇃ\�G�G�v+0V�XUD5�
	zD�gVaQ����m�4�L@A����֔�|�0-In�\T'�x���J�Tt����N>'bj��u�,u(�**aZx�����r]���4d�%ݤ�6�cW� �ɑnՔp/���Ǭ�sl�A���)w8��va�1���,�±��2�M΁��.]�.>�ゴR/��.���v�����B��2���&W�&�?����Ͳ��F��}�z�-Oh������_�Մ��ӕJ6�m���.����9����!&�O8�tZ�}!2�ޮ)���.p���4a<m�d�R���ni7��TC���;��g�n s�wK5��h�P����(0��´�_�OT}�{�TtX�_'������`�E��p��2�A�Sp?{d�I�q��q��h<Pu���;6�� �L�����z { {�	SN���"�߄w,��ⴢ$O��p��VN�f�~�vW�G�]�������?�WU�;��3�@#^�T?���K�/^�0SI�h-Lv%z��c$��ˣ�-mm�m�kA���yFd?�߮���Q�Fd�����\J���?���>'�F����{��v����R�v�Oi� f��\]rKS�կ�B�k�䉸f��\�2EE�Y��2i̔pI[�ĥ�~&��t��f+����` �ڀ�Ֆ���X�yUP����FPLp��? �d��y�;L��������Tw����X�Hc�y9�y����j�����GV�Ŝ��en�GE6��c�Ŏ��/G,>	�f�GH�ƃ��ӾPxUcB��S\�Q�dd-�%�;P�
�S�d�k�abX�����d&��hD
�k���(�}���.J{��om~[q�{�Uƫ�����GJۭ���H_(�L�q��\v��l��TKߍ��+^ �'�|Oe���yӿ��f�W�h]x���M�|�39Xɍ��u/�y���WNϏ��8B$�z�gKh��c�đ#K�֋q/ι�AJ��v���?:��08�(�뺃�������Rp����@C^�	nqb�)��h��.>F�(�b�S>�x�����-q�1T�vr��ѭ��Nk�|:�_ձ`_��*�]E>���^��+��t�&,q��F��Kl��,�����eq��Ơ�iT/3��m�/�� Qc�]�۱�g#U8f�W�v݂��0 ��\�o��D�`�#(]��r��+&��ܺ[���G���,4�(������@����7g�X<�^�a��e��"u���~Ɍ=���9դ��d0͔�gߡ�Z�Yk���WAѶOXY�����e�����r��T���[J���@$@�╾S\�H�ǈ;`���̼�`�y6K���3T}5]�[IY�G^��
Ԙ1�Q�6��!�TGC���M��b,^�3Ƌ���F��(lnU��s�n4��k�����I"88�A�e�`�G ��3P��Y�&M�@Ɨ|܋mMFt�,၍B��J#*��@��N�F|�.���Tc��1����%�*4����{l��:Gƹ�J���C[j� �rZ��yM"���g��Fe���_�1O�nA�܌�4�1�.��y��0r~�)�[�����˼��%һ4l��v{���U���j����*��ꨔ&��L���W���3ij����?�G��;��4.A��
�[sztL�M�t���b�����/���4�Io(@�găC�4~swP%B�ZA�`o��MS�[��HH~��v�
A`6\��n���������ew7�@X0��o{ռ�T\D'%tX��Bo
�v~b"~l����Z���UN�4���U񃶛��8�CAv�/�fc����.~�x|^�lfe���a�cH�V�ɮ	�E�%�5����y�����t�R���W�@q�����r|��E����rSq�=��M(�&K���&��2�v�u�������p�j�"��ǚ8��+�ӱ�~6�%pf���NyD/����w������|��`�*'e��Yu��cg�G����@w )�zĤqz��U�%��n�F�@�av}�h3�a�;�{� �r=5�3�@��ec�جգ�*������Y�1�驞\h����kt.��0aΩc(V��/�_u��aЌ�� ��`h���ŭ>(�\9��W���n�	��>��5����,����U��5��.�u# �x��𕕿u
L��́� u�\N�US���t�vw�_��A�B�:$����Tg1�<6�2#��R �ӫ�٤��ؠ��V�.�*�����a;��b���l�e�L��,���
�r����@Gx��FjL'��R�[كƈ�� ϴ�Q�k�h��c�=Y��ch踛b�&>� �>��Ӽe�\V���@"�m�Z�� �[�!�� A��q1#�?H�H�l�*�­����O���n-!�Z^о�R�U�����6�q�ˮ�|�+�3�\�<^��Ga��<�E2c�b;�#�Q��޷*�ɿ���A|q���k�:�J����w�@����a��qv��MH8�1f�Lܚ��p��p�'����+��yg��ؚI� �H&.��I��FӎJ�R�;맴W���.(�֫9������A�QK1�%��� lk�A�_[�t��%��j�oc�ve9���4~��ϸ~h��ӻ�t.���w�m�d��zZ�Uoz1 �{���dŹl��,ʁ'��>Nș�[���h��7%j�o(��x�GZ�w�` *[�@6A'�������y�i�ԫ��� �fCm���,�ܔin�E�\Y��Z���ű���o�.(H�j�ҽg=��5%
��jF��i}/n��
ךF���b��MG��kc쥉�q��� ��ɚLG����&@���6gMɼ{J}��&b�7Yc�ʩ���7'�6�$E_5@;Ji�j����i�B�+G�,Ž�,�ۥ�\e����B|��_/��"}��ܚZ��}'o�g��}B2.�����I���D�*���������ـ�c8����3qI�Զm4T�ر�T���Ê�R&uVo�#����q�g������	����2�U�/��0V��)w hkWQiI?l~{xi���2���I��O���ȃ�H���E��g׷k(,��D��<�Q�߬��X����?�_�8��~ ��ٍ�"�2�aw�`�j�⼥���c��*�]��1��Z_yI���NC0�/�خ�H�Ä�|�]g��-;��[��YZjwJ!~Uy\�n88)���.'����-�C%�?�+��]���	gH��|r���L�fu�k F������C���zM�v�|�f��	^��P͒�M)�v㰗�!4�5fS�B>-]�U��2�I�g���l!� G��Ͼ��h'��Th����LTw���k��r�:%=Z�L��Gz؏i���gk	���I�{8otWX�ތ�Ɍ�����l�L���V��$��=&��u/V�i&A5�a���_�t�3L�`��
��>���mW�k�����o��A��?*�����ǣ�hʰ�����Y�e����A:�)و㊖=^��qT�~��k��,I�<�^��1��3�%��ړoa��˕9+8���ћ�}m��9ȶ+[����%Q������(NV4+ws�j!�.�B#���ӎ�{�E��lnM�A[_����y*��JY̣�t y_����w���Kt��'�d����.� T2Ce��w���=d��R�FV=�s5�
�F0&�fN��{#5�rB�4�=G'S�unZ�'h��G0�u0��2�)̉D
�^K�J�0����.�r�@z�X�u�1��ۖXa;rru�Թ�!��2���Y�0�ɗ��ř�LC}j�*�4��.H5Qᚆ��gG�8Oa�jI��=8�3�O�H�� v�}�C�?#�k$?���Y��H7��m�@S��\�z���Eck�#���ؿZbJ�9����(sQ�1m`�i��l��0��;��^P��bb}�^4�
��/�?UJ�?��?�рpI��2������.z��8���D����,W+�<������9TXs���
����Y�-6#�b�ْ$�c:׵t�*��^͈�"�s'ʶ]mlM�SRf&P��}L�#�&MkwB�Svr�@�����͔2[�Ib�nu�<�ac���}��İ�2��'�iJ�����	����طߏ�RA�Q0�:I�c��ըu�p�2�7�����g�o��	u:.B�kwFߊ�
�)[�`���f����H�R3=���]�`�|�/@�/� 6����gW뒺u�OΓI u/ɓ�s��/��P���VP��P���xKm�ri�z�E�m	�|�8��(�2�72`Y����� \�\��J�X\�X��D�w3��`+ЧGaU����(��P��n��rf�)�{!g1��BVcI�IXI�Y+˨��|_C��e��\y*JY��\
���s~��Z`��}̭���e������+�'5K���A"��w\[����cϒ7K��V��9���m$V-���� 4N�)}=l�sd׮R|7s���Jˁ�I�Z�v�"�פ�nI�"��U�~�[�ށ���]%`���[�/)4�.�7�$g��Z���U����d$ҫ-���@t�~�LDS|�ۿ:��J,����t� �];O�m�lJU�*�p٨���l��0L/�Y�2���T���]�MQQr^#5n�6��>���,�c�psT��P�3�i����uZU�+k��� 6�8P?"�u��:ky��пى�b?ך����cD�~���4�	�_�L����E�*�D|�w.չ��^������Î�&��&��<dZSch���z�w����C��>2�0���T,��i�sʮ��9�NBb<�H`ם������ʘ��p���&A�'+��)�č�w���K��F����@th�h�ő����$���Գ}��<�O��T�Y^�QW� ���ɜ�H�"��i%�����p�株��3��;9L�P	9����c\kā�}ս�l� rv߿4�-��R�[��%S�e�7��*ۚ':�k� �ը|�����xiAX2����W�X����Q�al',��/���|��l;��ݯ���C�r[�0������#��rw|��F�-l7�WJc��X����,�^=D����E���oG�5���beُ%꟟�Nv�9�������a�P���_^�����' �7^��ɜwR��: r��s���"a.t�Ř�}p×LYmb�(�}�ي�܁S�-��K�(�&Z��oj/�ӊ~w��F�X,POȊm�m�e��G�P qU#^��u��56����(N*���@�ǳ�pCh�!]�Xg�,��������A�����0��L;��9GxkI��D���3��)�Z #ްF�lcУz)2T���<N&F��>A��`��0�(�>v;�]I�:�j$�붩�1�IS˖����@�m�k\����B	�U��h5�R�H�B�~;lH6V���w��_� ?QG�(מ���E�/UN)��S߃췽���sb�z?�U���@QW�|��Ϛ[�2Vo2[��j��!"�M�Wh��Y^ ��O���ӛ��<�������ѽ���6c�|݊�MVI32��<4�\�;�va�]R9Kzr�p\��x��H�7N��r_�*ou��T��8� b�T���ߣFZ��[��C�$͡���wdG���GT����7�5IW�`qtv�����ї�W�XW0'`�_rO{��^�Ӌc��g����E>��=^�	�"��q��M?
��>��L�D
�*����E6hߣ�2ԖJ@ЫXA��Y[!�=ҩ)�F��ݬ��2��4Y��"RH���xO��3+E�b��D�g�-�#�Ŵ��\���q�E�{:�O�0�E����m��⧒�Z8�"+jS?
��9����rjxY�\�}�K�#�%�#��ɼr	Q�����ƥ��dD �,��
�!n��A���`��*-��ы�=�KwE�r1Q��&�(�f�t�(:�쩬"Ŗ;-�T�`r/���t�D�5ڒQ�*����	�O�(�������h�>٣4F��o���-�C����z=a�����M���Ẓܝc�px:9��5=�+jG���Ø�1����p6�}ێ�Ľ�3W��H�7�@_�����y˖�>i������&�����f��.��ʡ_��|ܡ���@�J��a�<�m�"3��a��^��sȡ�P���-�'4���]��8S�舌�ӏ&��%��Ov��Rݍ��Y$p�
�{�ѥ(�|Y������Wb��E��8������Lz�#PC���@�TFtwΚ�8�)!���&#�#��E����Á���4|pt
��dc��AZW�
��	,�'���,�����tSG+MO�נ���_T���ӿ�Y�譾׺����ϗ{����T:@3D�zw�SSͿj(�D���5����<���go`2�}�s&��Ǭji@�@����/=>�
:�{iz`;�|�բ)�L%4v7�b=�[.����/���Q�Z]�un�;���:k�f���>IU�y�C�,,��5��1T��Z��|*'�,�T���_f�*u�T��p�X�1;T���
.�Nk�XqLb��H�D�P�i�Ol�YZ?�Q;5}U\ � _�����Iܣ��Op9��μ�bF��[OU�������v�d�؁�a1^��f���)�	��U���l�����Z���(L�؏O�4��%7����K!��Ћ|Ey�-&q�-�Y��Fv_,$�KQ�ȗ	��!�_:�����M���d��r& 9��j��/��A{��!���e�Y9��H��;��H�&����A�8�2�֝(�)q�+��ǜHA>K�⮠,H�$�C���daG[��>�[��(�0Bz�q����z"�Nc��Rw��X���d`���J&���\�6�a��(f��V��Lm2��U%��w�i_�,�'�Q�Y������<vGB!�U�ߕvt�:"�lg��R��y����C����i����$�D[��0�b,ѳ�&�;�aͱ݈H��5�<[��5RTz�ݝ�@�R	����@��v���{CӦjl�+��|g-XȚ�S$58Hj�:���I���̊�Pe�s�X��m[�	���8G�5�J�@��V�]C�	�d�ip99]"j�ϋ9�`��Ve҈FjZǜ]'�$��f<�9Z�y�sZj��hBmʭ��.t}W��3A*#�K��Ҝ��/�Oꦼ�`�/���j~X����"�8�� M��?���Q# M�ɯ/h�x[����̲��#��u��p|�����o+C�T�+����\&Q�=�oRQ�F��)^J��Cm���L�1��2V���r�� g���Tk��o+����t�ɘc���sp%�HqiD��� T;�bP��:줯Y�Piv����5L~�<m���2�h(�����������xS:!%�eaU#�>����C<8��9,��&ۦXOny��p�h�M:η,��Om´��;���:�y��)�a��b*ϻ�a�����Q�豜N�HU�2ԭ�g��2�.�:�PW��=�gU����BZ:FvK
Z:��uǚ�����"�ѲG�d�	����!��,B�
�ADSW����U ������4EAB��1\�(�9��R��Ra�Z��������M[#�o���D�`Ǜ�� բ0+�\J��({�e��f`e�P��n�4=�z������`�Xp�1��M��Ns�����rNQL�ܽj��k��q�|�G�}`ɋ[ &���*Z�K�U��KWe��(�j5��WO�8�3��Q��9tB���F�*ނ�M�omC�\)r�J`��&7P���a
xƎ����(_���l��Oi���Q��^H*��&�Kl�U���u��#�J��YdIW�C��t���|+�Z�sP��=���C�<mދ^����(�1�����1{�*�)��3��u�����5vϙ��e�b[d���>�T�ӿI$0B��;�����)d�P�%�"�_���5�䧰	��Ay��~U(������H�xс�"�B2�Z�D1�Y�if�A$��8�1 �u���z��d�6����0�?$�.�49�z}+A�[|�L��'e��ߴ�ܹ� ���F*`sfm�fI�O��MM�*���l���F�c�Hᑼ�;��z�i�ME52�|�. I�$��{��b��ۭ��J�����'8�my;x�M�z{a�6ԓ�^Gw�<�\�lQ1��&�Ӗ����r{R����C�����*xX~�v��>��xz�8�}�V�o����:�� Y��&9���Y����j�Y��j��=f�p�nq�W..����G8�F�~�|���F��x��~��5�GV��~��Z�����,/�׋c�� �2���2X6!W�$��h+�}{�8s���a��T 4(�bpE��HԯHˊ����\���!?�C�8V����v��Z��%G�]�d�p����-sJ�&�a�OW肀�m�1���\�ό3�WQɌ��p�9Q�^�j��[G����qїJa�����2	�6�Sx�/����,�!�>p�j�)4O[��m��}����hƌ��/%��l07[�B�'�İg5�g�?5:��_j�8ogٿV�B��{��nWQ���w�a�D���&��8�KȐ��F��c�~;���� �	-M�R"���L�|��Uř����Cn<��v�������Y�{ى{�t5����<� �
&�HY��_jR�9���1R$��?7���,h�5��'g<4�e���}e���..��H�K��ȶ�Ăb���^氨���x��xTd-��4(�3�lHh5��Y-��B�_<�TO�i+V������8�����ڥ��(�������wB�|�&4I�n�ډu��!��2tϽ�h־��;a�X0F%��Or�*(�����4���G�H���6��������J:��
ת:�5�!�_5���s��u�.y���[��#�S�j�A��C���]Ѫ�2Gt�Az��i���ɤ)=�6{`���}A�x�a��&+p[dd�MU��G�8�h���ozM����;��u�:���(�K���ኮ�3�$A�s�A^ǀQ��Q�7��"=���O�C���N��wDhd�,�Fzݒ�;���kls��f��J q����E���Ц�ځ��}��h6ё��u"`�QQ��T��q�vr�ءk
��;��lO=p\�d�<j;�0�Y�&��2wDゞ�X*D]�ɛw�I��������§O���@PA�� ��6gwSY�I{�	鐦	�Z)2V���#v`�5.臣Rb���]�e��Q}y�ߵ�q7��5ѯ��(L�8<�\�SS)����q�ӓ�L.bbP	����G����5�G���&u�1e��n���6W���t:�9����]���0�ʉ~�,Т�{8E��9��	o�?n��7{cX�U�[:�|�.��g,d{��J��CZſl���6)�uS��oR6 Q�
���p�s�L�.L\��,L?gbxҏK݋�#�@��d�L�<�4�l:��2 �� �D����4��͟�nFgDu�
T=��U�g�Fx�{���o�}r���2��w��w���N:nM��&�o��Z�kydF�%������A&�*�qT�뿟R�Scv �BR����_c� �s+I˵�.Η.��������o�į2Jy����R^I�$ؗ�*�E�K
��.�gn��y8��<�(2�C��k=�;?��֤^Yo�U�r�K{�nZ�rTi���B?a���N�]�|��L���6��^}�AX�;��C@0J�=%���B���P[��Z��CS���+���[B��$|�Ɍي^]�g4q
26.�����X�j�7�o0K���Z0�;�l~-)}`����	�[��J%vl���*oP��Co�5�3�R1G�b?IK��Nm�vI5N	s�es",�z�Ѿ&`�EdS�ʬ[)�C��
R�}cDBo�F�d�Npڀ����$�=�T�E�c�#�$c
���A��]�wc�DW�5���8s�����￨2J]M�������!w�ΆW��Ѐ&���7ǔ)��{�=��H(]���6R�J{|�<o�]�5� pj���w�1x3\v�Kk٢Ӕ�Ļ��j� �L�� ��u��(g�ʝ�Եj<D,���[P��?r�|�I���<�=����J�����Hn��u���ev�����_'��|�&~	����`O�Q�Vx��X� ��UHs{��|v�.���t �4."I���7ix�#�y1tw0y!�_s#��X�(�,nj�~�T���g�i��\|�jʤe�J��Ӝ����9�6'�� ���MKV�ñ������YNANm݊ᓎ>P���Jo��#0wP�j/z8�"����+ܕ
E3�����[�;4�ރ�8�i!�U1�n��Q �[]�P��8�N@�=E�^��o����n#��yaw%e�
о�?��w��6&��\�ԙaz���n��m�ˇY���(���y3��d�.m��NIs�K�q��M�l;�/DTI�c9�P٣$ԁ��7�(c�(��s��v����+�8�]Z@�w<?�P�{�Cob![Yь����!��J��(. 0t�x��W������� ��ӛ	�G�/��sAF"��c*�A�
^,�y�p��2��궄��o�H�|��oA�T�������iI@�ڈ��^&A[<�����J�FXO��O����2���vu&\�?|?����"�����
��Q��|��(� �r�A�0q�vt� ���f�n�(��*!�����R9�o��i�f���eH�dv+��8U#w����^O�����]�|\��Mݍwq���2������ ��|��g�gR'E���I6�C�1���Ju.[����ϼʼ$��H/7v>3K�?A��]���#D%4�L9��E};�}�l�)*�����H<vR8���*[�����?d�"G
��_Vk���	"Ȅ�����I��9�J���͑��֒��{��n�o��n�h�.#t�n���F� ���G��!Zc��4�v�Ŗu�JmK���B �g��Uj5]
55*a ��20oE����|�����-���
���gAu/2�Ǝ��=kq��d+���r��l5�������5���>��c{��M9�9�w��/�?I�0�;��:YI�v��,VM��ء��Ò�V�	w�4�\�7�<.�>H�����D�e�?^�3ϣ.X�3�{�e�����k޾�<��WT�d���%B?�����w�yKe�3��vd%��tb�[�"�C|{��q��:6�=�wj�3<�0��~��L�zk�mz��J y�h(��Y�2�]h��а�j�@���ɃA�V�"�*�����I~��.�Z�#f}C��*S�Ę�U+D����D�N�������Ǭ���'_��EV� �Svh�,��@˸{)�w�%�8���v�6�rs��*���q�kb���+(!�[9��� ,��}L�KS��I�1��}`}4�E���&(Hъe�!��}(�Q&�VhD��QoB��8GZ�(��y��$;���f�P���c�i�s�xn�&�﬜�I��KmC!��y�� Ɋ�!�����e����r�Q2�����a���5���-�}v7$[n.uĩ��*8K2�7��%M����	����
+~��*��1Q�A��^���Ѐ3 �u��z��#�}�:!:B�I{�X�ϕ⫝t��d+u�m�i-�"�QuY��jS�]oJ�S�	����&�_�l�nk�	�`�>���w�οˉ�+@If�P���V���X�h�h�=�,M��/4.z%���v��A���I��Y@R��6���ZL��F66�A5� ';��g�Xnϟz ���e�z��T���,�tu�+� o}2	���|��Aߵq%��]�l�Ƨ#vI4 -O֫�8�Y�>]��G!'%M��u�A��y~�Qܱ�,GA��o{�:�VZ,�p|�3J� �,e�0��{.w"L%d������PU�w��"���t&�*��:���2�^�T��T���уU#��Ld��U������	�eh"o}�}�ի/+_h�g�V���������>ū�	�<�#�^��ڎ�L|��h����^8�r.���ٙ��U�`~�d�t�;�_���~ƧX����`d�i}�9��tf�k�G�vf�A<��><�<�1[������@��I#%���5�{�O�sG�w�&�!�Or��C���EͳuG�UW"O�R\��u��7��;��:\A��Hh>��+���KP�mF�����X��QE�b�fFc<b}���0I��ף)	=ż�8�A��jG�C�Jht�(�s�Մ��"�
�(�����ƲG0��ʦ��9���d��;\c/H��4o�)�;���`x�BN\���K}F،' h�mޔ����_$Jy�����+�0�~�iIr��}k�1����R���AK�q���ܱ-�<�}ƣ�`�ڏ�uȎ�AҜ �wpH�!m��i��~G�wp�}e��}���0t�$z���y���Y\�9�Gn�n������1�+�Py
s�~�(49-�b69ʱ�~� ���b������!��	{V}�q��g�o\��/UC�9�*�L��?7z�I�j�^#&.6!�C�3�V�ƚC�����?�$\�?�:�s*Oָ�*5���qoU�Rw�p������i*W�lC��Ϟw�8C �H�򯙘�4�py���R�G�f�{[��M)�b��m��^�����ZL#<]�7���02i!l�� �ͳi�@��s����$�1�q�=�©�5R�
�s?6�;cx�?O�]��a]��mi��\���5HP8��j�X�7~�b�𲌳��|��嵄z�XP��w���=q��J��!m2/�'>�F0}�1얃t<�1���͑h�A�R���U�q����-���X��L�)�,�� �����>�(.w1&�	'���
�����̲VU}���}ɾ�O���j~|����+{�B벏ɠ�A�+�%�n��E��#�c�a{�\�����ɩ3�,5�ˑk�\�&�D�D����B���|��GRվ6Ǜy�� ��.��11@ϓlke���j_��Pj��)��ۗ��濥m�Mo��p�䍚�+�L^��/��Ʈ�-'B���)h��[��y.kwpa��ך��]cq�݉#�����X������}���H	��軫�\�
t�G� �6�瀣��Uc�1b'�	�\�����n)<Q�0�T�إZ��?W.TZ�mI�D����1��D��CU5n�Y�b��4��n�qb0�?�h�udcS?:J���G�]�^g���B�]݁���������e�<i�����QTZ1I��9�(t�N7�&�Xò��`b���j[8�L����ޭ�P��]t\cPsV!l�+ߩ��hy�D���z�珤���k���~#C�ד��Ф6���[�M:����$;<��B��ʻ���H6p�_�����/ةK�tM1�t��Z)���f�d�-v������@�ç����c��ƭ����O8�7hg_w��R�"D�_���I�i�|pc���R@?���و\n�����?OJtcG��p,laeM��<J!sf�H�{z?��Y&FJN�������ұ
�Y������1W�?]�x%�!�®~�~�@T5���NM !���'�'s�e��囃�oL�8=�J��<k�E���x"?�i�e�ꤼ\�X48߷������|�-$UPQ0Nx��u�05��IcͿ�Ĵ�iZ�n`7i��F1�S[w�9H����XD=��M՚.\h/�Ʈ"g?��T�
�n{)A<�/Z���ٳ���F����^僠��v��V�IVI�$�P��[��7Δ��P�F��YMgp��K�.����x��
<Y/5f�4�o�zFlp��k�^á�LuzԌs��l�5��2(mh���{�Mf��>��Q{�{=�5=�#��z�#�(6�\Ul�ut�JO���!� ��Z�A��=�0@uū^H����4#Y�,��t������4�����8�b]��5��A�O�m=!x̪�˒��n�\PW{�����i>�ܕQ��q����T�ʘj�sST4�fG~��&)�3��q$��WT���P��H���&�L��D�힀#�o4[D�脙(�<��C����y�4Bia���G�����Hux��Q�,������/�D�,LI��.yȡ�KT�Zc�}�Sk_P7%M9�D��/sÅ�d5���sF���,a��.6$���nq'@^�Z^b��o�)8C� dA�`��8<�:�D���Tu��h�����7��噫�M!/�@1�V�EA��Sw�,Em�V�O�A�<gI� ����ʆ�4�s��v*�~���1�Z\�a-��<��[U/���
���z?T�P��W�t�!f�+)�*���ހz�5O@Q�X	�� �#����a���[=o�-;-����n�z�����Ԣ��JyC3���E��-���:��*Sxʿ-�u���Ģ�Y�:%�Q�*Bp���US$���F�9�F��~No�O��ų�hYEw����PNء{�礌�y�@�ث������:�iO�!/�A��A5�\�ȼ�*�Ǖn_E��Q�.f�hq�O�H�`��Ӹ��T2����=�;2tfUȫ�ݔ�Iq��M@�i.ea'����o�~x���$�?`�籛��
<^���HP��Au,(�%�,�e�:iJ�{�N6�s܁rȪA�������������FmD�J�7i>Vv��^�-/O���Hԛ����*�
���0d` ��*q�
?]��Nbaa��B9�03�E�>��
�mF����**����g������D@r<!E\|p)q�#��@��������Kt���ҏ�P	;��o�Q��Z���d��@Q҇���a��}V�Ͻ�qk9d�7 ��"����A�ҿ�P7����9�b��.���}՚mP��-�@��D,7f��)ǒż��hz�j������MK�ĉ��oy̑�M�'WZ���t	;�T��4iP����3�C����n�FǊ1��)o��El{z�88!���J==�iW�1h�˅������e�V{�B��P�`� �Ȅ;1����V���������NV!��e?.D����3�jN��x��#)z���I�U �❝����%����ә�GV���<&��d{&�# x���)�v���M0�%���Z�r�e�$@lP�3K��)U>��<�&��8]��}m6>2� ����M�h���?�UJ-��R��R�z���_�{���$Q��b=[�>L7$m�㢐�\h��/�Aǖ��G��8aq��QW�p�Z�x2|\/�5j��ZHЫgk �[z-�*��f]'F�S�
��΀�̣��W	�Xc���*��t/
�ZWp�<H~YĄ�)3��b����ʬR�̜w����c[a֤ټ�'�v �����՘�d��rE�a轞�%a:�F�w+�����a���簉��� �vL�����>ٕ��7�g��=���?ob����C���ǌNVF�Ὦb��ss�B�6���9�����^"�裡�0��Q�#|[,�u�~�S��NK����0ZlK��Xj�Sw�����*ܟ�m�M���@��Wi���,w�B��� ���Cw����cBMp#qq��m4���m���ӝ}����$0n��*}��B�4A���7hv��	�.�� G�ەI5���f�3�\��Q
����.�[����Hقb/���*����רҨ���gY�]�zb�]��]k1@T�yƲP�B�������B�YBϚׇ��0��7�b��Ue<�xG;'X=.�l�0Qp�OHδ������wQMB[upT�c�av����/|o`��/I�ܨ�����U"�}�x����"���=�ALp�R^c�[��6 �������Oo���GO/�M;��Z���@v�UFW
DR���gm���ע�R����1ʹM���9G��xLc���	t��"r[Q��̜���=`��GZ�� �4̓���;3��R�hc��s]A�}���D����dI���W�~�������2�"��*���Z!as��*-W�`OAb[��n?�Ef�n@�X�#����&+��q����#L
Z�#kqgS�ֳ}��JU�J!#��}V���X��(?JɅ���|2�"�����H*�1R�"���;��Q_�D��QP޹@�^�����|�WV��b(����{�Ia�b����C��$ݧ�����e0��C�f�-l��N48�\j�^��g�����k�XC�mG�F"ޯZ�6(�����H��cD�Kצ0��)�jqh��'�-F�8�. ������0x�߇f���S���5��X�Z5OC���O�-�Ce�!b4�)N���	ꡙ�ب������r�2��}�a���#]�݋˚s.n2q�Yv�^k��V�������#����7K�I$�K��[pqj�0Q���	2�pW �?/��Ǜ���v!rjA�16�=C�3�z/A1��M�l�Vt�Ҟ�U��Mk:�ݘ5�  �h=�GҀL���G�<�z��U�ֆ���<j�z"j�;� �ߞ\G�LC�:&P�=�\܄鬳�| �AH��(ƥ5�#W�W�x$W��up�C��֑�v���I�8u�ۄ���ٴ�G�W��-��*��AP?5�y�
=��4�u==R�X��v�P��� ;Ce��Z�I#��Q� �<	���A�Iu�I=�M�B����S{Z1w��5y(j��ojl�ݚ˖���d|��ԯ�H�?��
�����d���z��]wW|+ ?z�B�TSd���W�
kX*(Gy �"5�)��
+�]7_c	AoY��qW~Z���4�2ݏ:|�3B�O���'|�x�{�
�
=�s��$Y�g�4��b����B'a̡٤8���̩��2[q�B���aV��S��!�����&�^g��&��}Q4��8��4m���r���������U�>��u���[$��Ê�oӜb!�L����с�xP����75M�t�^T�Ӣw��Sy��[M$ؠp�b<��j�)��5}]��*8��V��9��é��RP^�gx�"���O����eg=�8�4V�F3~��]\�����یy]�ݲ��'^���YQ���D.�XR��K���=���Dɏ�Ծ�-����k�r�`l*2������1+�ո)-y\wZ3 ٟ_��ɟU�h�2�>�-��5�^M{��`��}�� ��Ef�u�N���%(H:�c V݈+X6?��S�e򨞪�ӹÎ�������0>fe���PرD����Gu8�:K�4x��S��0�T1)� �6�@�Ȯ�w�}�f��GO4Td�!��]���՗�T�퍡�z�(�������n|����$��Ѽ�l�@lt�z���:/���b}?�> ��`'��a4$�=SO��XO��׭�M�����$����m��%�l�<�Ys֚��&�&{c�	)O��)�t�j���ܩ�m ��emJK��9j˚%��rG#T�n���������+	 ]��OI>����aI���$+1	"����M/�uF����D���u�jFD�ʁ�$�<A{`�ԮD���I��k��)uo��*M�~�C�Ğ?MN�w���d���5��w�\� ϙ%}�����W)�_y�s�;ɼ�2�6�Jv���i�9BD�D)LNi�^�_E3�?��p�YᠣĀQ�-��\'�ϓ� |Ħj��B�+���D��f^�t8����r���BgwB5|Q�T�	��;��KBu�Z��ʋ��~t�PJ�BF@�a<zvi̎�P6Y�@N��ͨ��4�~,��T�/��&$	��ߗ�d��h�?�g��܃T�Iui��D�"���){.��P��%�����9;(�Y�0�OD����E\��F�	�}\�Q�KA��C{vy(��x�Y���44\j \�$Ɠ dJ��qJ����7�R@���I[����xG�b��V����u�d�����OGN��w�V���F��%��'���2�IZmxB~
�{��1\m?�B�Kj;6���]t�cF8F�'[�O3���S�@m������B��i*�('���\ ������)5��a�,����R����gq��p?Ktoaj��1��w1�k�#ɤ��+��k�w,e-���`��4��y�_z}��m� \�'戓dm��I>�ᤥ4��j舽�+G�d���� �-�=��G�o��U6»@�W�I�A��.K3lJN�#v\��j�<� ��I��0�B��L<�K��|��B����W��dR
6}�Mܓ7Z�_�_����"��Ԫ��\sAxH3�
JC���o���=>���ɠ��v+�:������y������� ���j0�#�juGhQaf��.�?ܵ�v���?�=yd?����Gyٌ�L�
��?�������rd4�f4�5��%�y:���"���,P�T$$xͱ~{�]F���
�,|�=ϗ��^��2�d�8Dӝ�M��Һ��։ɫS�~��,u{����K
�⡨uN�}���(v(U=c;>|�/�a��}��t�/ߜV'�2�b�xEǱ|���f�B�.�!�Z �|�*�q����]�w=w٬_۰��Ԝo��V�9𜣇<J/gy��ɊD��m�Gv�OH$��c���W�2K����AN;GÜBi��O�o ��S�P,Ҵ^;�=yz��ld��%I{&���t��QΏ;�+��[��8�]u�Un7xW��qIwd`Jb��ߔW�|r�Z� p"�GO<�jQ����H\����I�견be��_PDK�[�U���_ڑ���0�K_���{
|J��P��^���Zn�X~M�R7
%؊t�z��*������U5��o���Q�їk�l�I�.ץ5���^��<�*ݥ� wF�+3���K�~hB=+�2���S�LP����2U����)i�@3y�8������EP�t-�zy-6V�>Xz#�:���	��`gD�vBbP��Y��J��*��YN�Ky3���w`��RG�(B�6c4���(��e�
�)�:�cr�D��kWc�C��s����,z_�*-R��L���8��G9�T�"}�dn��劾;��,�����AuGH����i!�+wJM0��(����q4d��� G�/7}���`���u�!���Ll����ˠl��x͠�=���`��&��1)����x?z�Yy�J	����P3@ktrĮ��r���f������|Fp�v��k�ֱ�[D�ƚDyJ_1��r��*�#PD(Ӂ���Z�Z���뉶1+�rR!\�ܠϿǲ)˨��2�� ��f��2� ^��oE�q4$�&8*�I�F�Ko4X����XH�b��PN�;q6m �;���Nڰ��+���V�m�GI�T!Vn3G��%P�`��.���M4{"�߱��|�����L-����)^J�VtB\2ц���4���ã@"�E[����쑱��nN�p��nZ~� p�z�2���*���휃ǹ7ݭ������Y#���'L�Z�A>�2�@XC���� Lo�����B��I����j��zPh+cF'��O�Ka��xl׹ǵ4�E��@�aI�
�E0�FNV#�!�&����P�\���������L��;�! zs�� u�t�!$�G)+�Ua��Hrэ���r���ݼ�}e� �l�9&�D���V��f�6���:����E��@��SEu>�#���>��(/�kaFϲ
�݄#s��fd�-^o<O����J$2�]e$�DP�c��\σ����f���H�G+fUG+�o�O����TIKW4b�w��Hy{r�x�g࿍[��߂�!]�<~��~n�(�	���j�T 9����ߗx��莄�&��)�J� �ru��Zf�v����*p� �{B�������6#�B�9���t���6��hY������~\�C|�n^p�#�Nb�z�&����殒,�wk�'�Ŝ���|(�$�}v��|0�W���[c��V?k���5 �`j�+�f�3���0ޏ����GN�shi&���Z�ĜU�D��a_�f ��=�O~a|5�α'Ui4>�q#�D�����-^����6��Y��[�M�Q�ɳcw���?�*y�c5Emyl��('��}��OnD���_#��)Nu	�Pλ�g�Gu&�v��_S�}^ܕ���Dp,�Ɠ���ҝ�=�2�!��u��NZ(��d��9������4�[vc�w4����`! U��3��R8SG�x�VnR@=��?��Z���n�k������e��E�we��y��I:�Mf�<l�˸��L4��w�̔�u�L��Q�u�q0�$�H�ź�K��.�E����v�ʾ<��D�}�C_�IU�x�p���(�It]�Z��-1��� �̙<1����TH
����hSU��y�{Jw! T���6�0�;�͛��rF��X�*�� :<)��Ǻ�+��k�T�eRS9�N (�:��Ó�Y��(��?6�B�����h�����͵i��[=.��W6�\(��ы,߬�2ãֱ,�������_̓"Dl[�p��S�x���	����u3T�Dv1��*�(ouQ�U)��dX;_ɣ��ᡳ5�ʢ+``8ٶF�,��,vzR�\����c��;��6rب$r&���ٞ�F�]]�=;v��P;�m��ݷI�g�M�<�$�4iP�����3.���u_U�gǎd'wŧ�hz��}��[��wFu�݂W������K�?5��-����b&n4]�˼u��R��!X=eW��T���v6�BF}�F�VF�gq��.M�͛�pJ�"����i�x��%��gTXKt�-�ќ�%��N�����3���X�*�;�o��OK�aa��LA���(��T�5(�<�	�޹l�M�b��NGB}���`��#`�5�ɷ5��t5�Zϋ�ѤD -]�7����	�st��b	Qi�V�������w���]"V�qD�#ڰ�4E���&���m��I;���mm�l)�߰�*�G�A��h'��p"�C���ʚ˶�WD���Zy5ۇ9y��)	� ��%J��.ʹ�j�,	d�ֆ_,1Μ�>�o�w�d�ɀ-e��emڠ'#K��֪:�������_:zz3qL	�ٻ�A?o&1�U�GϜ	��b�ʧ$M�1G���ɱ?���NI�b��Hj�^C��7Q��"��9�5�&N}�l�+z��G�%��ߜ�\;��p�@�#���J��of�oK�J��0:|y����'��o�{�N%:�B�V��c�`=<u��J��̝���Ҩ���*��c} @�h(ąI���U��}6�n�,Fo�����+�ܻ�W�@�����H9�C��/��bwO���g�#m�	�-�<;���O1;���B�ꬆ2�:������s̤ɡ��0W���|H:�0��<�<��?������v�%EX���o��ː=U���M���T�s�]�6��ŔO��#i���@*9�* X�4`�+n^�˕R0F7��VO���!�ɯV����98��IM-�������^E���鱒�x�W2�ށ�/[��>|�B�	�Ȕ�@���+RO�}�������!{%�X�����9�}��������h=��L�6G��͈��J�c���V�w���Cl!
7��k�k4v�h61�>)x~��V&�v�YHx�C�S�<���8>ʖ(&Z�Y��޻��.l�%2Q�����O����:	q�e%����$�����w O��װq���*�AI�l�	f\�s䦄iXG�c�J��w	i��)V#�jQǤ�UC�C������Cг�i���M��J,4�z/��[x���[>�W��Iy	09NC:��l�����]�DŹS�FPГ<��%?�m _���(m��WVhyA@=	R��yN��C�L&�
A8q����)�����}]�Ȧ@�$�l-���B��i7���D\�%����>��g�}n��[r$����-!uk�Q�g�MFCA�����M�1�_�Ū>
�0{`�~���0�l�h�$֐�F8LD�����M������;v�O����@�S��9��-�O:j�%x��R(}��8��bd�؁����f���Q���@d���}�mg�������&�6��`�YEn:�⌸M�4D�K�*�ƭ9�;\�N{�p�o2���j�ϲ�R�;�Q�9'P&uס�P\����]�FND@�v�-/��U�u%mp��5]7���M��g��v���m�vE 1G���1�.�%�ꚠ0��%���;��?��4��۲^�y�z���V�(�w��At�	t���Z�P7�}�J����ev8u�G�%�����s��RW-1Qr�'9��P��i ��dbn��Cw��OZ�̒�;&ukH�Ǚ���=U*���Ft {�o�z���[�6jy5�
ʂqwpM��d͇�����qE�T�3]��hk��di(b�ꇥ�m�����"��7�΁^�Ko��j��P�����z+V�2(����t���^�`TP੎�L*�}%�#!�@DJu�P�7����R�+���I�5�kH��q:�dG<	)�w�Dx\��Fx��X�2����S����X�D��=ݝ�dS��>�&��8��"�Z�j�E_���	� Ju��9`d�Nd��T�Up'�����ʹR�ɧ
��L�ޟ���-W�$%LF����PE��5�I�a��R:�NN/-x�&嘉���ʝ|~{7/�Lʟ�Es�S���ueO��w����Fk�gr��r`>뜢��P�>����ׅ�4��l\^��v����'-v�Sz�l�=�׭1W�&��n�$���7�<V A���E�	�g��z	�d�ΉBe���OT@�����l�?�y|�PK��LlI4R���;'3rC7�Cc	��סt����J"+������w.*c��`�q�"(;�~Yz'�X&Yh���PB?@�h��I��/����]��QZ��թ�o�g��)�l$���ϔ�����w�>̏ .���]N��:�k�:�&B�8'cS����\�o}�ɦ��]M
����^���v��T�2�oFq��oz>I��I*����n�8!�,����u����ѠV�>�W���-aKt���S�AH��̏%@Xg�b���Uʢa0�M�ԞN0�ֵ{~خR��|�2u�����@H�m�(�� Y�"z�T���v��e
Dx /E���V�r��O���@���<�0��U��T���*/&P�)�K���օ`t�or�����e+�J)07�g��l��ԨL�R�1��^ѹ=����I9�U�������)��^g�v&K0�'�a=�]5�>j��
���;�B��!('�b�o�:���˝���FaO6�X�����\
Ή�1�|�ٰY�J�ed��EA����U�6 ]E��HFQ@��B�A���k�#����4z֝��Q��κh������]�;����sUn����*<ְ�8eOh?����J����!x�"�ػ�D���A��F����Na�_[��z
s��k)̺OZ�Z&���(����'��!a��QU���o��)���,��ud��H���z¼���#E`�y���|�j�ֺǕZ�k�Dq�ִ��	ہ���?%��g��Zc٣p}�� ����ώ���EܪA�LԪxK��X�d�����]�X¡���t�Ծo�}H�7AE��\�� ��a`TP�C4��uشK��:��AZ<�]6�+�|��B٘��ϛ� �>��I:��,,l%j����m>��y��S�@Y_���!�qL���Y���n-�Ir+-C���ص��J^��{�K�G%-	��T_,�5!�BsQb`9j?���>���J�W�'���	��`��:$}ߝ+��Lb��(01MS%R�þ�c!���V�8�zB����j�'���� �Z��@�Ԋ�k>P�x�ē�xQ�Y�bT��X��SF�V��14�?�6ˎ"!n��g�u5�Z�w� �!�f"�Mf�l�/"�?�����ʑ{�Ty�"@L���[�rR������9ς�e�̿�%��i1rb�94��z�t˚����I[EHk޿W���S�o�4�B{��MPr�_��G@[�J�*r%=�X8�us�D�Ft�����;�x�9�ȣ����d��uDF���Hc�D��"Ei��"!H���I�ÄN�0�`��X�(�z(�=��Q�RŻ��UVc=�d�=E͗�C�fu}�v{���V�a*���Z6�<�EL��GQɚ���8��:�� =j�ƒ�':gW�wV Є̈ޅ��6�qt�l}�VH*:9��l��f0����s���A�e��|S���ʦX���/�}����Ӳ���{�����e�\��<�;O��8��2z����5���a�<U竔4�|0�/�����'�<�`����'���������l��~��qc��j;�ê��NR��(NA�F.R(V��?�w�V�����P9+�/���Ţ\\0���og��;�z� �?��uE�O$ߊ�q�ZYn���%�Ȟ'L�Ԓˁ<���r��-�'��c��MZ���v[����e�t^�?�0=���f�败k�gR=�g�[���q���個��&g�6L��3A��7X~���n�x[r�/p- ��پ�pE
��P[���S��}<Dz� ���ӆpf�
M��U��/� Ч��ڛ�΀�G�޹�H?�R�:����?t��#?��z��N����)ł�	����]@3��l˶��Ѧ��׆��ڡ�~f��$q�02�QH]��U�g��3Kґ�X���~�TbG�BF R�_��Ҝv�!�Y0,v�����+C��H��<�]t��l�K�@H��q��m�;�h���(a�#�}4�0����R��>�����e�6�Z��l_.�V��� x�BN2Z~B/�b�;������_�}J�Mw��U � �l��ٿ���8��z�������e����&�Tdcg�>�:R��#��Lj8V��)��
e�  W~���A?�Zt�����˹�u/D��,C��=S����ʟ��V�A��a|^0�<J�G�⍳�<���ܕ���\Ee}04�#Y�����*(�}5mk��u���v=(�C����3c5�ت�#蛪�L�?b@�%�e�T���]!���emGm䕧XC�Zݘy��x�EG��]���l���=�K����cE�kgS�-�?5ͦX=��ӎ�`�b٬g�t��dU 4�d,�u���?�N��X2�+jG#�Ln�J��A���H7T�x�/�E�,n��ͮ�z!���)s{�E�jv]�e�:dz#r��� ������?Ϯ|�:�^�Lejǔ�A�B�P�]�j m�e�`���=q�x��7�2:F\ ��C�5�[8 �5UK�}�5#v4l�������=�Lly-he�5%qaY@�h�<��Ѓv[{��+�f���#�0f�D��_�W����SJ�s��i�$�W�	.�ޮ����Χ�G��P#� ��xz���9�`�m�~��/� 2w�*�ۣKi��W�n+�u����1�T�'87x)�S��R�����"y긅�ҥ�#	��r���ʮjcg-á�����	wTjZ(`!��Y�=K�,��!*�Hb�cb$��?D��!L��톛�3c���������`��Z�����+�y�}02�R�н���-�i��=;`�,C0Z�j���`���+L�S��2�=���T�EK�v��AKvS�G���C�̖��z���d}EF�9�uC�Ui�Y�nM2��G��,1�O�:�Q����M���B�z�
)Ż��G��m���B!^������0q���7�M&m�o����
?�p>W�
b�� �#�,�T'־�|}4=�����? �vϣ%�/J� ̉o��w3�ׂ兛}o�K�S֭ė}�v��f�w �LF�	�#ރ���6]n�� ���|��X�i�a�����Р����hn�.&��kZŏw��)�?���8�!"1:��=�}3	-���/�g�v�ݨ��!�x����4����d�F���XQ�0�J��^ܟ%��)����ߒ�̷�m|gYFwV�$���`�)@�D57IH�S����ۂ��V�~�'H�J�Ҽ��@�
����l���Y�c�Fd�{�ke
��&z��,����Ȋ^j
/�xPp���~�� iEù��i%H��OG�\U�
�H:�y��oT[$(b�����������Y�6�f�X�$�t��z #��i�/h٣Y�� ��|��!:s` �/���>`C���S���*��K�}��{��� ��Ѱ�،�iu��۶�33�!q�shrL�F ���D�y�I���G�&���.� a��0YГ9:9�͝k3��I$�3���;�����0I��A=�yVm���	��I��L��~KǏ0۱��5'#�-:�>��C��7J��F$I�,@M���d��l!�@Ѥn�e:�'--��QW�2�	�\+m&�8Q���8��^eJC!����#�L���D���QpYv'���C��B�2�b@Uv��D~/���"WZNC�K�4��h�Y�J����ѽ�`Qf�w�p���XIi3
Է�m�k��$����Pugw%��F�D�/��*��
Q�=I�;�1'm��NJ t�L��!�ӐI�u���sb��܈�-��
�1]���55m�j�5�]�f���r�׃!$�ج@�W�lK!�����YP�����y[Xu���Ƅ\�֠�V��b�c�q� pg�l��%%�"�r����U��tE���h��/��4���P8�4���%?� ,�AGU �"f�$�.�h-U��FߌG�u��5��K�?�C�e!+즇�2ob���A��q	&=��[q�3zѢ����<���y]��J��WMG&(2�S���}h�*L��;��n�bΪ2�`V���c%Ё����o��~�e���٢0J�n����RJ��'%�6PSl�m�RA8n���kM���7�1)�p�^�7�w��yM,o�xm�Ⱥ�яn^&�Q,c�]�'�h�Mp߱� �͉����ҐPǻk^�i^{��j�Mth�K�|��ڿv�H��MI-Y��^ N�z�<�3�)�������b]���Ǻr��tO�D�+NR�hV��k����ӣM���G�;]ΟK�r
:���d����;��`��X>-s�s�k�樝JQ�A:���g�G��d\�9N�S����9W�rFri֛ؖ�]0����I�=`��?Y�7��i���z�CM��f��?݋G�4�.��P	~�KߑNM�`נ�&)}��e��w�*a#�������O�i�%a�Xs��.w}�'r�D(�^$�	�Z ��´Vؘ��[3=���X1ɜS�M�b̢$ᶰk!�7�E�ߔ�L$0�܁��8�c
=�2��&��d<&���ֈ�aVI���oZ]���$/�S���"�� |Dp�  *�a�6@�e
=be�t��W�S�$���P� �hھ�%�h�����y���d_�-љԄ��;���K�>hZ�g3z"wg���7:x04L��3�,`�i /��q��1���a�-vnN�U��7wr�e�}�� h���~�<#A+��R�I��~�Ln�u|�	�a����2չ���hC>�b�!x.��v��9��Y".|O�=��Zk��o�,���D�[�}C�c\��$I�,!���I���D��@>z���c�Dc11O�4�oU`/M�mWÀ��]O�60�#D����B$��J~+[O$�!W�~��kx��tn������.k��&g_��}����}h� �n��.�;>oB�m������N���1���g+��б���r*l�d���RU]�6 2��%���m��	\2+Ԇ�R����m	��Z�1��W�C������O�:5���`7�J��T/ٮ}T�^��i��-��`�{�E��\+��a#�	�$N����B��!�����p���H9q�V;�����b�'U�n��8"z���]B9�*�u��W�?�%sڬ~h3r@W"g�?(� �{��J�|��a�Cf!TcG\p�y�4H��sQհ$�t��, �gvv���xֿ����g��ר�Cip�I	�`����0w,��-�{�g���n�|5%Ց.��_��3�dbT� 
;�,�QE��b�a�ܩ3�T��|{
�h��Թr �܉P�?В2ρD�Ph�F�h<	�}������	~<��k�o�ʇ�[��4��Hf1�N�h=�~]�>h���k%Wd�9)��fb�;�_�Ix:s���9Fէ���-0���/ -����|0�р�P]����	BxO�9�	�$$<k��k;�"jv��YO'>�~g��g�����du���{�P(t��3qǡ����n��!�	[q-������{@�VZG!�8�/��F��D�/
�o�>b���f��w�����Fҿ��,u?�y;�b���3�)F_��w�#�h���7&�=�S����������".��/�>����=?��!����T�!L���?�Go{�	�ε,�j޽w��S���]�4���4'� G߉�!ã��0Ajc�V��a����-��z�؉u��]2t��ƃ���%�U��Z����sJh��3K�s�a� �˱�Il������z�Y��Z%�IW��Si�\�g#�硆:�/^�r�ZsZ&��r�0V���1��G�K?N��ɳ#x�_�Xx*k;!_˖ }����g���z\G��E`q�&cϵٖ��z���X���D7��J�����
|����|w�dJ1�A_�'t[+�`���VE�8r`��Q!��S���)�Ғ;�m����[�d���q2�)t?#b<�&��EgG��_�>�i��d��E&�O,��mA�l�������Wק�"��w�S�����zd�u�Cw1�k]���Fׯ����H�<#|��g�Ǵ8���S����U
(��(� �3��q�T6Rkxh��:R�"��d�g;���i��X�]/��=k�<?�UJ�a����}F�ow i�G����b4��$V�y�-�ƏC����F�h�a/޻�B�V�4L(��V���n 5!����	�8��15+Ҷ�����Á�������qD#*� HeT�<��[�x�sZ�[�V�uM�Q
�����WC|�M���{����ɼ�'��d��rb� �鄴:���`D�U!Q�yA�ݼ����菧�pXְ*�.r<e��cǛ�R��"e��Wu����vW�$�Ӹ��2m������U�T�B�X�3��(<v6h�VG�/̟�����za��O��17t����t*o�Jگ@+'����I���s��q�Gt�^�!il�@J��
>�������U)\N�1.%#E2�)Y��y�}�,�
���t�gH=SwN��wK��t��r'Ώ�G3Ը>�sK^���LIW��n?hW���a�L"���%���/x�hx��y����N��X���p�z��"K�$M���K��ް�^SL�z�֪�Ս����j�*�Q�}��)7��(ō{�p�J\� ��k/�B�/g����})re'���VM�N��:~�F�/=R,9�{�f����q{y= �H��f���L�nm�Cxl�ߘ f�IS���("][3�P���<]58����o��I��U>�9ލl,��:�f�����pt��'�Y�J�C9��c�iΆڄ�כ��*��K�u���w������sn邀����"	.>p�c�.)�:Y$xe�ӷN��@�^g]E��y,r���fy���5��"�8ژ�+�5�}��y*�,@�p�h����G��@�0�.S�,Z�Ƕ�e��N�'�NNl�r2�`I�C�
:�ʆ /��"L�}gi~��gI�>y׌?��YE҉��Mg�ï�J��f9|�*�:���Ζ`�݅\�ݾf�T)����������S���_ ���.��K*ܥ�o�%v���(�skWQ��&�K�?]SZ�ҏ§�GZ�Z�[@+Q u�9�C��zE���2 "���J��֦��8D~{�8M�`Tj����X�]z R��v9~���a�P�`����fUD��� ~��sN�y��IL; �8p�|
J�����WvZ?��n��>?;$��s9�G�壵47�ZB�f;��J����A<�|a|hZ���j:扃*��l�6!m�I8�/K�e���z0H�����@��)	�_��ޠc�5�b�7����I�ɔ
b��q���24�C';+�M��/z�ʑsj6`��f:��C�N��[
�0cmh�w�(�QY1�Z��s��������8	���+(���u++����ҭČTX�D��(?�ߥ�2C�P�� ��v9$}��%W�n��&)��A�R�G�-v���_����1���^�=ʽ�4��hC~���R3�����U,�h��:���`Ӗ
If�L���G^EA�!�q������d5��*��TD��A����}��*]$�t)�ނ���h�bp[��|S��?YmӾ{�#�����[gcO�>�2������lI��xm�q:����򾗥$�����������W�=u�y�jR%ޭ+U�M�g�l�u7�^̜�b5����m.�Զ�4���ɱv�ݖ*N�OD��j�w� �"�'@����-�F�=z�٣��KoK}U�&��|�oY�6q�;�}\P���#�����5�*v����<����\Ot�E'%��w���V��Q�3�rr?[k��a�a^Y��E}<^���4��՘���?8H(vS � �^�]\���<�7���Q��tb���eaz���:��'Ʒy�Q�3/ܭ�L_��'fL֡Ii�vD�G7�)֑*hfCi,b���6�a�j��P��=���|/%��i�5�����k��u���\u�!Y�����͕+��4(�t�_���?΅�� �\]j���.����}J�����$�y�&��9�]�,Č0ӷH��q�ga|��R������.�p$	�I+�IC����%ɩZ�|ֲR��0��=5���#{.�N���T���G.�o���+����.4ϣSՆξr��{z��f{�m�{-���č�Q�o�{ IG&�YZ5�8�;�~ j�&�6��<�	޼c����f��>-C=���ðub�8����%��y�}[�Y���Nj��\��-�ɳ�8��NC�_��/����R^ݖǄ�|D���FO���y#�GHV��Acb���ȶȇ@"3�sN���)1�]�	�P���k�'�ńy�`s3L3�0ԉ�v��UꮺfC!�׆�"���b^_��O43��+�=����&-��%lhف�(`cn'=b*D5;n�ȱ�#`W�aV�݆APDr��C�F����n��lE��ʟ-�.�=�b�����R*�_�rU��4�z�	�GAX
��Cء�K�ܺ�}ܴ{�D{"���р���i�)��
7w����������q��VL�i	gI?����;�N��'�e���T��]WU�c���8����H徼A}5�fH5(U+4��%�����G��M���@�N�N)���!����EU�)A?q.v��qí�g`���W��e�>N~,4����;0�O�#�K�Tg�S�_>D%������eƐ	��`ͱ�E������L������t$(Rߚh�A`�a��Ky�/��\oNb/�4�G'���E1Fc_��m��l�����"M�B�k��Phܴ�8�"�����Z#�����*����ST���gA�uC<1kB�jK�z��`\��Ő���b���ff9��`�ː"����������xnQk������+�M{-!�=�`�^�����U�ߎŨ2(3 @�q��6�%��tX,�	u���݁L+4�o&��˘�6z��6�L��fV>4:�,��?P��H�DO�AjїN$|\���W�����U��i1> W�:��5���&�}6���4{K������4߯йѫ�^���S7�R�*N��i���� �����%�����DA���A�<�!O����Q7��:u���UO$)B�9��B�U���D5PQ�ǾQ�$S��^�����	���ڼ�=2g���b���u9|�Z�+0��0���{ߎ����7u���6���F�� X�];�o&�z�NK��>�k����� �z��r+&��F�}�6�WUa��z�v~�g��r�_��}�\�,�	�<�g�;MJ`��͍��6�i��,�a����b7>��ռ��c�1Z�����j
D�����2_�:K7����y��}�_���]��Z�w���9RNp%)���S~{d>l�+�-���~!UC�n�T=WuKW;7�����&�w����c���� ��/n�E?J�� ��9�����Oh�Զ�5I�Pql�|#�R�k���7x���Ȼ�M�sg[��	:?S��~�f�z��w�˩�S4�K 8g���k�!�;5˘�j��;��d��Ӆ�+q��5̶Q���Y1U�����.�	�YWS���� �֟��H��H{j���T���;q�;̨�<�x_�e�*��c�$`����\ԜE��P~
X�	O\j2z�Q��G�eCsGَ�,j�`Z��`]Y�������IݼH�iD1�{���M���W��&۷�)��ID�ᙹ��m+r�T�iIt��m��~43Y��>�.��:M�S�áL���2�;c�N90�w��R���r�e�ϟpLta�F�isN�7�|tU�{�%�o�%�EOPIt�u������E�*Zd�:\�+R#$�.�k�Q��L�/�����E��V,d,cb��5���K��^���s3����H�=gc�п�n��d�yx�8W�GZ#�(���R2:	aP�"��%�|�9Gd�j��xW������⍄ucKh�I-d|��ި�޹�@BC��u�h���P%�e�x�K���a�ч�!�+&�� ��ޓm��F9Id���#XNR]���Z%�"�8A���CG��e>���l.���֜(Rem�$���
8�>�/rU�u��T�?l�(p�әA�W>���@�
Xϰ��/\�P�;;C0+�m&�����#�d��#��a����K_8K��-���+70�)ƥ]dG�`R7H���!q��I
�)�^f�y
��z3K��M!��5��{z�hu���seer��а+�jѼ���ŕ�i1Z5����[���G�0�������'�g;���6�����2��S��h|>8ɨc*�2a�:%�.ʹIN�&��y}���˷Z� �yf�hj�PZ��>v�kt�x�{nQ�o�Z�X�d�U���p�$8��D����4����V�$Nj2R�ף�5p����4)���x�F�[����L��8��Zܜ�)�IVd�5���̊j��ٿ"�S��w�ӪflY���Z��-sC?\k�k|�\5�W*��"�P�\��
��M��P�4�C��GnRR����A>!D"����K[��SK�^���S����ȭ�/���=� ��k�y}�UXq�s�Nj����$��T�:.£)X��i��E��_y1�ỎtM.	A%u�1V��4	�=`V�I���}é�*��4»;n9�m��������M��}y/Z�X�Xd�L��WZ���� �C8W=?Y6P�a����aU^]N�]#�w���G�Kg;���'�P~l0����I��;!�}�M�ƴ�{�e [�r��c5a��{�᪞K~	:���%6��A�`��P�����DƎڇ��O�n�J��X��ZI��yc$mF|���}y�7�'y�{�1��+|�X�Z
�Q� �,��k��W!�z���%敏������J,�[�7}m���|%���|�G�pq5ס}&'X��u�)�M'/tW���m�|�Oƴid�q��=�Ǥ��X��K��'�O�f�#�`�c�_�����B�,.F28������k�/G��4/���&a���9��~0�����:�1�F>���pA)Ȁ�\j�y d(�5iY���<]�?��Gu�B3�+�X��Ay�gW���qh�x�vQ{����4j߁@�c1�7�
s�����Rj�w�q���S��lr���l��ET�Z3UU�ކ\k�H����)����3K90�av'D+�LS�r��$,�Wq��+�+��L�U\Hj�X"fT�}�G:"�I,5���#3��I��^�
H,N�tf����a�LUD�T�b������z���!#���Ǜ߮�B<� ��j�t�r�Q����g�Vo8������@t�뒶�˩�`�9I�7=�� #e��pɫ�ag��f���M�G78��iK1=��$Hq�\cl$��G6~*�p��k��z��Ei1���+��C�i����7蝧�U�Lqjna��~�⩿+s�^-C�7D�8�����@\~?�Nƃ��\�э�򦕞�\�?�������?�҆�N��(3�=n$Q݁<�O'&Y\�F+�N��)�v���ԜJ����}�7m���KۈN�k�|3~�:�z�2�����hhBfU���j�v�v.>8��K-�b��z'���Y=��W�d���"��0��Oٵ=E�?<��$�1��g�����%/
�k8!�7�(2+���oEH���V$�g��#B�o�E K��++���S���g9z{��}]��G�����氡���%l������s�b��}4�L&y��Uf	S�9�m��x>V�r�u�E5��+7�p�s�<�4�Oc�����"��H�����z}�6;%�G�b�os3Z���[Rvdޓ1�4T0V?J��B2r,�Y�"�@n]�k|��Q�_�up���J�:��6x����8�?�bp\bM��xq(�&)B��a]lee��& ���R�,vo���j�`���z�;I�X�&<A���-��r^t��l؋��˟��ԐUV����$5���� T�h�z@]���Ҥ,�Th�5=�?�j�}����N���Z�����0B$U��Q��8A칏���Ob�&da>돕kC��E���z�J�]�=�fI�m3�Ŕ� �	��&ˣ��a,G������*-��JkyF������ބ�S���s��#&��깾�,�{ѡ�����kQ����&Sn�<{�-h��Ƥ*l/k���+�j����"��㦰*Ʉ��SO�CxJW�κ�됋������~^d�qc��β�oj^���ǀ|`�c��<)f��Q��OK&|7��U�c�tn~�F�wo�hZ��}���	�уA���x#g^���o o���nX(��n������#,{�	h�~;�[�0&CF�F� �*bH�A�&�:�l�=�~�
}��Q2�hK�"�`���u�Aj�LD[�������d�,�CV�[�8��7�o�tfL3���
Ag��Cү��nC�3��[�hE u�I[��J�vK�ޠ�w
�� �7ʧ�5����>6c���R�����`��T0��ۊ��J�`%~;�u�����?�+>����rf�h�W��,R��{dv���S{�f{�r'���kNs��dn��v̞��(�|F;K�q��Ҹ\E"
Qq��cV�Ţҷn�rOk���G�o�B���z!r�Z�
l�������������|� ���r�LxT$�O S;�$�Q�$m{Zѐ#���D�g���
��$T�7���hu����Cce��e��`�ٖ���bC����D�<u�Ё�C>w�mg�G�8�F�)�z������n��9s 8�۸�bCA�l��ٝ�P|42^�7�O;5QB5¨7�=ʒKjכ�}r�c��8I�e��CC�$Me	��C��z_���[ ?1���1�.:�-F+�u�Q��le��DΕr6�f���?T"�q-�M����||>EO?|ߔ��G65�؄��O�h���}TܑnH���>��)z[)9�g�F�ִZJ�a1�]��>�ڞۚy��>,O7,?ŀ�=�0���}Ճ���4@�	�
m�~\_��`~�L]�t�/�wv����~h[Q�o�}rP��f%�Um���5���c�TC�2����VN��� ;r4����/ٙ.=�#}$�*	-�3���y��C���S��^����l�`4�X0ZK���A�_
���z�qL?M#U���
��G
8�M�V#Z�֮� l�}�k\1n��び�0.B���J3��I�_(<��&��a����­f�:4Gh�������!
��tت��9�\��\Bj|u�� �m��\��Tu���yR�������[A	r����1��fI�|JH�f¼u��M��0m2����rzڜ�Ah��`].�� ���[3�@�m��	�޹�U�|ŝ��U-�r���j��}v1�(o��zC�8�22�O�Zo�����BY�Z}щ�~D���`C��?q���ۼ=扭�0�Hk��>¥0��;_̘�!u}��Z33��#�����R�|��Ŋ�`ڨԤ*/^�d��:���&+P���Ƞ8�Ҏ}��`x��������ג�Y���d���/�D�m�J9B/��h�AEʎ`���`$/J�Ȱ��h�j��A>��@��Ϡ���s��r�L�j�_<1~9t"�,�#�4��'K����tS=4K�Cʹm��U��kC���ж�55�Aq=���_�s
���I��Sb]6ʼ�6g+��65H�ȅ��E�ڙ�̳�Nʇ̳��&Ǌ7�y;�&IeQT��a��|���(���
"�� -���;a����zXZ2Pc��S�+RvN��MC���͎���zʟ�uv��k����D\���m�(#'�_w����L�B@���3�6�N�͸��aA�	�O/�?_������Z�?��ul%wػ�Z�'�2n*O�k�����Y�*��G�g��Yd�|Vu6�G�6��a��4�/t�֜���_���$fvp\���z�����/���q�=X�������}C#���s���OUVˢ�t(Btʆ�V8��+I�� ��r���_�*�l<�>�?15X��h_%��8K���e���2��	�؈oD^3������ʟ%�
�YN�9�lo�hŗ����D
��J1�Nb�$�*�X��9�?:�7&)�E�GL��J�X�fٍDy[� �w@�`��Db�Y��`z�`ʿ�E(:%�����]��mB��		���,t'V��Y�s/��?I�nL�Uv/�?փ5b�?n�g�����^I�5�?�6�$�G/�Y �}�_J���\j^��)��������ባq��Ύz9���(�*��Y�"�B
�����GnEJ�/x�J3t__y�|���&BP��d��Z#OV����ڦ�/\s��`��$E=)rٿ��r:�7 .�i3Ĝ+�>Z\\��3Xsw�O�a%����<��}��N�)��з�����qx��a�[�Y��i���6�IigxiMZV��Cе_Ye�9�ָ���1�}���~Ǜ��ר�c����տ����a��5���Mw�;��tŬ���Eڵ	7�[M�t�z�Y����"�4���	��u������no����٣���P9F�[U�'�si�]n���C��=��C�Q�j�����nc��E9�C�bk]VX�s��&�*7:y��ϐ���Σ�q}��eI��験�*x�H��B%�x�L!��Vl̐Q��g7'��\څ�B�ᬥp6x�C&���Qv ]ph�O>�[�FΙ���R?:�uL�r)���?����CN��+F�:#ۋ�I�d�?؊���R��7!z.���=w�hj�1Z&����"hͦ�j��+'��K�
�q�R���h�r;�J���;v�znQ���T��˨�I��?َȺ����L�`8������|��'�I����{L�%�^�^7?M�/�rl&*%i�/�} �? Z6y#?�Z��c�1�$��xao��f���p��#%����2�gK���b3���&�,�>h���v	���a��g
G��ܸ0!��2�m���� �Ƨ�C�{��Y;�0��&�^`�����_�ze����`j��K;��j�����@�ݫl�����F&����>[�����FN�9͌S�G��Mz\�C$^�R�SJ�բ(��Y;έ�B3����t�P�A���] �!�.�3m�Wfh:lR����1$��$Mm�z��C"�TQ(�FU��m��prR�ȳ����'S�y��&o�>
���$F{�nt���_�:fAW	��~sl��=IQ�<�s�{&,ܖ�D�.u%1�.�	*#��vF��ƴ��/�,���9�b��rf�%�I��,*+�0V^%��NI��e�w��(g3J�}1��A'JT��:��:�3]��O��~��Ĭ��L$�Dl�)�� �	�ɤ,O���_P��DJ$�N2�>VRFc��B������7�!t!H)Y(|T�� �p,ixߪ�am �4�l�4Ғ	�'TQ�f:K$D����<�	aK�1�ExxJW)�a��5c|�E(�]���;{���${ܞ� XX)Z0�M��>��C�����Î��� ީ2�!cm�xCtu�	 <5��F'�����C�AZ܂[�#}I��C1��$ܶ�0j�!ӭ��d�:!ew�r�5��
��UT.�����K������'ע�� �I�LLn�V�*-�D�!d=�����u,A+Yfv#/C�rI�t�ٳ�S�-�
���'�aخa�WH��NE���H^M�u����>3|P;�34A}[%Ar[)b��\k`���{�Đ��
|i�u6\N)�P)����F�'�<�d;����� &�V˶�r	�*���fu�8����M@������S2��:��#X����3˼���t?EAG��a��tG#�B&���H��U\��G/
��;�(�V��y@'�Tb�K
�)�����<}��1�%�.<-�����}�V\S��۱���u���rݔ��j1�`�ط�(y��ҩ�
R�`���ĒD��D1}��虒ĺS�p��y^PI��J���_�D�ƙ�h!Qz�L�,?iKsK6�{�&;�g��q�WG�����G��m�}l����6�FZͿA��rR.��=�nr�m���U!�Pۏk���ye���G�"��WB��Q �Ϡ}v�����K����=0I߹$�����1��XwL3t�r��J�w����ؤ��I/j�����\Gt(�-����_�:n��Z���Vpy�F�f�ZI�:l��6�viC�G{�{92놁q�h�� ���e���C�kq���kN�����
͏M���Ͻϸ=��I/�x��эe�+7�g��^:�;�+U�^$òj�,u�������~�;r��=�*8p-B��Ro�g�b�R�3y�N�=x�k'
�7i�q_�IZV��V���?�w��l%�/��\P��"˰���gjJ��ۭ����x[yj����=骜�$�A)���[�v�`�"����>�r���9���nx�I��乔?W+�	�#<�K���E�)�:����k+eD�N`k?��mDd�X��/���o:�V3����]��V+�2������`�GH���R�$rG�v�O���b?g�ˇ����+������An�|�>��T�Ab>���N*Ͻn$�_�RT&T�������.I�^�"J��Z\Y�F�1}�����_���p	O�����^	�|;N_�Q��գ����'���BrⳜh��D������)j�ޝCg��\2���.��	99�S�>�vӦ�l̻|&��W����z�k`5]k�e�^�,0!sPc���e5:L+�O���'\�]���Y�/(�@�( �;��I([�,�uҤ��{}�!g��>e�����ɋ{M �as��H����QDGkmUH��}f��ŦZju�b|��[�2�GC��}���jx53UL�b���z��2T��'~�X�=y�"q?Yq"��a�R�$�)�9�r�s��e@�|.���{����G��������f��`D`"��m���6L�?³B�N���m����qw��q7�^�-�8B������)n��H;�Qa����n�4<1��y�=.@۬�΍L�8c�B�jM3�:��p�E�ðbD�&,������ ڣk��̙�����GS�t���Iտ+��.n4<��;��eLq��_\6��_�O���e���,TS�]m�[[!Y��D~"%�zʹSȫ��jE������H	J��������QP>��&�ڤ��w�aȤ�L'eȩ�k&F��Q^��l�����)�eC�)d)c��n�K�s�D���QM^�F��8l=��G�����7�c��/k#ba�k=�C2�a@2�\W$f��]C�f
n�m `A��m�)҆�ND6�ld�+��B�n��O�MQ&jʠ2B�*�����Ơ�<(�2�p��2��E�?I�IxS��PHܸ�S~��������z�z;+U�![�n,M���g�i5�곭�j��g�Q�Ns�����0�G����~�z-3�Gnі�� 2rAg�`��!ά��weM�������<��#e�UP��z͟�6����mt��<I*<�'z���J��������*�?���~�L*%��	�0�є�͡r7{��Axڄ/l]n�\�V��\��;C}x��.U���\=�m����n���e�N� ��>ɓ<��}h����*�SRۜ���P'�u|��۪'�i�s��v[LA�M�Y���D��fƔJ[ ��t�]f�=��K|�ZM���!��]�J�g"F�Ud}�I������*�1f��?�AnG>�m��1=<��A<�WBf���m�6�΢�?is�������~�G$!�"R�ۚ��C���炫��%9�<l�y��qmv�~^%We���F��V��Am�3+�4�6���u�1�X !�pv>!��WU�ycw����Z�놶�bY��(��T����Y�����D}���kW�?5�a���r��mBfs7�e����?�-ѽ���01�Y􉀦�*�H^^��ڳ����q�4o�*<2sꗙ"�%~�!<�&��E�\\�R��[�RRu�H��6Y�N�s��D$ݕ��S'�!#i鋫�e65�-���%E#��W�39f���+�y��*J��=i&��P@,�EC�	pA�
y˯�0Y��]=������!~:�"�!*��$���i��=-�o�P@�k+'�\���Ѷ�_���u�E���.x��`��V��U=��/'3w�`��,��	P��� ���]	�H���(�4�h&x:�rn o���W vY�s��%a���R-���;�k�LS�h�O7�t>':�i��>�y�s�N���q1I4Gp׫Fi�$@Qް6ڣ�W���
w16Y5���2��x�eF,���l�&e^~׀�	(mDqd�%8 ;Ge���.'�P��Ԇ�q]�B�i�T�R�{����\���Q�s���ɁNL�)�F��Y
K%��*ܽ �Ho=���/	c#0`���ZʎG-*=�>XpK"bA�IB��ae����F���a����ҧ�=�%���|��j�����	��_�¿�G�_���%h�@S09�\��\5��|a��l����D��׊�=�ϩ�g�2��Z�+l�o@�jk�*��'��i[����^{��̀e%čDز�ڭ������ ���_���=���4 J�{%��6�����m���z0bh/�
��p��?q���u��9��Ƨ���P7M�q�[����y���6Xm������&J�bH�����o�|���՝R���\q$��t-�ߔ��=.v�!^�F�\��	!t�۸\�y�%ݳ����c��W�OG1䒻��pC��t�PWn%�?��G=k=�����m���R��v�����`J(��,���0��dwK�*S\�4�j���Α����|>E�t-��N���2X�o�g6���n�=LB��:�	G�ԎcɁ,�>�D���I��y������<S/��4��kZ�5(���#>�E�9�SDM���d�,���.�SI��߈	�W�5��{�lˍ��������AN�.�|�	jzce���d����gb_�\���9���'n���-kמ�T���w}j�+?u9��	i����#@+S
oo8���c�!ۥ��19r�3{N�>�k�Ih|����˾��(�Y�D���W�����H!��5������ڬ�n��.�9��ˊ�A#ׄ�
�uB��pa�'֔K���@f=��GeO��ω�-�TT5`>S�'��c�g���A<*9�ذ�������
��S���ƻQs}��_���ޡH�{?��*�n��R��>��D�����d��#���}R��h�@�%�Eo�XE|�kޭ)Y*���8!��܀`�����[b���q���^V� ��U�Kg�^�U=Q@�ȞH�� F�s����w<��ԫ��o�4��GHX�5��A6��u���p���n�W��o ݆yKLW����=��ѵ
)���@�/�qg����8� �b�t{�"�}BJm.S����o�A{s4d�5�[�G%[�_S�ޛ��E=\ׄ���Xn���X���������@$�ӯ���O��w!iy2
��M��g%��_C0�G��Ա.,����d�"��B���0����%�u��^�����jԖ뜺(�*�6����)}K��lz`�z�"�z�eᫌ���	ķ���L��_ݽra[�r�Z[�{�f#Ɛ؊��Nzk&:ü˓���)�K��&P�`# ��N�מ�(�֙AJ\�<4ﴢ����0?|,z��H�.�`&>�~D��Cj�e�"�o�B����
�3#� ��G�9�8��^1횠���K�V����9uvMD(\��P��B31�3.p �11���:��_d�`�C��X4!�r�_�x�5�T���jQ�Fr�����.'%ʜHw����J ��~�Pv`�peh��(�@�v��,i���L)���j"�LRX^���a���B#���z��^�^>W	��"E^��z��]#�J��G�7�#y.�E���Jr��n��"�<R)���k)��	Q紎lP�.H���5�5O��+���^�(��N��!����C�P�ժ�˥�d�ХW.������Hɾ9Yg�[�s������T�椄�9�`��m߭~�_(P<������Ո�$�
z�k����� ��.�z��}�y�r^q��mD�OH4c8������d�N2}�egY��c���(-�$(e�qL��`0��KФ���I�<!H�J�k���G3*��}_�;\��;Ƽ~u�Jv�	N����o�����FW@ߞ�\��Ry�������pت����.21�	w�3� 'l���&̷���4�}���������k|=5X�FFu!�3Rr_�%-�"O�S�k�P���/�ֳ�^�,�"���'�uj�GsV��@��@:t$b&�Ǳ{ٟ�
�\����e�-27CkM�F+�M�H�ŀ9u�H� �Û�S�{|^a]L�(ËK�]���E$34�[�p�QH�[(;�z����ۛ��羸�ږ�9tAGօS}���\�U�37���ek���C�[�@y 傦'M�B�К�o���i3f�LL<?�۪����Tu�d4����?�wI����V�gh����1I���S�|�K~�J��Ԩ���9!�v2��'��/l�ӳ�|�ڕ��?�]�Zs@��\Q� �����a�B�p�rZ��WcNX�c}���H�ta�sD����9���z��T�,�?�>���|GP���<W�������(�=��	oZv����hX��{}"�轿�d6�b����>P��O��K���X2Þc^����+�)b'����'�m�-��pϩX��&d�fU�7�Q&H�g���n�VHф�K�i�e=���ߏ�;����/���]eU���Y�ԎJ{���@�����F��	я�T��x(���x�}��xC��Xǃ%9j�͕Q��q%�}^F7X)�q�@�,��O�4X#��S�o����va�l��H�6=�� X����C�[ 1/I����g��s��T�n�����p����:U�1?���H�Z�0�V��m��b�<)~���ظ���U?%ZS	@x�����[��!Wr�@�=x|��s�1�>ާ��+�.s�8@DF�Ş���Z/Rv��5���N��I��F�u����k:sȂ��xCr��ð�����ҊCj\{X{q�����9�`����e��kn�90+~J#��ÿD�/������+�V��cu3��H���D3U|+��r�����.+�	�x����c��b""<���u,��Q*-��e��o��I�Z�@�i��e�2�T���nՑy����T���o�w���1+v���Hk8�Oy|y��v|����Fm���(�w��.������0�J�l�U���2���Z�֘t@!��S�s�T"-��N�t��`I�B]D��v��ցob����[�O]�U>����7��H+�s�I��7�*���|�&E�Hz�\bODw�'���C��P7[	��`�R��ZK�z+SG����ѣ���6>V�;�V�|�zC�"��l.�Vt0�^�Hj`��@�cr@Yg��aB�H/l޼h�&(���S��nyLC����)v�Y5Z�U4�	B�t�#�O�Y
�'y0���i}.���yud;k$7��Y1�X��U-�zc%��/D9�$�dl���":I��W���������b��2-b�`�b�/�X�k�+Z!�J���W�+df����uU�j���RϾ��
<���IC���B댽X5 ��?\�l�^�j�N0��Kc��Q�*��0��+f�<��.��2�挛D��u�y���`sO�)�I�����5~an���5s�]4>Eut�e'wļW�_��PO��=��4�5商x�>U�7{���Tں��V��O�yd�_g���@$�6H>uN+,RP��l��v��lR���?��b�����\d�C+w�Y�>G���Z�%ѓ�Ϗ��A+�AӀ�Qe�+m��Xt�/A'��P��|��"s�&�)��HG��$��`B�3���"��֤��'"X�/��v�@V�A�����]9E�U�њ����6:n>�c��R�*��?M�ߖ�m|��8,53��v�B_�8�eY���E�d��]:B
�`�r�v��ۑ隸�9��èa����t��N����WZ��'��B�u_�Vu����Q�56MD�v1A�u#Us�T����қ�sx0<�j}�8oܗ1��!� ��M��,e����8 �<
	�g�w�P�Ko"�6@�Ig���^!�`��E���t:(L5����(����)��ޓpH�;w�w��a#� }6��l8+CJ�n]0l��b��R�q?�G�c�2��̒�]�P�f]�HJ!N�2���6N$��n�y���[�yS��t`�t��,d�#Aoيg�������ԽL� T�p��(�$��w�����N�X`U�7� �S5K��o/e�H�G���0��%��.qד������.II�i�<i(YZ���8��B!6å�E�>NI��(�Uf�d;:�����f�d�<��gX�� ����~�Ǯ�����@+MJ&���>�;�t�mo�C~~Zf�Zsl�}�r��y!���� 9:A?h����0����� �t� Ԋ¿��u�T�q�8qn�L/`L��e��'7Z�h2���Qd��ԣ}I���Y:�<��_�:C�V�:`�8Q0����E�pz]���!�&�b=S�I���I��^�k|?��Usc
��$��,���M'��l	H4`y�+�z���k[S���Z/���ג �;��T:�?�]��}
�
��7Cׇ�K8��&���guec�x��֖�:���
̧��Vlw4G:+�,m������[��o0nw�zزU�^,P���J8J*mxd��5����,��#)8��+�
Ԕ��Y��EY��H+�N_|�l�$���N�~����,'���c��X�Ԡ57F�wt�"3��Y�J�\Q)O#���qc���"���/[�Q���bS�y$uC�V�_�KהY��K2>�{]5c!7!��,����}��*�b�׼8/IM�����ȶyn=�N�_�گK�Q�\�C�F�@ 9�����/�!g9�V�s~�a՘y�@�+���mxt�%��~��*���'n�Y�C�&�7��M�<�<�O����Ǣ�H��o{�/M��d)��2� 4C�S�=X�����~�e�R�w훯EϗP����j�^�b1<�ba�'R�c��ޕҰ�Us��]3*z�\�sgTؔ���u���2_���_��"�n<`T$�K�D���{���^a�
p
��)�OqM�V�c�$�9���&�bL�ǻ����~��w����O���.�̜�׃g����K��jKe���S�q�y�a���I������s�����2@"mRi�{h�4V��M�����������(a}Ú��,��"$>T,�-7Bd�D�I�#��vS�=�Tt��x��_j�-��K��
�:��TBe�����>��T�ܙ�-�MU��苴��O������H���Jf�A[Ae��\�oQ��sL���.Cؘ�'/#�.C��]�h/�>�n����.@��e;LqZ�;P��AE}^�r_���S��db�V�Qs;�h���JC��ɡ)��P�m�$u*��	�S���޲�K�8�(�S��
�0'"`!�Z�(��GaL�^�XN������!������۾�R��~�����c�l����,a���&�����J�b\E"����,Uh�y0 ����0+_�5qF���{UjCQ�%��i��;¿�AF3��y�_�y#1A�3�]Z�3�Ù�ɦ����|��c����)#ڝJǤ�O���l�^��<�6�Fc�Q��**��|�~gx`׻�RH�Tֆ1A�*,�z��]�<�� �	ߥ&��Ki��Q;,�m���]{�^�N�<�
��I�[���Zz@9��m=G��O�)"��v����ALÞ���]��_�x����д��"8GG�4��V��Đ��t>G+)�@�8�I4��KU�̦tX��"�C�y����ᘌAch� <�ҹ«�������m�2b�$���9-k
��&Ў+O�ʡ+۞g`�eI�[�������MB��nE(�'��$\`���o�=����{�t��8z!�����mj���b�BZ����t����)̘��Hyrk/eO�}��$y�fV��5c���j�`6l�w��������F���J������ZaG��ޙ�F��
:��~b~��}<�%�>1��z;O|3����ޙN@�U9%�#�'��3%���/��T���=P�K��zi�%�.%��?)0�l��swASh�W�(�K\�|�g��:��|�#B*v8B�:��k�ђ������<�Z�6cXe �ԏh�c��s;.3tT����?@�
Ϩh��:L<��Dn���zU����f8�Y��{eRHo��Y|L�<E��jz��o���^�t�ŵE���;TO���Z��[�`�?K�B�dý+����\�V�J�j.�A�f-����{ޥ,���`v
���=�ry�v^w��5�"��&��㑇�$�&��״��I�Є��N��k����GW��8�f)���!T��ͻ�Y!��s|��*?}�[�ܔ$Ih2�ӹ��C��X[��{AB�&��/��s>x����Y�w����	�W����E[@4�o�nP�u�w�5z�[��6-bN��m�(��<�n����w���#z,8���������1�G�P��;H�w��^���z��=��;�yz�מ��5�tF�L���3���Me$ ҩ�*��?�}��;	���ѧ�ǋHC]�v)d�*��vZ�4�j�o����	�˻w �׊`
ϴ1F���>����$^P5'�+�p��Ժ��f�C��&��,��rZw-J�/�/vPxǬ���T�=>�E���g:Ƨ&b�����?� %,2a=�F"�p{@�]&f������N2�I�َ��L�\�2�]��?[K�q��1IT<�TE�ڶ|�lx�NO�^����H��om·|�iي��>q�v���;c_鼯�"��ܹ'��L|u��!��*��-Hl[�ܩ|u�j���9�Q���{܉*{�i�>������ގ��H��Р���],���-��Z�c`Fƙ�뾱qDW�+�����1��F�&9������X_/I�������I<�]��7��!f�����r�W�����q��|y�.cb�[Q�t� �zu�2�&��C�3�UW�����\r�y�Jl�9�3f�2��o�`ZFP�;����]ps��x <��6cWh����t@��/m��5r�~~n�rIGZm�8�d������W�}��n��~a���rk�n��n�7w̓�S��S�w��RA����G2,�>�b@�u�܇��!��Ϻ4d�Γ�B�U�`�8$"9�����l}� �t��\X �� 
��0�N���e?u�&ƶ�\	��f�h��y�:��xh���.ˏ�x�(��9����v��o�d�:|'Ft� ;�?��t齲��iyE�q!�Se�x��� �\%�Y=���.	�P�F>?,J�ب��>�=z�^�>�Q�$�AJ���s^�i���AǳL��r:�H�������sE?%qI�-%0�(Z:f��W�"�03�串��D��<�K���~hQ*�G�Τ,�̲�3�l���¦}Yx(��nS�

کF���Q��s��e�)C��ЮB(7��u�"�P��2��mYקn�s~]�J�uX��dx���dcslʇ�E7�8�� 1����8cH��^��������V(��|6���l��E�[�D��m�1��,Q\d>�|'�q��y���-[��6���T�C"��)�2��t鷮�B-L(�����9�-�B�r��`Lb��L؀�7N����7J�n.G�����M+ԥ�`���%x��WQ��S>j&<C]��Fz ���悻��������Iv�v�?�z���kۏ��J�C���Ӊ�����jmL��(���V3���+Fԯ�����ʹȵ�L�K�O��-��ՆH�D��-ͷ������a^X�*s�@)4��bEr�S�w�����s��s��)��/���y�\���	����@X���Ƞ��#���
�=����e�h ֗[5������y�V-�0ɣ��� ���SF�}`����'s���#����7����9�_oX8`���7	��mC3��8���ʫ9��Q����F���A�o. G�;.��:	���e�w����rH������Cf˔u��UgM$����Y�&M�مl}���ۦ��|���Q&����f|�()E����m+,��>��$����~LG<���|�G���D��W]P��޻D��W��uW�1���;X݂�2�͗=S��j�&!�w.��o-w�M��
D�p�&�����J�PLu�=$DT������FpCr�m���|a���p�uțO|O��,	��J#��u���^�<S��)z�k5$��D��މϼ�Eyo�u�QV�%�lc�kH�,J3iB0���9�5�c23�ٿlD3#��K�Sz�=�&�@r���y���vhr�E�^i?��}���?2��!C�C_�3h��b���N��B@j�=u��(��P���P���"�D^]s7�Gu�+�x�#2�M��s��憿X���(X��=c\`ߊg�Ng�s��<�`����H���RQ q�W����m2��!�v�s�zۢ �]h�K��[`����4���wV�n�f f<�U���}[bx�y�}ZE���]��Z�q��@��+����a�vm����������@�8P���	���֮S�x!����l��=��U.�edބ5n?�e'�X~�~�պ�P���|�&f�{����p����bz_��@|7"/W��j���at�, �+h�L_-�9�O��hL}�\ݘk���/XlO}�ӯ��1j��\%6��qM�m������oa��Tp9�&4Bձ��iP���M8��L�i��g�l@�P55m�i��rJ�^̴ �ǣw�e�!G��0��h;���t'X ��n��%����BG&-�,�Z�K�YT/(�5lR�BJqQG3BMSǬ�M�K�]h�����+wr�Er�sȃ�aT���W��Il������S?�D�]�-�E!��x��Ј��j^xW_���k҃<A)q����;H�{	�/ZdA���[~)U��(�\��QlN"��k�<�Rj�r�[��=Ϝ�@�i�}ƄQ��G�)�Gvg7�f�۹AR�;�W���Ԓ�>�n$�Z���U���pv~�\U&$7=)��ϻ������\b�K+�'Aw����bp�}�x8�cbC�-I��C����}j�6_�/DFG;�g��櫘�� ��j!NR�X��"'�Q�!��������qP�o$2-�O���j���Z�;�i������:���a`�<����¦5���y�s�X�j�9�+�؃܅I�m��RO�g���}��0�������d�֔��G#��%94N��vG�1�H��Jhy@�����S�*Ȑ����$yF ��$L�%�5<τ���H�{5q*8� Ia)����B��4��MJ�V�����UC�]����uu��/�#65�9ֆ�\0u+>���׉�q�wV�z�[����Q�o��I�"��IR�ʦ�oC����!m�J�0 Weo�$���K� I ��a�}�dw��x�ngm)�G�'���ȦG}��[�L�Y$�1`j�Po�x)�K�6��m`ω<��>l�_Zz��˜��;Q��v!ٵxͬ�>�3���d|詊+Hn���Xn3��0��X�^�.�P����������a�0'K���'?��H�$�^�����pqN,)�NXs���+�����ۛ��B��)�`'�A+|�����*ByUK�ܑ[�w�(��<�P5SS���2��5�ev:RXZJ�g���}'��r��_O����=IA�z�(h���N��s�׌�h�D7��D?���,< $�/�4oT����<n�����B.+���+��T<P�v���*��=�aY'�#���>�MHK�ЗiA�O�4�Y�&��^��ٲ��tҕ=��?篎�ݛ%ˎ8m�@w���{q�5>%�oԌ�.���G?�ʹJ'�^n����8����j>d�@��%4&���֡�y8�([�Tg\U��rZ�"��^�"?���2�z+�Ɂ�.��~~7��z|�;�N�A�_��K[�J;Í�ŔOt>���L�؍�����"�c`����g,��}C)J���P�NK�x�?I�g����"<T�]3�
D���B6��A��!�L�᠔����<�[)GصN�dHp'�x��^�<,H_s���"�g��~@5vm����F?�s����Pㅬz?�ֹ��2`�<n+.�K����'['`"�)��(4{M`v�W�B\�:6�%�t��-�RY�^c��rM�m�����0�z��s��l�#����k@N�j�\4�LU	e�ґ���o(����X#��|���Y����T���9x��r�֦�E|��MQ?��>h�Ot�1J˙:���K��~p��%��
-Xl��R� o��b55�v1A��٩j��>����xmya���pT2a�*�;���-�;9>ho[͸�_�׸"�s��˺􇍽㦰�^�4�������)?����9��y���E=�I��8�mQ��J��f���Xx�o]Z0�zH�c�-��u�� �9��[��wU�V��c�}S������o"ʓ�%�@3��H�=������c��Y����J�����)����Pδ~
��V�,��̈�p�^g1�A��cٝ=팘���+��P��C�J���} ��Ff9
��
ob��o��5���z��Q�<������~�@�<.��$A�<��|�&�D]�t ^�5>�5bG�����l��G���J�og��Qe�%���|ɤ"�����\�Jı	�G�wd鵥�-�E@�-RX0����w�s��\���|�Ŗ��_*��Ka��]���K�"�����h��kۊ�����ڟ;��+�6�ם^a��A�~�9�-{�j�y�c�dcVÁ,2�cd���C�{�5eb���+9�)���������B��0w�i�>h�\�w�7���-�Ə��$m�D"~�e�B����pY"�v~����+�*��+��A@Rm�R�	OǼ�~;RJd
a���G#�'V�N��
@�A��b�,������rYt��5)��}�'9��/R���.����~��U��H	�X���#<ڼ��Y@���3����|�:*�7pK)'��,@k�{�ԁyM�W��݈�?ɓ���@�9\F�	+�,ֽ�(��;ٓ��N�/T)h$�ɒd��m�ݧۅFlQ���~����%e���F���[v�PJ7��{�yyr������o�ѳ&bƬvSKR�|���#k�*����-�hh.��}�����w��j�W��'�,�Nт�
'vTg
͚���f,l����8�%1ϹB�uG�C��`޳9h��D��D��4�<�!/SK�}Ҩq�qJ>z��8b5�����.�O���ku`���ġ�L��PEø) ƚ���e_B/���>D۵���q���o*����]�A�s�n�Mj�S���g�g�xϭa�9jD>� *��/SI:�}%�珩�')��[A*%�m`,;6�"�d�DE��2"_ZO�Xx�!G/|f����x^������P�&Bc'bE�W��F���8�In-A:ӹ��������%O��*��� �BL��d����#]Bbᨑ�4 �8Kη�Ԡg���;R���6�/�Loش�|���fP�U��;EArvf��� &Ҵ�K[d�Y`9�F�	u�M�X(	���Z��AH0�^:^�fd�����Z�ӯl�ks�yiY7]	4���L�J�vfjǮ+�2�n�t�hC����)�o3, ��\��B1u6Y���57*L����Q!M�h��B�X��NG��y�g_m�Ǭ��SY�f�������KX�f@�V�ݹ���oܗ�jQ%���/�����Q�����g��`x�|l�e%jm��O,|���� 9�F�n�pD�fO��'�)d�s=E�'ۚ	mBI�t0:�1��Wp�&s���7H�`1�O�J��9u�;2��n�I\�gֱ�#����me���u˓����A��=���>���ó�0�ѽ�ŉ�qW�5��ti�ojЋU���Zݳ�(Z���4����Y����wܟ�Agb�dB���̉&�5��z}K�I!�y�<Q#� �/ ��F8`G9���Gqzެ��pE��wbQ;ȤR�_%�C�*�C��!e��N�ԇ3~\�\L�W������>�ut��5Hך���0<��E3��i�����0/Y����Ĭa�wa�~h-Ҩ�\R��1���g�p��R����;�_�G-���uK�e8��pY�G]�g��-��H��ח�/H��q��>v>�u��q�=�@��T(�h�Q�Hi.�줛Y�5�'yO���<� ������S�H�Y^��g��X4~'� �y�E�תK��ڣ���讹�ηZy?�Psc�d�㲐��F�����:>���2��2:.�*5MX~����[�r��_z�����a�K/��e���&,�J������+��p �#+�^���_g]�̞��/isj�_�]a�Y�D��ns�>l����3	�l6�k����
p���0��q�Z����d)t)��w�]}=ĔSRЭd[�@�AY��K��A��
�2J%aبk����ύidL��.KОb����t�9-�#�].�*�D�Q�MM��g�w�gq�w��c�uE���8���Ѩ��g�noO�`��iӌ)ܧ `vm�53�09V�>f�7�Z�&q����|�8��'�?���U@H�V^>�=��mR4Ȳb���4�1v�%*�ʑF�C]��"�F����O&b���`AT��g�,�L����2�"p��ŗ8��S�w���_?D���-dо݆�W�#�o(�����ބ)��.��L���V[l���l�Wl��<���`gw��¶��D����.툏�u������Ei�!�p]o��#�t�ͨ�ߚwEr�����Y9�ޱ�F�-E��#�!�ǕN�F
g�Bv��4�yQ��i��:��&a�-Mw�o�Q�G���}��<m~�M�"���WYԼ�uŅ�hn�o�#�(l�!F�{hZ�}�1^6!�-;��Id������a-�8��d�n6���ɪ�y���������x�p���"���g&D�?���0�i��&6�M�v�g�r�5mm�#��3���qDo���}ZJ1�
?	��K��zQK*4�p,M���& �a��v�|����_f
׺�P&c��`j�KK��@;�'�L�E�tG�ظ�)n�|Dn�UʡE�^�K��_�}�����I���4hC��p}���q�:ώ�����g�c%�,����V��U:ɸ�Y�6�Jƿ�|��]
@��4��X�_�-G�8ݝ?�G�%y�g�����@���D��,���}��� /�M����6S��&�GŽH*hB�u�R�RS��:��L66��I�'Wx��^+g_�X�U.�+�,ml���ߚy�c�#�W��x�X`s�c��~��(���ʻh��D��/?�*'�%��l�հ��N���H�������*X�b�R�, �'\�I`�ū�[�+�D���'y ޿�ُ,F����1�F���.M���t��Ч����rI�soڊ�P�<&�~��OY���[��]"p�x3#'u�.%8	;檃��2�� �EJ��Q�!�{����FD�R�߻PFĒ,�*JJ�b��Z�e�6�7"����_c/a!t��sR(����p�'��o!����r8Ö(�ˮNC���Z��`�����κy�����$⎶�'�9<��7���U������Gd���)������L����1�¤���4�s|dh�Xc���29��14t�,�ֽ��c��FP,q~��^%��y�{�?��nM�U���f=��/���]����b����l�5��W<�;�q�ױH#�ެ��iugg�1]_9cLK� ����
�jOt��n�v�$�ƏRގ�胴	�I�<4�ϳ�O�+~ݭ�k�z�j8~uk�쌕(7]�'i{�=�3�{�"?�vf��H:l�[�WS޻�d�M^6�9��j֝w��mO7]����u�~�G��"J��1�\m�Ñ�ް������`�J΄m�R90���홦���\j�����E�T�N�w��|5p�
mHJ�W1S˧�7����:�.�>��07�Z�㩔�/�_���E]�J���uKv�|�ċ�L���kƕ܅l!V`x��)c
R�V�s��~�-V*���#�؟����Xۦ6�D�.lc����v���l��v;HՆ(���˩��O�������m�h��&��Ʌ�߱���Yf��	�u��vzb~�m	���G�����Y-��7Or�)��
�>���tz��oF^c=	�})@�$�1�t��5�<vV�)��7D���!�d�Y_�<��?0GT��ް����ɺ��*lI�V��mڝsպa��)A�-<��m+8�j*͵N�[�@h��2R&3g�äT�����kG�2�{,ˡ*��"�A6�%���j&��vH��3=o&�!��� :&��V�zߴ �~Y�S�I��qg�x�be�!'�i�y�9�Ḣ��m�����^�
8����<8�mi�V�������y`�O�"�p��������������L��H�qT�Sm&*�W�_�i�#֐�٥M�A��Lc��D�e�ֻN�?͎׸	=��<o���n�osT�� 	U{�*��ƿ?�G!��{��7"l���'y�l�W�B{���Eg�՛@�#� ԓ���j[��%����b�͂��+y�Ƈ��OW�� D$�Zn!�P����/5�zz�cR�+�l5�$���Q�vS��#�$ˢ<���_��5��I���E6ޢ_�B� L��UM����b]m��L���i"P��N�Tw���Z�V���ԥ45�/DW[���V�b�8x�A?�_�UbHfp����̊tX��(7יq(x�s�Y��a���aiJ�L�(B)m�I�|V�Ȧ}yy��R�:�*O�P�`��K�|���C&\�␥'
F�Y�z�{�x�y�n/��,≞Y�>~t;�x�3��2��U>��i!w�i���@F�fS��ى�����~�,{q6lUP�7 �C�{��s�)����¬T�z.��ͶB���(��E% �E�=�('���p}˯���1�g�_�H��䖚���iv\ ����_��G]�\��ض�Q`IW\"*����ūj��y,���A�owK0��C(C�u?I�L�?�K$���"���T>ң�=�Og�	_ot=��������S.9ߧ`,��� ��#I�(k�a��Bx�L�j �ii�)�)5 H�^~[T$:
O$y����<�'��p�S#t�^ۣ'/G+�$��r��J����R�R���egF�e��fݣ�G������IOe�7��V$���G��ay�)terp��@><{k�腭�6�٪���۴v��Ͳ���ZQ^X�0|�
b�]7?��"��.��{Ȩ��!�M/�DN��:A��[ү&	�b-��c]qͯ#�5�Iͯ����!�i|O|�a[�1���I�w�X3�t>{�� \Ҥg�ݙКNC��$b�>�p�I�p�ǌs� vlI��~$!�>Ⱦ���ql#W��}!��A�'D�UԂ��KNwR��ε
��L�S�0�*ۼ�Q���L'; �٠�W������ -(�,��yu��A��-�Jߏ�h�}d4x�ƣK v;5��آ
���푮�i��֩p� 8��ʆg Q�[���-?�w���(]}I^�&L�M�l�b ���O�� �Y5ı!�nAC�qG&v�#�D���<���f.��%h�w�Bb�-k�(|ʣH� (:NV>������R@0���u�_T�F��Ty)T�kU�Lf��Li�K"m�E�������ĥ�h���u3mSC*��H9fܤ�����J��:Ѽa��9C��
�jn|���إ��$5�Ǝ���6���ZU��H*;H�i��B���➀Qivϫم��aq����>GR�y��S�bb¹��^�|�Q�`HǾ�e~��Z�f�rS�<
��S��9���^�Y��K��wٵ�MסV���Q�I���5'0<͙�?2',��0�9��8��k�f�5딎�^2��j;w/�<~Յh�"�5q�	�H��@�aJ8P�?f	)��ЇS(� �MES h�嚲�i;�vee��ĔwbK���˨�Δ�U	Kǯj*�nО PX�>�b]d�,م���^*�OZi��ڒ����8��x�����^6U�:�{t#Td-+����ظ�1��G�A����
F���jK�5�u��K�?��M�K�A*�@��X�Jl�tr̓ߟ��s�5;��g��!¬dxd��w>��w�iA*Xt���*�1	�G"]��ܔ�T�A��}����#Z���1+��Կn�P!�Jwۍ�Fw_OraQG
��,�n|$��a�i��p��]?��S�&��$�EE912��rYv~[�a���2��R5��TL��2�y3�: K�YQ�m��v@��=�4=qz�XT�F�j�>�K#�p�%P���T��q��i�P��W��Y.��ܗ6윗�5��Qc?�ٞ��c�ݐ+�yb�Ů�X����F3�,�}���S���z��FN~{ ��B%zj���u�wT^5��8����ph�o��=�7x&��Ak���������4+1$���=e�����I}�0r,/����v�s5��X�C=�L_ 7����Z�aU!g4nxI0H�����7��|�ĸ_�,ˆ'��#\�R���$�1�)���/f7����H�ÈA8&gI�5ӝ!Uu��w��@�vl��E8�D'҃
aW�U3�������4=Obxz�\G�
wgH@\�� ��f��=4�\�]�*&�\��g0��Xo��:���G-���E[sZ����ɶ��H��p��� s�6^�/[Q�F�"�{]����$1�����U,D1�t��y�*����Q.1Cx��ƀe�S#a�e�!
��M\$��BT�vE�P�Q��ZD�9��t�o}uڪ{�>���5����չ��f���=W��ՊU�������l��m��tk�U��F��� ���$�j	�(i`�,�"Z�P\��k��e&��U�=\LЗ��\����s��.�[h��4k,�����s�GF�U�$͋	h���ErK� �H1ǯ��m�sD'��h���0�ٵ&���^�%ҙ��`)�Ĺ���1�e�<������'g����h|��Y�M��"�����yN��ǅ[�(T�{�d�)$�.61] t��QDu����g&I�D���T�����K.���e�L1����m����I�n�Yj`2�'��^���+2�q�ˎqx}#�����rjC��^T�nu��)�u�tl�7&��/�Tz�����B=
0x:�d��2剌i7~��|R�(�;Y[�P��=�u����)�ޑ!z�a�>g>��D�M�O<D[��T��� 
Q	�63�3\�q�S������ �7��nԁ�١ ����td"��m��yaV���rik
c��r�u��bm{����`�5 �]��ϖ]YfE��	�y�D������澏ͱ�{1N�O��E>I�����Yqˡ-��~�t#��%�-��\`�J�J�h'��QԪ���q�\+��\Е���":�Ml�P
�'���2����A*F��E�O4��H5�#�l�vB�0�&.)� ��<'����vG�n�`�[�ߎ���;����]�XvG��s�j4��������8YF�x�/���jg�0�E�C>�s�<5(�� X$cqa���qs��WNm�`N�*P�rlQ��T�(��i����I4�0l���[��Xob�����m^;��I)����%��!8��<���Z4J�K�#P���쾐�V�KH����5�֟0�j .Wl\�f;"��n�Va����7���x���� k�M�ۭs>>���y_�1O\�!���6wd��HD��(�%��6��t'����?�p�I�Rb�X�?W&��~CZ[_���0�I ڸQ����W��5��S�PUI��}��u�X2��T]߻/��^��' ���W�ln��eV$��6�D4>v -`�ϊU���pkcFI�pM���{�}�}x�l믫J��l˽|�B5<zd�Un�]�cTP���ԋ>y�-ĉ]������O��T�sV��U5kmi#�c��(�@'��7b��M%�a�=V��ۆu�R���nmyk��+���xE9犮����]�1���0��B���:�f�S
}W�/.�"��:Z���U��)��Jg�Ӝ5\��ޝ�Ӗ��]���P١��z̴p�8vTk��A��#M*}iY��Ƒ.)�bk.D���;q�F�܀� ��d���5�(,Mh;M������f�s�,���%�^ �T9����a8��k
Q��u7Q��ǚ�=큮�jj�p~�˃�޵��Ù��d�`V�;�:IAYtc0�����S�Pc�\Y�)`©9V����2��z��D���_x|��$ǀJvoX}a2��y��>�/0�7�{�U�Y��-[�b�<�>Mk��"S͉�F���2��	�rH����!��g�C�G"l��8�}�jgvu'��{�̄ˊӯK_֟
;T������m�+ؒ�o�"��S��k�%��A����FN�j9g���^'H�i��*��p+�_Y2L+��c�oV�v���΍!��=��7�l��� �a��H��Ȱ�y%^t�1�˰#���-��+=g�Ӷ�	�2RG���Z�if���+���m�g�W�D�z���91���/0�Ɛ>�hGAf�:�uy���ڞE�����OՋ�J��P��E����/5�TMdJJ#���F��3����lA�����ݪ�`Z��S��>�N|����Lp�
���O�B`�X7�@ U��\���boX�)�V|�!~�u�Ի`�����n:A�׮F~b�PǱ��LلH_����S�3���-M�(U�{?��V�o�&O����<UA���Iv���<�[�4��JW��t�AplN�Y���y}C�;6<X������%8��R�#U��u�;+�9xA1���My�2-�F����V������C�mpfZX$���}k�CIl��6҇;�T��^qU����?�畅��fB� �|I
�%VeJ�ua7�M�m��W��:A	����{�v�{�@S�]XD\`�uq�f��}�^?�od-S&�������3JÄc�֡}��(��P����8vq��rf$�ӱKu�l�@�+2V��$����Z�ܽ�8ښԲ_Ke� R-4��M1ri6�:H/_/Z��/řk[�h�k�
�'�>��?Ji�����2m'�A�� dR����#�����=֒��`bc�G!Łt]+1�1ǂ�c�ߪ³����9,�P�b{�m�/�%؀�b�wEO�6R~ �����`ƙޭ���|�д�B������XF�U��cMgĩ���e��V{ƞ���|kC�|�l�xn0<� �h�4l�W����(U���!6��zX� �[zT��;�/Y�zv���d�膝��2����so��ld���ĝ�(Gލ��ERп��yY��OY��F�>s{�WەD�H��〛�4s*ѓ5�By�r�^^�r
&AM��Jguz��;J�7M8��p-��8�A�Yq��1xd���ɲ�6`�v���	LS2C|geqY{�4��ݴh���xL��)Ub�W�y]@�ss<� ��!K1��?���i*�{ߚhA���JD/�u�~�qt�,��u�;�B�%�iF_�"���J�>�5�y�[���2��s\��T��ĝJ�sn��r�K�3=�rM�|��ڗk�nWX[�+��J^��H�-�R�1[@ḸQ-K��T~��Bb�$�W�Gl�w���?�c�+߳�B.�E`h+)W��*�Pݖ�8�#���kN��Ћ��8��JC����v���\0;��3�h����l� ����;����{X��j1�ndә��;� !���@���n��-��.0�hXQ�w�[U
����L]����������\���;):u$��,�� q#���Nr���3�Iy�r$���^o%�RK�nO��w���?pw���wu�kA�i3CXw�nП�R �u��}����u	Sj��R�ɦ;+�Ye��LxAiɚ��tˇ-t1C'��,��ϧH�tfk������L��a	
�H�a�3;�)���vH����J�޻R5�/[��ڐ�gy�63~5f�:�81K��dP=����2��)��c��|�9�Ƭ���".�;�)�ƟO�L�~GK��O�ų"���\y/�:�Gqm�ro
Q.kl�Ѳ*Y�:gR�t�m�$�s�a�j�k��J>O2{��2|�������p�h{#(��W���Dw��]��m������h�T'���e�H�x5�"�X3�$�"3�07���"A0`ټ���t���w�6S�������-��0y[�;̀5���`�r�Ï�e "(^����ѧ��Ng���RS�7o���%Z�(92D;`#�ط�#�.V
�9W�����u����:�>��.̏�{F�ejʳ6��،��2%�X���������}���]�-�6;��~���XI��,d��"n��46��%lP{�p-9���y۪z��B�Cf���»�'O��s0�6����9��<�/6N�g��q��-�?�_<4�0�7��S�5���L DTn9���!G,��#$�)(y1on�� ӓ��͡�}P��n�a��6�@3"��!����h6��Y���#�X�� rID���8R�8l�f>Po<`��<���$	�o��B��m����V��Z*ph��.�~ׯX�i���� �����ش�q)h��UZ��K��:d�H����&�M=2{[[�¥�q{'�L����:�+���k�{7���߸��9q�,�|��iR@��̵,�ȯ��MW���K��R3z�����R���֟Ⱦ~����w�G���Ue�@�B��r�S�0��a����S�������h��13��&���9>�9�QK��_�s�C�U"�-�i��k�̌ܫ^���H�uIm»�-,�R8���j�U�cc���7�tnɕ(}�=?���6o�*W��MO2�#�E>�<��q����gV�g�,�7M�:'AꨍK��v�p��pq�Q�v���3�Ư⭆4��1ɀ��2�r��
��5��<T��D�-�
���au3pf8/��B\��-h���ඁPJ�{��i���a�қ#�z�?l�9�H���e�1�ն�鹳w������Ǡ�R䵐؇�׾�@�DL�M�w���%O�w�Өv�F�,}s�8�U:�>��s^IDUA?9Q�Lc�œL�s�mxr�Tu���^�Z�ea�U{��	�k����h�s��pӼݙ��d�z����̕T���?-�������\'/=O6q�d�0�'=�sR�V2p6��}�^�os�{���'S����55�"%P�n���f�jFsI Qʟ�x������f�#�NJu>������i�"|y���Th�\jG�XRz��qj�u�����&��ũ��a%1 �������DV'�{��q��c ���sH��I��-���(Z�\����M㒟�ѨD���v�����ld�F%�Gwj������2y�Ѳ���l泥f�+�̢k�{8��d�TI��0Z	�x&j���˹�k���f�;=.΋Fg��A�XwN�0 �"�����I�q���N�SERx����l���mg�������7��[��$���=W����?�����v�Y�֔Tb���<!����x<oԔ�n�2�2��A?�M��r5��l����z��섔�t���AJB�Wk�6���F��A��b����I�%;��8��|Ъ2"ZR�OF� �<��C,��âa���{�����=���T.��v����~������8	hC:0Z�R�A�׷��k�Y�bV��2��� !�����=s��	��W��������(D�N���DL4�A~�����)�Q>V�%0�*;��z��U��&v]��e�.��G��?43F�F����Ҟ�8�RG�r��Z �N�m��@ jq\rV;�Z0/R���D�m/���(��$(m�iC�fMB��p7H�P�	����{����tUq>�G�'�)�[}�O1��$�R�3�	+��_XD(�뱺ҍ����
?"o&Dz� ���Y"d�=J� y�勓1t�$�f٬vv�$!s�u��$9�:�!���t�W�{Np�w3�h�I,+���k�.�q_fC�W��m���h��� ���J�(���7��'9���S��Ke�>�x�ڡ.Fl��DŇ��vF������7���PO18}��7<+jHv΍ ��.~1�{gF�����_�8��gA7�����e%��!����4��[e�3t)���&{9t�2j� s���|:x�����@�al��D��~<��"��e{�5�(�I�~�r�Y�R_W)����m�^i��8s��['D�88�f�
=�n���T�U��!�géC�@��Φ<DH��跻|ͻh5��T��v�VXI��$��1�@��2�0�IF�d�̺JXg�v3�,���L�P)�_�X��.r�]�:���MP�%)!�Z�1�7�PIXeA�+�jƤHxw�Z�@���ù.H|�/<� 3��&����ώM,e�b���#�g��U�CP��*����f�xK{���;�� �x,bm����|{���5(��~t�)���_ҳ��dC1_�T ����iR��p�h)�	R�x��K��
�S�W�5�.�!8���x>ªȒeI,v�$D��GY<��~�!|A��#߮~`�"�t=9�ʿ`��3#�%2�{  �� ��]�=.��w����8#����|H��}S<:���i2a?����h�~@1w�����,-)�<�����kj�����-��*>z����nk� @��P����=3O�L��;�x�rH�V,�[B�K��M�^6j��]b�r*�@�!��%�U�hwp�Ё�r�j��b�P�Q'���E�m/�;�(��\h�Sy��"�#"(g+{��3�g��L����>�V?��0x�a�$
/������a���j�R7H�6CIGH��H(�QO��	ɞ
�����/s�9���3̸��|�luss�I�q=bʁg�6O�f_�ʏ��׵���R��;=�鋧e�áZFe� F��=p�4](D����̒��e`#iQ��M?ͮ�N����C��$f���Z����S�)���E��X��][�O3SP����1����01ŕDFh(��ߘ��l��W��z�y	�6�{:\^���w]�Ӹl[�G|L̓\��Rݚ�E"Wh��g�#i1���D����hS���~���nO��s�H���.Ǫ���t���/KZ�\��A�$k��w.I��$�>��gAmTn�h��GN¨��6���*l�����/3֬����
���gG�kX�G
٠�����bJI�O}��eu ��K�To�4"�ıiȓ!�rV���������\���$������a�a8}��D�Gg����J�̵����v��iH�Y�r�72/�?�"�0���xA)� mHX�aj���w�I�RÐ��/�D�̣��pF����`��X�$�6��{P�:���cx_K���_�����;����w�k��zd�,03޸,5�l�.�]���7G�O�ƫ��!���w ��,_�@풝�=E9͐X��W���eyYNiX��i����ޓ��K�Z�5=�4�GS��D�(�N̴��6��Hh|���F�d��M����JB�zZϹ���ǿ��({�!�itg�����i�H)LBlg���~���Ý�9+ءˌs|yO���S&�=d��E�k�ת��x{������0)��7�(�ʼb�eN�^�<=hp}���r�lg�Hs���L��L2rGb"W!*k�F�TK�V�c�Gi��� �PD!�N���&Z�77��=n��Q�`�3���ET��iM[20���j��r�s��+�)�ι�w],��^x�MN�,KyⅩ]�^%��`�!a�]2򂗕���7������+&�!�nל]�S3��yeξ9���
���I�?������S���Ո���wO���h���2#W�,�%̐��:];t45,ꓮ�Io���HǛ�����:ã�����x٤ AM��nbH\�p4����/�d���,P���PпN	3}췘���z��5��.��n�Ӥ�����Ju��	f��C+¥��T�k�8����(r���6:��!s�y��	��4�9����[�-R��2v*��n�4!LHXCmN�����-kR'�"Fc���W:���_����3?�j�A/�V��u�	�|�k�Q9��T��^L^�UB�y��ǵ�o�M��Ton�[�]+�K ��ՐdH���du��f�3m��hd�]fH�hk"���7��T��z�T
�����t�d��"�pd,kG�[�˴�c��X|�Ի��D��[ ���E{���A�I�4��4G�d����8�~�����ԯxqGK��F3��ϟc�C7a{����x*��1Op��m�n���#c�,��蕮S-��EC�A�Fyg��%�~�]0X:zD���}%N������$Ll9�eת �*	 �%:����}�o�Dk� �*�W�IIޙ7�yK�
��\ã^~���B�k�Sw*�˨�.�H)G�6`F�v��w��B� ��7���sWd7gXE&�G@q���bg�e��]�܏�ӽ���S4��@�1�n����=}�R�p��)�f��+/���u���l��٠�3_k0���P���QH�DO����k=%�7�ݒ����焯-v'�u0�Ŕu&��k������t�9w�&0y�V�����r��x�|ʢ+FP�y߼�;݆�<�T�/;kyqfy����~w�6z�6{����߯k1ӝ)5�jo޽��
���V�T2��r1n^C��ݙ�8J7b�_%��w[=ƉD�mN� &�4F1K	�>U�:(�s[�<q�_�O_��N�Lj���(p8�³-6'������J\�T��RU"�Z����žM9��u�y�c�pT�r��L��ro��Z��2^Vή�"�ս!æ���B&D����(%#y�WQU����Y�����&�2����:m�n��XFsRg�}%����)/4��H��ˡL�Xu8Vv͚&�3���u��L�2�D7z3��eo�y`ҡ�>�!�Z]�y/V�?���Z�ugy�ȝ�UNE���f +����{����Gy,��_�G��Ǘ�!��z�����$R�qA�]�?z��R@�4s��˜�e�N �h�5�L:qe�@8%����<�.�F�������!�f�9��R�foE��w;,o�]�����A
=�8�u��Xݍ��bSj5�z@$���ő܆5d�P�ɍ{���Z���7���mg��-�C����3�@y蕸p~��6I�,���͗[���!�}o��y_!Y�3���S� �[G+�]�T���k�j�A��{�=��I�"we�~��Cs���w_����HeЪC��<'��PB��f�lE����4+\�Ч�H0w�?y��A�dX�L��;���B������Z:p�(�)�`QI^a����g�E�H2g�S��޴i�|gm�|c�T����<�x	4��fT� H{�?����C	��y2���A�j���$�#�_ﯽZj�o��v��[��,�y��LH"~�����}�1S�����q��8�\��+�5��' � ���ʀLcAT��%���D/��[1.J�P�0�ل���v�x&�Xv��ă��(6���Ǫ���VB�c(�W�(<�H�و/M� �g�y��1�Lt�k���Ѹ�h�d����x˪2-�Tb�-��h�`����0�j	sb:�G��$_R�N���h�^a�n5o�~Q��+��I����q�~+���9�H�j�<�\\�	��L������G��Y��[�x'jC��#�����ڴ"���%�>�)��j��
��o�[�8��:��q�t�m[ŏ��+��!��8LX���Kx�(���+�� r`�ۥLv�}D���'�R���Z�O��~�ږ�`~^&������5���@��v59�W��Ҧ�W4Z�!sh=[E&�/0+qO�F_	v#mk��GvTD��,f����Q�}�9���8oocoH-��3H�Mk�6�p�����N�ɏ�@��l-}�2�1~�� �ݏ����dG҄(��ZMV\�"6i$��s�	��9"��U`2�e֎��*��=k��ˤ'ʸ��E��l�n�y�RmX<eM���1=����QP�G~��^1����S]W]��N��Nt����g)�&n�4�[�IU@2� . -�)�crUf���^�/I�V��Et'��M��� �ʕ��gJ0���]��l��bE��65�cϱ�[K�|u~ ��|��/���ѝo��	���.}SeLs���l�����/8���}�jT�^���6�͑N�皃?o���m�Ùǋj�N�8�x��͆�����yV��?qBo����,�l�iŋ�EU<�"��((��.�Wv�e,0�9��@�#�2����܌*u��ᥦJ ~b�a�?sH����V�bS��%���l*����5�uwR���i(J�k��܅�{D���=�$���;j��C�v��}���Yq)$l�Vq��f@�G�����z@c��zh{k�`.o��(�bqݗb�k����gqA�(X��Qy�UV��F�z�ۻ�ˈ�s�/Цq�"�nЪ_1͓�6d��N�=��&U/`F�ݭ(��1��i���Bc��w7���d
�p��C^����)&~Z�E�M�ê����]	��f(Cz4��h�b�Z��T�dti:�@ߩ=@2(�Ȏm�R�G�i/�bޜ�����"��|T��,*Jr쾞|���A�l9���ddiO,�����4&����V����γT��.C+[�8��Y�[�kCk��7��;�g�g�T�L)5�z���r,�'j>nAa�(�p2,��k�C��������R�m�E���z�.���qv���}�s�}#^��}M�q�S��0���wD~�)�[03��|���5oz:ks'�X�n�{������`��ʁ!��A��xa��}s��-�P	%RGu���b�Ծ��V`5�7Z+� �y�E�\k<51t)�y$P�{�ˑ�m��'|�� �ڪg�z@1z�a��<�"�t��zu�bA��M���ć�?�D�!�_.sH�#"� j��Wa%�	e��أ17�m�g��7>�On{���$s?�f*/vRx,�t��V r���7�I�?9Y�8��А.���dS�=�39��k��w���RyP��.)N�uG�����K��y��7O�6�� ��58����$��f�yK��-#��NH"��x���m5�K�� ����WBu���-��捤��Q8��_�Y�d.l�����Q$����uDR��*O��oJt�D��rh�Df�L\�L�7 ����a�1;��kG~��N�&��FOg2�ueĊ��J�VVҚ���q^z�t��uzp�����e�w�1ί�`"�wh��9��E�~�y8b�'�l��ȺL���r�X��O��J���N8�&V=/�vN�#,�Rc�rl3t�dPN��AL���`����e��7z�ݼ��F㪶v�%`���c�l% dݬb�U��Sm�i��p&��C2�X�7�D"���^��q/5��7� ���ܨ4�$Z)ucX �p��t!��VC�נa)��@�!�[�T�~�;���
Gt������(<�*���4m�^��T���������uR�>~�6���J5.T  @�y�OW���� ��ĩ�xhtꃫ�X���3[Ja'�������-9v�*��W$o�B\�S�B�6v�V �����q4�J?���.�g�h����|W�E�=�YȣҦIkX`�\l�j��4y��%їJ]���Rv���v���8螒�ԍ��P�Q,� sPf�ڻ�)���] �e�7w�DL����A_x
��SE\a2����v������M�qu&Nr�J��|�K�i�c@��6�(�*�:����Δ�DZ�
P?P����Ko�E�"�ɻh+3[2?^H)�[����K|<��ҡ^_�4)m<���:&����8���%�7a�C����t�&�b<m��MLu�q�k�M2zp.@��v"=OW��J��_�Y�?y������>K9"7Д��T�z� �� Dc�^{�X:$#$�P�D���Y��c۸@��X5��ɤ�ҥ�����Ye�8tj=w	P-	�֫������ثN�?B������K�e6�`膐����;�| ��?�C�����I��{}X+�[���PL8fV��������L��� �o7S��/j7U��F�	����A��TV�fT�ދk�5� �)F���߫[���@>�m'�t�Wٟs���}B����ALO�WpJz۸�0���Q�ց���
'D��<&>�]t�p��)�ʇ_�����8��0��׬͘������ю�����oNE�xA�7,�C��5��Ϛ�,��:v��2�,������C�$������l�T|)����v.&@r�*��'���^�[-�jw� *����@�5,�����4���Y�[`��¯��6�a�睔�(�JdR��2&W�1�.y_�xo_���u-���m�w����s��+F`@5���*yP�z��}K$
��n8Zʾ��7��f[/� �����0d�,�7\���Y�	���!f�J߈�`�4�&�����]H�O��Q|h��ͫsc�86�1q���֯7�W=3�n�Wys�H'������=�~�Q�DN�hY���w�l��_K���Ⰼ+�Cm�C��Y����HI����=�*��`|�U�%Q���*�e�p"'qM�w�1�<j"�=����fQ]d6�Q�9�e4D�*G�{��^���$�u��ٓ3*�E�A�����#l�����e�z��IOW��4�e>�⩱J���vv�I��q,xcƛs�ya=H��|��"i�VQ���C�f �>�����ؖ�/:~z�BU��5Sn�0��л&E�o�����x#M-�ԁCK�%�?R��"jaE�y�7����b������B��{,)z������m"��>�/\,�0����ߥ��~¿B��\������,ϻd����	��q3�-`��i_E�Hf;�L���]�s�\M�,1`��~�˙艦W�p,�r��z�?�l��Ȁ��qF~��>\=>�)��k��8��]7{fu��ZS�(���afώW=b͑8W�.�l��=� C�2�/��(u'��vè�W�L���)	�H:)ֲ�(�ӣ~[}+�����H���M�8,*��S�,�_����%C�0u�6j.߾]�RM��lO��0��[o`�R-�qE��,_Ŧv�,���)�i`>�Z����v�o'����Iz:tG�r%�vݏ0螱�Q��|��({M:��F$��q���F&-��w5�%o��B�`�������~����yS�l��
c�;|^��@�.b�ŸC�U������c4�~��M�`* �N���cd�tPUf��_�7l\>���;�V���;[�]�k��[gɂ�{`G���I�d����bÙ�n@�NM�|�"��Ĉq��S���L��`����3�8���/���}ӷ��rf�FM0������
zsK������]�VKe�A�|��,e��9�� \|*�b�*��oH0�@q(=��f����I�����tLW=K�\��v�?��\�2j���H(�� �0gy:y�=��R�kܟ؁xb�)��u���ԭ�"���j�>ײ��o`��~h+c���V�?�c�#�����aFK��a��!�n8U������fI�+�>U +w.$.-���k�A���W�b�t�c�ap*��Uc��\��k���^n�G��}R����~�r��4�ô,��%�v}��t�-rQ&���@���M�z���h��Z��;�E�8Зr+0��� ls�d�k��~7��=C`k�E~]&�H9�r	��8,��:���F:\K�g��A׼p��phɃ�d<G�ƲB5I�
�U}����?��Kg�Y	m�Ҧ���n�i�!��D*�&40?�?L�\�E�#�
����)��3D�;�7�H*�jӞӜޛ��x��8�DJ���+���W���5ߖ~^�	� 	�9��|&�3�4�رЊI�R�qʺ���J,/?��dH���O*k����w1�9/�z��9Fꧪi�'�)���2w:�>�;Ɍ�0�\����7���-5h^-��)`���-���7)��&N�.�SЃ��2A�e�Ϳ���W"[��jE���*8�q%�)��T��D2�H�@/�)����/4|a.���i����Bow|f⊞�5�������!�ՉE�rŝB���_G��g&	�3��0u����D^���vyb,oEF�E��0����1m8���L ��a/���G��8 v��*�޶9s���n��xN��Fҥ����`����K��r4������>��H�q���Łֳ� 6A�2�S��8�R�peJ����3����Qx�c���	� �ڃ)�T��$�Ml��W����hM�xjd"�`�f�iBL�mAD����j�B썦��D��	���tPgU���g�G��X}���`w�К�.��M{�a��9�l4˙��^��sE�ӥ�Oܯ���-�/�q�K�O!�u	#s�ԥ��z�4`��yP�0�Iyu��.�����>$������L	���vx��7�3�D-]s_�D1S|6'����7�<�"w%]�|�שA���`����͚�8�\��KkH�a����<������|Ћ}oE�t��/`�1Wը�-p���
5(���;�����T�-(���{�ؗ&&�'ѓ�Q�AT�B�:(a��_�%���3{�T+�* ,`2�G��BO��
�	���Mw���P�����'H���H��m��	q���Ʋ��q���]���¦�,�*U���3Z�쀾l��y��z\��:$�҇�.��g�\�6�{Ǉ���q�Q8����|��_i8�)z�(�;xW�������_L{6b�=���Se���L�*���}	��'��yj,�#p<���6�o��F�D�$31�����E*�<����Ѕĕ�ċY &��s`ƴ�E���3��(�q��~�V�g$w�nV��!T�]�#�KJ�����o��X�}>�o4�JN�u�m�D��%��kg2�����Z�{ִՇ���tpC5UYg������E�Uj��L��y�.��D�Ȯ%�e.� ���U�͸����CCTf�<����5����7�)�f����,jX]�O0�X/�VX̹����J�=����Ѐ�+ r٢ż�+�������y(�M��E���W�Rt@�X�/�D�gZ�a.��l��{�*L���z}�B!��T�f���u4#H;�̺�f�S��l�^G3��fjI7Eb�QU��63�P�z�|a���~�yc�v�wI�"�'��E�X�����.���4*`t�|����}��	����-v��� DO(i��_��B��88�VaX�� �a!R��T��V5�9s���ـ�!|�P?a�/� tPAc�C�-7e15�&���Hb�=�e1p��uU��t� ���5K
&k�L	��qx��%>�d��I��~�L��c���}Ȏ;CĂ�xx*Qo�UdO4�ˇ]�񽥭�DE�k��Ewur�D�Q��!���7�X?ƾ,�`��
i3=��#���ĵ>��w�1+��/���>�C��Ҵӕ�o0��y��O�}���<���<�e�5�la���M��0d�pI��L]�x��N1�ɷ��A*/���pN�ҥ-�?��H2w.��E����~G')�7ڡ�.�iQ��ʮx��)��Z�RK��`����50g���!7��ٞB������w��_U����AH'J�d�6]`��:9d��ZZ�ʩ�2�_�R)�R�@��������,p"��a�ɧ�
�1�&Q�G�E����)�	~���>�ʲ�Z���t�о1�e�/�"�0g!H�n*���.,蜰j4��֫K�+��^V���:4~֦or�yJ�E�nd8n�K~bm�̶X����u
�/�<�����t�b�j��f� ���9�ty���(wU3��wi/?���+�u�-ؤ��pU��,?M 1�ܝfg�u���N�ƺN0�Ax�ռN��� r�ۖ����૘+��gJDJ�D�3���K��X�_�+�����f9���P�}��(xy�L�b�]Ⓖ%��?oB�*��_: w�B���Ӆ� ��y;I���#hU�ի��B��*��!/�ԒB�C7�t�H�!��:�������EM8�=d�Ҷ~faR	��s��㫓E���G�#�����9`�	��.^�v�#m
�<�۷�k����\{���������4���ݬtM���3R�N��&����+<�Iǧ8���Y�*���1f���볙� �'µ�;��e��wǥ��N̅GK7�iRP�?�ڰm,�x��hig�̱�g<�E�x�],�+ؘr����O�6�?F�P�N�x����B{{.=�'�ʲ�&��d�s��.�,<?I�]�������a�����W��
�M� šU)de5�UU�8�&3�,]�ߋ1&��۸�J�b;���-S�y���7汰vΫ=/�}�����Ol�)���l�~GT2Q�Aq���m���P5�fۅ�pl���U=���VWe��FB�ђIz�������(�3<3|4�烣q�} �=y��
ő����y���#Ѧ`��bOO�
�F7Hڈ���\5?��p�yEű���{x�\���ź����+�����ȴ�%v��l������XA6Vr�N������)+�2�v��S���
պt�VD
�P>L�/�Z������r���v��F$6��jT��;RE�­�!�J����,O/Չ䁯,Ŵ�R�EE9�>�q�lNvQ��Հ^OS���������b����@���=ۊg�⯞\��vO�7?� <�V0Հ��a�d���(�|dBb�GCY��t`|һMYLuR��N]�Jllb����� μ��'sjQF���n��qjv��:�*��i�~��{�/Ubn���t���lm�ڕ)��ⵊ��˕�Q܇+ˆr��<P�^��b�j���tm�Շ��u��˰|x(�l�#�&��Yu�Y1Ƀ�t����D��o�@�YQ�/��Vi���3ō�CV]A�_�����9��`"j�Ii/�v/�굿/t���"�>@�Y���YOZ����VL��E�#�܁;z���.�h;w��*OM&��nC��zm�!�/�> ��y�o�	��)A/������ZZ�2F	/�L:Rd.k�����scY2�l`�@���n���h+�i���%{i���>I��z����DR�N��/�|�ek<<��3ᬐ�D7�aJ=�D0�2��ߵB� �����7.���(��>��cL=��8f9��]V�D��7r�GRi)��J�k�Ls��� ��e ��h��ۼ|�\_=��a�=ʢ@O��b�(ˡ����/��o��q���ܝ�z5�ұQ4­���r�����h�1���^��-���KD��}-�+���:�x.Ju��[�B_r��?~����ʪ�4�5?r'c�u���.�O�-،ɿ�g![du�5��TA��Ε闱`��k��ykL���o�����vF1|��~&Y%ܷ-z�Ҽ�/}p�7Vm!Y3��Π�c/���۪J%Ov^��݌��k�t��nh\�x��:�_0�������
��[�i��h��
U��`8@�X8 ����K���q ��EB���v�qr=�'���Vp7Z��6l�,A�ĭ��R0��G{�s��i>�	�*�)A��q��c9N��/u�
}[�u}���t���o� #$�7Q%�M�p0�ok�;_H�^)������K^��"�4V��K�R1���9ft�'Ә@#ޔS1;�^9uOp;�"%�k�f�D:4�.��:k���mJ3�\ɥ��B;x`�������PoU��s�����a��=��C�q�K��K���oܩo���6E�c���up��N���O:sj�#�`�:��!�a|�|l�QBD��;�#�>����ĽA�I�n�
�i�8]k]hT���N�*{�3�5J�%(+�3S��yM"*et<Z[���M]���2���#.y��=s6\4x!���r`�ȱ��5����	}�Wpq�V,�������4�T����;5�7��Ĕڑ<�,,7�����g�@g��#�!�lf����H=�Hm�P��"Ow�o�"Q�a�xԦMRݚ51���������(�-2�.�ɱ5��翙�	M���+��7m<�N`Oe�}�b�#W�H@�7M&�|Ph	P^|��U�O�c"����`�0��Vά#���nzO��OQ�ޗ���D������Ĕ`e�	����s�_~��?O���Uf�S#�yޠ-���0�P�sf��ʡN[R?��}�B�4Ds�(!2��e��/��=�h's�Q�83�ꃎ�Nedl	�>��P�{6�fr�Ҧ~͋{�_~��8g�꺈��cW��G��S"�ޯ6�b��� U���������"�[��kr?���Ӵ�"��c*�"oO}Zn`iR��ͿO9���)�k����Ԫ������Tf/=,�z��F���n�nOa`��S+�؟������'�`��kJ9��~��V�@��}�{!g�ǲ!�T?:��C�I�˹���1Ä��)7�w����v%�#p��� 3+�����=�'޶��"Bhwϱ��_�,FN��,������6>;�X(g��u��&�s눖�N�MgČ�r��^���Ed��Ip��."�����Ph�Ϲ��g�F^�	�j��"�
�����	x�K��D��W�X9��'��-�E�A ��wV��éC۹U/�C�ow��<��ok��gm�!B���,�\q��w*�������o۱A��Y�l���&�v�v�ݕ��z]9k�=��$5�W�����*�O���+p%)k����q�jQ��������L�v�S�1:ΐbl��tS��ˬ�	A�i�(h��5qVJL��p�2���_�����iZ�ϫv��6fl�5��y*ƽ�x ��"�vM4�c%V�'A]�q�� �s�F<|dʾ��.�젗��?ú���>]��E���Oh��)��_A7�~���,�|a���t�����(&jb5�X�PK��@ h�;ٶ�y	;���a�C��t��s@��J@ԉ��B1�RZ��j�5�%�H���s]��_��%c��C�o�� 3A��%�:�X�d� �11�!Y����W195�Ql-�2?��3^�Vp��Q��nWU�:z-�iM��g'�T��k"�jӕs�w"K�;N�2��)q���u����7̓�u_�+`�:��S�i)�kj��b���A�VZT�sIoc����a2��� �*��pw^����.t�K��^���c&W�Y�:Fﴷ��as�&X|��pG���������a���t��˫�Km6���{�h���/X ӭ1<<� 0Y�3,���H
� [�'¼a�K�ᤧ��c���H76�����w�_֝�m�l<��Bx3d�:qE��D�;|?9�(��l��h?;��]sV���I��O"v�:Z6�z�7���g-SȒ��>b� ��#���f7�q�Hq�`��9��;��G:���B�o-�3�z��V��M
���p��p�'�?�A� �4�6�4���x)�Q���$F�&/�H��Q.�@[=��E�a����H�%(:X1������o�jo�/���3G�!�=�L̙Z*>(��g�)�v 8��,	`Cf��iB>&�8U�6�o��R���(���ڲ�;�>���]$����n���*��'�B��a�9�eh��܃ίm�S`�ڀٱ����P��ǼI@*�~�T� ��~��(�#¯�$�$���ը/����;-|f�_�������n�f$�U%.l'5����l�=�9���O|����<�E��nj|b��6��kG���Ӈ��mH�Dَ��T�C�G�.Hy�8Z;������6f�e&���h�B��o�WE�ZOZWj�̡ۖ�d̫5N,��N}?H���B�J9]��	�&��� ��Pvi�����*���d��)�i�[i�#�XD�t�mK�XS(�G+{&�ؾ7(��
�>a�)�w��M��4kD�l�V6��C@��P�����j�]��_���~5�2�/��ha<;���@�>��d,��S��}� ����Ѡ��ֲz��{vj�ۖ�
g�6�fV��6�=_�cϜ͹���0��n�EƔ$����$�e��j�JEoF�#[���`-���v����+�
ef���`��DY���A�K�o)Z7���V�Bɾ=bH�`��[G W������*!3�h�r�V{��l�Tec�����&�3�VqҺ$�Ӏ$� �5#Al>�jP�g	��L(<=�Y���m8D�"[d�Bu�%�G�����}c�nlT��iS9BIfт���?���a'\�F��S��ҟ��P�P#�8�@��"�f��"X_��D���Z��'�DE�d(]`�;���.7�����~�4����E�7L��0&7TV��l.���q������N�0ۨ�ӻ�',a����j��v��o�#�1��ᔴ�2O[�b���pD���F@���A�L���~.ߌu��qx+�g�_�g���0*�Cj�y�غ+���/�n�T��Ģ��$N���ʚ�{ ��G�M�� ,�
����E��Sç��S0`&��vk	��N��e���e:.�
��2�^dSGx\�4�j�ntc4{�z��wK:�0��#���
l����:�? ��AZqSu����:_� U���v�}�O���h�a`\(���	W�%��24�����3�e�BɆP�0y�2��Vv~�VX�s�����]z��uۡAR�����I�
����ݴ���f��֟�һ�>$ݨE:����e�u��Z����1 ;fy�B�X���
8
�vM�PN��!�&�-��$�YT<�g+�����D�:k�4��Ҿb��m����Sk5��,*}W�07}1�P�w�������!��B͗��Â�m)�񉔿ߒfS�����	�CY�{eW�1�049����8����9d�Wgn�i�o����H��m'Q=z�-h�x�F#����q�����V�"V�W�%FԈ��	�u��x�I6���R���+�$�(�QY�Ng͠����5�C��8��
dfIJ[[�_9䟩�jk��u݁�?�2j:�U
� -����6�,7�aս�":�G,���E�[x%;��VYS�!d���uv̫���S����B��gZ��U��i='!J������F�H��4;�������|��1��dGS�G��7��pH mK�,q]jՖi�?K��X��q.��mwc�M��D����m��9�#����pG�n|������oq6�I��pߚ�T�
�2Ό�|ŷ3��2�fD"x��M�!^��F�0F��M~���� 
�}��#�tn�ȁ����_CI��[O�`��R?����Ci7��{�9�^��T4E:f��C=�8��1�͋�?�PY
�`5فP�B3�i1�Tt���eR6����&��s�����>ο"bA�1��@AJ�T4l�yD���+��@��Όmq�7K�s(�5˜k��c��:�sc4�voH��#�Ч⃒�c�r@��P"#�?ZT�+�zk���؂KФ�8�1eV��{�Z��:K�����cut�&P����^����L|��������c�0�;Vf�(�!������76�g<�"h�X�jO�w��o�M�o�5M���+��΋+B�H�"[#c�Qku~�¦8�j' ��ZAi]S.�!�d���$�cE���L;�jbl����&���=���H�~�D�;L�d?�\Ȑ8�v����@�Vi�nx���OJs)�K�*Ce百�4�.��7�.�`��|���*��?���S�(�僸-5̨%Ѝ���m���u)#�,8��S�Xi��D�Ŧ�HYL�_}����y�2�p���R��Ĭ%	��+��T/"J�T�g�4��_
j����1�Cs���I]݃��P���S��M ��R�*q�,U$�a��Z �r�& ��8��p�]A+�nm]�l5@Xcȳ���`ӈh����T-�.@�M�/��O��@¤�E{�^�RI�wz\2�pKڹ�(������&���&Q|��H�C2��(aL1*���\��+�[)i��m�UG��9/�G)w�MV��n^�k#T��G��ϟe"$"H���;�����X�G�z���
K�����P�|͚P�k-1CU
��e��&jܢ�f�������v�Yr��X9����\w�÷��ܚ�	�a0YE��ߎY�Yt~�.��'��u�F���Ѩ��v8���rZ@H�>�Ӹg`ށc��Y���0'�����X�󞗗���
��u�&	� ��F��+��E�o l1Ff=}~�1x&� ��r�������6`�BI�����׈WRmȕ|e>I1.����"jj\�Ūh�B�8",�d/�7[I�!(�*�͋�	�a���P\�҈g��@1��K
Y�O�ٱT�Y:F(�52')��^q¼lpPf�:��}���`���+@��9C�LI��L�yda���ϒ%1��j�8@�@�.K�Zi��RtJ����Q�zF���$�Qt�xҐ�Z`K�#��X=��7�0���~��"��Ľ�X?�WǗ/>M�"��>��YT�Y�Q���C��k9?��09���DYF��N4E�����%��D��1m��:q��b�%�a�z|�
rKŔ�h>"ղ��Wv���^���r<��5��,W�RX��Y����W�(Ox��z�nUM��gO�5ܛ�4������ZNg%�&�"�ֵ�(3Z��cGv2Rst�Sk�%[�r�z׏�y��Y�x�N�����'VW� �LR�˼w'�6�Q�d. ���*v�(�7�����p�}h9/��ӕ:�9�O�y�QFĦ,7-��Hlf���X���+(G�CF(��rBs\���`&���H�P��9�p��X�)r@�m�|������١pӱ���
���鹑����>И��%�W?�!j��b� �W�����z���궚-'b�+
�Ԑ�<��9i���ho���EP���4ԝ��`̂$Q�qGf�kF�cڷN�q�j�ä��QfD��j��?����A�7HH�8� V7��Eo��7<�w��Mǟҁ�qM���#�x!��q�?"j��p����GN\Gϒ�+�k!z�����ea�e�+��U+�!bV-�%xj��pF�ͧ��>�'4^�J�~?`��+s��d�Î�|۔wA�l���F�O;!_%9��^z��}��y7>X��E-�L����ۼ�`=��r]/�)7"�=`13��@$���8>�S�kJ�H�3F<m_﫥�K��N�&6�V����1�S�>i�z=%�sΠCi�:�u�Vx��!�ĩX�a��>����r���������H��І��K4޼|<�H��xGr�Nӹ�>�l��kĦ����Y��H>[8FWe�0ҡ��0~��o�#5�-�tj�tꌖ+�->=��	����/h^��)��(��P�/�̉�T�.~aO�/ֈ�o�KX�O �'l��׮��X:fKw�V�'6�C�끪����9|ߑX����W�^��0w:ļt(	)*%�P�{.��i9O �.�6M?:}�Ol�繧���\�-�
a��_�1�\��<n�K1)����eY�."_��|Û@���i�R��Y���wBf�(c�_�E|߯ E5X��ؗ"�˅s�V�+���^�0+%ߋƴH�&��-�@W
��a�M�i�@ߣ���A߻�*���.C���;�+�~�Y������T��f u{:���<�sY�X��E?d�̸8g������)���ʓ9Q�����/��hQT������#�����|Vn�f�Gw����8���c�-�Q���ɽ��M�"sS�;�jU���PFN�`̶�����6���������7!��<�h�T4OǕ����H�R���X}���K�X�Z�}T�m�j�b��s�qY�n���VO�*7�)V
}���:Z���N���W!�;��GP���W&VwYnVf@�#ٿ!�? ���M�q�U���ܧ���](A�߂�^5< e�Ō���n�\�$����:�vɳ�!�.��Y��$�����h�&�x`�a��L���j��3��a��q��G�'b15t�����'�/���.��Lg����On��<|�����eg���ߚ���{/P�:P�v��3��IC�(�H�9�i[������0~���2�v���fM`A��o":4wr���������,�~�Y+ o��0AR�<j�h٤� �<���rq͝xd���nkƎ��/��x���;9�8_��ߛ�0�|F؜p{o�O�49Wh]m�'n�2���"����H�5g�5�mL�I�i��ƏW,�_"�Gͬ�e��ٟ��k��V��(�.�M����r��5��ʤ�F|.-C_8�EI~�)����bZ�_0��UU��k�%F%qL�{����,�,���e'y��_�<Z�R���J��5U��~�UQ=cݱ3���ҳ���֛��E*��t��ixݚB�vò۪}��}�1��|ù��Ͱ�#���{.�%R.��gU�(F��E��0]��,�sY��H�"�2/��S��~�J�~�w�>b�H�u��y�UG��4l�?"N������eBX�+O�3υG�b�|��z_����="��(�é�%2Жemy ����M2s=�$�`8���j��1+����K��
 ��%��ν��߰@�V9��W�e���^/ɳ�g���侐���/ܭ�PS�<�j�K�������8{-T'I��`�&]�c��ˮ��؏�k����y��8*H�HG_	l�yV�W���� E�OX$1$�C���:l����)Vڎ��^��
�CО>�r��d�*���E�O�~p�#i��(�[W_�����*�PR� 2��x��E�����������ځ��&D��#�ﶘ�,h�c4���~�D"�ki�t�^������2��[��'��;G�]Y�S9U�R��Hϙ�-T.�,+ �K��ۙm�٦���3�6�i|O�*,&I�����J�X뗜/�a�R�þ{ ��I��O���B�u=����n�}Mu%m51����P��Vݏ�'�=�Pcs*���$ 0�U��:��#�Ne��&%����@B��xgd�/Nx����\}g����܃��zg/Ԅ�/��j�p�`t��b�"�<WV](]X>śO��)klNR-oe:�C��o��WX���6�4��Y5r�7��נl�4�T�q��'�����%��T�U"nLu��1 +O���Qz�  &x�L����)���_*Y��CD���l\��L����[(�,����uU19s�U̮0$'�$yJ�������cf��Y=����ş3v�u�UAU�#�������,��0�a��ӾWDeb��-YZ����:Hf90����P����߳��k��.����*�h�����+����
������&���4�j���ͽr�"JC.����d#HP2r�u�s�/����������{�1�Xä{Ş�: �4�Z�5�Tҍ3'�(ڸx���,>���^��{W�Y%��<n@���)K魲��U��&	jO(d$17%x���+ъ�m�����3��!� �iM���5�p�6(띩�,X9����o���`ӏ�D�=X�{�E���"��������߯�i3'�{=:é�i�������ǃ��]8Jx���^*R��]��^��&LZԫH����0�/�E���i�Do�ԴoṇK$�Qߺ�rb��m~��I!Y��{��b��z\���hŤ�N�E�Ý~Ġ��U�t��88�&�SI<�mL�3���-�eI���@Z5��c���@ ��|}�ې��ĖB(�1��Pͬ�������"oӵ�e����.�G��M����Ű�c�mO���{g���
�¹����of�&����C��"4)A�*;���֢�=
:�]4�ũ��<O� ��Џ�e��~�W��j�ֈt�p�*^���><t�v��H��ͮ2��$6v~q�A"�*A­R6e��[i�Q�7���ܵ4�׭>|���� �ץ��7�>��VK��E�mb�\~!��e�{-O��*22í�ZJ>-"���f�+�5�}�72���%�T�s�x������M������>�x9޸gZ5(�F~:5�Հ����V[�潇h�ۄ{�[���*XOW��ߖ�������;�i��5�uF�O<��,8�|⧍��5���z?a�i�(H��aRf3*FtܪFt�7d(Ԇi��e�o+)���R+C��j��o3�]���7�r4JÇ?b�rX���hi��D%�o��lV��Pj�3�@)g�6�R[S�+�&�MaK��W���w�ͳlU�rOC.�d�Jd̚it-��4�|=��Rw6�J���81����=���e���Ę�&6FMl�C��-�Yy�h7�%�����!����$�RCT�k�8�Y��&�M�膩��g������OD�UE�꾺fh�����q�C5_��${�m�UF( )�!^��gM"��U�0�m,5�F�A�!Cb��i8k^�C~�ȬT&�5�)�1IYx�	
�o�.ڷ���:�˹Z����n-�ו@��(�< �4T�K1�U�&��U%�o���]}���?��P��8T�hD���-������â��������!���r��hlO��j�����kQ�y����}Y>#�ȯ-�����w5�A>1Lܹ���DM��m2������6ei�k �;I]�½�O_� \��Ez%�m����K�����K��u�*O#5�����'*�,��%+��c�v����g΍�BߞA�E����*������8�{�J�ن���c��Y�8�w�|�J��/����/�����4��Um�DWb�T��<���5���� ݲh[#��9S�# &O�Z��O ��f���ϋ/��ե�[��R����$�ԍ&Q����Ä�l��/�6��y�3Ĭ]�К��l�*��h4�?�E1�k�����ޞő�%%�z�-�:Sr@1��c��L�5�\Kk���cCnX���!^F�B|�K�"���� ^���6�eTI�$ú�*��[�q��5�w���b�y�7�g ���8hlܑ�H?g4At�敠���A��,A�_"�Aь]����W-����Z����ǻ��
8�϶�d�?U��+�:c{�J���[�jt�^%<��4\�1}MT�a�=FH���DPhq.
�j�!w9-�bVq�ɐ�T5ơ�a/�P7^�ę��K�O��y�et�="_��,�����@[�G��
�'�5���dHC�PMbg�ߜ�� �&�<w1�������ȃ@����6��(˚�M�\2���~����X�$��N �܊���k�w*���T��@��Iܻ �=��5ů�!l�:r啳	G\%���Z�����������L���z�1~�����f�m�:�x��1���"RhT�e�YO��B�#��f�+݄�$k�4ԉ�?��i�XT�s`>�����=Cs�ڥ���K�U��kes��A%������z�Mp��%��+?��Դ�ME_.�IY�]��x]��}����$.Q��3naH��nh���"g_s
BDQd	Y�qCv��d���� >�/�=�!1CW�a��\���h�YF��Y����Tp4�����Yk�@a�͍0+�p�2=��J�,m�����K�����H�:�6�,EB��jϮ��^�(4C���);��L%]�I��KZƆ�2J�Y+�M�bh�˚�H�T�r�3�>�h ~��U�w�^Uc���׾�&9���-��$g�ȑA�>���A:�5���8�^?b	��R�Q'��`
ü���T��U��������3ϩ#��������`�����3���ށ,7�R6$��²�[�A���X�$\c��!X�Qm�`�2D�/9�n4鯆��el�+�d�=61�G*���'�5
>8N�����}�dr���O�ʿ�mј ���SJ��+E
>d^zR��JF�'��,�a�Ea%fV)���V,8<�7T�B:��W4T��I���=��
�������
���H�^@`'��Wg���{�5?�&l[�1����K�;~�m��8�x]�8r�����e��>ԛ�$|����њ���H��^�pX�6B�c���JB�7�]�h�m�q����l�K��,�����B�gn�K�+�4Z�t�^k����<���8��f�;`����S~�a�-�����X|LM���Q	�:��v�����!��Zdm��U��-��W>(������?��|0:����i4�Y� Z��� 6]�ﮙҊoN<5lM����>���2��]���~�zbr��Ar����4��wŲ!��L�!U�8 '�-yCXv�`J���`�}���{1_\���|��=�����(
����׃�M��&j$v.�5�r�.��K����%�H .X[��[������R.[�f�+�6B�P����w�rbRW־jW�w���%d,'EZ�K �W3�Q�޽(��t��f�9`��J��;�O-P�b���O���8Pp��&(h�����P%-�6�����?h��.�I9IҎ$��t'7��3�%hwd�j��D ����Y\��t�8׽�4��`ho��HqW���$���p��X�9ΟS&��r����j`R�T?�'��g�k�~;�Y@[�8 �|�D)P:�8O<�{�W�IF�%p~(�z�8dr-��ߏ�� /���@;OH��W��85��9M�����L�,��eahH����1���G�0�I�F)��ɈZmr����xn�'��6�
R�x�:̋aF�à��_��݊hdaJ���X��>Y� � �ԍ���YDo������6�A^������O}&@U��*r��UZc�#�v�!�Q�d<����csE��B&p'7w�$��Ȗ�%�"�H������l�%��Uq���n01q�4
�w\Y����Za�ޭ��&��z�� /���MK�����e���v�Z�G7gIL�^����p^���΢�r�'?̪s9{w�a5'���@�ʀ���a����u� @y|�B���\�~��0�AfìL�![
���!^�e�ÒQj��{LoX�]�E'�%�	��p��/<5���ɣ�_8q�����	�H�3'
���+��ga�.YTm��\���*S�C�F�0�'n����0zR�H�r�\����Z� ���e���9x]-�{_��Wi^���jc��ϛ?�����cd��ݳ݆��~�mĹ���Rx���<1p]uKW�۩��N��W��t��e��<��:����d��ǭ�ʕ���'��4Z��XU��*�x*�i��w��uq��{�@��sٓ���®�{:ax[I�Η�[I_��	�v��u�1^�dC�A���I�"��	�Wu@�
��&�c&�n�;���>`+J�e�[�4P4Ǫ�"c.~M	9X�[ڧo=��(rF&��^P鐦v6��}��?���Zs�!?p���%�j;V�	�2�bf���ǚ��YO�.fP�<N��v}���
�MM��QX��&�ɷe�D�`� j)rG�0'ώ4�ŬF����n�#}{e���^���5�4�]����0�?��)t�	R-i�X�R#S�K_����7;�7���D>iH�%}��
�/Ou��)��k���R0�^ޠ*&���D����=+73G(?�(܏TP^��ϳ�T�6��' �u#�`�n}dtB�D
ýٕ���^"��yF�,���+�ҫR�r��q����gj�K[=�ά�R2V)a�R=���O�t1��c��BJr�-�;��P�K�{B-*������89U[��:�39��-��`@yEw����Q�+�]I�!������L|L�m
G�ܽ[_�wU%c���^N���Q�>-Ϳ�p ��<jS����I@M���9���A���bK��Dee4�a+��y�� Z��{��v�{`�����#t빤V�̔�jA�0Pom��ĉ��Y����rԀ>ʟ��ӊ�d�?*	��TW���ԳA��T��< 8he:�/N���'��
����A��;���ţ�g���0c��j��P��yz�x{�G������=(�.HO��)Sn�>R�1݆D�5*݃��c6|��Y�̵IJ��%�u��|�&�=���b�u�w�u�+����_�a�yI�� �2n�>/�$~xA���,ȗ�a�~_g��jw҂�~��c�N; ��B32N���wPS{5!��;
u����C��yM��ͼ <�j��7�-���~Y��|�U�$�@�y;���=��FbF�\�����#^&�k����ߊVqh�=�x!�qyU�g��uH��v��x>L����M�e!�N�kc �P*U�1"-�g��~�=�5��xN9���O%����6��G�>�W�9iy�V�>k��벃�K�6�4jo*2'����+E�+�Ϋ�b�$�����X��5����>���=��,[��kvO�4n��/�$\tOҸ��㊧'4�{5���=��v6�0�/0}MD����!+)��_1�b{��T+A�R%��r����RVY$�@����1��ܟ�j*֛=�?nN��.\͏���
������=�f�������#1C
є��x�M4��!5��E�ݐc�#�����f�x���<�Ms݂���7�4?�a䕝��F�*(�Fj8W��qZ�
U!ƅ���!����B�vJOK	���vq��#'�S~q��z&p�IN�f�o�$r:�i1F�'mN�b����;Ñ0F��l_�aM(��<�1F��W�ę���PQ�c����v:�������$3�銜���(��.C�\��x�C����9�����s�i9je@o	�=�[VuW�r�%U ��4�w�n=��@���b�h��"ﷄ�9˯C��W��W�.��LT��=0�Ɓ�m]�J_*��A!߷T>�nkL��y���"�_uNC6�����!���"��h1�#�2ŕ��v1�Uk�l��~�1B��Ǜ�\��"k�`;nt�̠�md"�P����cp����c�R+A,u&v�Σ��&V	�1 ��7q�O����)��r:�-�b_��SN�󪬩H�%������ÙE8b�E�2��	�E��U�y���8jHh@�׍[��/n��V����ה1RS�]�<���m�r�dlt�DC7q�a�'�%|�Q�8?z���r�~1�"F/r%�vKԺ���W���
�y��U����s����m =W���+>�3���S��l���q��h�/�p_Lr��$��@}F􃨉��<��m�T�5v�����q���S�������T&[�|����-��0�|7g����F ����2�I���d�6�8K%�'�����Ǩ��Fu�z���>��JI:��Ԏ=JEK���^%��Z��0F�\!��-Xő	}�.&�I�ܠ�/���_P��M�0�T~�����Y!����Öi}�9�
��� �o��>���ڥ�=(�|�t�P@�� ��CQs�VYR6����p��:�r� �vX�,329�-Ϊ�(�O�q]s��C�8Pxb�ӝ�F-$���?���8k�k:�vɊ��f�w@���rhi
��F�Bc��6V�h|��g��;��3.�uC���Y�
�a�l1K��VMqxh��Cm��[[��������D��y���G:��vh9�C��ʂ��z;����p�.��5�LD�	dLw�C��6�?Z��ou2�]	�Z:������%���K���6��9��pSv�X�x���
+]i2�0�+%4�M���0`e9$b��sBu��>Ž���?zB���ĤčK{��5E$}����w�?ѩ��g�k�j
"��ؚ� �����A�nzDkaX�!v_!�[2��6[�84P��t\���6����3�\"������%6]EI����ݥ�[7ȇE�Q{6�Ֆ�<1�P�A~V�l����%���� k���K$߈��_���u�1����李�Np����פ�!]�:O�p(�gW��z��T��U:1]��"�4�nz���]��y޿V#�.:Uh���[P�S�����|�劃A���(Ɏ�Ҽ��f�K���Wz���s��
V����04�C����*Ȥ����K�C"��<�_1�]�9�5O�A��������ɲ7�Cf�a�bB�C��b�P_���68j�>����F�g(.�g?ų�-ܻ��e���2g�/x���mzkrOj@��V
����:���g��8��X�׃��O�����:�҂<w��WN�m�*�".�� -�h14���{�o�|@_yـ(/��O�ݍ�I̲d�5���l:pM�5��wx/A�v7�#�՚�3{ЀѢ}��)GCaN� �5�t��svU1�D��i�ρ����f��.Е�1��W�%�;�S�LgpW�����Ey��Q ��3�p!�2Er$�$j��T$&c�2�FY���D|!WU�~���e�|ޚ�Fh��G�GdB��Ӿw�kv����������2:�
d��(~8 Lj����P.���j�N�%K׮�ާ��$�j�Ǿ����	2~dӐ�7B���a�:��P�2��{���
03��v�$Ϥf�r �1)r���F�9e2U&�^1ci��b�y�5BHƋgaPL��O��U��d�aӢ\oe��ݖ��� ��)����X6��^31;�%F�'(	b����J���U͌b_C¥cx��v��o��K��FKb��'����9�2uE�':��M�v,Dx3x7%�A��RG#��U�إ��;N��W����'��b
\Ҁ��}m�V�p������.�� ��z}J����@�Lr�+�+�L����,8۠��@e�]\t?ޗ�3��-]vT�l�x� ���:��F}J�̾�8炈�ᐋ�G��88]��cM�$�>��̍�x���s�^��	c��dO��M��a�M�4:�x��S��ͬ��6�|�(x<�K%��yч%F�_W�Ԓ#P�b5���<��u���������o��r�) �4L���38�4����i�n�5��?�X�h\�$�I�����<^���뺢�4�L=�2��RD�����[�粵H����蟃�.M��ȍ��׾e-�e�u]�f7�]�"�ޙ�;����oS�|�E��2>e��?&�uhDp��*�A儆����z3����+]�U��:�3 ����}sW��nJ�|�ߖ��,�X�>#�m�!3}lÒ>-'�u�H{�^u!S;Bv��)"�Z�l,Pm�UH��Q����ҿF��yx��e��Fڄh:���P7���m��9~����J���9�e��Zu����-�]�����YlAQ�z"�ʋ�@�]�rm�.�=�B~ա��g͘�?Uض:�L�O]��3E�2��ΟI�6<>�7S�g9�}��SEB��˕�U�uŢ|�J�v����x�=T����݊[�4J���f�$Dш|>�-*:���rVFm,vKh��gJ�ˍ�~u�_����r�02"=�`>�����]��H�"���Jt�E�zo�J��D��-0��Rۭ[�m���|�WL��O�b�f�9Z��0X�$ܪ��;��~A{o���{�u���R�y4�`�|`H:�1۽Ǥ��^��N�Y^����@�
�Kͤ7�KZΆ��peR*=�������=���oB �Z��q�tW�j=��"�4�_R"WSv����� W��4�S6A�wG�t�Z�~ޙbc㥀Zg`�`��_vɼ:&��#�C��}�'K7���<�:y��έ�0*n�2��������O��5 ����sMj>�j���&�	e-�?�9Բ}<��{�L�n��ߝ�U��zDL�pf�Rc��-���H'Uۤ�="7k��d���6��d�v��������M4w�q��W	~�ͯ�͌r:.�o��y�_��1��"�S-b�����4KJ$Gp�!�?+��a�U�ܖ�Ǔ)���9�G�MDabm�#lGe�����!*8:n�~���G��CU7u{����;��~q./����f�N����'ͽ�ֱ���|�yub)*��s�ρ��F����ǵ2#]ݽ�2�'��:�Ur�C�;�v����_�p��y&�t��#h�΄j����d�:�A� 1����hn�.E�A�_&m¨ɖ��n��{~����_]^p��:_I���.�i*
�*��&�f�	����"[S�8p�
�(��3ʷ�5��q�]�]]�?�<��v?y��%,'�1e��h� *�j�ymW��	�g-C��	?��bU&��p��}7k�x拫�3�/
caG����D�%bFŴ%"uIy��ѐ��LI5S�=Q-<���:�ߔ�V�����me{�P�̇�L����&2�U��G
��yU�`�#��-�T�.�3�,o>է�X;�+1�K]�'�5'�S�Il�	,1Y,�����L̻q��6f�? 	�C��I٩�y@mA���_���JFW�9��{�\�w�4�Ѣ�E	p!#h���x}��gN��+1cE�r��5�-\N+���ү���o�͟M��_���j���%���b��,&�f���?�u"Z���a�쯾��{�l���-�Qj�wj�S�
��j�R�;uC����8+��<�f�[�(6��AdJ���remOe�S�s��'%��TI����7���������8��9aN���'5G?�����׆,�4<��b6s����t�3���E+f�ULn
�s�O5��u��K�I��J� V����1!M�0��ә �<Ċ�0P�[��33p��߭��&��(��/����y�	�X�m��$��{ #V��I{��-q=i���О#��B"�S~��MU[�v[C�Ob^l
뱟�#2�J��][ea��l(��Y�нK�;�0N=���i.4����OU	Ck`^�(�<��c��Ej&!�������眫�Ā
e�[K�Tnh���Y�JI��M��{Af�&ǹ^_�cn�5Y�^ȿa��!��K�EE9�r�p-������?.�l0���Xр�����qɊu�Z�ߑ<�K�1f�y�Я�a�'���g����u�wBn��d/G=MɋI4��9;��h�
�E�Bp�����δ���|Ebkm���1�2�%�,h:�pcX�I��.k���t��^Xm�E���nN^��n�+�;P��$7���r<�nǌj^.c�:zm]��ܾTfv�t�|��e�:�#����3�-�o<��yQT#�\��dFg�V��o۴����Dz�:���������������)�N��ؓ�H�U%�<h�\���as��E\��l�q��%:JW�j�5�*��(�v˶�vD�z��j3��a�^<��a��=��ᾘ�A��� cp����{ہ��9���ͅ�M���f��N�c��[�4�(���K����D�Y�s�p�y:3�_���-���BC�m�!��ۅtuaq.����Y2|)K�2V��\G���J��gmR��H��A�A(��+�~��:2����P�6ݦhI�^&�je�g�g:`\ �E�Pٸut!kҷ�g¾M�}0�����aS���qc}��ZM�"<�H�@B5&��f���8������.SEUA+�A�x�;㨝T�4Μ.���PM�!�j���_J[x�k���|R�N����+{ors��� ���x��c*r�xĬi�l�O�F�Ԝu�v��l��H#�ѤВ�B2*���:\}�sut�{/:�U�n��<Ivo�
�n��*��]ƿA2l�51�es���]���b��
�J�a�ǁ1�����8�s���AȎ2$���Q@�Y���9�G�u&�3����.o��FY�ƭױ˘HH��t8�H^BwWn"`���kG�"�I2���,�B��%*�#ƶ���V�je�\�?{ß��O�cz��WA��y�=)�F�Z��@v�`��7���g9���*���+X�wԛ�Z1�]�=�f���.*(�� ���˵��P����Wg�R��g�9�Υ�����eK@R����,Z��qg��������X�A�xӷi��Y����9�p��6�'��h fɂ��ps֏�L���`���5KPS�nYPo(�;��r����Z��$s#�K
����=5"����q��Z�  �� r1�A��=;�V$���
�\����,�h[&��N�LL����#C�.�W���i:Ӎg��A�'�o ����f�)���1��]�ʹ{I�s�O��/إ�#���qK�B�v��Aϫ�Vԭr i�tu�2!��b�6��WW
��0�5p�*��JϫϦ�<��\C��]����:���F�[�^�%�Vt��F����F�������,�tSI).�H`�N��m�,�3:r��*��ȼ�m�`�tu���1鋟��;eQ�C��6��Q����Aۮ�%��g6|�٣�A��2����G��ZJB�}�Z��PH��<V�ޏz�,��\���5�1XXh�V�t���H��[^B�����8v%���h�7�UXYt��v�6^W����q�u�?���q�cW��g�r8�z(:��&��:��cAR��P��H�MK��
@mo�1�Nm�i!�~�V�L��2f݀��Lgx���r�,�c��JDD�jMx���.r�B��Ymd�x7���r��r6�e����윞���%=�M����_�:�\yҒ=�@�����Z{ub�8e�+[��rkY�"�`ewe���x�d�&��E(��u�|w��5��ɌFv���j��Wc�K:	��l��/KC&�V/�s�E^R�0�� }��h����� }��_�U�� k��"H.��\����e'ܭ�?qR$���s��ڬ�/��Ĳ�߆�_ߌ,��ٺ1{���E���3�p����H<|��{ll��>QzM�9�/Yx�b7N"����d�w�Щ­d�r	B���M�kޠ�5�w�(�1斮�B�뚔���T��(�z���[��! ,cLADd��;���K��1Dq�>YH;"x_t�L �z_[��zRЪ�I~�Nj ���b�z����S���K�X���_�/��i$ck�,Q�P�yk�q�¬�w�BTWW]�_�fq��ES p?�v��Q��=������[�}��t�st�)��eD��8R�\�|�L�3y�]��#-Ӽjr�B�k���j@ܲ���m J�z��Q�vW+��X~�Q��P����.VY��*[E~&�"Q9k"v`'O#��P�$u]U!w��C��E����4{�m��= G�VN`��I[���	��������1"�$(4C�Z��s`��X��\o����0L�
-3��JU����pQDF8��d_e �ʮr��|9"+«$����aN�#��_b���X<~t\�{>�Q3��{��)!�m)H�֖D2ns��7$��K��)���]����DP�E�J���Ҫ����8��t���sV��7"nu,�J�G����Ω^�\����A�n���������̣��-ى��4p�� �9�$3t�{���JD�&,3�!}W�|sdY; ���+�]6�,�J`tVQ(A�!5��7y1ܩ�U�z{,ؿP¹BB6	*;WYtz��Q�U5�o�%;��-�M��s�=�2�vG��� qY_Z7����95p�1�krp}����{��' DE��]�S%���R�!����Lq���r��k�XE�����_�?x��RG+��!D�f7�#u� r�ό>�m�5�şvP=�7��أ}��{����3��q"�i�qg�̼\~Ǿ�ۀ���v��(�m`s��\FI��*Ԗ���TԸB'���.�Y�*V��q�9q5�Q9a)���O�j�)L���t�s�9b�u���u(Y����0����Ve0^���!>,&����ϕ�P����2w�?4�3T��~���98�X�a�C]'�ꂅ:
r�w^󶷊}�/�T�x���y��L/x}�uކI	�F�Ú)���J��^cxS�����=�(��9��z���Ӊ./��o�8�C��]B����;�a��ʵ����OM%��"�BMq(zǑ٢��ѠC.�ϱ�������𙚎=��`���{�Ͷ]�g4)�����h���E�	��½X����!X�e���e_:��?,��w3S�J#�\1���_.�b-
b��Ra�.��4��M��J�#��W#�H"Թ�C��VK�B�X�"�l�٣�BG�9�0����V�(i��:K���m��Xv�~��5��{�[�9OKr���?�R�ٵ���-Fp��ǱSQ4C�>��>/��-@��,��J�)~�B����@�z)[;��IL骼aΗ��/*[�Q�aGS���t1�!�G~g�4X���2A�i/IЃ�}j��)Q�/C�l���W���Rnz�4��i�[�BԸ��J�fhhڽt��
g�U��UFՌ,�4����'�+�0�{�d�� C^9)���ϔ^�i�&b���-�x�1o�"_k�0,�;i�1����݉e>���?�I*2���*�����.AFpS�y!�?�H�@/�2�;��LҪC�|�p�d*|6],g�܂m�"���n`h������!�鈽�ǺN�;�M�|����čy��g�fB=!n�
�Uؘ��op�L�� [Z�w�\~qL]eׂT��(�\}��Hf�{B@�����Wh�����Kupw�n��u�\��+�1 Kƹ�&j�/HCE�[�.��]����{�<��E{���[�]�a	� �DL���<(/�����Z�V|� �:�s�7���[��Xƃ�^�Q�\�5�n����bM��j�3���+kC�=����W�����f��XC��u�Z�@o�Ӣl!2VF�}e�:�dw6��0������sݓY��z�dE�Z��*��er!w��7��]�B�A������4�׈�S����dq�T�
��4F�;>��L��w?�3ka�u�}�AIp�U��@����W_�|��!!���3(9�Z^��ũ�K?����]�/�aG����FiM�_\��#@�aYܝ�~�	��Zmk�l���Y��q�sP	����n��f]5�
�����L��}�AK`]D�J}J�d�f��KfQ#�^�Kt	����o����o\�^6�@�<����	ј)�[�W��֎/�ג�;<�����b��nC> O����H��ٷ����,6�n�>���Ŭ�����\��u��5Sq$%���p�b�@O�7� {(��,�6BV��EoX
E�i�$0��"W�N��;*����@�8�{�=E������U�`a'>���b���7����ѡH��4oZ�
`�"�O�e��� ��LG»�:d�Lͭ g��B�x��x-�c��No�N�H��=��o������ �S�r�2Bۢ�N+Γ#�Sqc�6������ubХ�ϻO�t��oub�s9���ů����#�P������M!����z�Ӡ�3v~S嵶A�{��!�^<�#��y�$z��V��*S�y�X�G̚v�uP<ūy�nwJ�I[��`��v4��G���9AY�3\��se�.6���(0��E.�࿣�,1�鋉޷�C�bl^'K
��s��� �1�A�@B�c�v�Ӈ䌞Н��pB�g�Uv��P+���pU9�G�_�ip��Ø���?��|��d�.����K����,��ѹ�����zYa�b��C ,�$]�>/�KH��g�������O��m�/k�V3ڸ������U���o�H��|ϥ[U���Q�Z��Ŭ�Ѣ������	=w�ځ�e` ��
���CfzD��/pV5Z)v:��.�K����hf��n�?K��t��i�h�J�7(	��"-����y��ы������M����!C��i,�����PA�a�6�0�C�R ��'Ⴧ��E����=rS�2�GM�����7?M>B�U�/�h�����,�(�>8�&ˍH�S�kR��V�A�NX�L�}�t�3Y���G�y�S������g��	#�l��7ç���m�#N ����8�ɺô��S�E,-QI�-?J3�걦��2@?�d��} ��B�:�d?�<�4��$�5���.o�d��F�Z�ᬻ 2e@�<0����aN��{�����xJ�����9�k�%.�i$A��J*�z�W�*l�
h'm�q:[b4�_��H�\曥)?���A�}���fQ��نe"�F��SʯS C��ߞ�?�FMb����|�B�K�Ks�6b�xH�"D۳�w��`[z��7)Uw����	*�ơ�a�vR�E>q��`��`�]K�q1_��J���K�E���́����/@`l�G��ڹb�dF>W��h�b�DN鲺2����w��=����'��.fU�	�
G�Mi�x��PE��h"L_Xטb�M�lS�u3`]��ˋQ'b
x��oZ?#Da�:Nx��s��rcIw%�:G}�RȖ��cE�5Rw�����[N]D�����F[�����Ff@��<����{d�6~w?]�����Ǿj�O�Ͼٺ���8?_��j`��^�;�����������`�E��}�n����~2�6X-?؛��77аt,����{7��h<�E�|��2*3�Xc#,�ћ���V��y�k&�q$��^�(����Cq'�¯�b��� �ݼ��x��(QO!��Ex.C�ͱ�U�y��/5D�<�i��i_=��B�; �٠I��u,څh���
��"D�?��c�\����=p7)68-�����0����I��
��r����ڧ�ժ�	�Ҫ:� ����ȫa�#� !�;g�r�_$	9�"N��B�S�^և!���-]fN�5�6�.U~郜O�8-VԪCt���(S�K�Li[?����fPv>�Z+)>Z.X(�����?K��BXFh{�&�ɑ�:!f��T!�KR�䳳��7W�	������8�=-�)�a.O���DTA�V"��z!�?�s���D�#����.�qh���_h P��=��3�+W��Ay��,aDU���,��郞'����3�'�ђ�d��6(����vD��z��ʭe���^E<11�Tb�~�� Y,�9�a��.`̓O������]�C>5q���@_.}m�l���R�p���R`�]�f,�69���̀�\��ӤT��,N��~����ڢYf������\19`+�I����%kv� ۿ{��j�S����W|���6�!��{d���g��;������&�= ��oѲ[p�?�+$%<n�P6;�H*���jK3E�Ā�G�Y��N�N<�Bb�8���G�uX9�s8��H��ф�uI�YW��&uN=^;�g��=^�.u_���6���"G=q/f�y�Q�a���"ˉ�C8E�z*��B�����3��S��]�p����Y2�S�;y�O��E�����6<�+�R�"\뽾��݅��2�[��,�c^��'r)��a&txH������reY��3�l�,�条v#�.Z�2c�;�4�@�;	&>b<]���d��Uu� uԿ�]+��L����=��x(=��NyNQ�=�E|w��8+r\u|�d�y;��>U2ej�����'{�8ږ.�پ0#��.��*5��u{�ѺL&�@YWe��gZ�G����ܘ�0����h��G�=�D��PE!��AG�C��s5�FS�ݑ�`�l
Q/d5���Bv��lW��r	q[��,���xr�pgs��&�dEex��{�OG(h�T�J��I����S�^u���<�\��%�	���Eq�/�AP�����s3VYZ���T��%�����@,�q����P�MI	�+A;oNmWy���������_��ɷ����V;�g2E�VTR����6�����	�I�����$]���JR�?�,�lΪC��XK	��7�I�WzJ(zЛ2[�x������M�*ɞt�ڴa���	?����J�ܩ���+�� �B�儳0���{*��X�7�}�B�U&��Si����?�i�J�D$�XR�q#�Zx�
�HL��Oݓ�RE7������
�KX`#�Ծ��}��"�p$��&�:�M`rǽo���f���2@�{�L�^���'�ӰyL�[�����g�Z����2rքcx�тX�Ds�W#�q��,�� Z����/��o(��@��#ph���:6��2�猁��0�0KWϦ4)�khc�!��R|(��0xg��N�@9����ua�a6#
S��p������'���hX�BM�%���-=Xz��));�.�Yz�v���u̬h�ݐ�{^���/ �a\M��2t�R��t�iuR�MZ�C)��$�Y��xr?VjܰLş'3�F���)	�p���
���)�(�U�R�2hbB��9�����zh�u�B�^ z4���A��⫢/��b|i��:�}ɫ�n��c:Z*X#��� p.E�oy��]m��������C���z^��C�%�4�j����
�o�S��������n߁U1���࿤ķ�:��!Fi��_�h��P �3W ����+�s��vuDpY^�8΋��wyA�ǧ��@1aP_�>J��+�V����}ZԎ��,�k��5�H}�$��ð� �~��V�G��p���e=h�\/0�g�a�{�L������GR5���l��8�	J!Q�#\yM����|[WC>����3&�;v��6�>'m�d/#�y=cX g�J�5�nl����$�D�>g'h��Q:�?&���#Sj�٢�69�9YDF�-�Mf,3.� !E%}�4�[)�*�:(���U�Z,��8d������25�4D/�mb3d]-`��R�(�CME���M��˨߱�����'�l�@D��WՓ�B��p٬��F���ܕ�*���d�H�wӗ�Օ7AgZ�~���u��ע���X�d��y�pOnc/�3��w�g&yԮ��F$�Anj�i�o��i@:�gh��8�)$���b>����/]�!<��m`[���ĘC��A�j�����'���)J�ޯv�Xv��X�i@Y��/��V"��:�lk�q4�M�"4���8Cw�4Z9�̺_BHg��d��{���G�Z@��-��44�ti������-�)
/
������׼���1�GO+1b�-옛,g�6e�p2TP|$HpX5�%z��۝�Xy=Ni�u���X�)�Ǒ�|,�N���^e�qi�8vޒ�9��V��E���'��>m�奠�(�����eQ�[�S^�,��<���r�*�=O�0@��M5pĭ��2�1,�ņ�R��
-|�N�Z2��wl��e��l*tȦǠ?��e)��o��;5Dm!=O����f��K+��Sk����?0�� �qh/�ٵŖ#��G�>����-`��[���Vc5�p����.ˎ`MF�#�ь��*�Ӌ�Ic�����.��!K�蛙g|���=�n-��C�l���5��"�7u\��Zk�Rq20an͔��<E�� �zD��ϛ�N�q%��y��t�������0�B^c���4=� 8SP�����(��VGǒa��F�`&;48rõ��\|f(	
m�=US��-��=��wA�H�d����R~�K�^W�ysa�tR�,B̲{0\'�[KW-��D�A }�d�D�X*��;8�������FJ��Y:����JL��j;
7ř��+h��x�:94F��v'�K^���w�!�tiX�c@���r^��r?��0�\@*
QFd��\HG���cE1�M48;�Z�nͭS�8�����x�1>��7�V��J�8���t b���3Zx��}��Hx������7�x��ӯl��K~����e^�Lf��&�m�,U<�����?�@��m.1��d
l$}�+_���o�Ji�
ӵ/�?C^[�\��TiPL���KE�,�Ƿ0�����/��GdnEXz�lm+C��]�g�5=Dr��G_��<���Z�gB���Ps�I��6����=<�Cxh ��Tk')��Mل �'F��m�I�,ߌ^��Z��c�^��(��!s�-��3���B5�V�^�^`�T��%�1��~}�9�{�wr&ԫ�`�࢖���`�?[����f
p 1�Z*I�=���[��.z�b�B\B�0��ր�B��h�����
0v�ƭ���d�}��;ម����l��.3裁0�_� Z��HQ�\ٸ���
4��t!��u��%N�^m��S�e�?[/��lG�h��/J]�l�!A"���,#C+�v�z|B���1��m�A�~�f>Ϛ$Kdo��vd��i��r�NZu"�
6�b��,�W-0�V��8$�y0Wxq�D�*��#,[G[Ɇ�9���-Q�a�P˿�UW��<\�<t^�o\�U)�>;$��sF�/��\�L����_� �V�0}6ZH��P�-���U9d�&$0C�@���,������K*Kx~"=N��I��.�g���=���^���l+��P?��@hYC�B%L?�b�}�}
(e��A��q�S��u7�mbT��h��ӯ��^&�~/�K��_M�*16U�KI`8����x��@:�o�nL�5�v�g~'�sܸ��ǎN�e������1�ҁo"��ǧH9�9�}N�wV��i���U��xr���G�j�X��J�L�v��U�N��,F`��F�B{��L�N!kh�)t�Ϸ�hH��=�+M��~�a���9����R$@?��]�:�ɷ�s����f������qa����Jߢ�Xcr�LPvG2����	ʴ��h��J�	\�9���x��� �����F���W�J+�#$o�����-w���۠O�?(h>���6w�6(U�l�ܚp���:e�^$���:�j���^|�)���!�?��:l��E<x�#��'�}��n�)�LY�b���xm:2u!����6Mbm������w����>����"|0֡�f�G�͂z�w�z�q�6&�	Ot��/N�������P�Jw��ˇ(��E.�8�C������/��t����}dc*ir�6�O1@Ev���0t�`/
8$�>@^ѹe ��|f�jd�v��R�!��Bf�3}N���q:'5�/��x	S�-��I
�8jM�OqLDl�o<ϔD1+��b96��y�!���I�'cgQ��"{n���t������\YX<Lu��oo}����9��E�vum�G�"���s��`�Z�Ժ�� {�]|`�O�B������ ���9�ڕ���w�G�\ope`(��
CXh�7��&�o2�d�����ox�ڛT>�dǐ"�am�:��#k�4���͢qu�_�
������L;�K����HNu0�^�����W�*�2ldL]�j�"���̽2�+{,���+r�4]�//���G����A�^�(Ob�����єO��ӟ�D-j.�ۡ;)3��p^��&c>S9�g���c�����oc��=��Atvj��r�r�j6v��޿�}��3+�<tr�~"�j1���=Ty��^�_�	��2f�9EGa�k��Y<�􎮨9A�����(P�{�ոѧ6�^�F.���{��8٥S��,�HK'{��������I��#�t�[����\UMX~�&�ꂨz�*gK`i�#���C�����oOupߜ]�F*�`pk������tU��^f��W���m8 ��<�S<��G���a�au�#����������w�sί�֤��T���ۊ�V����oP�s�]��`��E��L�o��xJ�{h�:���w"�2	v�i̮$���2%�"^��$�����¦�	6���0a�B�a�v�0�9���`f��#&d�'��0P���A��.e�K�(R-�Q�2 %�n`��+;��������Q5x��� =	iC&��\�ȗ5����q@;܇w#<3*���옍�x�=J�0(}9�Z|H�0�H�I�E�	
p�Xj1l�N�x���	0�����"c|��8��E��|1���u�2O����.��(k��:8����T��k�@�AzԚ)�� i�� �TJr,��~I���T�P"HQ��v�Ó������:H�����|�ih*�O*�iEq]����/�Y���nIzԯ@���,�P��gI�\�S�^Zעӊ���* F:T|y a��fL,C��wF�vK�z����QM>p��X��c�v���h'm�B�����g|z���'��������꿘�%�g���bo�@Gja&2�T�#ksP�"��@V�m�,4P�\X��=�.3	��:�-�]g����]����_j���z�bB�T��� �)Y��}����լ��Z�xދ����oU⚣���qz�	Si;x�yL�����7)ܾ�k��c��#Q��|b�%�um�.N�{�5�p6V�� &����lo��(+��X=��e?>U�%|�M�
S50���`�xY�X�]���#I�V�^�����>[����°����������-�Y2ʅjx ��m�pMoX'�/!7�C�WTC)Ի^)��9Rɡ%j�n�R������[:�/�H��x�Wp���5L���B���i�Y��&~}����3&>��~���|���y����sR��0ۼ�+�ܨ&Ȍ:B+Y�ꆃ�5��lUB��Fu��=�v��׬�h��,��L�$|�2�i2��F�T��Ί�f��Q��'$?�l�^�1Z�_|�Yi�0e�������ns�ԑn���A$��h�Ҍ�y�à'�����B�G���-J=$�v�	_|e���	��9p��7�f��(Y/i������9n͸/Kor|�}�)����5��ß#r�aZ�%'�c�Ap�}�8SO=#R��m����W�i�k�ó�����K�o=8kl�[�zK 2�������v[��bIɤ6�]�"��]O{�^��L��R��SH��wz)7
�v�ۤk�Q�&D+M����KSO2|����I@��I5Ͷm-�-L2��'�<=aSQY�G���QXҵb�#9^�;�������򴨕��!�z�'�v5�ۍ��k��������YL�	<���3�hD�_��Z�"ٚ�"_�)�4�5 �(SG���C��7\Ǌ�!A�ۧ=!�����{��qL��ÿ��� �x�*����?�/�9�C�FCa�� ���~a���j�[�81��ڎ^uv�6q��5<���Fh^�2-�[�2C�[fn� ��2ˡ�gټ_�4+ء��M!�~o|�%�(���glN�j[*uV�R��ϥ�+��Y\Fͺ�!��]�o������ѐ2�"��x䧰�� ><L�"s���I��93r�P�L�}m߉mr��w�{x�ו.�(����Hu��fh����6��2𪶪��f��h������|MN��{����H�ͷRoyQ�6�X)%��W�lS����eZ(��K��Y>�C*����H/��8ϭ��)��@�X �5�8xa_��JR��y�|?��4`ڑ�l���	��9�v����9Z��j��$��,4M�� ^{������Cn<J�KeaK��]�����.(��
=���ڪM�b3�����r���3+��ot�u~	���t;p�܏L���V�"����`q&X<��5
�7xkYN�=��������++�%G)_8)�]i��1���̠Ć�����#�J��d������&k����!�9v� f�� ��chRP�q�[�a��0���#��O�x?�G8�������G�jk$PVF?�ݤP��ZfX��t���Z�8IK�̤�N[��xc��P�r_�C�<��z��.�1�E�ysc��;Sv�{�p9���,�bQru���h� B�1?o�Գ�O��
MY�3�@��+X����j�5n��j�&����j5jC�ȫB@q��P�I��_���'$�	uC�{���R����Wc_\�n�·��e�{*�l��>d�._y����_�搾-���M|�A6�)+���:�e�Z(n��ewKp���1e�ê-�O�\[!��(Z�h P���20 
�� v1�ߠiz�f/��v�֤���ԓl��nE*����"�"Vk<k�*� ����Y-����7Ø���p�>��-A�������(����v�"/D*}��!,�D�e��C����T�Z0��>��^
M&���У� 4���z���`�'䯼7#;��&�14�A�b�aVpj�`9�4�=��|��s��얪9��!��m��}���r� o%}5��XS��&�p�y�[,K��"G���3��7�b>T�a�y�o���ҳ�̂�Q�5�������#���.�4�љ�$Uy6d� u��2l�c��'�,*$]t��r���g���X9�� �w�:��,��3,����s�c"#��!�ZP)`�~6o��f��q)j��D�f������f��u0��>� ;-8��7��MSp��k1��C�4��{8l���PYb�ʃ�Y���������Ê���)h���1�T=���v2�K1���P*Z�ۅ��'hvڤ�x
]�ӿ�l�:��T�n�*�mK���ܓE���_�d��jYS&�U}W��x���00��^�dղ��]���M�D7�o��R����}����|"B�p�*YB$E�w JQ��W.�@�o�U�u��S�P/�%6��"U�3	�>�dT$�h�����������>U&ٮB��)㜿�.ߑ�}�{���j&�Q����gC$�>6��iѪ,r5���c�R����<	8ܞMFp�Vb_�'��찎ġDꓤj
�ȁs�
C�q�B��G:�c����թB�]I��9;x��.���D�n�c<�U�2��ˤg'�~@⺾��U�\c��`a�VX?��-~)��#�^Ώ��>���Ŀ��)����ϬhI��]�!�_����gR��]ָ�]��(K��jYW#�-x����
�g۵y�h��K�r|����vX��آ�vY�$����_Z\M��������aFڊu�Ja���?=2'�EN2���<���'q�@�?��Z*bZBQ=�����	�Y�{'�8΁�����Q���TdHXY��iY�c� SJ���G�,S�y}-����g�t�a��x�g�O�At�'JD�r��ۺ��4�5 �M���8��[�/+���/N����y"���T�	|H�����)���F�G�u���L��c�vF���:��>��iׯ>W��V�~=3�ϩ���-�����O�T��� B톷;�����$���`W�Wp
C�YD ��i���2H3M|��q�:�|�v3�&��9MR����ǆC���j6yE̕'���!x���<�<ŭv3x�@&��?����Le��ѐߘ�"��X�J����^ɰxJ�@_-�(]�������I_ n~/'j��s�z����O8����p`6�L�1���(9�4�����) >��y|��5�;�_��U��\�����XZ9�DR.������73-d�Q��a�.�ܬ �_�*<atTɝ��0E��)��a�o����H��BK���w�m�)�P�"�q����Y�U�Β���"���n�]g�)�/U����4P(p��G�MYU;��(s�$��< M�ov?�ڙ����%1bl.��ĞM��b]�������4|���[�7�X���Ġd n�fm���Ȧ�\� }9��E\)j:�E�VV杤=@3��������g:��$��u&b��v�>�6�	�s��cӶ���@c�P�m�"z�7�!���${޵wb��jS��^(��Df��r�%mȠ�DLW�┄����<�V�-՚��b���h�=F!��W�Q���&�k��]��?�t\W�gC_����&���u,��.Ex�Y�Ђ��$�ή��wZ��o)U�!B�ݢ�,�9�;���+�gg���;���p��r��;7���BO������l@`y��s5Mm�� =�RWߚq��FK���j��U�vՌ�Z�ۦC�ɂ-iq���!u�� �z/ ����5�,��|d���/����r�w5��w��b-�N�{9��U �l���߅7�W�ә��RV���EEfۉ���U�5E#织��������7���x�n �\�L?�)jn�Џ!�ؖ��(�h!�\-n�gE����4����.q�OA� ���e�L��.\w��^Y����M�P�� t��e:���o{X*�_b�b`�;�8mÔ���z��bK�����=��#����
J��L���$�9%��^N[����ۥ����򅎢|o䪡1�_�=h����ﳮ��;?G^0��H;��XI\�ۻC� �%�����"ii��T�їQ���]G�{����6Ŧ��@NRn�,FxL���o�$�Lk�z�4�c��&�um�DuQ��m"8S=��"���$���|ꈪ��7Q7*������ѵ}�D|��
��`!W�p���ԻwX�,�k��rnf���ǳ5�Q<Â�����s��,�Q`��Ex]������Y��B�̊?�y����(�R��c�`h�����|� �_�Mz��Ye*9�e�G� ��'�//u�c�`�����I��7�_�R�6�?�a�U�z�5�VRJ��^��3�KH�he7G+������	9�~�	@%���xY+-��B�q��懕Z�;��crD�����a����e#e�� �xq� z��_	���[#�����p�x܍����晈�?.�YX���a��bnJ�������i�o��E+��)��\��à9��n\�r�)��v@(��|��v���.O�Ԍ�0�1%�7.z����n�
TO�,>-k��F���4�x�F-e/)9����QcB3�ڔ���O�b� �늅"WVB�y
Un����B'�˙0G�w}ۣZ���o���. �i����:ل���+k�#4����)�0썏�p b�K�|$� z�z_�g@�q\C� &��r�劮繘PnO��t�>�����>"ŲwΡB�s�6#i~2����$���B�r�k� #�˥������F\�T��GC=oR/.��#�U؛F�L�UN�ck�1haX,I�}7J�5r?Ų�*�C�T<��v���q\���C��؊o�^o�Vl5O��Iy� �F���p.�FOL&�Q���U�/(�A1�u��/Z����f-��BV�f� s���I	�-A�r��p�����>���I=��>De�
�\�2�z�� �W��6�Z���%m����D���b�]�%��F@�M��)���$�l��`DveX����v�c�����͝�s�i���9��v���+!�OCy�uA��[������"\F|�gp��G�dh"��P�wzؾK�N<��������
�sD9�reQt�����K��l�/�>z�Q����aZY�	"�K����[/c�H�H✼-� �s&��Kş�
n��@T8@�n������[�v<��y�ο;5�0}�g��V�+	�R\�ݑO�^Y���Ύ"�4�L�t����qN�:/���Rv���G3i�0HZ��ȉ�5ttߢ�Ҧ3�WAi�����W8m�� �J��%�F*+�@�;Z	�P�O8앏r\yr@��6�ih5���Wh�OG�x���Kq���h�B�g��~�Ոdߤ����#�/�ŀ0����,3��� ��I!�}�|����̵�
���R���^6�5VȰ���K<N> �>(�
�7�21i0�8�^U�O1��j�ۙ�,�x:�ڶ�8j��l��;�ux��6*�HO��X Tx�c	�з��*�����RXy
K�v���;��
�:th��(V�d�WF����w�NF&�Q�E b���Y3$�Cg���۴�캊�^��imNi��x�w��xfLԓ�$Q���'���E�e{���>>ڙD2z��!�jZ3��e��#��N(͡����I/(�9����|}e�j�J���'P�򳟮6�hj�&�\]��%����c�A7���K�Y��UվjjÑq�v�1�;�/9��CwBЗf ��M���J_�f�� &����{t�/���?)C��L��(%�܎��Z�O��w	��
T!���b��d_�T11���@���ea��˛T a2�����Y��B(P�8������n#���YsN
�af`q�	�tҖ?a��Ǹ�@6��x<��3Yi�fee���c�/�Η�����B�1��'�5D���͛%�Ȱt��ܮ���"_���*5�YXP������Av5G487aB��M0*�e2��s�@� -�����u���65(�*{�G�2�_���G�J	����Ɇ��u=�|g�&��7o��/���M4���1�X�U>�g��3�������7L�|��Ro`�'ܯa$�d1�Io���%ɤ�}��P�q5/�)��h|tC~��� ��wc�y��u�/��;~�q.���h�@��t�(�׷R�5���|��B9P@X냜�v=�a�����(�~F>2�9M�Jk(�	,Y�� �W�b|9g��<�p:I'� �]��up/����qҝШ%S�(	���6�=����T﹓+Dk����)Q������X���e�A��̉��n;��N�!M�g���cUH��;���3���3�������:��3��Hj�b:��@/Ke"Fk����"����$�0N:s|���P^��-��[��i�z�e(Z �O" M�I«�FiSkg�zR�GtW��h�k�4}Q�i0�R;3��;�>���u%8��A�l�۠|zv��*�����M�ڪe���}�V4���ϐ�� kڥ.1�+����v�B�lەA`�-����Òl�2��Q��|�8��C? <6WE��˛�hp��G�'0����M*�<��B&(ڈ��6�} �
p��) oL��$@6l"j�J�߸Y�#zw ��fݙ��&�Wj �o0�F۸�MZE%P�`J�t��c�k���P	�hu޲V��	հ�;�Б����ȏ��E��%�n=����h_��
��	Q��nku�σ���H������ߐwxQ ��?`(��+{Ղ���Щ�Uq<w��J������Ja��#r��Q(L�������y3M�_����Gp8�YU	�QR���9ơ/Q۞��&v|Y��D�W�Q����0�dO.��=����_ɛ��6�)٦T�i	��a�O	�
3|�[�L/u�oan �_ŀ���������:X�Z?�n_���7�[ E'aw}Kh���W��!P4�	Ǐ͂Q}�.�w�yͬ{9�,j|ƞwS
����L�ß+u����ʩp!SʨM��P�"����5�e�F�{cC�
l��D�B�I`�īк���TI�UHҕu]�4o�_�ƫ�W��`���1{�<%�&$Jҭtxi� 	g|���^>�K4'���[#�����Ң��F��	����./4����s8�?�,K��g�-{Ik y��y����
���������;��=��5�ͣ�^|��\�39=z�_��sh�w��h��?��os堅AJ�N-��.��^���d�G2���v-�4�%!}���.\��O�枘�||{��a,j>�~�O��_4�����W�[dD�2�P��բ��F������#9	+h�-�3�;�
��!Ir>3����K��߮)�|�|�)kb7Y�b_1I�ÖW��m?JhrH���Vb�Q̌�����iXj����V0�� �ǯ�^��ڰ�e>���R��d�:�<R�N-_����A��r�n�����#�Y̲#����^=�g�`/�hb7���*#�c6���x�[�k�Q�M<�3*}�7��D�&|������mj���$�+%}Bt�-��n�
�%�<�s^���
�ס�NW��ϱ�@�1)
D<w���	yU��?�o�fJ����g;�p?�0jV�� �!�2�	d���`�V	��<|���K�| )Q�>��/�%F�O�H6ῼC�²�U���A��,�9r�Ja��y�CN�V��	 M[���4j�h;�<I���<��B~� �h�4�J�R�x�Մ^ͼ1�2�F��p|� E[iC�s��z�="'��v�������F�SLz*�q����d+�/Aq������&���,�}rݛ��;�������Qyw�9<f˗r�_����Aa�,���	=�ZKH3w{��nS�Sy�Dɿ�w~��L�imK檪F&��`�[����y}�=�6&�7L���\J�����Zi9?����<U�y5��j<��as~M�d�|vz�T�"�ݝ�Q�:b��bt!���ɴ��Z�����
��?��H9��G�" �m�8�,h�0��XNm�l���4�����i��[a($�@sՐhu���Ҋ��Y4㷬( M?���5�d���p@ �m}	8S��x��*�I�r3��k�g���)*fat]��������� �c�af(�'@��:(~o��Խ�^���	����Rȥ��Z�۪2i4�5�� pM��q�[��q(���`����y���_��|/�@���U/���Z�l�W�z&�	w�>�e2�|Ȣq"Π�nGYK���A��h{�z�wLR&p%|(f�J.��-�\g2��2����x
���2nbLL����<*累�:D�jo�p7�n�����\�t�����ܼ`�h`폸Y��q�H����PR�������'z�"�?4%&f��j�ۏ�tx�������SEN�_N	7�.�h�9�d�42�>k/ԡW:`��^�%N�I~�#�yO�� ���кj]������x��߫�����:��}���\N�&���U�'3�44��Y�Yby���~��(��jY �v��:n��$�sI^��X��S#}�yB(*�Ń2w����k��B_�O]?R�h�)+��;�aCb��M�R7NR>�r�$�]�q��0]�S��5��g�.Ċ��G�`���lB�H#Zπ�^(%�K Ȍ�����,=p2�_�:���wx���FJ9h��Y
����S�1ݍ� �=-�PJFI�.�8�&A1~��İ��lP*DX<�R����G�!K3I#[5���Z����~��x����l����������cF��v�uQ��)�Ў"Z7zk�q� �z�5���K��cEI0�6�_�<jcIjR�j&�m�q5�*����s-Ï�j���$���9.��0���nB����7�,^ZF4'��GP���! �;��r�`w��ڍ\tT��ϙ�/'���Y��u!5�"Ǒ���Ya,P�XKX�u4m��U�D���vړ�豆h�� f�ʁ�}3�V��Ԧ�K�u�����H��5�c����Q�d:C��zMTI�1�4?pЋ�*��x���0��� ����r�O���5oJvz�}�%	�\Zն>�e
5�j�.3�z�E$a2�Ο^R�2���%�滔1t�V;H�.�f̰�d�����'����B���N�����$�ɻ^��o�},�n*�9�0�\*~?�(5RJ�d7T��;l���Z	K��΍�5�b�0�ht�~Fs$���;����/.�@���J�����6�B��d�%�������xKS_����x7�����ҥB�-� F=��>i7���ބ� ����P*��"��v�0��4��q�PJ���Se~:��{���!^gw�4�8~	�19�0�-H#7e���j��� M���+��Kx��^�Z.�_�K��2��xC�*u����!T�p�G�����h�so����e���8� �c��5k�y�If�, ��A���|>pln��c�R16:h�3g:���'n��h����CU�]x�󢆁�����}�b��j[8oP�nl���b�����zj�W��t![yx�R���x�H���G���iQp7sS8"���i��?���F�?�Q]It��~��d�τ�7�A�đ�ː�:}z�*�X��B�����]I=�-�x:�H�o�@^��(��ҕ3�鏰�RQcO��5Y��Ш�Vf��5�v����z�����(�n�NZM�h��q8�t3�+�z����XE�y��4)]{ш��<��[#g�������C��Z�4%2tJ�� ����W�wp�M�A�b��L���6��G�u�n}:�|�v]b(9� q��o�ֹy-wQ������b~��a��2���e�k�ྔ�9��>nw����DU�2���Zx�1L��E�ЛJ��d'�ݚ��h�9�VU�v����{��M�7�`b��c�E��Om��;Y��R��� ���p�q�^H1�^��q=2P�]W������I�e�zW�I&�>?��#C�! e��h��t� r��e E!E]����*���f��Xܐ��A �q�	Uq�;�{�ӈу;I6;3����P�2������*��8
�r�x��M>�>�Ӹ}�� 5E�a���M�6� ��?#�Tn��q�?�֯��	W%o�/����j�:�C,�ʤm��~i���p�2)�o����l`�A����[7 ��༃�׷xr��4e��_.4.=ID�z�W���/��yb��L�s�����J5���l�<V
�-/�W}Bm�����$��-.żҲR�i=��@����pg�$ߗ�M`�A:s9 �zcµH�0���@k��+��r����4�������s�`oH_V[>sv??� ��!�F)�P���^�Ɵ9�����o��÷W�k�8�c�dTk6�3�����>?�9�G�	,n��HP�� EE�ȟh�3���L����W��A��/����Ƌ��5�n�W��EK��]~�d���W9�.G�y��l4L((���y!��x��CF� ;p��� z�a�m�� �Ѩ]�����b�$��%��l4�I�Y�8�׊���B�xAim����eGu:�a#)�%�]�p0��+s�5v�μ�E-��W%��"����{\�� �e��l*r4m���L�����S�Gꕋ��V-?��{O��@��u!�F�v�|[hS�}����s�m�G4J{Ū����n6aJ뀾��A�80�Vh�E��\�����4�� m'(p{g�[uZ���gA$��K8��8�d.sh��e�����A��&�Ti��"�X�y��"z2~�ϼ%d@#(�ĝ"��Ct&�))m{cܰ&�H���]��7�l�0�E��Ҁ́�q����.%��������q~�5����Pa�P͜c�H��a��G�,�����N���>P�}�N"&̼ٛc9�R/�^J���	9!�����+��r^V�>k�{���w����������K��5GA�o�I���3���o�f�!zF���+�J>���	&B�E��Kmͦz��ls�2�q�)u�F�32���np�P��"\��E*�2Z�*�ˢV߫Ɋ�yޭ{V����rE�n�Y
����O󬊊v���N>j��~y=�u�H��������U�<xRʽ�\by�Fj�c�>�w�����MB��ˑB���ټ)s�Q@��/7�'H:/�Ǐn�����BqOV�s7<D�@��DoPq��ޤ��������C�'�?M�O�#�1 �$�vƎ��0��=��W��+.��ǅ��rC3vf�����Yo�7%c�ґ���-��\c��:ҹ�ǁ�/��0���A]�[m�����=��j�i+�,?�ǡa�fOb��X4�i2a��>g���E5)���kb�v-���̼۔=i��T��q�K7�_v����:�����,O6=�>uޢQ�@��1zM,Ԅ�xqL��dc������K�&��n�­��.ܬ�0T��:�i��S3�fdtڷݫL	�ǈ��Y}�A��4�h|�h
��ܨuMMn��s��#��"�H��AիF�?�*������>ƷU�!�r��I�����܀<�ӿ��{��B�9�]���B�(�|Uv�Ѿ̩�Vな�����7ǰ���ify����D�c��%�ۣ6�m�G���B)����E�I�ܮ��xDV�Y�p�O�m	�!u!���ى ��,ŉڔ���֗·��FrA�>{!�7�1/��s��a~!�#�4�ph$��ll�0��<��Q���I�Q�����i��	s�1�@�y��︿��MJW���Hq;���̫;d6U��zpb[7�N?#�{<��e�鶋���Bx��v�굺�n<�����
җ"�<T�����wR�Č����X��Tu��y'�MkQ����)X�'�^�k�6��㑠�8/��d��)��]M�A�����_Q"�8PȊ�˪��b|�-�U�*�Md�i��_,~R���Q��pd���"o%�涙ꦇ���c[O����K�'�0�t#���ܵ	&l�j�<Z�]�W�sq�`��`�ܳ�C@Ӈ��{�P���9g%��mK�F���4+F-S��C65W����u�X9`b́�CM���ا�Ul(���|ߺSVd�`{�sϤ
o��:��(�&A�xr�/t�lw�|s���\�upbP��faA��*�}�C���X` XU����ըü��gHN�ٗ.�xBݑ-'��I{�Y�Fx���e�4���lm��"��Lz0eLS4�X9z�`����%9՝�T��*������q ��q�/"�0��֔2Q�M��;��V�.�&�ddr��i ��<��s�`Ϫ�x�a]J֪�@�9��n2�(So����X�u?v��Yu�$-�5V�L�姡��9�D���Nl���V�}[P|$A&�77����S��b��Y�{i�a�q������b]	���!N�[���"LT�	��+��q��1��)������9�����`�~;�V$�ֱn��ت f�V��?�^صۅ�BΏ�G֡;0�v3UP�/�3�,�+�ol��r�ch�.�a�î��EX��.NTa���I�tt��+�'1b�	�p;3.9�����qL7v<(�쾴.6�y�Ő�/X7���H���8�Q��sl�Q����N���7Y��O�-~=̭:X�!D�3�m0Q���]����&ۍ-��j��l����Fc-k�Fwn��~�{��:Sc[3Ϯ]�Aӥ�����N��ڥ�m'SN�3F�'z���8fji�Ⱦ҉h�?���N�oQ��]]�l#��C�/���D&~˛1ލ�@�b��� ��4������s?��.�rn���3�����
���*~Uoe1�P��E�Qnj�����Ϲ�o�/Ԣ����8��cu����p�ȡ��K��.�l�Tt���ķ��xh�#x}"�ױc�&y�۟���˖�ݟm��F}�9=}�M�����;����!�Q�=��HVV���F����^�;Ƞj�d�����
5����N��۰������W�!䧾����W�H���O(���vN}cg�B�d����[�Z�&�ע���J�v�i�� �-Sx������8���!�:.��Q���hiϢ����_�:4�����!��a��b�<Qh�+�٣�-�%�9Fˤf��C�	0����W>�.xcAP������Y��6E�B�����K�XW}k���1���[u��P�W�c��Z�]�G-�u~3l�b㾪�I��ց�?�gw��G�������/_a���Y#t�w'!�d3����lR(/zI�ɜǩ���F�>�qK_"�~M�o�ؗ��4�[��s����t.]p
�0��u���=�;4b�\��^y(��k�b�����P�����Uw*B	�T�YEOi�hX$�z <l3ml�iw���<!Ա]�l��tn$�s!��I���I�a9汧 �K@M�+�1^\M�������|����_��U&� �먕R)�2k*+�,�d�;���-�#�>�2ZV��s����MS��d
���E�8�Ez�'���{hʋ썕^K4�b��&�l�#�vZ�Pn��ѕ��Po�uo�<��C���(+���n�Cq!M]������B[������t;xJݽ�Z�7�+Ӝ90�6��Tkz�}1�c0Acj�&�<�֒���}. A��4�@?���!�Z�l�;�Y�']"� 0e���JZ�#�(�/�2'����F�_C�a�an/N�`C���Ju؝�h�T�m�1�5X�1�kl�⑑��IF��_2�; �r�>{�]l�y\n�J�\X£裩�*#�}�y����٫t�?�6/�M �`<8����n�9S��(��ͨ� _� �)����X��7?�󌅋���ym��{��1� #j�9!��m�����]�<케�r7{9E�z����#+��s�p��D-��OzS�S���mf{��L�#U�%�G����+R���#�=z��K�&?�p��$�r�тd���bo{���(i�o�4=��5�D!zH��4s�ᘣ�ĜF�L"q�(ٍ������{���c����o������}0�&���z0�Ű�UCrݣ��vg�M߭E��ʛ�_J'�tkB�*]޴����g���<}���r;d���_�#��@�a�E#�q^5#�}h��]�+Y2�J�(�y��n�e 8_U̒����u���q�%w�Z�e�V6��9�~�K��|�ls�K���
��RiqWݷL`����#xnv�64���;j��j2��^O8IK���|���rn;�$�N\����2bҸ'�lXQn-C���lb�E\�>���V��5�R���%S��v$�;zIwLO�2A��Č��Eߙ@Eˣ�l�,��z|S��ۆ��q&IТ�����a��˚�Ư5N��$&]���;���l�po��Mw�A
�B�b��iA��N��D4�Q<�#a�:����(�ڕ�4������Knl�l����^�V�*�¦*��X�e���h� ^w�*��`�
��ʔM�xl�%�M1eױeA	�S��pq!����9��,�����R��#��A�V!v8��EL�qĲ,`����|�b]4���Ih~�j���_��?V�Q�@nM��P(TԺԓCiX����w���8��0S�e��i`�w����^�#�7���z1蘛���)��9y]�ƫ�� ��+�ח��?�}��.��������������\��l���;~Ld�Y��B{�Y�@$�4��)��>rs��	�UDE9�H2��Zeh����PLH?>�`#�'NS�`�B����b���~�t�X�n��r���eI�A�.�M��u��L���.#q+��A�t�\�D����)�p͐��A�5��yRG�D���N�k��a������o$�5Ӌ�=/�MؓVW�H�W���6Q��%�[@2�}����dg��("
9� i%xY&��;B�u��If� �f��e���lǏ�hCV��Q4�4��*���?-�g��oG�⫭l��I�=�9�a?{(�eZ�.�UHl�]A
e,UX	e��Ծ���:dH�L8g:�(��`��6�?���Es�����e��wTɔ�/��j>�h�1As�e0��
�$t�"�~�����~��a��N_�N��϶�.�W�ԡf�Ƣ�ǻV�|��U�F�ܾi�畕@�G2H|����@6Q�^������5��Y�v#�@Ϭ�NyQaW���E몱VA��?69�>�-�d���G�s�
^�ߥܑ�d���e�O��QY�F�~QS��F�Ջ�Ñ�D�7��S0l�]���l�'+D��1̻��O�#�O�	W,������4Q�NC4 �6��D0��T�U)�qAݳ�+����|4�L�R���gd�a9W%��mc�RH��X��N�s��"MX ���W�����DM�Jb��o*7������_��R�����%��ͫ�����u�������b:�+��Е�j�0�[���;I�ZCZ]i:B��P�^~_�k�'D���e�F��t������z�j�0�:���<��WZn*z;e~6��$�P��?f�����C�i��,��o8�X�x��6���{�/���"�[/���b���4姥�׍p	P.������d� �e���-p.s;5΀�<н���@��z���p�?�r�?�5�z%���x�<��=����oH�>+����[?������V+��o��i)�٤M)��R�,H�Q����U�����i�[m��+i#<��X;�)i8ڸk7N�M�8e���I�^��_m#�X i�% ,W�w��y3.�Rl .gb����40a���g�p野:DGj�u��g=�R���ĻKv�#�֜�H��s�K�.b��i3J}����=���N5a������	Q�
�ɾ���5�B++s��Ђ�l�W��N�ᬀ�v�x~k���^:.�ȶ���5��)�cب9'��&㌻X�������w���\��ņW�F�P�y
�_eA�-�*�#��^&�����,y^ba������33%�-@��U��r����ݞz��:�T�#�� td� C=�D
� ��:l.3WG��Wm��9�� �p0�fM�n�ԡ�7q?�������,Q|�6�����@Kd�f���Ml��2�«��'aGK}�o������SOߌ�5'���^b������}WJ�2��k;�bJ��@�K���
�BC��^i�&��p*��27!�=s�b�ϼ�}�����e*,����`w���J�C����֏�\i�%�u
'����h���r�C�v�H��]|'�Q�9���UR�Ƈ��@�樥�( �]]�����ﱍ ��@�[Hg�t̼z���$c�'�g���h0ؕ�ѥ�Obo,��0�J�xUKHJ���`P[}��i�0������eT��!ե���h����i`J��]/!N4s��N�|�e��[��dcx���8�~͠����;o�H�!]�Q#�8�#@���H�G}F=>��[�On_�X2[N��8k�(��+��^:�z3�V9jLخ����8'>�ŝ[�1�x�G���&sY������}l��g�2����M,�����J�>&(�=�W(�+�i�y���}���V�ȸw�ox��|hz2a��Nx�g�0E$�O�O�I^�W�)��^÷\*u������J@q����<�o�E��5Igz Y?��@���#�:'�X8����8�.�5��8[6�C����j�/p:z?�Q���V7�����)!Ŵ�ѣu;��O.�j+<C�ՍH��>yޛ7��C��zWX�é�?J3�]A�>�ס��&>��hT����y���U_��~���܇I��i9����,�fK�� ����yL�}�;�3�ގ��W��� Hx+>�_G������I���	d��� |��ծO��s�>��B^�njSd���65mz-�N^N��$RŢUy�b)>]����� ["AѪ�f [�X��B�c@D�����l���'�c��P�%����`��yPC���遌B��@��ҿ�S�x�g&��sފڂY�"뾚��D�c���"�:�+���"3sd>�h%jfOA��_��V얊~R�y�g�ҭV��\ж�Q�D���8	wT�_�x>����V����!g�i�*�f4�5��K8K��3o�ֲs=�N�҈>B#ٵ��å��2�#g��%���5�-4;>c�M0�p��B��r�Z�<Cx��I�V9-����p�!�@c͊LsJ�fI��T�7"ᬭq �3t���/�K��Pɢ���H��6��GT�|��$�ܭV���4$$$R;��[�A��= #�4��9�"�.�u��u����Ȍ;ͨ��x��j>C �u�d��I�\ �_�Э;��L��=���
���"*o0�>�o*ޭ�{J�x���ڸ��(�u1��E�0f��+j�%�|Ϫ�hu�Q@Z=w�T\��"��uE%C��J��	�|�`�nfz(I��ag�첒���\��*�_��J�g�T�_���u.>���B}���1�d�8,V
<51($�&LH.q��:9�7�-�O�k3��Z�"V�c��k��|A�d�	���" �ůL!�=]�;�{TP�<�����EcA�`�T ��P��#Ԋc������5��O}�U�0���5)�6�,����A���B�ӃԪ�*eO.�=�5�D/��N?P��t��3��B�
[BA ��a�����=��Zr������J�r��� ����
dv���J�3v��ƻ��Ur�����CK�����u�f�H}ك����RG �]��fbU_}�ᱷ�{>�l�ݯi�U�i�3aY�?�i�C�|��|��OM)�e5r�o�	��S�m7pQ�?q-8mB%���i�fVŬ��N�P���)xs9��7&�d����6����/�O�PS�';�qs����-�M5�9}��h���݂�CPvm���1�����<$��J?Y���a�d;������!�9*��/�g2�S�pǔL�7$	���ph�Y�v�
Ѭ�c�A)qvs�Cѝb�Z��lb����p��{`���_I�ŤS؊�̈���ĳ����4�ݙT�E��Z`�S�S;]���X�C�#$���t��aC���5�?�jް�K��.�,�NӦ/�7'���;j (��������H'���c-�&\Rs=a��|�9���<�FưlǗ�>�R�'LHҨ)Ƌ � D>A}V�>���V�U�b*�v�4oj�lF��V3�o�ժ��XN9���#��2~�2$�(��</g���柆sgv�0;��ӣ��z[���&Ą��X<��E?��UX��;u�d�D��g'�
�k��l(�	��Q{l�g����l[�qe$[�2��?��P�d��R��s�=1Jj�qح"8�4�)oj%����!���fYi���)S�8��<������_�X=�ۄ
��F�Fto�?63 �q��nǚ毓���������2�xi�N'5��+�;�l�D�fN{�!�߼k;� aۚ�`�G�NND�]F���KQ��C�n�^q"��}�� ���CH���bX�af��<�A�4�򏙽!f���f&?���T�SAkLſ��f=��-�h���� �s�X��F��g�l�X�)u'��:_��{�Ў��(���.��
����̧�]�Ԑ�~��,�*�;�!9��%��P��B�įg�E%�hJ՟��RO3/	A���YLԽI=]��g�H8X��������uXn��Qr�`�Q�)�e�;�>Lxi�w�\���lk������b��̕lS�L���^�0��	$@LT`R{�8���ŒB��jɓ���] I#��ދ#���'-}<Vi��t#Bz����9��0���0Aj�L���x�Q���l�KN�ϓ|:#�%���~p���ink_�8f�H�`�8Z��
鎗q�|+j�1K�%R�z��E��[F #�dX��p�!lj�����2&��}觔���1�ִ}H[��6Z���r���\~xa��h4��V����[ڶ� =G���Rԓ�DK7�G����s�Fb�S$[a��a&<1<c����*-� 	t�#I�����&弟T����^�@�b�����\��<����d!]"·��.���s3������!�ggEfE�L���C��\��q=E ������ۡ�/֨�(�̋`_�-�������a����<�c���T_&jgKٽ�:�iO�8��R�i���(��ʍ�g�gg��!�Ex������P��֏�vcG�V�f�_������ ,#�]X{�sΎ�MoNm�^^̼��/͗[S�rg���9�J��M�}�O�A��O~�e�L�ѷ�O�Ұ�6��>v�Q�r�;q�♽#
��E�T/-�����;BoEUo6�]�B�)�#_Z�'���r����Ă	{������Yl�|�;�H�D���&F���@��4}�����x��_\����Z!�H t�F��vG�'o��n��df�b����\-��,���H/��^�s(
hr~���`��ve�Q��!�qq{�����r�\�وY�%^}�ޱٛ�#��R��a���xB�ݾ��r�q�gRx���^X�Mh���X^"�%��̝Df�T�B���Jl2�/�W'4߮\�	z�!��8❇�*@�:�d�4�#M�ޘ1������w%k��"�	k4g�H�;7� ?&w]ˮ�LX�#��J�Su�'����e?�+�B�f�*M�2?�ӟ�*SK�CQW�<G�z�&���p�nc�N��t���ʟ�x$���R���dNJc+�I��nL<���Cxd���:�A��s}��ڮ�W�ٍ.�l�w��t��3N��5ߢ���Xy�v�}�G�k�^���Xc�W�(��F�އ�Z��u�?��?y�މ��P|8k��9G��ߨz���l�bPh�Ỹ�~������)mv�z�z{~� -	�b�kO��3.�9�(~�vy����1�����0Ź�Q�߶�XԵ�n�u���N��C�JЇ��_-�;�̝�͞����Tn1$�L<9�p.�B�g�:_ۦmp>0R"�7�?XW<�����w�m�J�J�뮓����f�8of�ʪ�(b���E%E�qVPQ�jByV�8�3/�u?uZk�d6�}��k�����@jE�ZI���IIHbV\su(3�.�w~6���7k�R�G�<�l�qt\�G�-��v��9�+A� ,�;~����.吧��R*O���)����H�"4V�P*�Y`a��ĥ]�[¼���A`���8���񩧓'Z�{��VF�f�?�BԵN��9EȞ��⚝*FU��m]B'�^��&��ֱ�e��T/~�nٴu78 d?zI���4��S��ZXz=��;簑D.�[��y�O�0Wŋ�y4���2X�_{��� �|��	ϏBј'�/~7kN?*�4�^�s�dgR�ԨD��{�Z	7�[I���o����d9�5���ZCeP?�[M�Hg�A�ngZ��E-(,MRde�?��L���:�u���:v� ������t�c��	ѱ���������=��WL<f���zkYf���qc���1�'�ZSKvE�mH�TK��n����7�^p&�De�s�(�q!�3���k�5��7��
.��Nu�g���X�1��=|Q��2�{����f)
�nK꾸�:8��4B���|ܶ��32?O2�`��2��.88�@� ȗS��K�u�h����I���:L���2'�#?��L@SaY�yf&Q�rr� x�ߟ9��	�R�s@����s�Ш��G�xl�V�$���`�����x]u���#nT�������Ck�\����0��/w� �l�Dsh8CI��!h����Mt��$"�<�ݞL�1���E~�c	�ӹ�0)�Y���ׄa�e�`q�d��)�f���tê�:">��!�C^�I��� z�0ƶ-�#�ɒ��	� P{[�d���<�Ŷ�QK\��V��A�wU���^��)b�]׹e�X�%@�C���s^��-��0$E ��XJ����%�wؑ�[h߉�g�U
@x�KזD�'}��>�
��+A(?]�Q#���e2�꒒�"�*�b&�M��pJ�O�-%2����Y�4�����ہ�D:�1�l=��[/H���*}q��#�_e,f�a_�����\�~Io����N��5E;2�70�c*-�X�-�����'λ'��yۂ��kՑ~Mdk���\�Z��{��s��&Z����F�q��mY4J<�:H6�`�,X=�b8�̜L�B.Y�|���#�|�s��`	��u��z흟��bH�
�R����G��4�T��{��L����)�Xfkv���y6L m<�V��FUȁn�n��I�
T�}��/���.�7��A�������}Js�m����,LI���,��
Xխ��2��P~��f��!���5Lsg�k����'�<��oUe����0(���P�2��Ƹr�W�ů'�����cW���䜈ް�&�]kN[�|���4+�����UD�Ek��S͏X�������$!�o|W�Q��FC����j�}��{,���r��	���노x�lyGBk`���Qݮƣ��yD�n�q�[ᏡD�&4���JrfX�S���so�=���Kݫ���3���� v��7=��noFE#���Ѕ�Fݦ�h��f���}Ź\��Kr@��PНY������ R�S]S�@���m�B����GL`���{�*G�]xX�|��*u�ف�c�$8t[Q*�SL%!��p��m^��R?�ӌ�e�����cS�U���	���W�o�·,{b�]�FJR�7�}1N��Ir����\q��򣹎w��~ȴ��`a} F4��1���S��E�7�B��Z�i�}�������uwsL�E�A)�}z���XZv����{�}�M�C�8/�zh|Y��������4�&���wI���<���f�I��P�_� 9@�w�c0����{��L�D�&�;�=9W����u3�+�F���Dp���J݊D�u��J|w`�UR�(ѸM/�D�Bx����JBa��D����謊܌,ǤS���+�!��.�槨�4V���˽<J�-��;~�;��"r.bG#�C!6�*<y�����ղ�f��Aem�]�R���5�-j�����t�o29�����ָe1�\NʽC��$@���C#�{X� D�ck���:��Qh���b)���A`"Ox���6�δ����p8�ZL���g�Ý��`�;�8�EN��A�sl�i%S�����cf(�s'��=�+**���:�Iˆ������G��S�1ߧ#�����-ۤR�s;U��y4�(52�Q����"-F�!@�џz?�3ԫ��ˠ��w!�l!����M"��6�S��G#K�=�=�"��΂*J���q �<hk0e��n��7{��>���z2�&��O�V���&J�8q�Ȑ϶������,w���i:�%���!y��[�S(ҁm�������Zyu�d��^�5��M���d��p�����ajQ�?~���r!\<w���i���f��)��2[b�[��c��T���i����!4��}`��t1��"�M��C�XQ���N�(�z$��y����n�C��HΣ!x�b�u߆y�yd1��ib���Q��5~2�������a�a{q|ǚg@����E�j_�/��OO�+��Ȉ��Er�?��Js�T�]����.��Q��n��%�l�y3�e�3�C�3���
�w�@ؙ͗j-�[��w�qaȰ��PVD�K���-��&�l����j�DV�K��d��3��((èv��ĕ��NJ���$1!|#����T�����C�geK�Q ��g�8i�)���qR�/��c���M�@�֧�Ȇde))��Ci	hkos]��k˄���t��7f���
��@�:��h[�%���B�Q֠�G��h�I���2h�_�9���E�Fw*���"Q5���=w�*�i3j2ͳ���� �����P����f�� �%����7���3���u)g��ʝ�J���WM%<`��8�����*(4+k���e�6���U�^ ��A�����'"$�Y���Y=��"[ʒY�]�wF�b3��4���E�eI�����C�bQ���C<,<�}lC	!�)��F}r�X~S�G>v���H9p�%N$umF��8"|�X&���
�ϯ����3g��E;�	�c�h*�z�����B�C��;峋Tk�w"�[T.���Sh����JAծBE�[~7�qZ��A#������hs��uU�:��K�\"��V�C�.=W%غ�y��:-�io�ͮ��/����P�0��7��<��qw��	̹����ȉP���~[O\E�	���������6���5�C��ɣG�a�4�ί���Ɍ0�r^-6	� �O���c�M%�_��")K:�k����ǆ_+�����$��e�u�n�����As�Z�m�!�0�߁��m,z���Vn�/�x�Sz �F�֤<	ƽ����y���&���
��_t2~ӊ�z�6Z�]:A�������p�
E���b0��$�fF��"jhV ���U-[�"��t��T)�@ "]
���g��7���r��O/P�Ԏ�M�Q:����tM�.h�p����D��o�z* :�/ ���i�x\�()�$�[77x�;��H�i�_K��I2���f��W�J*>SGɹ�����2�9(K�ќ�\a:�K�_��9�/2'���cds��H`��~�����Dk}��VkJi�0O�?FL�.��?���-����o���d�+b�FR�x����I��/ ���'��F�&�����|�ZOeC$�-1W8����bK�!gVp4���3����Ү��g8��Fav���>��}td}j?��X�l�2P:�C4��W[r`�3��杳<�gT�,�~��.�g��K�2���?��y6Q:ɤ2%d�i�؝'��l �Z ��p2��hI���F��r��`;N)�/~��}#�2��?��R�"ﬖH1��mr"|m�g���G(D�n�	M��r��"�����Z���q� 8U�֣p+{	�Dr�h�2��<���Q�͛#'�3�Q�]�$@Zv�|�Pv�����HQ}����\Ը� �>��h�r���|<�m'�N�g#V��ާt�fxp"���pd��s���Bc��`s%QGM<�t���^���EA/���G���2��('Ob1���܆u+�_���*�0�[��K���ٿ��i�X�U:�^�dzsy�?4;-��n�9�S�:��J�yB+H�\=�V!�9�m��iДͦZŀ\Dr����ץ�f(eꭔ5y�u0�=�[MJB�b��f�nӊ"�㛜�ƻ���_d#5t*:��K���!�a�Xѱ�������U���gZ^{M��á�F�����<@D^�u�ְ�6� �X�;\��{�;���%�צ߮Hv�a�Ò�_՘��ƨ4P*2�R:UUd��%���!��4ܻ���0�{��궨�g3�z��%�f���u��m�ϙE����JO(����^�d�%�������Q�11��,dbӣн��|D�:%����ġWnlN��ԎA���nx�2L}v�z�f.�.����sR�O��m�����b3ņ����<�%S"���;�(?�F���--�u0�{V��xa��p�Y���	U_�{�vQ ���'-��\J8���0��W1��:Q�+$�vc��|G���BI'O-|��k����h��r�#����D� ��~T���&~������P��O��cӯc��U�����s�Z��𘷂����~���V��!�zD%�G�n8I� ��43��a�о��	�\�^����E5<��&��&�D5M�j'�ڌ������z�.w�4��A<{5Id�� �Fi�S_u�n=�)	��(o��\9�����J5�@^#��
@�(�e*N�&_�.�a=C��8�É�}�5�z�p��,�Ny��>1�^�s,o3ɽ��6���b�t$��!� S��o�2l�i�OQ���-��J �q��~�����4��������F�`�c�@s� ��<�r���fH��+��DD��G����xz(M�;�j���ַLe�Đ��"�=�O�/��/F��H4�d?�dn�ǌ�&�z�f���t����ѧA/?�-@��-��N=��/�AOxv69���>��.@�t���m� FF�{x�{=?1�qN�����v�� ���C-���ĀF�P�[,xb��Gۥ�RJǳ���aE�6� re��u6�vsW� ��Gp��A����[O��-�N���B)$i�����]d6̎��R�4ǎ��ܢ��]���Ґ�n���O�����>����X��ʜ��� �M����js]�N�60��(?1)
�32����P�(-<�� ��8���p�*�q!ڄ�̞��]��r�[<efaT�����Z���p���}��UM<�<ı��pp̓�*��&��t2�m�ˑ	�BH�ҤY�4Kn�Uו�_����q�~�N�����e2����nI�1�Wb�j����s�oy�CO��𰗪�d��`O 6�T�^P����G:�����K����2�Ϡ+$��./�[��yz����4$�|`8���T��kT��ح��������0 ��R��e&�G5݆����%;6TA����*���^���[)��Tt}��Fh'G�UxƯ�njz��>c7K2�����$��x��^a1]��Ԕ��>��$^ �'�P�@%�R���)�����ɪ
�7�_���fl#���؏o�7 �c�/+����I�8�\�9|��)Gr)��]�4�R�R�J]���4�F����ޓ���`6"H�$�˃��o4��EQ.���J���RC$c/8�U��0ꥴ�zz�����G��"��r@���A�v.98F�����#�LX:����S$���{�%l���e$/���F�t�Sb�� ��i�ofۭ��B��<r�'%v��M��d��ǿ��1�}B;��虬t��#��r_�0�u+VY_���A=4.�(��)�scF�R���T��T��F�R���x�U�7�<��c{���5���+.�oH�h�d�@b�<���SB��t��5��Su����Q�Yc��e~�;ӏY�P&�0R0�$�i|��Z��~HZO;�\5�l��ni䊥P]���^g���dU�Z�&�)jX:�}��/��Pq
5���W�&P_V�L�o<
�6n�q�q�����F�����+cܷCS���CNV�Y�"wZM/h��?� -q�p�`�P&T��cI�*/1�w�5�:�{'�Lpo�Zr��8aOY�L����\�`;3^��9�,C��ԟ:�qa�<����=���`mg�S�4�XT�HL�00�b�j�ʔC�A?%0d��*���x6���?���)4��������Z���~q���]�ju���ڛlK��O�`�"��G�'�1���W�66�:��v٣��xf��4*ザG"�����3��]It��Zx~J�����r� ��:�b�Ӊ�6~�4��_��z��Lj��*[獏�"iC�WJ����r���3}�����3>��������4h��:k)El�̯�r�58E����[|���m�Zݤ��& �AQ��@;v�	�%D&��Xp�z�Iɨq�����u�+��n�(�e�}O?�2¹}�>^BkFeEڧ��'�2���m'轵�U&ÆYX���^�as�Xt�Ĥ��
A��)����t2%&-��P���o�S�w���w�7���S���,H�����ܥ���1�T�dSC�d	7��5��7TL��҄�,�8M�$(hKc����*^ΫB�@Q�_�__�����-SM'+E{Ao�GP��Õd�+�tV4�e]Wi�xO�hB�x�M���	���q����{�M5z���P��/	,{� ͧwϩ�ɮ@�P�~�O����&MX/���fEI�8�Z'j ��Q�#)�M�݂Q�r��F@].{H�������% ���G��
�=������/$����w�V|ߣ��V���$��r�O	X^�5c'�mP(4�A�{�l��]GTqɾt�W����%!Զ�O��}����}ޯǫ�LN���!"9D�>h%}?���/�	x��� �9��f�L�o�v�5�O���i镁G)���Α��qHg����c��֚�Ni6�"D<p��������+x��/���kP�%^��A|I��Id~ �T�oӑ}�C�9��.z7�AxgHi�s|<��vwG�tP�����l�:�28����ҕ�����5�H�W(�$�b<����V�5�X�+)ix�F��D2rі�e>���,�^ʎ��Rz�-l����Tw��9 �1���H,9���k�r�W�@�`�y�d@F�D�wN����%�����y#Ii0��R�DX��[�4���9P;�ЯA�#� ;��M��@r|R!��xϻ����o+-Rډnۛ�(���b� �#�誼˺�E����8��7��L}��`ݺ(xm�
k��N���`#�%�t����ƊhJ�j�jh�$�>1Q4f�]C@%�^kU���N�qC����H>��e״������|��035�?��]Ǻ���K2�Y1�N�~�滓�=#X��KLm�7<ތ�ݦ���̒	��)o����$H�X�k�r �����tV�R��̓y{\8��G7�I��M�(��'���,p ���ɇnoLO�m,T[�'F3��������ˡ�W8u#��}f�M�b�\2e�U��R���,[a���ݡ8�E�,~wy�-�H��Z3 zaI��2��e[�=18��z���ࡆr7�D3�*�P]!F�F��pO� T��/S��$�wr}g��D���cA�>� |<*֭��|5����9�za��2TZ~��R?����;��W��	�:/�)��;�Mu;_w��;�i]b,f��&_ �bn1^���iM]�Ԇ�[�7��b��ixA��)RE����e�r�����J�$�q�j2;�{fV�n��FH -�+v5�Q*�Dt�������M��{eZ'��ly3/":��u�I�w�O"mb 2_9f�Xǡ�E��c7o֮�LM�����Y���#ͦ��Cm� xb흉�y�<X�,@���,�YDx��a�}ʽ�][��P�Q�sn��3�<V:�kl�i�`���f�/��S1��B�2ٸ��[��%�@;i]d8�GB]ƽ�MR8�0���-	�'>b�^XT�0��ْ���b�@���t9�
<y̆5�����~��7u_w�}O�T�F�WV�#���U���T���:�~8|�B�Ztv���ޥ�\FcZ�4����Os����X�]lc2�$��I�t����au�H��i$8=�xY�PO����
N���07��d�����+1�\��z�ow4�M��&6�GU����(Ȯ����P�w�>�+�)���y�^�Rr{�Ծ���[����J�8k3J�`���'�תǉI�<�~�,kEz�U��?��;�����';��P<�`��C�a8}�_N��g��?'��E0uF05�a˵J�tt(��Lv���3y�z��%;6�_DZ�1JMH��\n�N���U���W�G=#�JK�c�����",R���|pu��\$��x�[i28M�Wx��=3�k7�,����0�o��V�c([��^���6|�����.z�ߤA���C�WR�Y&�~Q�6�w��� F��4�E)�"�m��>���wL0�G-���nu?a[a�U��q�۫ek�*�C��^҃Q�@�]̷��;;WY�f.�PT]P&<dk���7�M{�̝rBd�(���;�_:Z�vK�Dr 4�v�T �x��8��Us^j�0�<T�qíe���	��V~�:��O�I#���vz��i�-8�wje��;���k(�z�%�z����͐�k�q��6��HJ����k�TQqg
�A����R��$2�I:
!�v�#z���'��LG!D�8���2��?3�)�ͷ��1r.�6o��Pm;�j!$�Y���n�ݾ 10�d�A���r��I3p�(��%S�9�2�ؽ��φu�u+x�,�QT��	�萨�Ē���^�u���(��d���g���D�<�Д,�Gv�JX����Hϴp,f�6�;�W@p���
$�(G�j���2�h)�d-$�ʔM��)�Y�tڥ�� ��7cj�s֘�m�5s�ޑ>�������t�(��֯�B7~��L�*�=�v�VWi�0�Ġ�N0U�o��i2�!2�;UB0ŌXWno�� �f�ձ�>��o⵿��� 6{���Y����WM�C"���r ����=�+z�6Ȧ˯d`���N~��r���eI�&9;	�3js�ӝڛ�����VѤi�s���F�����a�!CEz��Tq�s!O�Y$'�}��Š���|7��c}��DzT���i�c�@v�!]­���I��
5h�^M���
�UZ��k�)ڪҾ��*E���Rl�B�4y&�o�Ԁ�t~�\"�i�f>�b �����%gv�8��nŔ�L>�B-|�r�c�#��u0� ?$풝T���D_W��ҋ�Tk�a��
���rk~U}C'�z	�aε�它.�.�u�5 ����ְ(�IG���� ���`>|�����,�0j!�rH�Ӷ��5��p�{.쯏Ͼ�̨�}7�*
�6D4�M������@�U�~�g�"|�g��`6�~����2/��
�'^e��QM�ь��eK#��s՘xת5 �~�\��7�ܧ1�^�c3�F����O������Q*J�f>�� �H�C�#04��q���4�L�+VM쑻vҐ���d'�+��EZ�ELO�	@���.��V1L��M��W���%��{�	VmQ�dP�46i���#()�HM�F<"�����첯��/��d@��(]�,F0�Q)3��OڲG,h?u�ip�p~�DP�_H�W�c� �%כ��=�Rc�|)��C�u��pܽ���)�X���	;tP����l7ݟdz�#*G���f���rY�K��˽.Wy�ל��|]�*����OǦle��v�hA�i�ܥ��$vrS5*�4pj~�He�y5,�W���{�,��u�I�侠I7�e<�����i��j��3��Ex���0��m�/:t�ia�&�bw�fb��ȺP3���K�+k�mYE�\n�,�#d����^w�2����K�W�)4£�Ńs�L� <�������r��0N9�"4O�1��v� �w��)���܋�C��ӄ��۟M�� z���4 ��'\�G'u�sA-����
6qP�d�Dx�����VEh,i7�$8$��z����i���ff��F�s\��LY|���1������ƈ�g�0�Ȇ@J��ț|c�ؒw��S���$d�x�sϘ��r~�ft���͕�N�w.f�m2y��eYN�)	9�a�n�b?�����N4��٥4̳��.j�L�%�*9���ъ�������ӆ�4}2xN&xq`����e ��x(M#�Y)8ݑ��4b�iU7�ę�y<)^�b�ղ�Y��I	�l�k�c?�-�'�8�T�]��{�H!�74/�t�v�BɺR��)j-m4���X��s��ބl��j�� �u�K���&.��N먁D��p�t�7��֨%7~wXX�}��OIt_�;C����)���$���Px`5
A)��� ~����F�����.��U��@��[�SK8�J�</�da��]��B�{`��x�O(��]<������/S�K3�m��#*lqS�6�Ks9n#m/� I&����Z���:���r��b���ض�c��X�1���%[�D.! y(C.�XD]2O�vН�/Ԙ�"Y�%�{:��O`��G	)��ʓx�T;t¬�� �r��}��C�[#q7B�z�u����[��+��{JQ��S�)�p��f;�������xR8ӯƠ�9���
3�+��Ś�b���0���H�%U3-��bH��Nf���A0Y=�B�T;����T�D���)�EPn6���kȹ�7�~Kʄ':~xg��>�4�G�G��z,�9�D]��s���S�V|TH���ݯx�p}�F!�(j��͌���T&�w�h�8�R�W�u+�5�jO�ˠԷ@j_g��y�Z����C���b��6��B�X�]�l�,���)��70|��;1�KA�Gu��?��U%-�`��{6��.��++FK,K��u �P@ϛ�Y�QL�P���	X���?N�������i��=����:�G{���A�˒q�sI�������i@m��x�����N�q�mP1`�����~
+��.����'F��{��T��2��)z.!�[����$lyw����#Eɶ�$�v�����5w�oޅń#<g��^XHy�nq(+��O4�bϵ�tx��
�x-k��H�:�N֑?qf1��3��'.2��S���/.��u�
�*���P��@CK�M�B�p3{'�vZk�E�ڏ�=�J\&m��|:��o�b�������ML*�OBn@��v�nA�i�zx-=k�q"�����F��ޙBwxL���@���k�U��4|q>$�$jpl�!kIw�tyH:�.�LN��]�{|`�9�>��8}�p�\ ;H�RZ����G�d)
��n1��|G�%�K��>'�G�u� ��ڠ��&^
�����8�e�����©.���tv_��:?yl����m擇�S�P�bD'�5�7S�Hn�< K��*\�l����0��.Z����!�����Ǵ��A(q;
:�V���8l�O�v�Y���J���ˮ� g�6��k��>�7�6��JM<l����I�*��������	�+�[e�nܕ��kC+什���F�j}��_u�7�`�S}g��D�m�ܪ�rW�ግ�q�̓�����N��WUwG����_f5`���v�W�x�Qq(��|�c"K�J��Ĵ��a�,��6m��w�t���kJP�&���ŀZH'/��Sbi�]�y�uad~�̆Űae֥�L.�~����B{�"�|/��_�h��>��������"ї0yŅ{�5�<�9����^���{�Uο�Iԯe�n�TyA�1n�-��}U��B�E����#]��$:��!Yz��t�t)W��9����[�K��`���8I�M��	���.����I��꠭[��O݅�[��^7G�SJB��� ԝ�a8�/I(1�Q����<���,��c(�ؚ(٤O����Dg�!�{czHA7����[��6��*�/��b����aVʲ�+ڌ������_�H��T+��h�ci���3 ��aV��6����XO�m�*.�������F���2�}U���-2;$���/i�M���e�e���{�٫y����d}&��z�@Ne)��a������`u��XzIi��@�`�X��7x�<8��Hs�w��k��,$�3�<`��PL����J��$A	����a��U�kڀ���5&,��jT ��toѯ�d4:	�\�d��J���;���EHg�����aĜV��b�ݷC��W��� �W�)��!��T�t�|?.�\�!�.	F��Fa�?n��a%Uu$k1�#�M�G6�o���c��0a��s��*�����i�I_t��O�O}�����TӁR�7ZF#��&��x���;i���3�oF���[D�c����C�q���c�5�d�*����o���W������HF�-]�MW��0�����^�@~0�5t�>�t<�^Ҁ�I]!j�$��~/�%?����b���Ƨ��K����i@G��y�Ź�"b�1���b���/����v@��N����������G΀5B��~�9�a��͂so�R8-���Gqs��3ba��
s���1ko_:U�g�6@Ղt������\gI�Z���I�&u�*������>ћ������g4j;Hd�0ץ4Ol&g��á���u���K�w'厇��ֿ2����o6��hC� ���ح|�,(��7���]|�ԚP��Ex�aF�Ʀ/��u��D�Ap^�%��5�#{Z��h�˜Kĝ>��PM��v	����/�#�1�&�
 ӑٻ���j�����I!��yf��8��F���:!�ܻ�����z��q-�?󳐈�A,�j��D_�>�U�/�p(θR���~I�����p
����o��BB�_M��4pʚ���p{O>\ ul�Y�����ݔ55�p����&�MjA;�*�;m{��b�녫�!Ի��R�~��M��� f�#੽T��+9Р�٢T�Xg2�x|��t�c���[�tŃf���~z�Rh}�,��:��Gs���}X~�l@u�C�$r���FY�&���}U%�
�2����n~&v��a֧�&B1�"m^yK*@h����naZZe��KQ�;:`1�;m�⇻��	��N�G�k��>�Љ"��E������&��y"W�|�>�A�+�<��ˤ���9i��)�4ɽg`�3�mfi/�@�U��-�9���������z���n��1Vw4i^�l�ޚ��6��"�,+%=����iz���bZ#Y*��l�Yk�X�L
eXCx�o�7�܃l��2>�o��ׄ�{�������A��x��v\��3�����ͅbi����`D�oZ\pF-D��kۍ��<rU�z��g���/S-F(��X�+�˫	T�ז�\��1b��cS@�O��*_!ϑ��O�B��c�ώ�RDWnr~��tv[4�cř%,���Ǌ�+������wY=��q2|���G�o(� ����L��y�h+)�J	eS���G��85p\괓��xo
ߑ����f�p��}o�w�v�[8(����he<�K�3J�����-�Kvw��JB��5c,wm���q�g�za�Y3 ��zq��@1v_����dB�9u�Q-��_��[�*{A�fD9��^T�$3�,�ҥ>�����I׵�����0�N�gd����Q?|���v���� Rv�/�Gyhd8~a="��;C�ѕ|b�w���q��Ẑ�Y��)jpl�q�K�>��ȋB���w��]M9�#���?^y�Pp�0��Š�Pa�D�Q�\���^=���@��ؿ���;[��D��<�JZ��ů�r�d(Ll��E�3�r�/��|������Z�N\�@�}�!WKW�gw�<;:#��>fA�ǣ�Ӷ�����,��[f�?��Z�R��*�`�������/�e���V4�(��5h,+lM|�^28h���efˎ�'9wՒT�g�Q�̺�Gh�؎b�r�m��π�~` �J�y�_����J�QW��/	
ZVg��1p��D����UGf�����e/d�g��*7n;]�j��ۡ�.�4%��=�@c�ŀ�8ܬ��u<8�&tn~�L3��~�h��H��C[�T�.h~�����;&��ẽ�,�є7�Ua×�����ȇ�b����3�]P�a|52f�Z0��x���ꅸL�2 ���/�26]�N�{[���Y�4Ι� �)�Ij���)����ǘP��:��%��iQ�r�=�\RÌ%��)�Y��iU��bu'w}`?�R �H;3�{;�(�%Z�^���G%�$e����I��zle^@����[%-���p~�_����+v���
�a�����R����u�m4����,�
sbt�J1_�x�eU]WXQ< @�o�j3�vF#=��t/�Ao����@��/�����?[!+�P�=	�n�*~�fTYt�K���v�&_����ɤ�Ktyu�>�Xx��O E7ʛ�G���a�Ԇ&���اU#^�U�e9I�hN�*aHu�=����H�a�
���x�T�T�/�(%�*�ow�t��F|�Nݜ@pyrA�]�I;�!� % �bD�+�P���o>b�����C���г�Ь�H������Z�a06w˄�YGo���8�,�ZKqSrZ�&En����z�њ�Zu(�\2�X�]�+	�f�Լ� �������b�F�]}�uC���V�Q�?�ۙ�9_V�C0?@�z�O�j9-���T�?���ϼ�pZ'���K���1������*@����1NM�ɼ��h�wP������m{a&��XQ�,�T���?x�NX'��F�������pr<S��h��>�ݶ|���"�?�&4�Ԏ��T3�&����E޺�5�&�K�6#�Ň(�Q�,nt��7?�f�ND�v���af����t"���2L(	��蓮��n����������?I�����k�\�_<��>>A����*�]�ss̛��{�*��L�wc2��nu�|Pa`��I����z�`JJ���H��?Bd���G���w�����u"I:{�1��:�� �9ֹ�d(h���QH]t���>���0c�Z>h�6���q�>)�\ߜ���ֆP�u�J7�n,x��E-��R�DI��PY���9�����F�Y^����A�.�j���%��8?!��U�Hc ��xU���E�����b#��v&d-�cu1�����x��[�6��I�|X�0�O��P5�~<�]�Y�$�ؼ-qe�+8"�D�솭��6�	���Ӽ�k�<q��ńW�>���U�z#t�<	c����/<�ٔQ�.<���RBh/_��4u���v၏]{o=�+/���D(
v���See%���F�RM[!h7��7����	�P��w ��K:��Z��X��F�T5r%!Y4�P��&#|g<�o�}��)J��
s
;�@��h�� �ʲ�w�F2.�g�Q'P�|�MQ�f���h��ؒ_��@��,�P� �8�pP!d�T�ien���������t*Y2ݘ�Z`Q9oUS�#�OÄ���������Z������\f��YX���ʺ]-�T����0v�CN���Ȫ/8g���#�B�����zHz�?m6��Dq�N��F%KP�>7.yK�:���˷�E�F��6Ɖ@E�%כ�cz� β�$�u;��{�p1����\to@�U���R¶%�y���3��D��y�p[��YM���W�s��#�WX�L��B����qy]��m	=��PuC��D{*� H�3?c�5�@��	��P�,�p�(��T ������9�ݬ�l$�1���ɂ�HG���#��Z/ GS�J~y/�6��ȞD[_��9`I��*)@�b��}�/sn���j��P0��ا���NK�:��~�^O�~�U����qz3��i��ak���X? 8��i�f��,\�,D})s�?OͿZfu�F�B!o�Bݽ��);K�$fZoV��`����r"���Pl����Ԭ���Ќ�Y�U�18�.6����0z�'J�w����^#�2HBe(���������k4�?v����q�kj;�Ts@%����	�N������]h �4���ʳ��₦qc���6��
�T��?K�1:7(�S����wШ�f�Kd�aR�i������!��X�`��(�ڎ�n_�J(��p*�M�ۢ��Z�3d�d��s*��;�| Q�^%�6}e��S5�Y�4��8����|ѐŲ�aU|L� K�+��G�X\2�E^��k�Y��n�#d�
�l@������ٜa x�����M�j�ՎX�q�%����g���Ƴ5o7aYH��PӀ����ִ5䳛�;8�IPj�v��>5�YG�o7�T�A�B���e���x�{�Ubix�M�����g^�5�:Z��`��a��`@Y���]���<݄�"�+��e�Ů}Q�s}Sfzk�aM�ٗu�1�'?���0����@/�0h$�x�H�W�_v���٢��>��os�>K͛�l�L9�Y:h�OP�����EZ\0uYbf�^��$��� &��7<	}���2���Y�%C�p �G��<Fb��+Q�ձ �u[�����;�_�j��~��/�j�K��b6��)��(��W2ӽ<.A��u�����
c���ᇑ��%�z��DyP������}���!rY����"dǤPh���W(�\��r�J�w��n%8^�_�WE��T^���|Ne�$¯�e���<�ncO	( ڒn�~�"�J�Z�(�L�O��FUE�����w�7�i-_��V�(u}rI�Aӡ��c�����?e��Չ����XK�ε}��/�غ"��h��-��z@EV,��`������]�1H2�S�!�g9$toͿF�`���_�����j�`W�b�o_ڂ�����p�b�W��*
fg��1��QMX�,����sd1��S���%���Ëi���I+�-�����a7�o�:������/��x��*
���3������K����1Vb�K.��
e}K�Qϓ]��G7�JQp��/6]5� ���`��ѓ�k{�������@4�3�ڍ�6�m{�*�*�L������ҧ%�5����C������3�h�|�CI�?/q5R%S�orOWr�c���'�`G�	���Qm�S(�!�||��
�,��3����.<�peͿh��-L���x���xI�#:w����ޟwPt�����E�yl�T �L͉��'�oz����};�EO���{A��5EbK������\�����N_�O�_u�>�(4��u|o�C�c�+�\Ȉ�ؚh%�Hd܎��4� ap�z�6I+�X#�>�L�+�m�H��;z�b
�m�,������~j�r��V���SJ؟�Ph� c�R�
��l��"��
��>���2���CnC�nYzK�	�La_Dn�:P����q��p�Ve~t��j�'?B7�;)U��F�G�L���!�3L�,UU��s-VQ��^�5�����%�C�����˭K|��QT�9-�'���_���u�����X2}����MF5�t%���,���p0�P�`������(��AB�ܫCI�0k���	h����e��{��ְ9_��,4#���q�R��B �g!u�h��b������Ta܏ۣ��'J����N ��CD�/�L��<<���)�,��RY�qjVr�!7��%�-�(q�d�K���[/�?�@X�^�����h�c��`���BX���N���˷D��qH_�A�,��[��\��
��iD��?"U,�7�;�P(�������?a�aJu)J4~!�r|%�0� ��zҎ�y���~����Z{��cz�fAg|����>X��"�
�J�'2
���ΏL�qk�z1{�j_?j��ۢ�!�Ee���FpT��[����9BY�He��b����[?�������:�$�L�ٌ}��X�1P��U�,��.���
��O�O?�T԰ޣ�?����ƙ&�5�`fm�p�Ds���E�kE����F��b����dY8��Vؕ=��/4�"wm�5� ����}���67�niޤ�p�a�ۍw���L����۪=9m�t���K�5;4D��%s
E?gw�:L"�Vb��i�~�ֶt���2�^C�M��TA�۝!jG/ҴF�py P�x�2[��إ�;�s�`�v���J}=r4z>�<`w�7o4�������4�+{X5�IDc��L�]+�2ƂJ�j�#cT<��J���͒^N����W�߷��V�ed��.��������A��V����r. �oIՑ����v����Vz[76 O�^b�dt6�J�൞5w�&�D�(�-J����MLa�f̻����6f�v�,���N19�<\�;��#�o�녁�Zu2��ԚPr����� ��/�6�(&������5��c<�0:�j�H7�U���ԕ$��v��b���9���5�`��)JF����[��<Ą_�E�1X��&(��0��K"��*�ǫZ �@�|]��k��1�Gw���Ǉ@W~ԱZ�j���P<���$m�a0�+��r�E+��wa!�0$�j�@Z���M{N�O74����Q�<�C5��,6$D�7ﻜ�H��������g�s��-���Ӊ&Yz"2'�ȴ��m�I":�bi�z�4.[Z��N�D2��_�ڠ���o��R�pr�*�J'�.^}�i"��(����m't��T]B;�b_+�~��z=����u�Xf�	NW�l��ɦ��o� ��Ԅ�m��!�I�	r��Ȑ-��:��}#l��X� ����_��L�� n}FG�=�a\��B�rʛ&5$.��=AJ!a�i���?,$ºe(���	k�2��6μU���9�gjST&'_��t����!@O�v9�+�g{��o�����Uc����g�Q2}��m�Df���Qn��`��G���'d/�����9��9��1�"�QFJG��T�W�]1U��,�/r��c�fv�9f"39OdX'LDJ�j����o�`KQ���)�����NmO?���,��9�^3d�4�q}Ʈ�pE3��;ͯ,*rM�S���˳pz��_\�F��hKeH��\��pp�G�!�"���S���0|���b"�}T�N{ĉ���~YAXg���e��Q�	�KdJ}�n1��S��k��IL SX���c]}����`9[h���j������w��g-8�O	�yÓ"�Q��R���3��|YOF��/8�n����T�|��,@����W���p�MJ)G�#2�XvFf�Q?��G׆��1�xK��ӭB����7� Ȃ��Q����(�ʅ�f��Qy�a2��t0�m���o�X��[�m (S��V�D��^���astUܘ�̽뜐��y��70\����fr)mib��x�ڏ���7&(<|#8|��K�2H�[�͐	Ut�bj1�����.���h��ш3��
���`g�+�%<Ӌb���\���%`B��z���+Ę{R��W��T�5��x��ֿA�W���C�*���ڮ�Ϙ�Dzc�=WJ:��k�	v��
7�p�0-�����$*Z�rB��^���Ҭ�ִO��z�=,"lv���6���w�j~�⯪E?�q+]uk���)M#�#;�w�X��AY$�R��Z�Ik�4���5�P��+�J�q� �>W���z%s6�]2��-QI��~�I�*T�8rT�%�Z���,5/�6q�"�j�$��7eX@���]_�^{i�����E���<��˚ί��d20S��,�*<���Ӹ� 3&{�h|��D�Z~�C|�;&�+�*��Ȟ1:x'�!�`X�~ZLb4
`��'/_����n��m�7��(ߧ6�?����U���c��5M�=� o�-�R�߄��2���H$�;�ۈg,Hj��c�+���YK���O%�{��6~���� �c,Q"zb��Dє=��}��I��w�xi��s�q�Лvu�w�++lb��3VqBi�Qr6�Z2ϗ*���zB�qq�y(Ӎ]����+2�M;@ڜ=$␺7��1���b�!.{G�5RD���@�	����@�����Յ���DV���ǽ����!&�i�� �.<��-ƞAa�;�r6H���z1�-��bdTa�F�P�gȢ���:����vJ2|�"���^��[)��ThzB�O���y�p{Q؋p��x�Tv��zps�K�ÿ���43�L���|`n[��5K�N�m��),���C����\�K"\``�G�a�sޔ���^����M9��ƚj�Zd���թ_�F����5w�r�u�7%�
�7��y������)8��2�i��ș�m�ץ؝�b��[0�Q����F���w�+��C՚(�� ٣� t[?L�\�1�n ��s���n�l"�����+2��ٙ#�Z�1����=ӎ���:�Z��*.S�+F�|�'�R�X
�W�Nb�������r���Ӯt��r��8l�;9���ΟK����!�02N|�o�b���tyYKx��� \��#Z�~#�T׽v�]�8Y���9<5��t����LO��Sɒ~(���|���7�M�P�1�Λ�\�G�J=�Q�s���W�.��evT��h�wO�h��'*�C�񨩼��H3�Z���s�!td1�0i�X��l��u���a��_O��<D�h!1B�2�b�+�S���ߴ5x�>'_��`��o����U�����Ds��R���\�`(8Ө��ĉ�G>/��d�N��Y�.d�H^CS-NqДT���?6�{2��F|Rd�᤾w�D�'���"��4�%�?Ϲ!��Bm?�1��# ���>*�E�!a��풜w�o!�����ř����*l�{�t.�%��D��ɵ˨8��~L�ϧx����ԩ����:@H���R��൤t�1� h�����3��x�̵���O=߸��uf�͌U*�r��l�LE��[+�f/�pwuK�@!��`t1��4�|�^<A����?
Y���ψ��m��x'M�	%�%B���4����-ă&��ѓ���k���@hI�8tQ뺰��{�����{;{/�w���S]�j��2f��vm=)`xf���ҥI��l\�d5��pi�b�#:@&.0#1EN���}M�W��4ᘆS�	j{�Gϙ_���ї�R�G�X�����ਙ�{�� �*�R�q$��jԇt>��>����(Gǯ�ĜF���1$��Ջ�F�A~/骦��v#���ݽN9�<�J�'-��� �E5��(� ?��qϬ�]@�]�^lZGo�F*�
���1�����J�&�;Dr��\_��O������sU}?R�=�8�����I��oS��?#����	�ձ�*������ա�T����Q"b?^H�Xֽ�l�д4Ɔ�����Vl�{�+�P�Tr��L�o|�^=*�1s7�'��}�gA2��(��v+^�Ĵ!���.�.b*s�-:�^Y����7��� MV �T-�r��Y���[*�ak���=0(ɦ�u4Q�Y�)B�5���� �@N��t�.��9+Ţ3ܮd@8�Lg�A����E)ز�������i�.%��6�쉠c�Ӓ��aX|׼uɣ i���G���I���_������7��$G�e��Y5<4�V���,�0������}���L?�/a�r�&�9�����7�|���`���	��@������A��>L�4�C��:I[X���Q����x��&�
�\��J��<��ܯ���I��V��tJ9�zF�.���7�9A�e�8I�;���*��в~z��p|���(�+�Y6����w��p޺��"���%�6�a.��f� w�uN o	ަCY¢�a�VL��$��!�� ��F~ъ���<���d�{�@؟��@�zo�E,�V/�k�*�T�ATw�9V��jEI;�}T#������� �ן��׹�MÀpQ���vҩ��6�X���I�M���|_\�ꓠn�NF@ߨ
dDqv�l�^�_s�y�JE皥NThL�ėBg��D���BP�����{$�L��]�as*	��R��L
Ϫ��3���=�k�T5H��#N�U�K�t�x���,��b�V�֝{��>�	0A�bM_Ec�Y\j��W�		�_��_<���:oe�[Ob˒-�d�2!W�{t_Ai�� ����戥��咐ZZO߂���a�n��=1��(��q�A��\���Yr�C��	-�@]Im�e�|"t����O`Q/$�I�X�p �D	&�D�*�-�D �K��7s���������4٪E�����MҒ�����H�.Hy�un�u`�C��+L��1������$��Du�����жjKU�����_v��v����#��椉�|�	s�.�f"wH��e��n�6���n�kƑL��[�Y�� ���}���z?<�̷���1����l��h���-�E�?�)���a�k��@C{Ͽ�-�%V��j6P`Ru��6�ԣ��Cn�n���h�>�B�X�\��-d=�"9���Ű�M�v``=}�]o
���8,
�r�Ta�\�7��N���>����6�:�htxd��W�,&�|˨��p�ܓ/6:��|/֨���nh�FZdO[{gen�[P������>�]g�''��n�2�w&/��) y�6e�< �ʵ�M\�
��Ş<�#1�R�x��sF9'(q���ŏ󮥜����^h뗡�?��A#�b��U�i7C��v˂׬fI*��y���a�oE�1c7]U^�-�t����6�ʽ�-����\����4�f��d�'��gvm��=G�W����&��'ʤ?������AV�����,�s;Κ�^L �׷XM;R�5��-T�6��
[6�>?��k���/P��WC�^
_6G�(*�bwt�!0�����O�b����;JV'��zay�5|��_�չ�9n�������oʶ����q�M|���7���yeN/�@�p�w}<�G��\��A�y�V�8�9���w̺uA�I+!m뗦�\��ZUB?��;˛�Y}6zj܏�;B�Eg4Ĭ�Z�1�-QA�TB!=Ye�t�����Y�Ne��jA�F�
L�=��_y��E��/�e�X�<ū`6JUm�؉"��<}�l�����u!2Ǚ?s8��o��Wq9j�ylx���V$J��_�5�o�'8��[���p�'ES��U��)��w�6m��)*:@.�O�o�T�ذO��_�L_"0v(w�j|B�h��
_��Q�2���������	��'Rc��<���/qb��?�>P���/�0�S�vi��u�1~<t�k7A�g��5����M�%Dt����]6^l�F[��!��r!�����Y/��4��1��ᅏ�2k�H���-u��zI1/܀�ƣ�f��Y�G�4��6�wh,�{�^�&���M�E�K��9*��`�I��ED���;!�d����c�ıA���.H(m�Q�Z)Ě��΃Vl {lr4�}�.�I���3�*��m�x�in�b�M6.\%S�%��Zc�!�w�(�~�8��:�	����m
L|,s���8�g���qB.$%�]�^�q`�#"S�a�:��T��8��>CUh��&I�Z���.{����^��d+q��������i�Z�#�]�&h�+d/
���; ;c��1J6���8��ջ��A����D��&��~h�������q���.x�S|$۠,2���Λ̂͜�z~�8J3�Y-�dEj�/=6l�]1U�������ђri�Q<	(�>��đ��ַ�'��-@V�M�w�z�4��G�Z�'Ŏ�AK��IJ9��51���M�T`b,�H���.���',��Uv7���}YX�,�bSm~"vv����W;�@���q�r�E0���q%Q��D�t - ��(Id��1(��z�g�_���(3��N����<��[�}���H��j^���+m��?��5A��g�jt�i7D?{+�E��ɷ?9�#K�K{���b9Xj3�LG�4��W��@FLj�?4�m����8�Zς?vˣ�����ǥ��nJ���Vv3����Z����χiS��e�I��
D�Q���E%�p���k��F�#%�=X$�{�<
���W��]�j��u�/m#�6'k_	.�CH���e�N�a? ��u\҆ӝ�4g0�6F0c����W�����E�1��H{�O��B֎�S�Pa�{E�4�Ǯ5��n�w���9��Ú�)�+�NI�ָ,h
������R�+_G��Y*Q �����
O���*�[��gq�}��h�A�����=�1�"�Ky�=���'E�!o#84�ι/I�LJc7^��,�*p8&�*$����P6c�]�����JĦ)�QJ�V���՚,������H1K��Jc�:�-��\����N�{�������r���
�Ji��@jL�p4���c����A��A��Q���P���M����vG�<�Yk��TS$>��}Ĥ ��>D�	���wR���E�:R��j�?���ՎU�� 2\�{|vTsg�+3l:T�����ư~zax"0��+���o�
�c���e
/����*?.�e���v��1wAѾ��(��y��0<{u
��_
c��)�{M��g�
i�P˂�|��e�j�I�Rle�R��?a���:U����_�,��u�e5�_\^��F{bh���,IhE4B@{�����ѲYɥ��j��Puh��K��@��W�B�k��]�:J��z�e9��[�?"���I&����$���|�g�qHEb�1� �Pl,c:BG>ߤ��ra`� ���|���1��R֫�P��˔�@��`�pl��F�F�fC{gm�~$B�L+��^!�W/��a����/�Sv��2�/��;T�}b��8�^q���Y�R'���fr)���<��M����Sڒ=ް�� ,�<�jO���XGF���QI#>�5a�zN�kڷjK^�3kW��}�N�b�{�9� 3�;�odnI�_
ϡB"4b���Sy8V/��K൅����x:��V�%u��p����ʚ)�*�M��YX��0�%R�M�L�l'�܈����nw���D��T�Ij�?���h@h!_��b�����9�n��;����������{������2����3�.���D{�9���>>�wM�-
^����h�$a#WolAb^>�������{/��b ��=��������p2�*C�0`=Z]؉y��O�	8P�L<R9Zl�i�Ƕ@p��)�|�$� ��r]��@���ڰ^e	�{���*�*ON���l�$�"�
{S�%wP����D�<����沞�z��_\~`��M�=bK?2	�b�x�>�d��6*&�����d\�<�aP�7�z0�s9���|��j�u�t�)�0#�:��79�)�'�b�zWP��؍j���\b<9�qU���򉝷�����>h��$��\�q�����p�nŽ�7W#�M�5y�`�Ԟ�ӫĭW��&��W��$���:�>WQ��;����.@ !��f�\`����9x�FO�+�ң�4�w�D9������!�_?2�(���\�@iB�4E���o?wt��.�l� k�a�T@���y�MR鏽��O����"�=c��
̴�z�G�9�"N����/B6Hd)����c�dY�1zS#��� �݊����~�2��4�'��/����rN�!��2��`��".�G<�U���~E:����^���?��"�PٞM�U�t�
ya����3W��i�x�BK��먺C�F�4ٿ3�,F���g�a��q/;�����:�%���[�,~�e\�ߍ����p��`��Į�4�ܟ=񥅀����*^=�n�B�u��s�H�1?�ե:N�b�Δ�T�KjxY�����?�б�&\��]�'�g��)^�L%�|�f5���-K�`��9���.�ژ̀��-����c�VO�"�Kx!f#�G�)p[�:5�ph;�si��PP?�)�x�*�����N�$MoD��i�Ҟ����3|{^��ڻҔ����E� �}>r�Jݴ����B�������Bz7+ra�Db �NM�	Y|��w�� ����q&F��y=��U��~5j��x�q �H�p
4���rK���2~�|J����8�8��4�|D������9��n4�\�J��|W1.C�:N/�+�H�8�n�Xr�E�~��w��Ag�d��5��6�AMځ�����"uG	<?�R�l�Y��q�+��G���t��/���d�=Bz��H�ɨ���ݓ���2��S"�Ŝ^+��a\��I�7���bt����H%w��5\�W\������=ӗQ�6'	��];��ݍp��>�8H��pݿ�z,#T1�8|�=Y��RlH˰��++�H5�y����6�ƙ��vF��
6�R�s��5 Z&hwv��-����b,Փ�َ��2%��U�1�hq�ȖH�9E��F��$7p�����U�:-�ٙ8�-��{I>~�4�l�za��(�����"�x�������W^�e.��@�צ�`r~V��S/\-..r^��=xwl/g��p4F ��f�y�����Tok�ʒ��P{y\� �>��a��E�_�.(P ;�/��%�c��o�wO%��؊i�}�������&9�<��k��r�Pa���&��I�>��/_\Զp�q���7��Z�Z��(�oCl�tS�p!�z)G�o~^�<�:�I*�����x������{��|�&�҆�@�#k)�#3Y�k�(F5|���T���v;~?�r����pA�A�5$��~�� ܔ�g[DJ��pT?�<�foD�UU�GR��3� ���l6X����S�-���	@ ����'@�&���x��b�Wv����k�w�E��@DIN��u��8L�~��8a��F0f'��?h��bb+Ը��h�� z\0\�6�,lh~�P%��Hɏ�v��ɟ?P��4ْ~�\nM�\��-K$�&�	h,ʧi;y�烰=*k��'�EH�=��֦
ը�W~`�]���^�W�4���%܉(��KCc�C��*^�k�j�X;p�ѧz04A:&�j'�:g7�'���A�c2N������¯���S�(Vߚ��O�x8)���SW=�_��[֎o��Z$��%��XM�A���Fq&�W��Ua^� U��y��!%�8��%6�g��}u�r�}�֗>&k��:��P>�H\�P�9^g��k��V��F���hpp5	J�F�w���|q\�s���RG�h�� E���n��e��Egm�� ?���s��c�C�Y���y�B]��@������v8	�����W�y�ݝ�)U�ÁJ�Ǘɩѻ��Ñ����"�]�]Ѵ����j�WU�����t�Zh�z���A����*���s�WO>El���6N@����m���IdNU�bxZ��uљZ<'H:;��4J�ڵ���σ�m˭�L��W�O�����.A� -�
Ģ���׬+����5I#n�5�o_�f�o�!����y\:հ�s��}����O���Q=�T �ݖ�Z��8(�=��L��B�|���w��҆2w��(��,��Ϫ`"��'�
���`S��A�+�%����M?LXߡ�-EH���r��}p$s[i�+�UR[�Ubm��O��(ƾ�����CpJ����V� YVp�I;�C1��F*i6|i։Ɲ���5d�JW��\.:Qhe�#Ɍ��C9�.ɖ���G��W�n�v�L���6%:��Z�˜��/vҰ�
�F��ye��t���OI�J��M�S���ށ+�_�tX��,ɜ�)�'�RB���/��/SV�r�,��\��ͤ5i�)��u���s�'Q>]I(�c������_4q�Z� ��M�I�K|./)\c�)��4�9�ÍE\�ĳ4��4D>ɭՇX���?�,	�J�-�+�L�
_A��(7�k����=5-EWB%{`�<�3C^�K�DC
^��l��Ytw�W��Uȣ��]Ok����=����������s�ٯ�÷d�M*X�մ�vM�eg?2Z���^�(�pbA���}Q�}����nٮ0��!2�@�������X�����Dm��� Φu�T�y�V^F��*�>G��9~����Ty!�t턅�$��0MG\�qſ`���d&,���<R�ds~HG�F��b�Ci��)�2N� ��T�z��-i{L��7�T�X�;� yR�tr�C����H��,��e�-�j�QۢZ�n������8e�W��0/^	�+��a��Q=�#���M{�pI7]���	��_.M9���Qx����р����Չ�4��X"��5h9c�|x�_W#��周�$4��o�fA�E1�����ڝ�(,S�J��D�/O���&�%���n��}��-#>2�)0��ê֠�u��ެ���qࢸ�����a�>��,S8;ﮄE�ڍ	Q6w�}=�� �Jit���T���X�$���1XE/-6q���'����Aq�]�'d	��[0�Ջ�	A��xg�"גܗ
_l�X)�/�>C��f�<�hjH�K��t�s��"zL|i��������|ן��~o�GeY�$��9���l#��A��3�Q��cԲ�vR�22�qe_�>�ȃ'!�X	�2�n?�ʺʥ�_�:�	�1��Qp�,7�{9�;�9X�kݘ2~a�2� �:o�֕-v����@Т��+��p&a�wl	?�b��};.��`꒲M]\�e\[��i���)�Q_���E"(VK�L��
�Z6R�����R������~	�o����y�͸��z|Γy�����K�2?�/b�D�����J߇��pfdt8 �.���O��	c�+�l,̶w �ʳGg�	�������WO!�Dؒ���'EY�H�����]����m���ܑ��Ǒ��#�����*p���fPĂ t�6\�!��Q�����|{\8v����O�	h��.D�tQF]�#�R@��aaе���|�D_1m첯����Z;2g�U��+C�UǞ@IE�&�-�e��wG��(��t{�?�D/w>�$�.�ƒ=�\K��`�����j�Ue;	���������@E�%��ҡ�aүOPќW����&�q���խ2	�*<���wQֵ���{��2U�H,&��BG �5��W�� >�]�T��ϸ�B<�5㻶}�=��]��Q5�ޘ��L�~��[����w�˦u3N��a�r�t�c-n�'Љ�c����|���:�Z79�-�|�*��մ��yu��JS�Qͩ�V�K������c&�n�iJ�/���u�V!�N3$Cmg�uܶV<d��S��h?�il�vKI��y'�^x#��|�aK=R"Q�'���˧�̡��մ�>�Y���Dle��2�E��L�VI�+ѨTY����B���0���ue�����P���"�l�M�GS>0������՗A�k��G��7�ڸ� �f��9�VT�T��A���3t����
3���P�F�&�8I��*(����G�u�R���9v3қo���S����g�?�C>�<�+���\v� O�A��HQ�:)Eɭ	�b� ����k�`=n���׍�.�,��je?n'4?^-��Z&�0�!��Ü��A�[{��_ӛ��G]�_�Ɔ��!R���2�},��A���o��K�:�ٶ��hpz���{�kmV[�zL�p���M��S��� ��!�&w$u��g^v��o����K����D�<)l��k�E��
��!1d��ԙc�I�+*�d�J��H�|ŝ��SX��f�.H��P��Ɇ���e3�籬pV�K�/����i~���������a�-n�ۿ�����;����`?�]��a+,���Y��&�����#}�Ub�n���� ���Lc��,I��!���R4��F� �7(�9Ѯe��Co[�)�'���#��;N�>�zǏt���(�]��;���^>	�i.�?�#��^�J��z���:(����q j�)~𿘹��%F�{��wD��w�DV��z5x���ou�ew$Đm��kq��K2	����-b�d�����i4mꏻLq�f�e�J�~��%��*��TV��tYji����;P�G
����@��	FP�t�V�h!�����tw�bڹ�L�y�$E�3��@J7��Y���E>�ga�!Vy���j�I��,��;�oy���|ޣx�ۋ��*����p�a��6E�S{�XNd��^��߂�D�$��#��$@ �\�x�p�F�Z�˖�㟫�q%}N޸$O춯��ڬ�� �7�"紓ĩt�k��h�^�q�ߊߌ��t�a�uќ����tB��/���\�J��G5�KJ:ZfW2G�{F�T�q~]ʒz?���L���PK��Y��`��q��ֶ-ZKl���M:wض\�PtN��e��y��l9�zv��¤�ޒ&Z�F�g��L�y��'?9�1C�I#	Ӏ����{��z �ͥۉ�-���������%��zR�d������F���dI��UlS���^ ,��B8���j��S��]��b�z�׸��Y����^������}
Q���2����0��w�^v�n�f�{�훢P�K�R������Nd6�i�A�vf�c4��B�~�;?��ɡ��Z�(/A�n���G���s�GUo\�[x-<�4f\��!Kf�U�KW��נ��}e� 6�;߰z�e<X�O	���h�m
�P�zo�5!Rͺ��1#[�!�``�h#W/���K��<�A٢~9���c�?�kC��~-������!�H)�C<6����K�HpXʹ[����I�"C+�y���z4ܫ�q�����ë�%"M�L�CV.�l��$zE9պbI;�+����XP��3j�"�Y6�����W�������Ί�_'�&q#l����/��I,ҷpM�4?�{e��;�v������Z�� �̾!���t"a�����x�ˎΏ5��][��(O~�R� xN�׿���f���ߛVG��C0Yv�^��I���L���N�\Q�S��
���Q����C��R�2��ː)�U�s���%��S<�Y���Df)�+ؖ�>s�2������MO����;�s����i�*�m~����"ѹz{*� �T��������[,}D��f:�5��2Aם��k~��1,i���y��jv��5Q5�&l�
���vmQφ|$ P�v���d�.��?� ���Tȍ��hyY�y�e�ʛ��=�C�Y���/2�9:
������ �8yYYJF;��Yx|o��'?�p�N$�h�RR�n?�o�	� q	ގ-.��_��*��Ne���µ�M��Hi������C�*#�A��E�����伽s8͍>�����t�mKbR�<�w{��v���A�eB�
�B�G�����C�F�����l��C:�<�%��-��}�U�g|N��	��p�?鰍7� ��(�s�z��bL.�S*`�_��z�*�Z���%5����N��M���-�5[
��W��t�R���	�VC�{r�y�������;�<��*������E�����O�#� >n��Θ|��ή�����{)��D3ڊ�XF��1K>r0 Ż����NS`���OJ�ıZ��(�ZE�@ 3i�6��s^�n��4�qQ�Cb-�fi߸��=V��b5w�p0�X@ͻG��>���F�i�A�Ƥ�L�j�ᝪ�3v[Q�_��|�]r��9(F2�,�\��WCKV��Ǘ�S.��r�m/`�a�ѲV��R/[�P�H�#�Y�3hQW��@o@��q�9:n���H��M¡�CT^~�V��<E��4G�V�m$f�"sႥ���&�L<Y��������{�ZR�?��H�����V���&̉�V���A�@��@�q��\+�v�]1���r$�|������"�JN�a h
���t�y�7y��m�L��k4�$s�ho�����,ZO=�l�s��Z4A/;���ؒ�m����o�g2��tY���/0��kt����A���`�70o�>jq��I�gS_� �[�Qp�i����郩U%3å�C������l	T�k3�y:t. �"�M��BЁh`���3��;}juS�g(p�?�fX�5��.i���R;v�V�3��а�l��4��/��遇T��#��@���;y��h?K����{}&b�.���$���@��[�T��#j�V!\�q&>�����Hy9��)p�l�O�:jݝ��jF%�'v��v��IX��FaF��h�;��r������(;�����	��*�O3�N�V�-j��	���C0�k歕]+�-��vA���":���XUc�I�t'%��sb�`��{�X�^�Ƃ�7l��C�|_���p����&kJ/X�Ÿ�⥍2�.�{��0vz������8x`2R�4O�:K^?��M?r�1
��C9��w��GcaOK���5���F;���@�]V1���hk�6�.�Y���OS��2ނ��}r@p��Z���N�ל�p���ۑ|;ws�|ţ&v�f�G�B�qW����b�d~�U�1�����G"6�2��3KB�uS���(���CCg�ۊ4� �� ��c{��|�P�B����&& "_.�;!DO�5�]��tXF���Bp�AWgz�U̍�7���.;����=����**9���d�j�.i&�;���r���{�8^�>Ub@o�9.�p�����
w�Je�Lu��qKu���	b��ք�/P����1�봽��Ba�zE?��.88v�5��/6�R���t�4/��:������H�|����*����HȵKe`������+^��1�&��)�O�J�j
S�P88*�f͜���g�v�I��Q���^3�5�4���v�0x�-���h1 \��ˀ���a�Ǯ@#����㾳벟�H�Oc �)g��P]����q�����g��E0�
��ҍ\%o��@�$��T��M�PHYJ��|�j��\�������/*��"��x�x'v��apK�O�B�.���t"�����;~�3�y�m�-E�3�f��S`�1�l�+��s��+�R/S��+ڮ�R����n��4(���9_��4K�C��<�JtM�hl���ѯ�TmJ��fz�H��g�*��cp����*�%z�oM���F���0���9-�<<��2\�hd^գ�ǘ8x����"�1h�~��.�+ys=�EG�H�P�}x�d]�9�dssk_ָ���Z�(�"T��N�ky��C9a����LV��GGT8u�N�t��'��;���w�NU�6�.�G�,z��ʚR�B¢�&$����;~��x֍�s�n�^㗛��F�Pj2�4m�&�Y+��-�Cݿ�T�7=շ��z�z�>�_ү+���WH�<^*~�,)��M�<G�C$�{�hgWm����9EȼP/h�e)a�ۧ�i�Ѣ�[��4�np�+|�my��	��r��0&f�������q}Q[��M0����s�b�A������{�%fg�Vv;�oң��&��(�Wi����T��w�`���Kt^w.�[��3�ݮ��9��=������ڲS��5�ie}�nS~ �Lx��j�I��	��3���p�������o+/��a��0	��M%)n������w;��٢Ĵ����eT�v}�95{�a�C�4��)�<� �2�M(~��5Z�F�,�L��:,ܔ�a��-=��(d�D8�Zv�W ��+uS~��M�@�By��ĭ�@3�A�-��dz�s*��ϣ�3�I��{��G�][g�Kяঐd�"?�c�]�?���zc�%o)�뵨�ӊ�a[tV�Yoj���s��0Ս��iq:ѷ��"�7;�e#�(VN�k�W;{p�i'�E��䥽���L�'��Ȫe��7�GjOn7�=%�����O12�K>�b���r:#yJ܅����A.~��X�2�h�ev�D���F�+���}��:���voޭ1�0�x\�CJ6��aC>�|��oh����Bl��	6��b敘9�ݟU����!cK���ME}% ��f\����|�NE����� �"F���_OK��@"D5����h!D�c
d�-	�x:j����.x�>�π������R��~�R}�M4"'��@�;Ђ�#ĵ
Ě@�k�����$����e�8M��H�|�L����*㯠6G���agP6��!Hr\�l�a$��i�ʒ��Ǚ�<'�)��ڪ�G�J��j�l	�<3��V��m-Vd�!bA�=c������n�h�o�˲��8�-���d�Д1�)PO�`��L���uBsC<�elN�Mk�F 
��ۊ�8(�K��;ݧ�-���b���?nɤb�`��l-�'����p� �2�@y��/u�_���`$H�!hR|��'-� ]�L|�tA&�dX���O��mZLdE�o�kF�Vs1tۯO� �˞7��?��W��4��l`�д�s����5�s�xQ@T�����=�f���*Y�X�C������˘��Oq�2$�.�����L��삃g����������(�&�9g��Ը�].��P;I|0��{wg��;o_w�A�0q����-�ժ�o�k�+)=3&�>ȃ?��S�i�n�k)��@��2�t�ے���_�	��ی�{�r��e�b��SW0��`�5Vs��TL%(7ך���+�'GF��-w�kE,4���D��7�I�$`B�� '7ӽ#�g�'ϧW),��s�d���#Lw��e��g�PW0�a
.r�r�e�$Z?
�"�J����h�:�fb�350:zs�#���
�����&��s��0�M�����_��4֘ev��5{�LSB�kĂ3��@�C��Y�l�-�L�n��U[��z�� �P
��:��eɌbtUD��r����[k5-)�˿f�#�y"��WO*nE$_�F��]s5���$�ߔ��u�RfI	����p	%�_�V�||k�,寪y4���M���22����Y��9C��x��F3��³=J���Ñe�5��6v���,櫣|LuE�$j����E�C&��!�����ș���+h+HO@t�����p���bq��_!(l#���lhMo%�WzFp���)�ր�
�{��fZ��[�ꤟ[m���璃K�{�L���m�PL����Tq�C�������#դş�*yc_��>�_#�GB}��-_�� � * Ւ�:�U}�V$�0J^.�Q�-v,&�� �*z
-֌��fPJs��m�)���������8�ځ���Q�M)_�䊉]`���K�zq����?>îЧ�렼R�Q�{]n�����y���z�F�[7,"��P~�!z�*#V@�Wb'2�P�`?T6A�<_��-XI�BQ��jf�(��d�O?sc"��Z֍u�Q��"f.
� Yёh{ʛ���/B�,{s<3?e[D�����^�
�������0��6%��ڵ󢵇�������)���6�7����������6��[G9F$����	7s��������a|�ȫ=���J��rC�I��Z���{E?��p��Bsh���3�������PW:�yۭ����X3��l�È�sf&2@ J59���'�5R�&���+��p�F N%oMo���Tp�Y�C�%��ڈ1�9��V��#
ޱv� ���pݢ"KwI2�{&�+T�~�+4�r%���|-��J��Ƙ�]q��<�kj�7�XhI���F�W!����T&C�z� 4�UC|�F#6�6v��U �Qn޶�C�i��6�D���z��.t�ٴ�7^�F�.ش�wu ��;���>:~�T9�o3�N�/xW[4�W#`���`V�*�vqDߐ�ٽ���}�w(�]&��T���}~�ӘR\�l����׶�]�1$8����`T@�w�	m��Ic��q	!���f�q���^��v!��u��g�F,}fX)�M/��]�d��ff�:۸O�2�����K}Xʈ�ҹwMz� �u����O�ě ���rRL+�y�xa	��{�7�1��)�z���#���ẍf��`z��Bу~~˦�Z��R�
�׶�QX�6W6���ڢW�k����
_5�k\�Q�)?�
Ħ�8q�iO�2"�'����h�tY�O�o܆� ��Z>"r�+��7���"�ipIGK=���%�e�h�ͭW	��T%����D¤��Q��H��/�Y�
o�m����� '�;��0�0���6��k/�#BQx�U��b����^�����x{�9ݾ�4�B)��܉$�}ƛ�ϜYY6�c&�D�4��G��-�ro�ʄ��gJF3� �Z�--̈́�|x6� &�R����j�E��u,͙;h�ڐ;���g���-�H�vJ��8�y�/v�)w������10I�* v�3ϔT�����6$9 V�o�Ѧ�j8����u�/7�%�`��
��m��[@�u��YM�V4E<����o�!�q)�H��W�Ye���ߦnv�3~.��:aݤ��t�P���F��z�
��z���U�}�>'M��>c�47�ɣ��x�Vh�t��;��T:g1�D��t$�҈	M ��ҭ���N%�'�14m-y9_R��V]���K�=<?f�)?f���H��_C���0��^  ����Hi	{�e ���R��;�3<����U��"{iL�������;�` �f)m� :"� v�o�;�i
�h�G!�����o�^�h�ɗ��O��S>6�-�;�s�o��]�$����&��&$:���)$S`�AM�9��3u��ZW.�}���=�TD�H���9��\��� #?����9Eb*��~��Q$�v�9G��5%�����(�?��˅�a� � �|,Rp��*DL�qR��0�I�'N���y�S�������e�(��\1lL�#�0����6�P�!\n�W�P�*�8]����	= �?�h�Q��,�!�E�
��͈��h6�FaS	�=��2=�qX�P��x�$�&�4 ���͆�Ø���T�?��3�ig7�w&��"d2�P�^�u��ou�ALՇ�w�f��%�a�����eҒ<�$C�uPGV�!d��n9¨UDE��'j�(�ݳ$�B_���W�#�mG��w7�1X����=�Y��y��G�`�H�0Ȗ	a�V�F�4�42%bwEe(L�ԑd���?�ѠS��>�	�[�1J��X5*+��֧
��0l��}��vK���np��R(9��DT��/K��YC������@k��T�)=�A�ܼfuo�!���c�����{�o���a�c
;��*&�1�-ۺw'�z�@�BO��(��m�LW���qwn2��V�����>�mZ"#��qqc��{���m3��,JJ�`�ta�Y}�vN��3�&���T��n��E�,ç���b��;==/�ĨX�aYrN����%n��M*��V���+x5=Ec�P��t�֒5�V�P3��N9�������1Q̩���c� LѰg9I���m�ky��/�#4D��ݦ�X��|-_(�7�<jbp�b.�+�k׳�J�,}n�ʻ맺D�1S��H7ċas{x�J�;�����L~����<�~��4��H��>�z��.�F��Y;��;�N
}KuQ�$z�[2��PssYc���P�~�Pq��i8q�H,V���Uq� :m%|�Ì�u6���ʡ�"��y^V[(�.��>w� o�*��p��>�j�71��G��L��~�U.q��t�_�ӯ�!*�Q��D���|+Vxa!W�g�K$�,M��O˨�]����J��^*Yߛ���]���%uĊŘ4_�������1N�Dt����Fb	8��G����[?G�h�H@E/H�ӳ�}�̀r�Ks�����2\9�8Y�����2y.gJ�@��G}��F%��)ʷ�1���;;"�F��(���&i�\E��%�L�@`�4Ny��iZ!px��h$�� *2j*T��{H����T� ���+&�g�&ħ��:�Rߨ���^"��P@�^��	9����Z���.�6�H�RT���v�>_�'foH�G�Ҥk�"����;� �ֈ�!�<�*}	O,�I���RN��H�wc��}˿��������|���:#��;,��iZ
â)�p��K���dke����lx�:B�گvӅж��C�g%�D�T'���!��7 S�0�$"��'�t�7L��P�F�����%aY
�#�Տ�v����!r� ��k! �i~�Cc5�F�Ut�V��_<B2�V�{���1$��u�hrv�Q3�I�8���3�r�*���}�"3p�;�ٿ�eX����A���X��1�i�۶�?��:L!�{yWL��r��Κ�m ������ju�J���\���l������F���|4~�7=�*v��t�=��į#��kD�E2�aRU40����A��ݢX� Tf��{��.
�w�\r����\�ٯ<�&��^�J�/Oh)}��xjx5G�d��yVad�n�0�j܍T�7�υdc�Ԇr�(�MB��H4E�&�����T�*�
��¤
9�P�b�-y�+x�c�F/��0�N�*E��;���ъ^��u;�u��d5�@l�@����'@�����	�%������ ���L�aڲ��i}�?v�����/({w804�š�G~�1�ܡ�mu��R�ث�'�|��������e	Cp/n�=�7�W���_~-m�iF��i�&9H��d�^�?��4{9ï$,o<��[��41�(�R�΢�̣���`�5H��tjl��%PP�t�-A2V�������v��88���A�mQ�նZ�E����,�Y7��n<B�c��9�D�B}cy��~��4����dB:�Qj|����1�,s��:��Q
�{���hE��次W7�E�΄�9��2��I�n	�37R�G+xi�������72� 	ni 0.Xh�qF]R;M�h��Q��YY�-��C_�[7��n�K��O^k��n���	p'g�܏1-�zV�q(h�uRŗ��(G XS�Z���?�g�i9�Ҙ�/�Bhi����h�A��~��y��p��r�>	D	�4��T��0�#'�j�B�W����]��X����1�A(��n��S�Pb�`�5{�l���8��7?@ڋS�_��v��䧋�2�Nq�� 4����1�۱m]V-���{ȱ��k����x�Ⴕ8�K�U4�����>���<GDK�m��a��J��.�IĞ�����A�,M��}��{���� ��b��"�n'������:�}?��'~Yy�)�����u��N:d��c�D�xN�@��-��6���.��qY�E��n�,/7����+��h����m�'��z�'5�|i�%������{�b��(-Z�8��*[T5j�56O���~n�[G��v��ĸ�n8��{d~���@3�.�J}KYi�e��J�8:}�_��9��ę�dG\���r㸖�%ꨌ���G(�����]�<�+B�_�xX���F��:(�����̦��[������\�g9x���ވ���մgݞÝ�뾛l$�O-�% }ܛo�I�G�]d�G?e�([p�}Q���Fz@�\��Y�ҫǅ#�j݋��2�H�q��)����0O�DX�k�{yo���rA��X=�gsþ�j%�����amJ����qwb�|oB*5u��U�-���I��"��-.���ֻ����'�cҤhj�BL:y;y��5$�²;��=�y.$#�����LTx�lf��s[e���T���m�Ѐ�/�w	�\Velh�b4ZB���t�2E�
�d`�L�ʙ��$��Q���,�	�(4\�2z�z�Xbvd��	�砹z�̭Y8Ly-��C��-r�� ^`-�2���C�І ���iZ�Gf��^�t%�@�i��i�,5�vnH��s�����t�]��5�,�j2<����Q�%C8�&e��ktb#���]u�0��%s���;��*��{\̱G4@2����l=9}ˆ}���Ui�C�S���L�������uw� �=�ZH��{�ӜL�fÅ%�x���d��"�2eì��M)��		�y�L�#�C�Ŀ�Y,^�?�u�I������m��7��ݻcQ��R����IM�5|:��E>�����>QAxM�>�`ʜ��i4��+�l��ύy.#9�ga{)r�q}�	�<:5�Հ�Y��Ҧe\ -�+1\��>��	����y�'l���Q�|�����<f�.�J�Z:*���x[M=;��O�K�Z��4�gD�'!��|ſf�����F|��.�w�K�}�/�fv�"jG���%̔,`�1��"~�׳o3��V-�\<&��`c���Z�D���TO<w㖾�~>4�wZ����Ԟ�������{�l1�fc��F�i�WSȉA~M}���
*k��+'(���m�F7�Tu�L�)C�TGS�
��p%�p�BY���J������)��N'_ar̄���ܡ@��M�1�'�ɡ��h�];�[oP`���ڜN���k��@pzb��J�}X�&y�ߥ����Yρv��Pjz �� �,���4�$؄�q�o �����Z�:��!�Ut�O%Iy�$=���=�SzJ}�T-�?�0�� ��SP��$����h����F�Ȣ��RlR�<��@�6�� ~�Bɽ��N�w�o#�{�+<!�����$'�"��y��d4�B��Y��M��7��ʳ���t�q��R|CeR�?��Ig�;�[lD���|��4���O+(�v�*VCQS[���a�~���)1���\���e�'%��,�{s.���UH^�Z�S�E?�CY�8-{b?�yw���`��e'�o���O-C>� Nؾ�@�zΤ�E��@�-i��T�JW�5ژֈ3j���?��U�:��<b�3jn���up�\S6;{��G����B�гe��iY��Fu��|�������`��ݬ�P�W?&eS݌�G��G�04%�u7
�� �2�����;�H�ř��ke?� ��w@���ɜ�;�Ql�zW�F�%��6��?fD̩��t^���!�	=&{`	|�m�PQۻ����O���mr��Q�7���!�	�
�ڣ�v��&���x�}�� ӑ�a��c��f��V{��C��F�ׅ�;i֍T�W�Kx����|נB]3+	���"-!!�9I��5M::�m�l\'�0�kh�gWTFB��5�@~�j�wt!b\�i}�ӗn��ҚExt4��d�{l���X鱀6��Z���B�C����*��J��Q�31%�[d�s��a������Ɓ.�/���	G��p �B�I�|�N�� f6�[��B{	w�������꙱Pli�8�D�|llS�:�륪Ǜ��7�t_,��F`�R�J4|�����m���] ���Y월P�F�|�qN���2Y�q�֏(��z�}����]�R&g��?`��8�(�u�)-����+JT�ZK]k$��d��,��5yՉp��S �Š�Wp9oy:n3�j����ԧ�B���uXn\�̧4;����m�&�F*�UrV.#֊�qO@�[]PgS��@�#ٸ���qK2P���8��b��k�j��%�䂊���>bU�B�~�~��|9�`�IKO����n7^[�۳jh[� �a��"�� ��/1Uz�Bu|��:��p������Zf�9ab��ŽL���'*6��C�CNc�V��t+%�%d!�c��&��re�=��-��5($�^�r���)�V�ۼ�R��`c�Q�]s:�@����$p�A��׼<kd�iNQ��D}��,nc��񉠾�h'���'��u������:.�j�0b~��ܶ��w��o�3�?����(���d9�"RڊTSv��*�����poY���΂~K��|b����S�Ԃ��4��TXw�D}�L�*�R�R����F����GM�M���%�X!�y�7^Xo����6�K��v���`�S�g4R#�|b۴W)I1��B�G�,�&����J����-H���Eק:8�5o�.��֡����~P�[swCā��r)��-��dsk�g"xF��r.������t@~������*��s�� Q�,�WRM���1�z`���T��9s�P�N���T*��wsj c�,��S��VƆ���"�u��[7�������ux�s��.�}B���-։n�g ���:S�ȃ��t����:���]�/�BH,B=l��m6p!�� s�yӮ&[�2Pb�+t�
w~�S���O5��Cp�j?� j� ��������a�~����%~x���~2��\7Q-�?��	&�ڥ�2��Ӕ�|�ü��fY�,^s��G���!C�B><�&�~FѠ/g�|�Pv0�đ�W!	�x�ź��|�IO�T�+_�`Rf��~4�&��&���<���JøC�-c@%�	�h3;!�������c��/����L>�\��$k)^���?�l��&�d"QC��GAR[z�o$�Xr��o>A2H����峒����w��=úL0�����K�ѺU�%UN��n"WX��%{�,"��("}�5��Uʦ�\F����+���Ϲ���d�7��{��k$pЙ���L�}nPլ��ɵ>d 4���_8����b;(v�@{�Fp�&�À���u-�Hd۔n�N�"�͚$u�\�p�G�r{�>�y�;us#k�"��&�ʞ��/]��`.V��@%{u��1�@IV~0zc2�{Jq��+������e升v���U�;��?�D�E<A^��E-U��5S��"�������0iޜ[��4R���2�
Vv��#�'%]0�'�ޏ��}EΪU�y�p�&0|����q�
ޘ���-����?��� e�a�B8�<s�ysIb%�^�Ӂ`�ؚ��g\��U~;~Y2-L��D�Uʨ�nØ^�E�n�^�yV]�vdW�y2��(�bL5���t1�ۊ����d�1��ݝ�E�3��7-ߊ��� =��#P��q�=���|�<�w1V1Җ��$�;su[ 8�O���zFX�|c�	Mt��;�Ż6A��� �Q����@)��f�Q%H�m���A�ı����C$�� $�O��,X�;H��{G��AmI���=1'c�`,�'$k���vi!�m�\�?�Op�%�c/�gU�}��pN(��/ϰ��Ꙉj̩�@���_0�XKD��,���l��x�q�l`�|O"��@�ы|`�7pK�X��,���69���o��G�@���.����*{"�JgX�g�r4riy�l1�
�U�(%�{+\���n'l�\lS�� �=�j5L%���H�1�u+���m�v�z�}�J��e�A��QL�fJu����|�
�������v��j�����<�b,��+�h��0"�yp*�����ũ_k�-\in�c�3�=Y�9�� �Oȇf�4���4��4/&ǎ����؟FnA�.0�O3}=�y�*��xZ�2w�8�{/��|@8	(�6�Γ@��`��A>�4i,6Ή���!�/�9aF�:Ճ!%��Y�uƗ��� ��hZ�V:	��$q��ec.��mzX��vҹ�BJ�������>�&�~��/=p�k��e�Y����>�Y"U�(/���z�
��sS��An
\��1�:�* /,0
7���f͊�;?Ty*`23�������bڥ�w�Z:�~����˘��I�i��-�FY�rU���'�=X��l3�$ן�m,�F��@(}�.�A�7�������I�Oԅ	T�B�V��������+C�;R>��V��TN{���[��p#xY�c�{Z��-����N蘺i�(��I�B���k��2�<�#�7���w��
��n�B��<�v^�!�*S�>;���^��,�/����)零=���)R������P)�/!��M.��������$fE�1���P������<��B�L�ξI����[��Ƕ�E}��"�_�Yc�����δv(�p,n��vH��{b��[*�V42�rcL��\3;G�NPXI���=�bCc*x��XTXI�WO�4��b;�y7"���5R���wm���%��e���ۨyr���`�{��u`�Z���{�.�}�LQ�Tk���l�i��|~�� �{�^1 ��g�l� M`6}�09i��d�؄k�FZ%s�Ln�W�Y�`<o�������d�"��0:�ԣ��g��
����S�\(�E� $�ۄb7 /��ќ�л!��3G�j��9�\y1�!�?��er��$� ���"��"dC�:
 g)¸7������F>F+�k.=F����`-zu �-�+ysJ3�����=�D�"`u�L�8�'�5�$< ����+X���ֽ����l�L�Ǔ%�I�?��崏즗���W�W��9ל�v�#����g�9cDB)'�w]�0F#	�(�S�a�^�0�ΘE�,bO�rjU7�_���I��Zx�N��`�l�&H춶�1;f���?o���� �6LE���$P7���%�{�C�!�rI�:���rn	֍��`89�+���]��{L��Z�V�>ek�b�F��o5����K�@�t.�u�y`�.�:�޲��� J3��$����?QP��S�����"����.��sa��5�p�@��?�`5L�c��#�
���ϛN��o�3�����|.,>u�H�2>X`��X�1�o�8`S=�R"��;1��#5_��{��ow!�FBJ�2V�v��`���g�`+0(;���˼�6��^��{��XY�ç&�4M����B)8���j�#;�O�{�����Q���f̓P���baJ�4���?���(�k �ݣ�vJ���gO)|��d�d�: �Q��My8��VC�)U0���0CL ��.L2��+9��(S>�T���КC�)�ZY5�a�FXP̎蠇��**�P.�E�
�:�G������u.D-iyT0�v?d ~��:�J~�K���=�]�3u`��Й�G�}�V;������l�oĆ�tx�#z���H #f�+QP����9}_z,&��5���H��~��=�ɕ��@�����ћ���7���F��m��Oі�Id4���®��<����{pZFʒZ3���"�w\C�+5pz�+y�+O��j���iHmO��Ҥ<<&�c= ��{���{��x����K��P��� ���Jm{��}v^�fKC�8މ��2`dRr�M��T'x}e$�����d��<��4��H�ݼY�o\[��c�@vk��Rg)M��zA���B���ZO�Ѱ�h~�"��WBJ�R����q��C�L�pO9je����p;JH=c�;/p�UA,bk\�ɍ)�u�|���!���d���v��O�M���D|�e���Zq��.�	z�1z�OZ%t�c�=�y��t�x\�mfz8)�?y`��MB��٬>V=��M�!9��P���'By}f�b��ё9g�
7;8�� kb|4�R�jpx'eT�vJ�6��s@m�iJ�I���7��̞�[��9�5��Ώ����5=��嬹*l�')yqn��1L,�=mWKK�;Xf��9U�}�X)��/!���
�&�=�.�7|r ٽ;��6>IɄ���'���4�a����pK��x ܫKPR�[x�{ז����X���j�8�q{ݫ�p�7g2(E��U���z�G��/l��'5�w��3��ޥ�*��Z�id6]�j��5��_�%�K?S��dp�����^"�KdH���\�;?6���}x�c�3������W�w*~��y�F�Š�ϛYk�ۭ�o&���n�A���w7-ƽ��h��]r�0�W�ُ'�Hk�sٵ�#�{�;mP�`�`?I��O�>�fiW�g@Wr5%�8�S?x��N7On ���V�F I��A\���x契F���=in�cz�o��[�tnJ�,�I����%���m�)&��J�\�RUX�E�V�W_�Z��G4��[�i!D��/��N,�.�� z��o^	=�KY�g��D7�����oy�&7*���K�/
����`U��9���w�f�m	�A?]�s�AQ \���%���*"���#�[�P���]����]�b�տ�]���ŕ��Yn���(u�z Ȅ�cxe�y�[���-�u5+�
m��G�I�)@�hr�Z3"���m������_L��\I�mr��>�6O[>�N1��JjL	���&a]I�7�{+�J��(�$�DDy��Z���t���{�aنE.8%�ݞ+��,p�("Ez����@1��ᩞ�p�-�Q��Ў1V��1׀�B����ꂉ�p�� ��;�qf�k����y�S�jO�&�o&���Ӻ�X����d���8xPN��P^H�߈צvD�Dr����2T�&�������>��N�$4#�y�!���m>�]l�8:�>�T��.��/������t��%�RN�
�x�UQ"�/�r��	���ڳ��{�J3��b�3��| ���F�_��Lva�@Lw5o�=��=���]�a��U���Ң,��¤�/g���"+o<Y��ƪ"io�����<Oi��ի�@�V1cƽ���tR*�xsf<ہ�$���ڨ�f�j��?/����Ƣ#�� s����`���g�M����R�����Ǐn&�Nt�.Wk��1A�W���R���[�$���q�D���,�&a��o�;z��f"�1�F��_6�F�1��Hv�7&l�u�-���Q�\�P��:����(�wqIk�(X�O�=c�=r e����s��h��{r`+W�v:����;�A@�����Y��<�L�K]D���A+� X��^'/�Ŋ:�'k�瓽��Gx�iL�_e��,����{얗j�
GP��`�Nֺ��;i����a?H�7n#u������dx��C?�g܁��w0r1]Q� �o;�6�Lq�i���S��\�L�D^`I�?E�
�n�U��!�PY`^�������1�%�d�'#�@����S��F��^y�����G�#�z���I��c��� h�ԟ�k��.:`-#��d�1���Άnt�|�T����9kŃ�-N�t�ؔ�I�?u&r�K�'
�����W4�D�1�5ЋV#0_#H����;�G�X��v�}l0M��#���l9B��pTl��J�g}������$`��]:X̨�5g-���z!�)fb2��;h-��z-1�&��y.�����u҅��1+UnRznő_��X�(*�p�u�l�sQ�,D1k3�Y,��gz�±y��8rgh|��vc�݈�v�+R��4[���8����("(����
���^�m�A�ǖ�m��Ж�뛙�n+?i��-)M?7�^��VȔq���ne����[R'β�/���O�~(�7M�<��X�z��P��j��|�8w�Cv��:b�%W��$y�+�0ڽfeq�L�Y�Z�ہj�|�����vd�Q�[fgZx[h�Њ���Ȕ�O͈KA0��u�-�臐�ʲ��OO:�P×�x'�i4E�Z�(y�s��4 K̻_9�6]iqu��k�X���h�0�?�UF+H׶y"�d��V��^qy1;���=({�f�8�U�t^n7>K��~ő��R�>3�?JA�ꗅ@���,Lfƛ3���a�C�Ji�uB��CA̥HL��TR����J���0&�&���M�c��@��%O�+��|�����j����X�h$)O�2[� ,�Z<���Ϧ�-& I���4�Z��$p�FQ��e����7���X���e!���������ȩh=�T<�z�g �����=��L���k׊C%�.��~��5���O3x>���v�Z�T��'�[e�6���U��������ՅQ����J�pS@إ.$G%�>ni�5 m���0c1e�*:�Ү���b���q�t\^u)c��i�r^��Q�Z�뀩�t���,#���Q����Y�\��#P-:��n�fD�}��Vq�g�L���b�N ��	<��KX��ꊃhY(P��vu�`�:T��%VC�3���h��?W ��X���}<S"�h�1�n�?�q��W=ԧ|�P�A�����jTC&�ONAOŝ~Ih >�������4�
�ᆈ�F�WǍ�R3m�a�T�<F]j�[����hK}�@�M_K��g���t�U�)r8��mU]t0K+�G9�ߣ�{�R;h�e8��[�hi�t����	ё%R�ؕK;kSr�Œ�����Z�d�ܰD��l�	�_0��)/�|x-	<&���'�@V�G�6�/9H��@���y�idK�`<��R]�D��/`���>�]�'ZdD��(V�$�$Uw�#�0��f,��b��e���R�?|]�&�W�����CF�~kle���e0^>-�*U0R숥CuL���u�y�7"i�Ş_箻c8���W^D�M�����F��FT(�`Ҧ�uy���e��DJ:5W��ד��u����I�L��k����:g{u��͘>S��E���I�,�/�s�������flê���:�߁0�T��b�O+�+
}�㡵~�9�����L���ѯ�G����ax/.s�](OcIw|Q��'�<Y���	e_l>='���7#V/�m���}W�ӿ�&H��Z�nO�\�K�~�4����fo`��?���h7���;1��-�a�Ϗr߯��O�99��ޮR��Ǝ'&����v�h��R����H#nИ���&���a�%�G ��/i��j����߉��48��(�K��BԎB����N*Kn����aֵ�'!㫘6r[�'Ks��/9����Xi0����� ���*�+���!j��v�Y(�ZC}�fn���_��M�O[��D����臅�_�jPߛ�Gx�]dn�%f�V[c�puA��:(Հ�m����e��\Asu�k=	�';�^�: ]��t�@��eD�Z�+�|�f�7�E�Oz%�Aݷ/I׋���ؤ�Zˢ���-��L��H�z��]�����ɴ-��0T�]�����&�i�}�5.at�C!��%�%s�{�Áz����8%�%䄳�=V34�������(U�|�`��\+�2����Ya�-�_l��xl<
�>m*¾n��Z�N6�)�M�|���FN��zTE3݊Ï�8�D���6�˲1�`~ _��#߼��U�����c�����"�����\�Š2�j=n?,�n?�·Ɍ�sd�_m�òK��66+&$�eh���Ը�8��!(�W])긚���8�]O)�}��?�5	u�*t�((e��#	R�X��h��l/=}�plcX��G��A4-+�et�ë�W��-��� �ܚ'f!R��t�v�@����J������t���SE����av	J��o��&z���j=+W��kp��t�M1s)�kX��R�?!�!���Jph�Ɂ���&�GSt��T�Q����NW�Q\�����UKc:G�����"v��AOj�ȱ��k?�D~ ʽ y�gu�R�MV��%V�D��O��*i��+��L)���}�ϛM�A��[�䬓��e��N�Oi��X"����7K���V~���q�����j�!��L���˰���0 �EZH�Um�9��D���!�!�q�mf�"�;�e!K��ŪZx���o��0����.�V�[XIw��H��Y�	�9��}�c��:*&�"ŝ�G�~�a�z1}�g��@l�V���8��J�Oϊg%i(Y� ��8ש��W�Ȧ%�a�W*��J���6o�S��Έn�i�H�NF`�m��n���R�S��؀�+��&�k0,Ͽ�����eS����.�������8 ]b�h�=���g�5'�6HB�ڠ���fͻ���6#�Ҍ$�TK�d����ۥ��s�2����ۡV�u\��v��ah���K�s���A������_L���!Oi���N�9F���m��Y�̿aԹkq4!�ک����,�6CY渡S���K�V^zs��8�&O�5�0�� &�.��I� �� ����xa���E�"��4�D�l8BC��
L�:达�v�Y&mQ�2���ҕ/ؤ��9X����� `iA���_Ͼ|�}�����& (�<���!V�AS���n���#�u�_'���@��Ռ����N!(Z.���aC�[g0�^?�'(���e���E_�G-�'7}Y���h{��J-bU.7j=���>2	x�u������aP��Q6	�6˖��o�u~��0��>�Z���*���_ oX��X,�E�:7��ߘ����Dj:��)�Ҏ4D���o�@�gm8uY¿�H$��C�]7>9�>�dd/k���iCK��"�R�,/_u~��:�˥l+cA���s�D������IM�_R���X:+['������	M4I/"'�s��V�7z����ͽ�c5��q�T� ��?�9��Q��2�.�*���˦_���"��\Ec���r<Xa=B����x%s3��hu%Sǀȭ��x�D.L,}[fzJ+	�M��mxsk��)K�W[�\���]���0(�?�Ŋ���_a�'M2��u囑�і�_�jC$6��]��~�Z�L�:Z�RuBU�$nd2�n)j3�.Uo�����|�*}��,��זV�|q'
Ju�lj���aM�8�3�)G�����N�<�R�!b�����5�C\���c�@���ӌc��c�g�8w��y�1!d�>�B�(\�Y;�<s�J��~�RÒ��M�߬H�@�["�}�����VM���Ȁn�J%�2,�P��p��ä ꎨ$�`B�$��%U�61�Ae�$��v����Zr���H�x4��/{};��M�՟����;�xXb�]XL]���m����۔Q:�3Y7�i�MWx�ؗ�5�����+B�b��3?"��?�S���{'��n1������8Z�2���d�����[�{7і���|:�����N /�߈����T<��\�24�o�G��m|�@�?F���~NmaI��YbmC�R�m��}r?-J0���!,���<��cvle�v\�y{<'ğ��o�I��K�	|���=h�����J%ZՑt�����Ý��QC6�+��K��,.�Z줖��-�^�u~���s����D`;��.0x�
j{H�G�u�,3x���Ǎ����޸�
�7lZ������>P�3q������#���av2��0{r�3��{�Cޫ�Wc���W���#4r4<ٺk��Ɉ�fC
@ϾZ��N�e%b���Wa����^�D��L��6���/%�%j[s�1d�56���6��L���������o�{�ꛠ�SA*���sK�����+�����4p@�ߠ�p�H�-��y�����T:�Dn��Z*
���?l�}�J�	���^~6-�O�j��7�<y�xw	�̔�UR��BէR�DyvC�n���
��D7 cf��+�X�k�v�f!<����XA��� ��4�<��˴���ĉ�V~���E�s��{�L��Ƅd��3���6o��ڦv����җ)�0����ac�1}]C/�o��ߪJ�D�7�7J����?�_+�h��Xn����K7����G�����=��kp�}�/�*#|)B=����sB����k�>;��-�J�� #7����z�F��x�1a�i�:���6��q�`�1��謭v#�;�c���������
�<}�B�u6spY�n��*FQ��}����-G�_�������Z��z��{D�;�9.���Y	�Q������~,�r��kD�p�7c��b�}	�s� �C���-!N���1�Y�R����c���'� %����'��.u�n�*�\IԮNH�,'�<?�c��	��.����>���Gc/y��S��$E�N�p�Q���F��i,�?�ſU��p�z���x9����{�B������| �[J	��?	���`H�$Ζ�L��E�.�L��vb���r������'�i�o��Qd]��~12��?zٛS�����&�' A>��R%�
�h�b|�N�q��pΈ5�*%��2�&���#
B��-!�X�X��߮p��钰�ȥ�ts�\�����+N����!X�8ONr8/�Qp�����q��q60л< �4�a����9������u�eb�����_i��/����k�[���n��ti$�'�h/M,H�"]�����R�{4���P7�ͷT@�z��P��y⛄��K���`kWd��P�!�b� t�}���",��ْ+3��ܕ.�65W�q.�Hg��O�q�_;���s�	�\Z��u""d����+VRUĒWY��ME�d��oxH)�J��P�|w��3W�h��0�����H��l~�+�6:�:�c&A�s�@����;�+o�bh��	)�͂$��-;����6�p���)���0>��K�驯/�SRg�vR\���h#>o��}c�ܒ��3�����w_U�����3�0��#n<Ii�5J��_�A7SHe�&�>zZ�"�B���n�+�vݜ��{!�`��T� �;{_9���D�y��4��'IZpػ�F���1U�:· �]�#]��8���.�Bc�X��$�Џ��>����z��:�.&���F#?�l3����J�RF��vݎ}Pi�M�;�y=,[��v[��t�9G��nm%5Ȼ\;9''��F�ƾt��`:���j���Y踥?[5�k�t��L�S��f8�ݿ]Z~�����RhN	�����nr�[����r+U��B` ^x��V�6���mA���l�^Q�	��>U'/k��XCtN\��␨�v!o��'+�p1�Mԝ���f�������p�La��o��]3�x��TZ[p�?�|�(k�+-���9�)#۸��6@Ȑ�ş��Lj��<���S(��dT+�Ն`(��G�#C��5l�L;���[���#C�MCb��Lڝ'da&?%�^[Q��i�5��/r,~�