// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
gCLm1SdMHFBh9kWHj1Tyh9pqSLrrKlXIai70o45j0Do9EviCGCN6YhillV02L/9MxMuZtbXkshTM
oSC2cEws7voEdiVPUhyB+XWj0XNsWGl9lbUqAZHd5g+76knpRT6TsWkn3VYcg2J+bbV1EsuYzeI3
2Grfg0pN4/7/4FaS4DRzPZRFFsD0KMlg8uDS9sGlFhBJSRD+nZ8G4RExFwfzQ7g2CkSkMIsNHjEx
KUcg3RYMJDkVWpywfgISXpR7pgN+rH+z7TsSTWFN2VVOL51ceDPxY3s780PRFyZzFqJTeGXVcdsy
YWoAFofIA6riHcDwHAdS0Ohg015W+pT2VB/DvQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
OKMXDZL89GEGD23g3vBWT3XgmJm6KKtcGCvI8BWV+LCBsc+XlUBQdolKGChmAmnpLuCzAoDg4aNc
6dYjgNsIhgP9LgYog76o+JkxGox2PasNa0kTxREaeboS3ILB0kznROjCnw+ZWzWGfI7Axol0+yO8
mEjNdhcnYP9vO6FSiLWBcGtC/VEW0Rd3OT2YkldQctv+8PmpdKuW0S/vjbtveLwwK84+z7u3kNes
yuGrLAnDoX1YBOQHKw+RJxQfIW/b4/1rofzJ4ehutYYdhBQoOdZ+Z/jILilkgi2qrWQcr7jS2hc5
cHYeRP3a0oVmLXhQ1Qy/aRITTXpxCWwVqHL43H0cYwtoHgZJ1K8mG9jhve2B8x9eyhvPvJfst865
76s5ZyWCTdAmQSTywJ7Jxsr9LKcaRk7NsJjoJAJjmiqn4bSfLe3GlRbfwBpFXsNM56zKwx00bSCK
Uu/bpwqyZ9gMWtu7O7sVwpxMrzPCSKRQCq/ko58LKlXwXNMsD8+w1H4k0WPvrWTPwpJpW8oAdxWa
/8JxToU/wBwINjhy31JPk7QcYk6zYyaEBELmO8L0IZfUFSx3mzVCHRGG5+EsvZQ2IEMu0kSGBpFY
sy2QvHrhfh1yx+7g0eyMAh/ocTQhWsPkSJ4I14oXEOJQa4agOvZG5tKf8MmZbo/sanLZIrnzolpY
RH/g09PVswjWWs+W32X6I9SRpq9uHX4+DMtpRBtw4rx8CKMS9/0bTM2qFXIHKhbvnKQmaNaXn4qa
6njElSx6UduVrOKygCs3eyRR2JptVc1YN6WTSmdGQIB2Xw3do23BOCZ6Dg+bU9HA4+BmLIlzMle3
S6MAPumjwu+kuczOzFeAm0IcfFQ7VQHk4q+9G7C3yM0mJmaoS+JnVA7yQ0wUtY2vVc4c2+HQDI99
wOqBzV7YV7XJI2pxUu/lN04Igd3JMNFur+h9/tRUZwDXp7+JHplU1VSQhhn8JDUrqhX40idz/Yve
62EDZLRFM+deJcvyE4c1eXXpaHLBkAhy0BjBR7MaBck7ZRhEhyKlS0N6YH6mfO+N+6a1gQ+vDnbR
VQfdToQfuTyk+tSmv5BLGY9xQuhdAW7peMws8cmpmLoEomk2DvgyY26UGXZdJdolL8CtbY7hf25y
uoT+GRRjyV3krj190gSB/ZEClJwwozt2P//lCinux4eq50+2U0EUto0F6IQmVAbLu17rAhGTditX
0Jn5UEFZfVV27FDLgfq9ggR4N5NRvAweShF0pQcEl65Ohvlp7xCn19CN7B7VeGn8dZ6tFR/qI0FM
Hcz8EL6/vqiO/bBVvynsA7Bp5N4dO8kokOmQ95YoNAF8uhHoTEQsvki4xw6KFE2pydGgTEGrzttH
QAqg2bKfPKK2JjU2SNx21Ce88jocMR86iXRH9uWD5vs6aHoSxD+GIf8ix/0kxxSsCqUFmyy2IChZ
Ifhs/p81X17Gx1FLWy416Whp3bwjRH1w1nT77DoSQIkbUJfVf2MgvJSc4qCBwdn/K56+VKKDe+VW
5DDTFxVi5LQ/bCya2W8fGMg3/u9bX6fm664Wpe5o8Tegk0m46zLxZL1HjwlRg6iuDD0QwfKUaGRs
/JwbwRYeVX1D8ydJpssIv429QOLowuqWXaB3raCRMo2LXu/lALV141fIkuvs0qdKDrYe43B8xvR/
wD8KLPjArxerk9qqIHYlA5c2vdxdOhb8/wE8FvF3cQ88r85/AJq4yua1n7HlmRuAD77MAbZzIeCd
ctOfTRSKICUmGQ+HrZPqxWo48nMbRrkoDkmz6iFUpWERHYQmIqgnWS3DvRxb2ucUsR+bqfQo/E6Y
0+G6gWgYgjRToK79oy8/Bv4QSryQlUXN4/vC8vbmFg3frEFBibcv/8/fzbm4Cg8cnaJo5SXB60RS
HQWcV6rNAVFM+S1XKkBf3gx8N8TRBMO8QhR0YVDHx0vi7XA/PPDEkQoGSsAn5DkTagnDm2Ewsny0
w/79jQHmxFzZoYEs5OlhfjeLFefxlJxdtqvXEN5azhuq1MtIOqwSMC8WJu+WHi9bR7zRkizhyg9e
gkzuZl9A2lVXJ3HSKx4il+SaR7wYsl5/aU6O1nVz0PxA2Iqs8g8ygFSg0r4nuCt7bAx3Xuoh/85y
IhNkWpaR7L2oXgchdpMf4Ral7yDyUYssRDyuNFHJWF6ftZdnxzKiQEIPIoXPGPJ5fHyKiqsYCX4G
DtZh3kf6XbCDlU48kRf0oS+UU+XrXsPEqsoLWFdU1FuxiLyxBiH5g+yk1L/+PugR3lPy9PY3vVKU
lsYBuWCZOF9VjQ63U4HWX28/Rx9n1JZJV4sdRhXZ3PYhh5FzpI8A2gOVa4byz6JiDp1QCrM/1uOH
atZtvfjTNj7C2a6fgt7Ptd8ytXvHcEkK3nPQA8D3Nlk4koW1iapmiquV2IB0ki9UMapBUneD1JfS
Tb7VmbQR49Q7uz3JUZ7A0tub/u45cAJEhmdF9/VMkWfEJXd9anf2czrqp93Vmbt95I68wXTZX2BS
gQNs9tZumJxdp0a1EmniPIjSgMtwnf0LYZ04sPK/sbeNOPRwqmjzf22UEQ4RBK5//6CugYVh6JEb
fmxx+UTqFWqa8WswrXKaBWXJcZIL4JOf3y37UBseVUVKziK20zYidQlMgYhrJLH0gQHfP3C2iQD2
xwfjVyhlQTEu2sUa6ratuMvwcmsiYu3MNLFaVShhjMR+uTCNY/csdpgaG2KBQTUh/GC6MEWkL9Lm
o0w7lohZE3OfCQqP3s4NpfZJyMQm4ZwDrIJB3BK3pOhZaWOYPd4PgzsOX9gl+QBSDLdwEZikSAKr
V5G0ZIp4SVyRg94IJYBYlbFncebq3aT3QoFnUWQ0DMcfDVPP0T1lL8/+0tHQUWjJ1kQcYxx216EN
IR8RtrPO+/OZvvRW4E0ITB/IbEokYzxeQqkhWaM2sQ/4FBrodZK86Na5y91ZzNz+HC0e2elFR57U
z+21DLVV/PpUyHplcjN+mlwOwqI4CM61XfdZ6rO4DRYUlKWcrxzE0an3f/tE0eexC/6qfvhasatG
Cca74UQTQqZHA5gRT0oKXLbdVKoQw6QcyUXodM0kIvP7/d7ttwNOTKn1/FhIjyL0oUbL2S0xT0lJ
puwzgfPUCbfjac4TCIrM2fs9pUYh195xMhZLf6vORwvQpE+oCe0EJlPkDwfGEPeicQfmfAmTPPU9
7m9Tn5zy56tekQTr7KPZKv/MrH9jAM3pV3W6Bin28CLNKz+KxHFhNZ9079jBee6UdmLjkw80JRgy
captb3vBir3aryFPKYAfSc/Fm2TUjpxug6sOYtgY9JiMAVxKtds1ug6QTJiFX42gwfXo8B9hrhBa
cu0LODwThNatfpFr09JMho1U+7q8duw5UbL7XnW0qJ+cHdow0Lr8TMXGb+8fxQnvF+aANtGC/jxc
kdUvs7yTHKsBOmXCz5fs5MGt0T4d+eM1FklsemeE1sSudkSrNM5AcqhHxRbL1wMOvomXW8cd+1pv
A30itUlTH9HdA73Uzjo3oBw+tqjRi9wI8IHsg5WmSdVRplJohHX+9xPKkfNU6E98O5mLDEHRWQct
cI+HhgHFlrjcClUrWzHg9/CLBIaYnelfEy8H817013C+ZG9lxujNlSF6zDngi3DO2ZPwmvd2uRfk
yjRciXazHaEXUO1rmkgsbxwqiU82QsrXqdx4kD65Hk2jCsKJaFJI/HnAtzJIhlQ8cfqsJE3olcjT
BwGWQOIXCTClWcg3ZsVZLUxUxeuTQ3FaNAKQeYinT9fXGlrKBK/kco7khR4jXbgeKo/uCvbOohz4
2wl61z9yJ3ys5MEO9/ScyOVdYo+FCkyelnr8BNVMuoGDNMOTYDzvKZp6vmhm2v6NmfkqG+ZjE7OC
ag63VQR4bQXWKOp97IbZveGFrm7Fe4V633OkGgIys5/nlbQqSFHVyUB1OEM3nFfoKpXwxzvRFE+L
Oh51kk7xfmac723HRt6lDw6zpMJwRBTlGeo6fsyTcC/fvYy5GRulGaLNPBs5TFYvKSrd0o5SOMci
zFnOz4BgBsSUiF3IAJ52vhADAIy57XWBHRaHPHhpLbO0OdX4dQTkPnJVS9HBFkI4As2DA1AnO9YI
PQA/uGaKzZZRIa8eq+f25v+Oxbf4h3nxSMt2YCSliBS+aswkFc8jWgMEaKzyma0Sm8j5G0JFEQNE
EOs6yhAh6fvGa+x4zYKlhIVBk0+2hmvUZZvZt31mP06mvYUzhh9r+/oBnI1s1uHwotlu+Wwh9HHv
kb4B+tg4DIlaTHIbV5BbnLOyN+oXJlqcT18njUIQEF8GJDRFpSR+LetBtl/Z+GxC7keykzsKyFoU
G7UVEXPVTCnkn7jy1LNDjMJ7BAmdbmnD4f+akPYORcUIYnA1xj2u6pq8ws7T5JvYqfZ8buXAIlnP
R9tgSd0T4J0L23kEGttZ+MADB8Aw4eLK8hnro0XxsiJ3Huc+kPC4aWCpc0k8M7ijGjdaJdLGDCl6
0gJHEPIus3jW42q6kgcWHffF4THODAZTbg3eCyVOEkEuivAExuJnQ9VKKN5jHyWWLjp52munlUj7
eE41HWPMoBcv2/UH2MsiwuQBwdCiLxs1wxX1BTZ4TA9NUsjvu3TSG3sc8vZQu5K9CTBKt6eHrp/9
D4l8jCJZ5csplqZQEzJDRYNAgCspEcCbodnbvfUSViet9EbkvLOCdHJK4pDhnaCcA09mGDlVJ8Mi
x2Ux7GvEO54BaTQH6cDptMAZadrkiKzJ8v+kSOQXpJijj9H0ct2rbzLTbD7J5rh4Ip6D+chpLJU+
x7cvJ4F/JcUO3V4TVLhUSFU5fyXH4EcvIotMADDIxLC18aJojLtoUyzkMtsHomyZwzIK2bLv8dhV
ty6fPwkJ9Zn/lsRDTeJs5UuJVFgPrvOnTTUMRaKpGcDIyUpTlFXdW+DlILOeM8YhD+3vasIn7wcM
xW7AJZuLx2VohEGLIr569JTtUO6WweKPeZiGSc8aXPnXi51bQpA197ifrLbnsYoIJAe6lYYSZdhQ
3zk6IVdkirQpTKEk85ghY2VPAof6NFwA2WUR843yy/r+9w4ef2tJWBKT5JqDkKzWxKFpqDkrNo+x
0o36hnu2/WoH0ZbIrLUhtJa49tetIcuHXuYle2FksGXm0Bn4twZy99bwy1LBZU5+NGuq8gYCn2Df
zaP6bJoUOG3G2wjTX1Q0CnhthWVkXEXgK7I1RS6GUPf4GetN1hpErVX+4LihXYO4/s8OtIQ84bc6
L9CHoedL9MlzKa/wWthJX+OCFir1HGxdgUKrHKokPFUII5igYkEgUNN7vFiF4AT7GvNKb9GFlo5w
i9pObE5Z4Fz6Y85qdC1Ekv0rIEnr6RvCAaBvX36EfIb7JCbObZKfXuqAougP+qB0cUEu0zfl0SFQ
xUNo6EX+Wx6OrryYS3stn36bxLBfTSBdzhJ7Hm3//Zf+GYey0OsK9iW/W5kPdM0I3BinSbXl38Ud
cluj+xVq8EiF4np45jCSKK1Sk1IPtCuKIPD2VAAZ7FYsVyeAsbmtjANA4uLgxK3Oj8jElK5PmBK7
8+QmMFfQ7vIFVQYeWmMeRxejOZ1xMrN6maJuDHuHXEvTgM3YeA0yRXnQ1eAkI9RKwTx71dUCKhC2
fcOQ0tj1QKnmMKuFzzR0LEjaWgHWO2bysbfcTG6WfiD6w/zYwONxfHkueACU8MF7bbUWmwomvzis
LSPivaga2x1ecxILCoP9wLEWg69HQNHoesGBlIrXhIdNHILIVI2YjjvyXclSz4mERQWBfm646Oem
Ils5dCytk0vi0kPNf85wRXBL72jUIOzYpjFd3iOUF8b3ojhElDlXzlqFixcDRKtuR8ahKIlX8v0U
Ll3ff4jSb3dNsxTdeyPzi0JF6P6TUXskaY36QylnEYj3tktL+tJJ6p0e07dR+LEOocU6hQV8TDn2
m+bhJTjQ5tzGuMOFs7aylYwAZGgD8hfqmdfAnlw6DM05Cncvzd8pGgMe3XJyo/JIfXpi1zpZM4uj
LdnvnSoQLRr6SqkIn2B549Qo7SSOHp8eagiCme2oqCO2X+o+hfu7R1wW3N7qvnCQSVTtmFmur3Js
NkB95gB1c4GKJYVAN+2CQ6stkV0AuaFMeNwt7hYjYcu4weFqEvjbeJV6slaA3p2sbna8KZbVVeM1
fAaoQZsJf2ktdmxkJu3wzEPX0XgBjGOnnKXsPOkrX5/13hY2++JIWUkLcwRjV7QYZWgRjDyyVzIw
cr7E+P99IIBqW/kkOn0HcxYgj9z6p/wpUCduFVCNtP9NZWFev5Aa5CpZ6SChvETGIdqSEwKrV8ol
e2gGRiMK3c27TEHgMvOThSkuHoh65ujpwvufcBdqzvlM8DqVgdjI/IyA3UJ+ovFGljlvC2s9REfy
Ub2plzLJ3IJbuS2SDo5hg8RT9Do9TPL8FN379MeP0iSx4ib6y6/O9WkR5A9EuWPIu7nPcoUPckD7
gJgL1UKaOfAy9Qv8bYezgNuee2YKZHFNXsf9DjjI0cwVYdIHTPKi9J7+bPbwsJRdHM7i0CFT3pLa
GHmkOrqmYoxb3gnej/3/lvz5ordIwmXCwpePasBSVIUVgfP0C8ftD3T6CTaYsFOZY0H5ZH8QL1TM
ZFfoyOmvOdmgep/UDvmtofwowc6923q/AkUPAjxl6xtmtsYXWs8TuaH0szn3Kq9kB52JYQ1iUaiy
5NFVZoEz0/h4/IRnEBZYzRao9GmqWz/aSuUT/olFWVUGXHtuOjD/LydCBOW4HQWKNzeaNRUjVFzN
NQrll4FlQPvAL5lp1R7xDMXmQg1AmUdMdXWqH5RxpAKFcuUkXBrLioXJghgb31RtyJlu88gcokNS
cqFFYW9jete+AF1vdMVMGa3g0lljn4EAHUOTQWZQAlHdqQ9+p9dTszv+Pu9EhBekw1ypFhbsZjd6
vb5hgoG4AM29Q0KYqVMtLCWPznSfdRiDNmz8kJ3dTJHiHkOWaGDizvV6m/Yvuc0yYk3YKAGrqPbQ
4Kq9bC+1u9vO3ZXS320bXzVXefNGBpe9z78rZHO4IU4cKlLJBfgYXwtax7jEPjlG4GlYsANhaKew
x+RnkQsn+fYmlFPdHURyTskGLRU2CBdtXVAgjsbzbWdPCN7n7YL2unjDG44Ehu8DwcOtPhw8+SKQ
uAq1NNr4uKf43Lr+oblapb7pbvdnGVEDCrYW0CV8AR40yqRen0np6ZOsh308orqfCD/1IeVoo/I8
/07/xw41jXLwhBhxWAeeIs4mbYAoWCoA79sYRguXKliln8Jj8Sinkmji9eUmT5AwMDbRbNtmqvMZ
4SIVsCCcVOUiBs/rcT8vPFNrWCT5X9LRvaf17NQghG7FWW3/C5+7VP+ZfDW37c+mDTI6GopUxAGT
WVG0XTd3Gng4Kirg17XTh3ZXklRRxjvWwoM6zAThNc7uDchyyK8RB6b/VyZa30yk0Ls8TxKkF0Il
ptoVmQF9uyC0SbGkH5rS3J5EQ3hPkR6cFHLbNCUYBeS+dzqEvwqyhy0IP7GnE4jX7qipFZcDT+Of
BU3MgW4Hsom88ag7j9Bvon88TaOQu88sElsSgSKtE0mnpnnVpTWc6eIOfodEbLworJ3C7CSw+E+f
IyEm8gBZuU3sxdWwtw6c1kEaTv3AH8h7FBCfYogg6gB87w5bEKJvc0KbuZEnlfZJxLuqNzIylp3s
pWZKugzCWVWFZTn5h+y4SbhSxpX4A2HpGgw4RcGMQ/d8K6MgRfNsMW2G0B1adePV3RXwqQSIcFsi
XiH22SLJgLaKEleWoqVB3+rBETiGqm1COWRWQX0YOyrG9OVUXcx2P63LEFCm/1Iw1KiC/lmaNri5
oCQRXJ/QzOnNG/WBllGy0U5PG1i860MRChX0irqSHSIdnv9cTomeqNjpWG+ouMqkqgur0kZwL6z8
TyU/AKlVdfsOc5M+rKLW43u4FzCH8rsYKX2rTm5rhBW++W5xi28aM+Di/lM4KthDtzG0E+aFDaWv
qfaRiFJl5mSyXQ8XenStRfhT9E1ySRVqPF3qZuKsbi/kN/+OfmIm3WJf8j2bVQqyLwMl9xe9pB78
gOltVcb5C8D4RVfXaJNz2o72SUAA0R8vKx5UcET4t2iDBhiHI/faokAR4Gbv0umRExRgQtNj4CMS
t2Gjuo1x4c5gVZz8rpIbS8tyuakiJf3CMgLpCt1XxA9f71Nt2m+O08Gk5rG4wUuYrY3CA/3Va0w5
SAturvWj2NjSJ6TRBneYEIqM/aKKCkpRaALLJd/qR65UdfUSBA3TAJnmURkjQ3Rw2cGqoX9chL5p
VGjmVXZmD7/h7LrIguJ0EyeMuCdVU091V9+ma2+d8cwzm8g5ZgkUUbarFh9HajcEBGWIWKw9Nd2r
StrAHkdvgPBAEwOyVE5JHRF5qPl0xodsULSxGPwrUdjh9s72RKQaBAQBMZ5syszdFKwn3PAqldHo
YsjdedhMX3INrloNvml1pB6idYcQGatV7+IVybTBuYdQaiYUjpr1OkLqOHSofh2pv+B/hQhE12Bn
UVgCTEfsk23Q/N+LxIGz6WRgh/OMrpQzZmfnW8LbMRYulimEZs9/hGCnYem4oVXPZHyJO1AxSd6j
lV2LkqzBb6gvHSOYptaZpl3bjNSvy5EnjVrLgCuFdv/BxvGOWGicCimiwS7Bq1/OH7uk75i02JgE
b6q6Fms1dlwVdlM3zIfy7PxdB2W9nBhSzp4y5eLDQ5TpBn3IrnXSDPNc24MHnRS2wwJeQRGlP3Lz
+KICeT9vvDYAp5Be6/QaQd0HjyUmom73MIcffRLRhfTZHqguQsJzBWE/NO0l0rN+CsdmBTvgiOlb
ijqBQErrnV+S1sIiubNWQRfuwj+MHR3l0FldNlFdiq4sY8y8TqD5IGURoPiRuBlp5e5TqfPxigHJ
4ufxlNE/lBqEbhaU8jNPH8NgN+kouMs40to9FJuY90ExoDbupHLK1lROM1F6ap+4TibsGClR9mis
E3AcwzrzxlsreYuTSnux60JLotqS7b1tLsTqdjEQ/b/WLCLSnGkDVffiiM3xrO0cbzhtjdXjuU1/
2jAUg0NKjITAZahNgxeT1KNregoLm0OcSbFYjaMNtEzZBDI6QJPISY9HM64BIhnJEaHMmhLQ/2v4
vwwMJBrbOf6fDGx4Z8050mHrucMetS/Ni16zLATvR/Ne5IT2jLuav2pf1wAQZKmXYz4GnjvsQ8iY
b1SIGhlYZccknXG3LHY1LG8gVWcXzWfr34yc3814z2pzIX+w5pxaaJNrspjhYwET8TBIpux6ouqq
hjO4KwnAdLRAjzQJCOmz8rzSYjnKrb/b7evbo8AffQtXQxo91U/TJevNLRpe4NUihrELV+bVmPBg
431hm5VRvQo4aEgZR67X2OcwSjhC0fMXStYwIIBg3zwovSThvbXnSZ07xSPIIMHE11jeykXONXK5
0a8KAJgNHT5JZK+S1zTIsGHgImoCcVZPNvQgecNoSranubo1vQY8aQZcctqWQ7rb6yjVJNxani5t
pwL9bmhU/j5l5firWWiOUOIpHUvMkjK8H7Z1Hy5/p308CZSXFHbbHcGJKDlsE+6JJK6n1HFKuVRj
M8/Kgt2KvbZeOKAlLtMezZxTo/fjscHiSPQpFH8MvFvFgDD/C/3F2pJAd2CxhKKiVDIutb5Vie8C
H8DD3bpckKsSYnZ4uxLNv3/zOutOMFJmmwZEgGpk+NcdG0XP/rv2t5e3K0BGR2tMBC8Fm8qMicB0
pwa/DWREEiymJZ8HmDkCB7nLDxE2zh/nfBJlgJbna54001zRkRKdTXefin61Q5VHdE1l8ro/ycvC
TsKjxISFDKkdSRTinHiRvdXfWh/kfS8+lbDjptw2zR0kjUxIvGJuIply4iYO5d0tZ35CmzpC+8rW
iEzw3eqHvji0AkWr7gKh+yqNx0Kt0bpJT/Fbqj9SBsp5nFWQWQtsdKNW2TBkgPZLX4Q54vgSZ1+O
wH9T8fwKmMF/OkeigXoa6lRsbixG0nCX/XEjmYFMjJIlCAw92IFNNPVDjlsQ38ae0Y9zAjXapeI/
+taSn1ekeQyNcdGeBlZBPDTBJkv5jAQRhEOJeA8W9ROw10vpL8xBcjhY1AdzuH6LSvrkCBeAXFY6
na6VKgYuuwOT7e+WSCJwIDniPlE9GvrJgo+aNqH7Fzq5kz2vl/jRn2NG2YmfeYbMXfB9PvZyg9pO
QF2e6R3PoXz3gq91srLFslyJw+jXSdbK4e9lHZXUEg7AtwS/ClA1ptR/Ep9SIlN0/3WIDYIX2Rk6
we1oFDKt6DG75V7wEziON7V8gh6LiRSGH9YVmUc6CjqnNh0wfPEZg/DD4bmX07IZgSJK0wL5K9WN
asYV94uOZMKiM0TXXobQ0JfAFW2nGvS3qczIkF8ucm0qajnnh4v2GPnCy8jiJEcNNhIY8YINWSXP
BZotOgd7VuhXgEb5RRrQCdUemMbe+/b9C62gC1/TSutWf+Powpmc6/DoNH0lkaHYgWfhrGdRP3fY
P3q0C2Oo6NFI1n0SrW7PM+vj1abh16fv9TcGM6rAVfeJ8f0ylrNYCT9P0ayG/DWGwtwu3CpCVYkX
yIwZgti4x32C4+jaBhQDv+UsbDEGJwllZr5kVtDetT7hwlG4D9wiH8Eme7Gfp9l7AxlbMEd5yJi9
yx5qke6FWGvSveg3xYt8Nk9foDmiAnWHtYAigg7NALzLbefhS/VQlTYDaW/l1bHQKEfrRRTCamdV
EPzJqTMpBltvBcW1mro10XpD5Fj7opJ+ecJ+f3B+bcVXKl9ln6dw9wpIkkx8gjJoWYSPIOV06gAF
VEfsPNLCxjcUcgiVbBmDyQt8WIIDRRda+jpKDO8x2ee1WnNHhDR/EReBFx/wZmnBFd0B17N/Q13v
qIwtA5ANBwVxbt2m4k/ymdFha79uXOc2a05tyosXSjwqWFkyREz73iYq66sGYYWXYagHjkZjbypw
k9Otbd+quXKiv1ylgj1A4hsPDw2J20NPROqOeOQdv24DreYEK2yV95FGBYwHCdlIteaDTLrzf43G
FnroDg+SjIEc+HgePNkPC1I8b1c7ZjCfvC2LPF/pDdMyKj+2Fq/JvL6OzzFhafJTH7xytGpeu54Z
o8dAD4O2GQR1wm7bSWxwx094ZWwCM88HI/5FhbhXMkuz73RquKHFa2gc0b7cysILkX+WvTEWzba7
lDtdXBQsi1fqtZ98DRR9JIYVfzScUPFMjlnN3qIt8PApVPwpC6YU5JH3eYcJjmP5zLVZ2F5zvnVl
b7emjWR5eeKekWdhm7e3jkA4CgKnB5szK9mHWHI9PF+urfbDscPUhXdq6UTGsU39swLxLmpgBhsS
dqxBb55GJFKRYzaKV8NKC9Lb2kHfdo1u/rXtLuR6e5X1amyT5mkK+M1aQsTJlEPUD6h+QGVAxtyz
vE1yY66P8xdNyw1EuQupKFct/0Ql3sjaUEyb78PD3Hwf4QpG9ctGcFCkiyy4Nfu8rfrob2wDCljl
nOvoXWuJrFDISNtFYZG4e63HMF9VO2PctPe1WCq6x8cEJzDdc2LioQNVQuBPS8AGSZgFWwTW4ske
j8b8iKNQDNMJqy2tZmHlV8uQcKv9QMMWzUNnX1B13a/i9+STryiS4vIa1RVQCVDEHc3O7x56niht
PV6GIXEYPlW9zGHwB1/JDnvsfazs3mceOJJ466aubx1BRrJ5Cdu6Uah12nKnfptQ3SY3y52385e+
WcP3odstQyzGq1tIWa8SbQMtERORyWx6XRsaaTK2t+qTV/nazGPgYo8krEB6LrVLwUMnmQoxwJxl
zQwsJ/tcMoCud86SdXZxa1gJoKzdxTLbjvSz/c1vScrYriPRVr0yp5s2xbk09wOjjBsGnsJrhbYP
qP6n7T8xQXZAs+LBLS+QAc1gtzyvvw4m01TKdYkIBiGqGEguHRyJOwW646NsxMC8DP3wWGcXyEG6
LbaBKJJSMqaI+lk04ip0R+BhEn52v4S17bZ5v1GOsD8cfZw24x8I2Meh3CMbDmZ6At3Epa/wjb6K
j9+qxILWjK4AP8tUyBK4mCyPhhF/pyEww5sCzXc7b3d7Z3TCyfIsPz+6aCd6g1qa7i6AOC75r9hE
RrMzrsrzdmwhpcDwS7eXXR19BGeSMJrZfjHASGs9ZgwK9WW+0+aIbQ7HEfgnRB5/ymGoAULpFEqE
eGbmeoXqQjIk5E0MTlCGlv7JWW+L+WWQWeek1gOmUd36/BlEHJx16aBDJX3kQf+LJbkz6zvrY150
ze4t3dwydPJasoBvQnAI/haL8kG3VoPDUH/5HaCZhMpoMPkNSDZRZw6SIRkn87f/xRlBuRJ6nNIK
B6l8/IzmlxmQsbwi25/+z9Amhp9ykflaOL3xmI97he2Z46aiQpXncyMpTLKmgV8tqm2fLH+S6Kxt
FWWNSUgQD2y8sxnTJlqhiEy/zNkmM14B7vX0Z5sFhjiGHLYOFx75hsLLrmjMhCUMQIP0GbKeGhMj
6IEQZKxF9o4ENSwTWwwOzv4D3Xx2e/OYWyQohHO+gsTMP1Ne4p8SVcGdYEUl8UYFE0x8m5vegyIm
j+fgXprIVhozlpyEQJ3II4b05k6crJdG+5qFldpmQb0FEP4Ne+6cj8l2DsLXXczfrsvIWFXUFxgu
9aU+fZ1Cttjleyj7tw/tIsXZzV5UpWJVdA6kS8ZYYICgKEH9UOfxleCH2r8VzVc7kPCzRmS+UlUv
u1bqP18bwiWyAcJZo6lqapH6gJ90ZFm2szFw8Up0kjYMwplN085eqXDNppeLbyWzFFqJnD0MeOtk
KPhAto2fqH1sZ3h6ZBcTgAC7CeJv1PrqhpYvKaJ355C6F787HxK7ycbWfzrrsHsEjPLBGbIinRM+
a0KF1NCJycZml00iMT/cupCFsxpsRsbv9gcPfyZ84hPaR1V+AoakzJYa+Nl8wfSWW5PUjvj2nXp1
EknB+ieRZ3yDHaOef3jv14Pzs6HaUh2LYUsNuCzcij33vkq5eQMMwdEXr8EBuMDlq5mlmSKiJiuD
CYscPU/jnf4UKMVgMoASg5juum1VgcVMjHkxzm9WykIMVE6NX3G2fPiAh+fNl5grHhx6B3kagWyL
JCh1jGFlhH2RthOoxpjX25JWDdKR0TVbCgqI7QTcWaZFMeHeh4vHWnT9zn9PQ4COinc5LhIdf39q
57pVhMoAIVMl1Thks1p5TEXk+4JufMTD/Ryy+ZkLPzq+mOLAaFJbTWWt/N5y0uo48kp7mfLbDxdm
W4hNYsviqqwSHebq8RaejuSkVNTDfqzuVAx3bLdBEh0/LB/+xGiPfDA1BM2LbWyWLzInSZ4HjTMO
AVwOX68QbmlYgaqzIm1xE5l/jTKusrhPNtPx/rpPmsqFk4bA8ttmMG+yKxuxvJTBHamQ1ipIhEM6
21RnuR5K42cYb0hgupsE/07IlZmtILF6uJO+vOWFvbRBD9oxWHr3BqGXmCPCOudAilwGBMy3FaB0
SCbSb+rdIIFTv9EooVBdKVDiydxVNvoCdeUDAy02MhXNRxUzV9AL/ynuOetWiS7wq5h4GeuQmrk+
9HyZ0Sw5r8ck8YJjelpecCYlcwDLRGePKJ1kJkqCj5vzUkJBrb7PokFqq9zvyY3QZiTUVE/E24n3
yhGHovsRBfJyhDKdZ9XXSF9IaxY+yFpFi1cDouBqN1HQifXp3lioxkLAOGNT6UsWOzPu4vjZjJHg
VXfWVp1vD0Y2JmUJEgI3cAU4sCokLtdR/wmObCyya57KVvswS2bcZbFs3vTvfW5xXM+LMUiGPOlH
mR+rkceReKVKdRF+oExTctwv2JVtjcBd+LBdjDA0nvxckZ0FaJF5a7gvslUI6lLhCg6bRv1OhRXX
pQKDVYhKGlj1BIXT0Bzal4ZBb7cirMUJPbTdgyuQO9ayAzels+neEvPEoS6sGjH9GIqg4wwlYECZ
P7FR31/a9P41MMzlEXFs66rfxqIhdq3bTC/YwVzS+Dtg7v2C1wWM3JBbCF1ni9k6kCs10RAQ9Duk
2BMUTizQlrvAs7BJSV3CoVY358CdHRqThG01HiADbuRqAhH9Df6CnUPgxo7XwyEKw4zibG5H//O1
2FZJUXu3kCosieRDxkOxq09v95PeYKXpl1lxBGU8otvZMiWZHQlgoOvLIVsK7R4xADrT6vCETDWA
1pJEuW4mhF5/raOzLms2EE5XJ+JVVF2BaShJQIAOaVxlMNUEwNSh6qcdSZlYWHhIcMV9B7Vxoix9
3EBOMeWMJBMlq1NmF4SGeXUHCdAEayypp5BwPqEtS1JBvVrMjjgMutpqecLLEZz+rPpKO43x+4S+
Oz3fVvMCsykFRrC5n+0iPqrAIIYKk3m85jtnZzLzFCcnpilnxEv3Gj1LLh+1ulaPJtqEceXf6HTy
WJqEhxHtj8t6FRnAuWVZttDk5VirqZol9fQ/xhCXsXIjpe45sd9od62T5lieX3hURaahEaKIwHf8
e2meEtA0GiUmpVBsfjfMLLX5fL+R88MzmGSEOGNlPwSAtvLVPI8GUCF38KD64q3Q4MMPf46Li7sD
RbM5c9NuBkwwlD1txeVFWdEuYf3EADNOxMyTLVEjpJE/O0DMlzUmMdjiCaORNyBTwVylQo/wugQm
HJ57wlzpdUKZXS3+gMrnLRiMS6Pi1vQR8b5FuzqLTj/dVMPrWM2itWeWlSynKtBCkvCd2aPdwgn6
FKR01f4XO42tiaWjGGZ9WGlbdO2lz0itpVn1TwSrnLvXkFKZ10p5Z0x7a1izuf5Xmy9YUUN/B8mW
CWnolwFQMK+mDSVTbp9tCijwWR8OkNmsojH0BSVOHQfSpmy0GIBfhN6dZ7XMqp0fkz1Ht0O7S7bf
ux8yItwquuB2D7UT1X5/C/xVOLrsIqLaBkqmEcynz/DyDv+7cR3utOM7vTM0ofNrxQu2wBHOIl4u
TJd6c7BPcc1tmWna565mM8ZqIuVif4tjsubqF3HZ3VlcZe+1C7mBtz9u/ten7X7efqHbhGSvFiPb
pqtQje5rbAwmJLFcluTOXEQ0yN4jX6yB6z6YZfMerATVdR9+eFsRIk0RCO8/StYSotmDMB9cjLyK
0Vu0HaGJ0utspxFrh2Ck8oGl2n7/MwO/7WKJXvNhrntG+Ntd9yfIPNjrVOgIXem7eYAE0gpTtLpf
Z4Q9PYKlu+ul0iZAhoMDOU/PxvBpWMnd62QCpPGz1TSVkhPoEvlfsadB5/r2iZBTTcKLzs+ky/eU
njKlonzR3Yn7jPdarmuSv0HSpvJ1tZR81zWa35xS3Qtrzj11IVfDBmimD71T5XrWvkG+/KUJf06l
96ESQqmVGWi1bM3EqLGZRLClJVo25OSDv6t0/CidJVAMpe3CMSEd7XZdtrULsIl7eMBUeBC6jGX7
XK9AwTKYjOKZfiNlAxRXvcIgIluW/O5oKWx/BG9Q6Rt7uEeYKU6qhTLYRkrXKpd6uBUokoo39Sxt
0In6bIWlD3BvUAOZIK+KNkkdyXUwVZuWMD0PFkD8HcP2wukugX9KNon8Ob2MLO0pc1I9dU69xDOk
J/OJnfkC/k9mEF8YpRg/bk+GKYQUj/gFfYes40/K8A/qPzYXyZlNx1E6q0CKRKxdaiLNVe+hqyF8
TcSO6rlt3J+MErCibCXK0QlKtpoBUCwJ1WN3h5nCnw13OX8gawX0XsWbHsd1i6vW89FQ6D6VpR39
rMeB9ywAH3edSV/QhB6qYttIV/K4qAuawwGmu0jJxpPKtWoLeQ5gzAbj9Q3d429K0NmzdLDZPRW7
aaLPa1/axrjfLEMTpvgXzbLNgQe9afUIcSjzV6CqzjpK5EjvMGUL76Z+a+coBg8iLS5ooBCGzkrl
Ed7fl2r0ucfdN2VlNpHh/Uq8T7tkcHO7IM+RcgMDfKKhTLV2e6zaFRXbA9xg0xMzMbHk5NQCaPP8
35PbEJufSnHG1N8ORyCy9WstEbDtRhD1DSRMNzBkQ+dKAxX2uXAihH1tApU9QRmsvyE2EcfYAHrW
DwW9Dnh5f2OSNsA15y7syxjsl53dJS4qv5/SPAZQeCCILitqyH78oSotEdmb3FI48yDxIVE4Qouu
9tdyW6nK2C2g6AU+ntHXCBfZWMr8mF9d+HD3RiibvNnYGwp+bkzY8JT0wVAoQahSbQLaT4zodIwy
PoabT2/1vBk5n9YbFBYQLm1XQGD0FtXH+KetzygGFtw9kD4EjxXFPJjW9S81pkeSQkZKk225KqrV
O4BGnTXrq/v7roV4JNdRvtTiNOZTcyu8Lay6Gu243BrYGNWrflar8Lc67oVa3ZZGTJlYNWfjSU3W
GLaJC5eWP1+s2/9d07iJ3PQiWiXE/N5b+4LwHcaUx8FqAjKiotpoxx1iqJNcemqNzgIgzteOfCzM
h67suXMDbw4Qfc7yixgEawT+r2wCsUzHHF1sjzBmZlRImWdRG4DO0QcGURS5IcIWuAAH0FjpGuoz
sTp8B7egMjzN1k/qkVI6IHqPg6ElBMvsSnH8xa34Bemyxh5vV3DI9Qp+N2Szs6hy4jdFZmcDUVM+
zYfT0APRM35++VGxzBwVyON9KoNS0xg1Bvbr53nYAEF+4FZb93aJReFgaEjhDND8VAcA2+o5iirc
dQ9kavd957rjuC0/SpSU16QYS5UUbNWEOnmaBfCfm4L/K0ANLu9r6z/bDxf7Ts8Xna2kkDSz5NfY
bP0fguWOTTkY/samDrF5sSUZyjcPuoxuoMjY8EJO68n1EsSY0/4FH3mGiqP9wGnw6iNzNaf2pMM4
BaHif1949ZyzM4g2C6GKAPXBErRIcpbvgO175PIhIy9L9bL8hJqzofgirojI/6ACXEYIMvKHGGB5
VJJRkR0r09JCw0fuF0cba53fnlwQy3A2S/PBef6H7orvETszp5/yku/4BehHWY2OERXfdUrS3F5d
N1oWCvph7dR2fj2Uab3XS5pKEGkp42Kqc5Qsh6+UqSoLxUszzqP+A56ROsLX2uP9W8Q7hrAL/ifb
yaTjqWetgeNMYnS7UZ/zBOpJlFN5r9h34r6AGWGLiq0puTIy4GoTGv34HpNiSBbCtZ6k6wjvnO3s
DhtDMi35MEBqGGXl+moLcFnoGcl4AjQAUgW8kX52qk2kpeXOTqvZ/RAs6int08auJRvVxioHd+Sp
UkA/3QJ+q29HS3wakY3wAH+ao0yezbe7Z5X6H1CeQTFhvV4+UHunk7nZSZdKVT6cBHKmiafiaM8P
q4UVsaGgUwdlwo9BplUukveZ3NdDKQASRvuMpdSFIYsPlU/dqgVfF4+PZ9tx9hn2+aramLttnLNG
xg8GPJVPsA1BJGIu29dG12gEpJvC9TADPsB0jdfi4FZ6roEaFsqNAlFBuNYkLH8v19gyEy6nmHFA
HhxQnNloingz+9wuVT/0neAVu8AbfdZMbItwlyB56umgAzjcrM6Hce7GE8/yUtAJ14fqLsPHt/Oc
aD3Qe1MQ/W4YywRHwpthPG0d4rpDnnVg46BkPSQqm2Mc8or35gxP1BjWSAeU4GMn0QZcdHGRgNV4
Fl6hP8zwD6Ryzt4oWZt6TxL2uiHhpOwr/WGL7TUmfk9wNMDgC8yvftmF2LYR1153DcIRFDj0gkKr
gTOcSAxByDxpJ+ElWEEgRu491NbcUQXOOtyZCntEeZjrrPvD5eq+tZml9GXcIcoD8uIt7anvj9Jd
tYJ0VcJ1nhRperA0pMJyrzVnoobp5GAchRkxSZfJOw2y+ZkX+oiyRoO0fzXxt0s9A8rx6Y0NUWtQ
rdI24+CXC1RyLr1aPz6mVSvnqzaJP+Xe8y4ndO/iR5ulc4RCJLHISmUdJSR1QBc1WtAVH90rk3tB
gX9dbkYe6yK4CMh0KPX6vtulqa+md17beIaITM2nH+wT31JksALRjQ8xL+x4MvonQjEt5q9YvLt7
uiUNeR4uVjN6ZzGfVB1rOOrpJAxJWLayAW4vnyNhF0S5ILoK31gKhaAvF2seb8FNEJTUSzsNZnc+
hxZa+k19+WQtmXVJREor34acgMDXtsugTYb9dQPnP1e7C7c2QpQtTN6YVNDTwMuMkxFGq6J64au0
bHA1SNnMI4WLZ5Rp8LAkeQSvFygvvRLOQLACLmIwNIxbEsKDIvSF9NJor18JA1JcSt8cxLxPOkyv
6x3G526yVC78LrTLxaGTjH86OwKcfcr6TXfm+ujUJfVUDjVds+q5lktQhunsHkc7nf/Ahb5n41qr
dxCuTTFD1+d02Lm88xp8QGOvHmxHTbx6cGdK+QHZB/s+CspsvJkrGqjVaLeik/FjSszN01KQgVF/
/hjZEh8yegR+kBXGoEZe143J9G4odJsHhGiVNZPYHFZt8hC5KZhg+4XHvNbi7hsTnWG64z1+Dq4Q
H4Vu0zPfxHIJgL+tQ61F03KXok4fuTV4U5rSeJwAyaK1BUa6YqdjVV2979Rofrakgy+3GsHCBgGa
D4IbPmOyMRZA8TZgIDp7+x+SXHQSvxXWPov03e3CoKAPj3PocZyL76uCAsFCcpT2pEFjy4/kdwtG
12Cjghqd+vji888TwGS6hTwWwtNIX0dvN45euFGUwDk3r/6ykzY4yuUiXstIsxn5trFaCVb17gLE
JhOjiJuSxm+0II8SRNHQ2yG7TNpujfRrheyxgs1/4U/vR7EpkXkB2yXAPzsxVRnv7kpHm7MRLoMP
jv6OL9A1a1/Xr3JKtZSH+nN4jKqgIvSDEGqS8dEb4J7dlEZgxcBUQBUap1MgTQKCnCnRC321ym92
Mw7E1bUd/kmSlkrXFwcBEZJzh2FUISqWQNTNtKwfT3nguzf7dIhUc42Pzs5Bom9k42nKkAdSl7Nn
BHU+dfdjEWTT3dAelnlXpoqWryVzBpbq/LWbdbDAyZwhqV8raZZGUgIIWXD79ri8iIqXzvEVpHy2
B0gJbV9En3GduKjgutmRriGZVZweo2Bc60SaVNHt1tOYHljAXPnL/esy1hkwhcE4110mk/VATtX8
nyreGOPFnCSzgeEU13fgY7Ndf2eX4pdt4b5UKTrL0m+GEASeNvsJPQUUJwASxkjGmnJkWplxyJB0
axD7uMFL1rg/DymMwU9nkwUBk/kWPcZ1uSU7tVLX44BTammRNMdQNAjprYr0szxIhxNJLrbQLBap
oiGs0339RHRYv9WBqFPNrqmdbmwOERzcI1PG1mHk7bn3Pi52qDkAXVrkdkiw8ajFboACUG1si2Sr
0zkMPMDflejOU87ARtMYp2Ozv7w1iq3akfnE36Ebfsacy+cYHt0+qb3KeUnkIHZQvDByg3SmCmAf
WenmfHprxKndF9qq6NBaeIilijrokR+HeoLdgrAvrEQibWr4i+XACTFlw4cqSbnEIKSzOROGuVl0
So6ul/enPrqE1otJ5wpBH8dsuyUBSEXRfMmxSakAslXCzPrrCtD1R5CN6HLJXmtGYz/1OUY8j0S4
75EXzo524ylDdKc4nSDeFBqh3su+9GIrG6xbfWou7KYq2fDgogyLlEHacrPVLFj8/0014AGAp+DI
+mFVNPn22hgi05XKK5DlwkRwpkWAW4mlHtfwwTOxqwfUdxnzaTR/VZtaWth38enWQRDgJ+ul1NBD
MHAaGcLarsdFQE1xwRsYUV5oHmVvqxnKhxslv5GcQLQ4R3niJQumoTgILwiJQdeXbMfsHJu+XhFm
VWXuJgj0xHVlGwV9jrOKcHAkpOjhf7Tnx0oJdvlfEZpra1oL+FjBu7zdO6SjVLk/O1sjUSRPeIZ3
O81VIG9fGGBdOqGsbZAVAC/OeJGDDCXd3TSMLr6BLEN9k3Vrs/usaMjDrXn27iLt5wEH4z84knnN
yg9VHdzWZyvIB/XpUSUJ4fgcbL9DECOBv2s4oZWksRrsGdM3kw6kIsGbsXJNFl+Co6HjU6Lwuwaf
1mb9eeQCWFu5qQJ7I6NoYVX7MOMWMyJqKhBY99qLECmEZh0RHkQGuglWXpXx/4YKM9KYVZoAIAY7
h+Hdi2zOQ+wnIzYo/4iHWInOjK368nsokNSQ0VGIbxBkhDvccmck5jY3l5g8BRyla/I+iB3nvZI5
hFyMWriq3mAlwqRHsEdLjqIJEnnQR40DJDbjoFOUfniRFRyZE2FhjRaVM2aRN7NyLRmdylfcMGW/
ngIUuajEeK+tucEpbk2IQPgbb2uKMChCo/iTwzTTLBkes1o8brAcsWzctXoja8fFuIpRjgSjgDud
cmCyOg5XehgVEpaZvamuwTpvZ5KhWp677yG98Ga5r1x01wy2IxvwmUJxKpSD7vnbh9xl/ZYNYUVl
Fy8PXbGdZiSbWgEx/mmbQpDXim9poKEoR76Kh4oihJTltW1f4F/dR9lADQMj3Z/KxaUclHyVjT+a
G1TdSp4AJhT7bap6WJgfxGw4kCVIbx3JyzPEkTPMyMcPwLqHgCXrLFpawQ46bM/u+Z4+jIQtN6WJ
LCnPeVyjT0Pq2Q9bnzQMQugpaZTzQFJ11tq7z6PEWsjuUxC+MPDcFa2cJ8EEwMiOTp9uKTiZ/uA8
VJDQu4o8SHnsO/+KkTSsgP4L5Juti6QnI/6BbbRYY99uEyURHezH1+lcWrTKuO75+2t9SyoW09Tn
a3Ztn98TjsawTrUAxKMICRt8u1xx2vDXC2oPI9bOK9AHzyOc7QPYJqVzj6UIahqAU1D+gOh0Z0Lw
APofdLF2z+yI8eZ8xFiTirAVESDpxyNLUKBy7EfoyrUY+yD1ZREHSsjayGrA5eQLHL15Xb2G2rFs
rHKzPWsFvCRtsutMDHqmGi25t83WFIqEOwvRrW2/y1DzNFjAQI17kGuSPIVcDV1G6gH0epa6OegV
5u65rhaHtK3PvfZfV/vdzZmt5Tp77pvpkyd0TuFHXRTJI3kqs2PTOr3UVIqaGYbt3r0gopHe6ZwU
cJLIr5w6ZvAGR9H0Yh4Eu3hzhTb3tk2o6F9/KHy8sN2UOovga98II7XX54lragrsfDH8gQH4XY38
HdBHyTFyOVNo4uQLMerOyCUiedH5Ce1WTPhFfmZuWacFqYpiSI7soj4uaCCwCAVSBH9hByUjY/VA
fKZtZN6Rx6PSGR8vZ2+dedH9RDS3ljRkZdTf8CJs70Z/pAh2874xPS3Vd7dmt5CbbZq4LmmXSlvt
NMhZjTXdssyAsNtgUkRc2FEtBsPU0IP61yN97566814x/vbF9g5JBitT2kKQdKBrE2dxgtG5mwgY
Bfv82cvT7LAEprYIG6GIDbwDOuh/lP/LSsQgrvgOOXqMifKCRESIc8GT+8tjy1jFufNvWti/CVeD
q6YhoLuqE9lJOX4b3BqF8hoDYEu6UUXLoHijatJwrUJeViyP10NbGmKB16Am3VjkV1naHvP4FxJu
VoKT+VA5s9bILUMpJOIeLfJnRGlimNtynPca61pSoUATJ4y67WyQv23Txo7wugj3f7PWANN2UDMQ
FmTwJTZ853zun/8doTtxxD7XUdVH2JVTg7iM4PNCr7dzUDY8fnzHE0ReRE5DLYYAjlHTrLLRm/KU
f18fy4ZuLM/+2/351MmsVUYXgVpyCYxRDcAV7Gbs1HAmHaZl9ohH8aKQX+6i0o/NsuD7NWrvdLsi
Wseb4Ri7T5nNU2CEjLkMzDzG0zaVgsj9TNiN9IbPQSaYKlpu+CrJJik/IQof7W7Ndv1yD5dnFbkt
N8bIfv4xcj3PJwo0BXL6iKV+fvqclOOSYwdf991HL6PiZidqrpYRq3geMdt2EChfduAplw9U9cD5
vxFuHxWodBhDEJQisCpzpom26iftzCHiWGVbiB5agHekg8dECQUSLpRZ93TqnATJ7g5rzAMJTtdi
8QZ2l+jqy1IlxUbQJwnYuKe3v2G4icDRmAOWPGBVYK0XodiEW4jslNx9rT3ygPziqTSccAPG2H0A
bVnFmpg9nCZ0HQp7q6XQp3Uq0fhpy57DHP3PMW6H9+VzPWBsAqcxoARxHDMuHzAUaIsngMNNKHI7
ZsGRDxiWMhmIYFvHPertprG21jBXmKbMsS+RCFVIc53jEkn9u4F5AJSDRG8arEkSoz8cfRiP5YhO
pKAGIXEHIJOCvVNsKQmNpwO42ZamOLQE8tGMtc0Xp4NzK5NpLtowteXWbc0MAmSzzOjHjftJVE6W
+K2tKn5k5MWZ7ImSBvj9BVMgC3QdWY4UkdI0MQDU9+57vK2s5vbSlpa34zijS4prQdtWVCoupDhr
YFHhtCEeYCPmNNNGCqdkVM50ftdVYtUBCZP8yWK4ZwbHI4HWFssSv5CsNs03Ty4tzCBiwOPlLCB2
WMTgNoo1ONbSxDxaV+4S41/0sUceLo+C/LSBJXFQnyh4l6fAvr3J3JUM0WeFg5ji0MCy50x7r0AL
85Mz7V658uYDGl19RLqwF286rGw6LWYEO5FVeUpBd8kIQW1Bv/hjHnFWrzqIQOTUIfbnOOHNpL/O
niiLWtfIwI8UsV0LEZpUac0ilKgOQ2A2yCSyNTNwEvyjoNv7AH+vJsohXH84xVhmt9o7/r2nbxUy
40sS1xsY0ESeaWj7vDQZynGw7UADT6cFtiYhBlUs56ukMf1E+B87rGln48Ib/tKFZG9UHjf3ohUl
Je0XOSKWQvM8f3HkfohXF6AJqgO2q+2mBGeC89byZiGZeGoioC+ymDYk5ql11iaFJbOQhYvUgmTy
A/4dnNG2qADM4N9HsfnnaswKZGOEKhow0PMPa+BG68PQ4fOK6GZW3O0naAs82SuPK85W7phAD0s1
4IWVXZdkcvJ1vpjiLjxjn0Dh849pPcxzHHLD3M7+682DMlPDwJm5dkSnHWw7TtYFd701H3gtD0lj
f7u9PJXXfQZEWVTgt74acLXJl/i3BcdXyyWZZcr0uz5jDuFS01oELsqzCrx7AyeYorhT8FdygZkM
KVqJ/iqmJrOZyDXmt6ua3CUrPf0Y7xLMaq9oINAqaLqMcwJHsg1Mnyenff5dqqYTL0hSJksP8d3p
VvPYxSguGm4bLRgTQdq0dyHaBnOsWqZYrDcIirG2FQIt1El5jRkVW3xTs7mwPluIISvs3Cp6o/nW
jttKZy08RjdiowtPAlFk9f12Q7qAlsn2R1QwDF1brVjRUGMhk1YnziYqboB5C+pBj0+XeTkNXyqb
8sV5x5qvw65wBwSxa0r6rmcGimKPAJdbXIe6fCQ0+obyyjB/VEnCLH1GUuUre04jQVUow/e1lTWt
y5NSiVxUMGrSO+cVyE+4UHiMmOpZ7pxWTsJbN1spirCP4JcGzMrRqwMAd4xKmOMEskfOCzDknYHP
rfJ/G6kjlkqSDArURr4kDFl3JZNk+gU0Q+lojp7ASwef0MoBwkDP+F+yzKFDK99no/gfecPpnyft
BVebzKq/9stP5GW/Z9UDwzEYiIgonNYhb681juivoFKAVF+MAl8KMjs8BBpM76ueImlFZy3pkrIK
PkQXu0mS5+8qSoDEVy2w/QbaXgRoib9Reaarj6a1s2yazD2gFnFia4uCJnXsJm8uawzccp6Ht70Z
hzUE4EhM5X92XAfmxGYvE4CgEcQYVzdHuJxd4hdTg1gpwn1wqF2NuWF8xuR9pW63hpXd6Z+dzakB
8DQl3+utQ96BRuir8fLX/n8gI79NJXd2x2wX246ZojuH0pHr5uJNZy7ZfqMDhW4nyUfVCUwXXYg2
6/VA9jijlx+H35HgP/g/IySYZxlX0nyCyo5y/BcMdP/y8JeI9oNyseU1BfenYxXJdzar1xBCcJd9
ulYanxtbSPhx9WbWCNdiynajl98Bgtrn6HqaNqFpEl3/xKVN5/Tvckz6BknCdO+SM3SZr+VfHq1h
4jqHlfkEragKvSKddrJ3pA5fdxMrSMBKMWZJVDJraVauihXBa7NoSvyTn4uJA+TQLEgzRFY3Vz63
uTEDS2R/pHeygpn6MrdFeQ8Z2aB1xt/4G5hdvwNPbAIni/ukAqd7kmHqlqwhKw+5uFqE3mC73Nle
Ta6PJ3IPC5ykU0BMJ35JN7ipQOzrd7fWhGdOrogdK9Uyxg6kNB18FLQ+5/NOLTPbJLOScQI5RqRN
HoHzUweBCdGd8ooWvzBAIi551FavfWiC5aP1kupdgMv+3aTBAZfTcVdUYZRwemS2Q3utEq1sqO4K
lytUsGqlOI0Jp4vs1U0DjB0V4Q7wQKrpUT66bgRAns19ONYSPthjljnND1ZvF1tDDuUToP1zmytB
dLrsFdjQzwiUlxkcKHRVQKdxNM7HalvHEV0qmFUfrKyK350B17JrSyeorYRLzqPQsCN4Vcme6kuo
CwNZ485WYCiCp7gb2KklSiDgo+fdbmmMw8xxv1wC8QcPvuHJQO5qJPbEZTsrvYPQ9C1CTN4rxxnb
6OpjoeC8C3aziyHncSjnrsGyEX+fiH8sgH9Qqk6Eu0RgUddGwdve/UJEpkMVod3o2CbQVFJ+Ban8
IZBF1GqD19dn2eXZCqGSMklDwsfgRLT1xAaUgopaExvAhPvk5CsiaUecH5qWsrm/qT6imB8v1o9G
idNHM0s6Yd+2kV4E138uhiqaqBU3CVGaoxptR1R0ds5BgJKPnIfA10bRolZNq8KsfcpJXVTqWTbV
WeM1p3kicQWQnhBk71QPKMObp0tV6U4q4XiLA6wexPv3mYzPMuqZXd6fLHBHTVh8ks7ZOB7RKco+
BYZNSH+O3/78CW3x8OP42/EpB59MmbiA5XHx5WTa4RWENGsUsIpmDG1yjW9oOEtqoBBsir63zKwt
tP5/dStQH//nUprwVBqrNgFLSqnxI1hH0QZ0SM61hMuI+NfgO65bClT7ly5EnBtY1t+Hyl6hYt9v
KVwF8ne1xs9J6H5xwMIy2733h7zv4JxlwY91XhyONRWV1s7k1UZ3Bz04W7PF/QDala/f3O9RhSEo
vq0GpdBmBqb3IvUgud0Qyc+2GdaLYBcN6G27fHpoWkrIWH7ZXD2SGC2k6yKBBy+TTumFKRw/er0O
xqk3y/I6+63wm+G9I0NQuRrtzRGJEvLpsrpaoYi06w9hB5U9OJYQqt7iUoxtnKD/wL2hfvlSszAu
bc9iry/PKph9zuW9zCMijzDR8cZuTwPwW/Xb/SGoUrWF7ej7p6UrA5vlIuuybNvK6VFGY83uvSA6
lxs5xAHB83yhsPicTx3Jkdj04ooRxOl7g6vjaXni2c6NUZfVKYAcoh8GD5JQNLy+t9PHY8g4VPwf
uGTo1YDTWKCW7KNzXYLT3LSiAKv+5t5tAdUFJJr8S25qDeWkwo/hy2EMDcYRnKt5gNtuBUaWfvz1
RojOPYEbyrfj5PAQiHrc2KM3HKjvqbM2zRQ0m8AlwiVqo1WeWIJjeEGC9g8oGPVPYSxsEhSLXGJo
l0JuzIwBLybCPTzt6Y98tl9c2DZSwRZZepYeOavOCTpdA/55pURVEryhrPwFZJFpwT8swsX9/buH
kdTGBrBAOoUj+5Akli/T1ST3vqjAWZUytGPWb5bGc8DS0F1vsh5h8aGUW7psu/BH+cG/HQ8fRAYU
c6p9Fw5R1LesDq9gr/MjmNTNaoE4GP8CAfsIRcna/2YWL+IuB0oFJtp+VXh4NCnHokvxkG+VqIE7
NEKNGSzqXDTzxxcvhsHmC+1cI8hNJFt2P57S5RJ4OrEo9I/yelRTgYJpT13q341t9FwSdL1Plr40
hsbCJGAo8OQ3+K4E4XJ6Qa8apokm7rCevtPAFVnUWEdq1ubDW9I5E4UHqNol60qEqlsHthxGIwci
b1kvxaCpgi+Wny7U0RS7dElwx5yjsmEB72PsAUvRsdTS4EUTnl9/e7slOZ96yqYtH5OzPxGAZqIV
HBEDYII4HagSzB9riKVc2GN69kuOak8rVIJE3TGtqjlQ1SbIhsR2gC5KADgKa4YNR0d2KzJvgUdu
1Pn9LzeCk57eZwasvi3JT3Q5V2LCJCNule/EGSff36Jtp+1DTxfvdMd0Wk5/5sLHsRvRX9H2h2Hz
hX10ssYpr2LMJZFEHQuJ2uAz3eMkhFb+O/9jcwNrxiy2EicTa2YzxEomlzHWawct4dupDIs9tMmF
rGtYynHQ86YhMldL7jmxEqSQNcplgXfCY8H+LNVZHgIrUq/u45PMftW/WWb+/yScOmkvMlOdCv1y
hFmmaJii73udlLZWeTg6dYZy8xxmZfMlMIdbgg5RifrqhjD0pppqnS+V6L6V4XD6RT0i+j4MCjoY
nahzq7yYFa5AFCQnUhiUMGT372ZT/83zR6mEM2CmGdk3tOD7wJTt8dsgZAvh8+QFf3Xtb50mzAR4
KYODSQOItMDU2btzTSOcdnbqUTuHg1NCP1NzLtPXDiJWW1tAXTd4QMgditaL1PZdUM/WF4GA/1C3
FjPkQrJ/r+pk5or4XgDzGSyqfwUwFRRikOmTkqBTDzE0vjDXvD5kXOv8VOyg7PibdkiVXym+Kazs
zgcLZjuQu9z78tbq72IulXclzNpvYFAXXzfRzjS8TLSRnNrqoavdwf83NakEeoRQ8knzBpD7mHhg
5aIO0N28isGTJhguNZah/Gt/IIQObKiZNnUt0btUajubsgWMSXZB5NmCdkysgELsZUU8Jz6ikn5b
Rx/5Bpy0PoyzxrA3o22A5voO5D//wo8EuK1pZ80WUF4Cur/mpRJr1swIALn+emFBExSTAtXFYil4
fFvT+SnSjx0sDZzr8xrE58pBsGBrOsenHT9YI/G+QaH/I/0LNisWaT55jDb4w54O4ePfY/ekP1tf
zXSxh5l1ZFNpV+yku0mEM0mTSzu6XGjJnAqv9c3Ddfw/2+zQhUpA+jvm/ypgTkvrmSfdv3I4jNW9
XQOZtOF2ODm5/wnLpfcXTXjKsDcwW5yjweSLZuSLq7afKpXK50gBT4M/x8ME5C1gZYjZ/HJRwg7M
Mg5MSi6G/AYGzTS5lP3y/YqK3WMGIKT2E0VOav3dENJvdAlOwiiNdKP+hm1ODHUf2vH2gm1WEVvc
b/+jl1oFgWLYyferLUcgpXnv7WgV+mKkf/OT/rm2sUE6cEko01ZWZuH9UoHJmky3CUosqOKIphhe
wzYB9pHfajTGDiiVjWJuVOJGiN87uWQt1bqkvmM24mb5HsWLoKx2iVy31zI4woY5Qd+vLOQAGFlS
J1oTusEAEoarIH5WQUrPlf6OF+Yo4adu4xG8H7EU3NQwkkQKwWB5xgicybtbhF3vrH8anTReOBYy
AKcGCkRh/ddZHGsXsgjz84wmOCSTvDxgqLoAxq0+NuI+jV8phvYDOwA3vSc4xviO5W4UzqjL0erd
LjtiyMTcRF+cFExwGVsSULtO04Rk2sZDLNEnfEctGsSodrgF3WodjoJ76Flw1WnhSVtV8+VsFXo3
4dn606OIjPXisGZWtWWw/vvxD2tDMdLxcSK0JmhpB/fiNsP08kJMTJs4E7bVXgL9Xj4T+85rwnlw
dILsFK7awbp+7oq0kY2SEmwpqajy9b725+I9WttIxpBhuibROTVoWx2ZxYwf/aJ9hz/TMGtISYxA
d/HxQfXFpuKzzAXTUdbtRJWgfKprc1vaHFPjMIt2REvDWREieevFr6Qa77YDdUqcD41BT3rsWehA
sZb7bIbh2dTinjKDkBaMvO1ajIlYH7wEjm0rQ7gQriDjYZE0P0rX9AhPlSRzUT4BwW5KHt75oZR0
/HQQPRyBoTxun++s/K5DE8thPA8WV23XtGgW6ewiWEtwkXAMBYrt2KGJhPyCmn9096CjUdMEW0YI
9t4sNHZTeWMwbfyzQZSpxy4uEvlXM8jXmH7j+rYZHLzmGoV3N212Bg3CA8vdAguVryWxFAoqFkT8
Ja6z5xHoJolET2byjbWdoAuoeZT4tOLEjqyw9GSWO43hXle7AaIcvPsKim+aRwfM4zzkS8hrB0rG
z/cGSPBpwIxEs4636LBBFmgIZ1Nv22Gq3SJ6iTPQrCElv1S1BvxWO1KWELaPp4K+KpEB7h1CB8UA
xoFhFgVPS/q7a0FSHlysH4TxGuD3Y/jBCEl6my9dV7ar2VnvlvSssPJGHqs4P8O8EjFZB48EQN/d
J4qoG2aLqM4Fn6+I1MKqvd1IMKJy5XqiwyODxZcq1uO4s35rNNmeDaG3PhYDaGl/BAk5S2QCf/b6
dJ5TUf6d3hIz4S5m+JqKuUUJl+/T4cJa56EVsBnsw2cMY3qXmHXPyo7KAxpoIJpIG8KU4kbNb3QD
7wx6jV2Ar0mrpyhQR4eM8SfJ9AllqI2SrIBOz3lQN8VF5tSGBunfsh/rXZjDC+2+w8ud6Wjb7piN
wXUnokoz+lxoNR0BDF2RhEswycFfRzB348VBaMoLV01x9qQjNiGUwILb/MiAnXoPWJg5msD71RxM
5VOTHaVQ3GWBrysrQJpf8rt8++KlkVFgKer+8KVu7WSgr5z5kqddcaErkI/a33crkMkWBLpu0bdh
2Xex2lhXtFnmv7wqP1N/OytrCxpHxyYuGjl/7eZbB+Tv1nE3VNy0nb+iYJ2Y36abB7lqEeZ9tH3F
Df9MXHcJqsRgKe+oX4KN2ZCJpsobnyYeTTaIRt8UdiHZ0uxl0js9fbqM+mHH6u/0cexSp0LxrRY2
vc/+utHYpHF3fFgdQiEZh2mxHiqQtXVE8ia8m/ZSAArVr4RjLb+uruRfh+DYxNGmVqGQED1HgvfY
oNG9IbB+tejnA9DuTeuMlEiFxK3eH9XLgrbYXjAQwyPbpBYjglv5NIs/3G6iG7mRHUSGwhJenW0A
lB7JM9HgHc0OcOFUfptSSgceDd4ciu0676dF9Il2q1sfsJDykIx7H6FCS8qSKc+MIAj5CzXAS/aP
cH0qItl+E5zjPFZyR0uvssWfiJeSXWeUQyxUn+6ORz6F7HA/53YgCmqcgnea6iCcIXZPI8BzqCkt
S6nWaMWz9qukJX/4viDX2anuoHjrSqYKEuygWWpUY4u+9k+aBvw2ZpL+dQkye09cAUQlmFya9iZF
p52riGIFEE7qMhlGrMLY1QPMwM4FBA51UPjw3oxtby6vbj28LHbV104KQx3/Q9kMzuyANKFJZniC
oXrHageh4pXN827hRZvWltuxkKh8GhPXqSvkM6RXIsvRI8fzQq/nBsoyBEWgaAaHdtmPx6KW5yC/
/XouR35vXLU7V9i1WK0QgP9TESfXyOfZ3BKVAz8a2BXdpVjAE7ZICEXL51zBJLuLqQwwO27hYEoG
wZazKYTAIeRVXQm5BftXxbUYP9Yy74gm+sbnfjBWrobAn903QlWiFesehXgZ7jQceCT5OGCw1VA1
OyWHuYBceEWbe279dzmFdeY7TJzq7jj8CZZn+fLOPBGF+HO8YKqh5FI+3Y1xGkrBo+EStTZ5vrrX
z5n6ymLVyzwKLjonbacDMb8D2ZoEs0Ox4V+W5BESQ/l3PyXLQPVjY29ZJo2pFLhvjoWFidtNRa1a
V1crvt5mNOGdgQISSo0oP5bYIg/Koq59cvjAKw56OZuliO1wKxDjBOGbGUANxHZqJzYtpZPHDIEG
kP/85fkyoXP3AJh2BQmytZPvzhTb7kMw78P4Egj4LXxv9OY8q+RylmHp/6kMyR/J7QoZVrm3S3Qw
aIJMUh/fiHO/6+FW1cp9acQO7Ib6q+w2bWAuc5sjgJbKufPik5lTn7UulQSFbG7fQWMlyPEqtz/f
XT2hz7mfKIfcWW1fBSmnOn21qA4lqKMCtQei18wIBwh5WXuADVPny9AYbkYMuJOClyA+Fi6ve6oZ
7q6qqLtmulmRTYrvH3Qa18HTupzNOvDM6CflseaOjA8I/YWxX9SNNfiO77F2zEQGr3NFHDTmu1rC
T48uUR+kNm5d/eCZpC+/L4QV6RVuvE9jMarPiFWcSd5vQb2VfTD5f78Nz+GnDEuuixqvjxkEW5C5
dbcmRNWuhj2Fv3sPWvqnZLuoa6SyPg9GcwHNfJqNjjIYNQ5dsIDdaaDWe25ZgJEZkzgMgjmG2fi4
dQqNy1uwLr5KFuFLKrIHRUyTqsMvsgwK1Lv9opuVbFbeBOwU/0KSdnBSC2TZrENMxxkbXZRDGl2f
NHjWfjo9YVJbcZ1Rsa3GUePQM6ag1lvHcuASCTJ/F134mYoq7BqbtxRilbX2LgBDjFW4Ay1W9SCe
LQKKtA8Z1iJCSPvY0Lr7mwIjJuhb/Qo7ewHJvsm+Lrh8U5A5sBQFNjE6qHUPDek83GGq/MTeSBLF
1cqDDG+BZ1ihRYI6psz0ZawGvbkGJJShDFjIeVm+jj5uX19CzXu1m9e9+TspNBM+yDZPYUL9FSQh
XhjFZpFDxO4earNB7OTwGjhYWA12jRJeCY9xOIh3HhydwQZqqayvO4JIQK/V+ZICzeIc395gvQDt
ri9uwFk0cvwR4UONfKf0LTH9tKfathnY1VAgOMZHR49GFxRPaJZ2tUmn3Pm9LnHlsS2M+HvU89L0
CDPhmHOATiMv5E5RYWOTHGe/A2qfsbCVxIVyPniBjZAjSMsDVlQCwTpqiNnn48jMhdBOhl2G8AYT
iOAv+OqHoCmdPsac75kwzA3gQvTrTwQThT6mrdAjwBwS6UfqnR8KgyD4/MGlvnDCdNJDXcwRPv0Z
Jp1+D+gpHMfypdnMIeewOQVuZXSLsE974NbNF1WtdHwJQ7bUPraeDxL/T9xhxySlxqAorXClbur5
3U2xo1lLlbwZE+/XE87k+rC2xXozcM/uausZOpZr2YlaN64nNCHo+IHSyN7g0A+XxyaPUDvX0B6s
8BOrbEoNUp2C+smVlxL+2NU69xffyWws3DFOmNJse2brvYuK2fZsy0M5LnAGlkjMIJ9rXofm61Cs
Tp3k59PT4NxU1qa/jxKaqqRDEQbsxLsDfwvqBu+FoPS2+khzCIBcYwSIJL32NxHaCzTTqj1iJr3T
3NnW39bEU1qVWzNnUg4e1MGO+xfGXpcdQSlNfeaOOq6khonWW44mgzLggs/OQfL8M1/mHnAOgDDK
Pk3sp5gHd1TlmJdq9qWNWaiBfk2z/8gAykUEJ2xkm1aKirFUCfrCvxKeIlLpI40/4AZaq19DUsqP
HbCHaZHYSqPGHq63JR6/5msfyULt9p4+7r2xEXJ3/Z3xRx5j7w6BYb5Yv8nGk9yi0fr3nJRRVAn5
1F4O/OaKuoMwfAYWbA9GLEmmKE8qoYV4trhUHSFXhWQE6fAph7k2sfZDb9J1eSlMeGGy88NNT9YT
Ys/kBaQvt4xVTgRWR33OYZEBPKzhtVG+UzRUrMC1Q53QaVY0RndirIiM3yLpYwd+tsi4SgV777yx
26kVkjxPhhxMblIxGz5rBisk+m6ywGCrbBhwizYTGzGEAgNoeuanMz989LQngfcel6QlD6n23j6v
AZSlvXfWrdrR4PbjktmKa6v9SZEcJKxCSrSGd9Ugs5ldhEUvvvHCQbVdPm2qGQh2r9LZutGf2K7a
4okTDIG0ZjDLbGLcFBJBBfjB1nvfaZZsJL5B/AjQZdfoazR9ve/WRmc2RiJlYd7V/vht87E12QAU
DVlhekRbOe9SsTeZXOr+USWWfFd2xcaZWcyPtUF16dWD3vE3WrJe+cCltiEHMpO8DSqu+y+qKVMM
+hWMtoJQ7EJ5i9lXlve+Px/KQRtE+57V2XEKEcPrzrYN5PZaTUwcZKelbCvHAyvx4Ej37XROTCzl
ebQgoglcoy42U8SzhiMwERUwr36wsyU2C8w5ocd+rp/ymGv1Zr4/E0YpEe9xo8erirCsxPRNbCJM
BOeThGCVbVXoc9k+MztVteOJwdxaOg9Ex7goVFIwfjwYx3l1osvnYPte55UUuq8Y2QYxGi/+Qm5h
VRAuzQYDhLhg5GznliaQy5qV2zjpgeuvmxr89q7atGG/dToIhPT5+pTHpaRwdtiLtkxVAJEj1ucn
DzLQBOLx6Uop97ojx1Q5Elo3Vi/iuJa/DymoW8iagDgZniDVrCRlXSW5a1BgKErWoTqhI49lvnj+
hFoIt7Bv/gBUanAm0C6f6/pt0LzokTmn5RjbP89Cq8SeEJG0ArvwPBjlD86UiebBKq6uUH+AazKP
WyvvsdJxsDa1C3w9k4ocjunhLkEKdTzlg58pJy2tWKAvbjHDHCeNKkbRB0J/5hIDFQ/640NrY6zr
lKf39om9CTiHKLJTbl+kXeUMPyBJ0hldPlmxvPuJzMO0puXAAE3E02U8i9LvgQ89IChzY8mSxwiI
DpbYySpM32ymuhQQb8DKWlY4C5I17yLKuL2laXekgcKfRmf0xy4bAeD9PJ/AA3btCCfIVwQdX9QP
YiUQn0XZa2FlD7sWROnOI6w7kxuzgAz7zPe3/Dp+qMPszXjoLceGPaKlbgI1+0u7WkitWfubtE2i
2yvRJbkvUX9iZpO2FOKzlq7HAtsQOZenMaiznAdQ5z06il/of6tyMYPQ+2VZtaNtPJLyCaF0Uf3m
xEC6/0qBvsMargHqVzQtMG5ZjhMVFJNSiNfPjSheTCWNAJRLUlwiq2lCKAPN7rH+RTI4i3EZXGIV
x7UFEbX6Hx8lgouSo8WR7FiEp/m5ZKYsbgNMrrY4or0M/mnZbyhc/mqbUVkcEQL4iIWG4MkmABWo
C/2GjuDdtJiZJ+OF8CWEAIJQbRI4JifHJ2AJrDIyPOFfo6nrRrvuOow1SA+xSsRf78WmRux+n+gR
5dzDunsF5iGklRA3wjCmYyZgHYZxFrOSEP7E7VKr6VACQ1SsyHtWPLaY5h+PJ6qKjZic9y6le0j1
ZTFogUmf+F2vQVNqAnxtyyRSPmpwcn/6nUlNPjlPrYZTWGqCqr7jWqEd5+R9KVD+AN4eGt0Mo98i
TygHlC1u6X8j3mgu89WKFdtF1hw9hhNq+/rOrYZi2jdLrdM7C+AKEk8ARLTSb9UUtcTVMXQo27Yb
W3Hgq4+tXggrRnhVdp/HAOB5U8DGaI8svRbfJmzFX8vIlKEOwUqb7pGd7bZ2yArBoyZrNCS34qJF
f+ivYo6C8W3BSZrdyb0rzXTP0y8UWf08iKteSEsGCdg9jZOKYQ/eIAXe0p4zjPoyTf6gThaeHnWv
5oDV1AAszN78hfPFW24esBhe4jBdMlTCfE5LrmTfRUZNMCY5fhk4V3gtkAqhdsIXuBZXadzdXbmj
xF398Oxa8yLlr/ZEG4uEhRSanYAiDXvZlAlD2gQyw7HE4M2z/VQynlrAUEcDYTeOjm8wBcRUeHIM
tcYssUIr4XCmQpEeb9CJ2Qv6+3cVm04IL0l4Cnoi/75//Ja6Vz3iXVp0tYtehYWhXlJ4sjZN6Tu7
EhpUBNvllV/8/jLkQ2g33qTCDv9FiLX6N/A2nKlM1xHD5HuoCKbFHDrI5XegH/ei6RESwUKiB49N
tEYVnGx2WpTjjMmP6LtHqlIhYdp7Ic57m+WFca4zVfCkvjqSpdKvPfuiZeBpigy8sexGBxGs6fNE
cJluwF5P+djL8XL3PAwTb+nedPIUyxXuprYppFZF4VM8gT6Shir6gFl7F0/1z5xG++ATKm6vPAFU
I73u0wlkx6poZChWUi0wfwZguSsimHOC/rni048L7jITnViR5dc6g5ibJWBnrSV5mDgDD0oKzrJr
KeZwX5lH6p4S4kJVRj6o4azXPPCAHaD3HQ0V1xpdo5oRCGJ8a+go8ygsj9pRepwVYPEPTVtwJC4h
aXf5tvvPoYEwh5zjqMFW8P7jrAHXk7cG/Cqed5Up6rPK3fewFwZfdBV+bj95t5aI8B65uBMWbmOr
rt5ZU1GcnE0AzxCfHZj9FwrMP3jO7dfM2DqI/f24OQEfLfvhX/21qbVmk4Raf5PbolhrsKRp1/q3
/EZ39vP67pyz/gKFEgXvNrW79HZVAYY5M2u0d9I5eBz8QzlKlGGRoGHCIuwDlK4ClXiU28xNOWUi
yoBKUjL5aHSeAl1sTX2U62Ef1HyqVsDolfE+oIP01Y5VbiU/az/sOi3lPn4PpuONZNy0Lnjqzj9V
FozoY7/Cux8i8puUabN5rx0T+JnTrwLVdg1EGqNwDBQRqZiZDhGn8t7PpWxk27JbDNWN/1Soe7/G
tRQGE8p9427jzElRKib2VoSOccPavEMIygGK/Wy9diW1rC7IQDYgZrRJpRrNOuwyLe5OVTnPIYH0
27LrSWgxLxQk6v0FjbaIaS4wGt34lZ9mNS9//mmOCnREKVZyxSf0f41ILob0Jjh3C4Gu/n6kYaHH
WpsrnnQMMqLcMx1Zy7Op2tm7/FlIUp7uaNz/qtrMl5HuMpxmcgTza9vBZS2rUcK/eMwg8lM9e+UY
vGsoqcU4Nr08epxMY7doSSOdi2OYffyNI5gLubWeAhEGKc48aBu/81imZBdH/lJ43qylU0W96zcZ
KyEtOIR8VD8zjTCs0GDd+KkkF++5MG59lfLhM3ATsyBzoKeBBeWz6+ilEwe4EFNwtfSXC3UhXp3V
mPYpn+tNZnpgcbwlZU9gc6H8H1tozRgLcoYUwlU3YRuesG+/Rz4T6zLBiuF4XC+yChEehcD8jn3H
ydJgbEyFKuzEPEl1wWi2/52J8SB/p5d0h6OPrYdPb6FQsC1lYss1EL1KLB6Zt2bfHPzPaZlErpa6
mBZKbz8AO1vmUG7SxzngzcT76DAYriodE3CImI2Vbw0cz1pNyT/RsA6EPp/pxfy73so/MIQaCX9F
03/hlPnAlcRQAy+bug0Dkk9miacajfxOJdMdLMHFH3YWqiNvTpsu3D9FUfXwTrkwi+4Ka72WTG9m
F2TKxDJvDYqfaQblkM9yufY9yFXvKiwa5w3PpsvL+CxicRdK2SmXkh39TRzzrNFEJokfyTuJnYL4
ekhRxyXaBbPCRrLWdJ/uoqso7FJ76hqyVIG4uY6+i9vTYoYs7rrglhPE5bylQsmDHoqGJ3obOAwb
OpRdWD4VBSiznGMg+cov3G/0gOBwXAl2ERLFiaS18cPoqfcmhKpzD0Dk+u6lKbRwPn+isucXev+9
mBysirGQWQiyNWYgKSOo2zUt4OM3JUktDYYX8Wm0Nq1DFStaPP6ZlXO2S/nDcZrauHCSCAqc6ijT
aXrR/ePSZkmWeGqzXKA+3uhF0GkkaZkGRAfQFc1cdGUoIg/r7qlIVEXEdUMy9Wt5Gumlq6jByXKa
qcLu7gAsmERwcfqeoKklmm7FDy40u2J6gR53+CK4LatQqQvHTpo1IlnSQ6kdaTQbz6XP6FGhxzfn
CwZObe1w82b1K1jW9PE8FCHbTr9sTtncY/5rOepJIzETTKhIpt7rvVMtlT9jmBDEzhPiZ9uwN3FF
QxLgrk8AKWHAhm31FC3RMnS6KjZ7sj46vW2seVoNG1Xl9g4llHa5MYFp+yNmVfvnskU+5TSI7wU1
zU6pPWhXPnbFI7cSdK2MXR0kUmJS8Vwso8uw9nEMcAxvKZRx8lDX7iEUVxSOFYd82QyjXi649OHX
Jl1aXSmOpSc4QHnWvz+thVlFLDXeQ1DBGTHPuPNY5X2aRzaSdWGxoWJ1G/QUF18zzkUwgGk2y98b
sG42yLX8qjNavq8tyNQQGRIbSIvNy5TQtTF1DzSK8b7i93+/GwJUf0zRyleC8afxkCyNlXbBR6WY
RVeNBDTA6jv002nP53Av1+pBmC54cLOBHJBzkDTSigNMYHcfEn02PzlCdaW1VOUdDh0gbPjPsW4o
yM/eT+GNyjP0AE5RYX/Vgcuos4v3o35sG1S0P0asPCa6uU2UXc1zALyuOECrGREYiDkpZgZVG286
2tF+UlutBMyDIzpWmHFu8Y8CaEmScm6P8sjoz3TOvDAGHOybd6I/TE3S31fPcFg53V0W0V+XWS8b
d2QbH9SknRgaLtoD3dDCdvXpLZHnpgWGPY8KT2Fm7KoJ5R8WESUYMwphjLIksba7u+yiqbYHTTOz
+GlsSbsIF4NTw76NqwHBfPr1KebHYqwwR7Ap4xxQKOO1CNvvxwY5BnjqVRoxFS9xt10VAsOM/oCx
7/hjPdB+YJieyLl4ZsXHyETrlKT8a9CtW/RV8ezmvbytztizJuWpy+2U6+NWJQ803z3K708Jjv+M
D9GXSQh47rXY+54AM9H7VL9jYbddwZFt8npGeNfW+Ha366/rXaochtRKdi1fFUGHA8iaHHZfYsvw
l60qlVo5gTFUC0vBTe5R3Z7/vMtCiwMkk7Lmhs9XmOGaC4TgPEs8c0Y0eyHYbDelL4HxUXWne7WS
6ocVKUT0Yh0x8Isg/krjn7ajVtFt7lOFTcbqmqFzuY1+LxNNr2BEhQz5Wumew3RN3nj8/zPobXuA
UPM/iv8etD+i8IMzsUVOPBFjbe5TBW6RWUIgWa46U+Y7DvFW3fDW2U+cqzVPSEJzKw8uj0V16l7J
FZzEFlqmBSGp/OJuahLU8NjH/t582jsF3SKms/pFauCsurwju2Bw+87ULwNlHEfSM0sVRmv1dmpz
y2rVEt76ljsHo4lbNcHEPrfvthMVCrp8yvfzgDvo+JcUxEFG+9HCorfuM9wy8IOVFFD1tAPdHrLT
Xbap8kULvASs8GDTdcbbJvE6MDtw4azX/KLoLjExKH3sCDvwbk136VMjXAmV5tCGLL3HOpgyGp/9
RJX+nCjoEhatNe9pWOpAR1Ba+s2bEdcKp+CoelgqXo/rkeYMIYcsm8bXmYp18D7dLfGAwZfzQXCI
VWP9U0NB25rc0lJtQs4lsWPsE1BIaSvqvILFeK/TQMoTQtOnd0/gLxBHiMJzjDIH1L1bk7xvuVU6
pyrtHtg15ZRGMmWATNayGke5G4PoNmuIZiyS5oZhL7gfV6vBEybfxQ8Rk5Toi/CDyPwkf2ovf3kJ
c82CfR8vrX3imLp1X5dEZtJvQXkpS8rOnGhbblGUcviVPah7parpukShiEdk1VO+pCRW8VLuV/zp
GO4OTQAMF0iA5ZLaA75ESJHZN66PGCyug3BzVGSkrkxeuJcjkMBYQvlthfc5GeZFNBMbv3ai+/Y+
vuvrAVeRSbPHvX5j+C9x+LccpCvU4hrX+m5kivkWTHHso5EDJmdwNDSTnaaKz7QZOWke8E2nRrYL
Mf7y9Gdljr7f/RxToZ3q6+QO+9+B4MQj6hEYCm7FJInJ5e/eNXSKuCGCyq2QXITFeDVRuhKvOTY/
aQRWtSPoUTBdcg717FqvFXP9VELbzTolygpoT+5RkxuykjkP12mdyi5ReNM6i/WAS0O3EgOHZjAg
/J//O1NBWIwRpjTQwkzkkIsatMLUW7CSRkDr9Fzdi5G/Zs2tIA4jGqugZ75iMuICcMOM/+RzPVYk
ykDxAPvyM/YagrlHtpmJyAuUsk8E0yBurWoWcehKlJ9/lFjAAHmqQoxYXmUy7+LtaP0CdWF3dzLo
Yz/TB5cA2IIeWaE4tLBULixz8tVQKnN3y9QN4k5Ab6IV2HH9T7aIepcz3XR46q66hXNnKgfjNnUu
TvepvUHcBLAafR5EcjIwcgsBJoV1V29saC/t+mWwSVy+30lAbuyCAZucl+IS2JD1VyLX+29GFOwN
zgXD5L3oXV4ES3QlpfK893zb63hgJuzhq17jyNyyBcA0WVitIvxwgdJntKYqACjQFUE/FfQJ0tJT
5rl4iBNWCiT1oh8ds47I9A7U+JzB4nwdwpFwOHQPD9Al6gQ6zbGnuS6xqVPSRTJaBy+FdV255t18
6YZzY8h2th5Wt1EbBhS+M+DkEP4EYCsQU4dSjMOCrA893i2UwYWstCzb9HBIdEhquU6342E2LrtA
PKdNmqITCx8cp45ukF3T1GZ5YGMvfSzxStpXAK42Ny2TcmKVAINGHgONZDoEhBf5vi+LWLwXxCEw
2K+UdqvW1siuZS4AcxHbsulF4Wqdnf7i4SjpLR/0iRzH7NvLMyhI9AQvbE2pQvVzrsdblPJQ/svb
j2l5WNsdqC1W6kYpwMXzY+q0NjuHOuugzJRBAU5XdgnZMkb97MlQ8QPuJffuRb8eIKHoJzNT9u3m
HpFRWaOS2TT0oukoYX26iSFdkI6nJpU1IKB1gjlkc1LMn11YFgEkBne8Uo3u/qUOfh4qrIerD3FG
g3UMf6sXHp92EqK1jiLF9cUAXmjhNDrG/pe/aQL7IFRwdxNTZK4nNNh9G4gxmgxk8jntRnzdR5I+
QkAt2dyc5rbV/Y3m43+b15Sr4/w4OqVgb8kAzYxselzSPyn8aePCmQk0kGsQNNiE5877Y47cWN9h
Ksv5fAWe3N+GCqLQRgpw1sYXK5WxhXDnJBwYQQ30zOs2i1WdsFdTPU+u5NLNBcbZY5sA9jLEfz5p
RF/lstBqNpSADXJ6vQQ4UhDoCbGOj82o6A7lhSEjmf5+sk9/AQu/+M29e3vuhqW0F4cv+cvGsBBc
613KArfESW/IfCwhyQsUSsHNerOAEE1DCcpNDt0LySgVeGsT7oHTMmgcC/0nuXl6/mVXQdNm/sEz
73D4q1ukEUOTKjDy2MqDyWaYOsPza8mxdsh1X6+n4SCEK3WrAGno5Kp8p+a1w3S1yYsdtS241DzG
PTrl6XV8jHDMe46XA/qllDBEFdle5vBAxOSE1bOHF+uzkrx0r38OdxHnnPqbuNKYdrsaY6f+1hNm
wGXhuEn0Jw712+Lp4mzFvZJGcb7CmHMgmhmmZiQI1aQ+Vi9n49t9kxUG5g0DL+8CpdZ/i8BSYYHZ
SRDbhnoStMk1mRHkNr/wFa9tZwxt30atg9Opwx7lwQkYlDX+HDkNlfhkQ3Gz/90eLaADMwcB42/J
EoOk1jfTskDMIFOdhJ6mEeigq03vTJFL+cwFfEuzHAZ89PFgBBim19bSiemC9uAXuZfpBJc9cxK5
GoFBG8QOcG139d15pdf2OIKtiDH4I/VDrHk/I2PdpnfHUMMcA4R22XWTho/EtKZVDBLyDQmGf9ku
ZJNICzSwlszud+skzrzmSJHrosmVzzdQQG9kTpVc//ryb42ao/P54/miPHVmVTd9VGOkRV7OTT1h
e7OLfxknUSBbIHBE+39iKVL9lm4NgwRtG3HDabvmz39zWKM32b36FP8VUkjc/D1NL8ncO4RuwsUJ
ARXEOJuilFAWhqBRYHs7NM32TMJxX16ehd9nIX3NocE/mN8k4ofa56+b/7B/m0Vz/R4FMQ9qvkgz
izbt91inJX40D14XWlHQRBy/RoeFkncSHZzAbKVz3AyRn2QJdKK7jbtRY8DDLsDTx3JaCqCa2DRz
/A9pSenhyj9nFJj+CLhhxS1hW0NVvoCxfnbb+APKDeszzRKDz6QsBe/vhQ10LrK9VtKbmos+EfnN
RoohVLp2UTr+cdiJwO/udTihxqCOFlD5qHi4rCByNoXlenjQBoJcxYyztmoqgBbC+EOpH7mUc2Bp
rEK1442KR+Wow4MaAdUxZLd01exBY2ZkJCF4spErWqZs1MFhSDBr2OfH4SU8VcjK16NuBHlGxAkO
S6tcW+6pyUjJw5rMK1orq4SXKcvyMV+fi4QrIweGX9Zorms4b7/Q9STx8GMkar/zEK+AA/R45VsI
h+EvYHMwQ3X4jT0XMxtT5YuEz13Ewpak+hopLVCvZd3Op131GWyIxjlBtUO2g+XUDo/vD8NYz01G
f+Cp+6G5p6g14v5tkOydUes+vMrD6fcqMUpqQIVrSjVjXtHInU+KRFkyDKO7YXDLfXtz278NQL4U
wOq9QVTqZz7Zji4bbkJtYAoT4nxpImu4KO8gSo79QCQdEkS5/Yj6eQSKGpTsCmOp9MTcguNp2qGC
ZlL974Q6W7eWqCrDN4sr6TS4kdeWkVm+p5RpTk5M9o5ZMg2MoGzNsGaHYUw/fpS+Td0t6fZTf6m4
xBJXbo4MF2ryQKWCWi6sVAXp9vD/pcL6yK/KIHP7iH1BIwBy/TEp8hNPqYm5yr0b8zMvXLYVc9wn
BVQ+bn6f+nDBlmvtQOGtO6M43r8+EoOH04iR2982ROdX0hV12SOahXJjG5rMXwmhY5rEK2uPQJRJ
C8j/XUwLkFWgr8G9sV3WzPEoSj3/rm5FRYiPWRJnC3kadpzLWDUN955DwYXunjSkSih91cFSA1Qe
PJj+Wlb3e0SkkU0goJTaxlulIwD/xMIcKdd3iZN5FCohxvRqJCf2EWOtnegVCbTip78Iosi/E6vM
YBgqU2maE1GZHPp2/wyflQV3PV7ev2XwtE5bCSJFO6a0TveL87a7aL4qccco5LpEOUeaEUIm4j3q
Kan9LKx6VCVhbntxWhbWxbnNpG8dC1CrvaehgXS3MWUix7cZsIJ/3IbhaWt96unJoYoTA3aKBP5a
ReJ4OQi4nrDCPT9RKVcBwPdt/AC/F7eJXvssHI10B3HeVrYWQiRMUkqJ6EOsxGFF2hgWZixbZEqO
/IuoCRSoRVxieV83kGFckLEg37+pJvnJtGuBF4+NBwdewIPg3yRaQtjdg+MNhIUygy3rhqafOq7r
4iwVBlqV3NyKxphGE36g7MjJtn1tfQhAoTPDiPBrKzri4JHoQptfqK0+cWXsyGA8f/iNHah6XBNo
WoJBQA7fpI/NRn49bRjb0p+/NDLQIGJmnqWXQp6BPD3tylpyfa2Gaanx2TuBaTR0VCr6WEo3uM2X
oMYVaxOMb+f2s2eScR6vEnmvYAiMhphwQMXqm+3VdypaqUtFm48T/pqk7hI9jyIfb4TpLEmrjE+F
KRO3+gPhPqKvuwDEa4D0IthDMEXqn8fq0TakzGRb4T226+Br4Y+mc0voYovMy03Kdq38JB7xgxmS
PMJ8T2TN/fQq90+2uTlgFrS3s8oE+8IbzT0+Kw3hxYwk5msSnybcwl6gqjnLci8MNxXFFwOG8cIM
sOjF50poGLhkRiE4tiOSYkwwOltAfepjxT7RtUbpfZEc67JIAIU08gOjbmNpg41BifJd/Y2J9LJC
9HuRLZ3bfgh49w7w1UWqnZyqUDa6cfwFvaPUBfqVV34Y7u60MAPXAHLJRh5xHN/2WEffXVPcueFc
lJevhAqOz1PCZ61ss+y7bAJpCSzf0sxKnrOQfT0mCrBuJwd0iMEueUPskn8RrBuE/AKFzpvtJ0kR
CbVtg2lIEKMMUYoshnIpZ8Flc4YR5nYxgMu4Dhs9k3DcvjX+uP6A6S4o/G3pPMeb+LEtevZ+ObdM
y9I8n2FePczVUaKCCYmzIKJPJOJTJiHY7SqYNd21SK75ZWYsM+fR9jMbj7FGkKG8E2Li/6R+SdGV
GmyOnJhnHmoosLSFwVXtOMjT2OYP/TIfLLiK8bEQxFurj9x9q2ZZD6Ww6P3pm7413OQlWBsQSn2p
tA7JOKOBAOPUIn/6kcYvT/rengHmSCP7pEKxHOPTc9llRz9P6DNRa1B16QTxyWjhwIAmh83v8qa3
NvQ610eC8NAbBXkooMh6URqtldKpBZfB7inQDdjtUybWB1Mash8F74Y3Vv0RdCi/8JxWNjgr77Wy
I0LaB0FUclPgGa14ma61y+hUhstGRB0F3e0MEXzLEtCnJb7JgWKmz6eSmKSlx4y21mEoM76l9mmc
b2TVqdRsgQhDSdL1HZ9KaOxWuBKY0dGozY6jqw9m7M0pgUKFPVp1oCZOqqJ5W1oWLhztCxpRkjph
76haf82jOjhE1ix+3NJ9K2SGdYnID+UMREmi6BpZ54oQNLNFDP8RrWkZ3uboNtuO4oOfsS72y6J9
PIm9m4DZ7jUbEs8Tcazh6adgJ3XrWUfk3O1SE+jYSdK1j3uYdZUTLUL2BJOCMXpte1922TDtgicm
Vbnib2frxcGVoTZA0CKf60ddg0xK6g4HILAboLOaK8a0zeVO2lQLEgD+YBdcMXURkMpVuQBQBwdP
O1VnSkEn4dvvg65iU/vfmEGAMn7v9p3KdixTobbZf7rKNjvv+/5JLRl/KxysRXX5Uvw6z4h0eiWz
IFMjnLdSttqZxgoZnJa0bQE4xpMxEm6dVonENSxZY9ZMxvvdSXy644bXLKWPHzVsA5WR9QCc/QHf
fkzw8eb9B8gt8szNj15+O9spOUNizgzqjsv1V43b7WFkT20t6QxcvYPIewbDMwojk5yP5orBmbMp
t00exybOv64SYOtWmzNJIOYci9kbNFKdNO6fF1nn0KXQXx1HajAALkZgLx0ZFgYbkQOs6iyHqPSR
gJ4J0/PZvdVfgIu6JrYDQjB8FIXcLo7GAmxsWRV3ufPhAWxaGR3M81I0/XzTXI9+zCTSfFt4mS/x
tcIbN1aRSEIjIdhG4Av2G5zec5neZC2aVK3KTjseFCqJ836sDK+6Cca/EQgRd0BY5gjzxPkcDr9Q
FhbFS69HmINPJNEsGIVf1Pq4j7eFc6pucTFTorBekfezCwaE0dnGRmOEDE4qSFCo2wdRxI2hzYgd
uF+kaYfJ0MFTHLWViO+OcM5HXvlxXLIVof96rweUrUf/hYhs/zHxCKMPOAkUNB5Obx2gNoVTEm6B
3t7pYfCh7Jf4cdUiYe4gz2lQupOBeb1ZJgDsFi0Y6aq4edgnsBhxjsX8+CzEusfneluCpv8ChHsp
jYeCRAGsmOLkbgiEojI6h4YE3AkuO5E2wf5bNn68uEYD1iZWpgnCiRg+maeS8vlPxuvPtU2eYhcl
LPvU6UOJ+Ukn/dl9xvepbyOaC7gRNG4/8fgSzbiAlZ7nNDi1Mscp7jMnCZF9q7ygRNE4oLCVVsAV
qngWo+fuWG1nMjlWpgP7BXUhvy2ZHEsPfooszvb70+PP3yXG5hQfRPhlpuUiF7c4WhLxiWJVWN+n
1O96/QN//Ek9criO/umPUQTrpCHTL133gSVXKc4Isq7qzO5iBP0M2GstKq7InA9c3SS5HiaYxHfc
1ktJU1Lswc34ugIRa7Bl1VnBK+KxrXAz9AKC19Eszhi1sPDoyljVxP+0rzpLdXRltnb/tEKPRTyT
9qvO99LNY9ddE7A/AemiXWiedecUFhLyNVbJ5sOfWCFP4Mmd+69VMq35R2AbEKjfWFrfXBkZ8z9K
O2C0Js0iKaxGh7c4xkLrT7k60qi2bQAzfV35aI6CBN83E1YYlDwDagW+zAYx1NAPh/D7YxG62aRG
R+YG94mUy74xzKB683P6+gQvttP7kuyC6BAJ7PVbiUfeHmqM/OePzJ/z0wesiB1m/bNZ1Wd3s+Ru
4hkNz5FKKihrmHsMYjois9izc2LiO4TAOipo8+tRr2rLy9+FFv2nLZYNOCoN5B4lZYMeuaKunCrH
vmVTrNqh6y7YlfdJCeTAotelMgG6rN6MVB5+k2F3zs0E3bvvSS6m8kRxmUMlsN5vG6jctrL8JAdv
WUna2kehU29bPLXShupoqLA+siYMPdarHo7jeosbBQVDdXYomvCvFAHiOHJ+ZX68AHlPC1PpNdGq
M/1sqeNzr+UZlweVjx/gDvEOrFxVVZ9VfHjxNFMyBBCmEllhulXr0LU66CBdW1jZ+iQBIvNYUW0S
ESrtJ8qSsubFutkO+tjpBI5FG5QP7e/vJq1hfyNBg9EzDHkGvgzSkpUlc7gl0g6ZxjJK8VS0+S+b
4c5Cyd6x7v99AcHLX0IAGzn++aE+U42ZSn04Ul42F1CO4e1EDCr51eDYjyx5gQIViyXpB05kcEO0
BIAneaZUKtaKzWxLGqHAlKwx24bbxDW8hW/qxsIVHxy5qZGMB1WqUi/2w1R4Y5sGfjvOh2z4dqxE
uEAZFS/LHcZwEuDFW0ULOyzhDWDnVS8fHPrw22Cn/sQnxv9Lm0V2GuHS1FxnWvjsFi4EAvjP7J2R
7r/Ys0mxm66G7j1BzBEoVgI1vIVWeJqwhj/ZLoJDw5zUW4QfPKmqWwBEGGLEPPEdT9pkqQJYIaeg
PS3Gl8ZmoNkcP66r8VdiR0Mgyy9w/gbii6gykU6ZBGgFhbfxUy3buKrYSDhT1/n98Fb8gPDTXnDI
Q0mKwFHDmoD1J6VR3z9vo5QEfqcstb+0CTUx+V9IKK3VYgzXtfcw2emsgZZQZ8wKe4cwBwMiwmT4
Nnkr+4rcRq37IHjm97ukE+LKtn5HkYkcCvSDatlVU7URSuMXnLccTP+U6f20RP+iWS0M3JehRx+r
ZGJ+rkOSCP4Tj7VM/QminMnD0MSWIYKeQjeeKxS0fKchkO21ft3AM9EWl97u+5Zk8IGA0JfVZE1P
4xaq1rtFNOM0/gYz+TW2iCC2BR71DWdcgu8NZ5e3NKK3zzytBHr/fGX31bcl56l0EtbK8N9qMy32
NJU/qQ2Mr6gZSoQ34Btb40mCEn8Aa4QDiTkO20Px0Ua2dof6umtZlqLWkkN3Yd8AhO22tYVxE2wb
2531ki8Xb/gMXk9WN2eq129ZeW3vLsACIJJBL6z5tfptUPDs36ALT0j6vF2jhh+pTruivZsnP8+t
Yj/mitvwguLlbTGGegWHkF1A1g+63sBIlwKm4bKeBpMzStbeFjaru761+mHfTSCFq7ppmD4w5jy0
CJmFGgYuwF2O6mpPvVTPceUtANRMBy20P8zNRpE2RhIoY/q8GtudrXtIpYWDBfTRlA3al26nwb+u
AYZKh20ELd7tR5Gzf8/cMFf5RxeXJ7RM/HziGrSwaVyKu27y7Q3z0d4MK6wNuRkyWErvoNypqf3e
QFQ5cUgZSfBnJSbZ12QSxSvM8FBxI9Q5W8ydwWoI0SS/STB9LADrmcuelnl4iqHqvLLGE57bsBn8
Cvu/tu1xFO1XEMOlCGavIKTmkhOBNGqJqJmTlelYEpH4XqWdFd+QRaNrcuWbZkUMfd+E3dr3wEXg
F+BOXkWRYHtXnzcLMzzrF7LI8A1JYNcXHYYCoEN2NDeyXFy/J/b0f1/CwegCsQlthG+m5sCo97ub
qlRFGrckZ/6bCbA9JHccuGo/w2fXaPmQf6u5Q6Jt/EU4XqJzfY39XEwUzBUS6EWXW3PVhEuNnTs1
1OQedRbtCSyELTE0CstrAttUtm0c46MqgZbY5h8yetfhOCJyHkwRw+EQKq2MLFnZeYN+JwtScNL7
Y86yq/W5IRE7AmqdJnAHMQ8cYEWJMzCZYiCI9uaTtrqS+KOjnpNDXEJIJYXxLQQIwwcrQ++UVcQh
X6dpzCqLu6ZgNcIahRgw2nIHzAVhgHSE3q+Z5gS+R3KFLO/RzjVg0uMUz+NHuP8IedF4TxBN2UXu
jrOiQB0FnXuV3KmXm0ZY7tEN6kBJdnIB52K+ah+fWC7A1B9coMFNO67BeZ+wfViX/8MeXBEgTvjL
QpBj7tJfQDPam95XWsmSLXM29Wz+oe3sZg4n+aFRfdUIJ9+9OiV7CGw3im5lYQ6O0Wkt87sCNw7/
IAkpOsrhb+kIen5LBcg1KOfwyKyXblOzEffDaEBJ7VEY9vJ6mQ0EnouGI9d58NBffso5dElN5cKo
BZntSwoQ18+p/nbkoUtcxN8HApDdHRcsJ3TFvkG0mAXY7eunPPw1FW6yTJTnzwfF9UyPgGWxB/NQ
82/d/s/9hiHy0JQQGZ4jLbjRSSz4F30smaUdIpSJKkQsUqOhB+i8nk+6tVWJfWAQRtIL4H4Tz0ZT
UNaUkURmCj5etUvv1jIv4OpNpC8KefxCB8X6b8RttUz59rdtACXIr0rmTY+EI3P3sCpVLLZN5Qkk
YzMNX/ytKW7YcYLVZQ3DbUUH9l9LtAviyKu2q6l8oSoVMb7A4zs+3UnHyCmyFxYERxTm+rAjXmZU
OZ5mYBfoRN29moq9aDzsSaNRKNz+vkVbgTMUC3ATDYqy2He2TjEYf1YXKROADyNvWLbNA+CDQR8N
mNO+RRhNHSN5AEl8b5mLuecWb43xIUJIEhxfIAyUcKHFkZJjO/HLt+zQucdL9lEX/JSv24TZDUNl
FKG/QPm7yOah1G3dSNmmpXJPzmaYygHnMXAQFOYJepHE+3+q+SAvPpF/ANZ0SqRxwI3yeDjVRNbH
DnqG6d310BoCr3k/jf1kF0imtav2znO9U61ifDshYiC92D/mPcQ6GLEr7a1HEOVBAhkmwhbG3FyP
fsjY7W5GLORRgt2SLug+jC2kEv/STHEfOwZV/S1habTmT8ZwwrCD3GUWCXbAIgZPfcvcuMTsFqLW
HBs87noSEK+c8yO82eY6klbX7+voAVldNYcURBfz9b7sk3eUPNNYUr4IhefowVSaMhMtFjcar7EG
XAeFzbEAdaMSVa/DKQbDfpTYPkgk4Qq3U3KQOxrY+AIPS0DSqnYjMRmCqyWjaJIFIUe9hO5Tal93
gaRk3UN2nym7fNwni917XiALyEDhJhd7b0uDFpTeWOtydG2XMRfwXFDM2xtfrZuoXGkQWiEIuTDY
jR+64+4RtsJPH0wNLtbAyxCkGo4Q7Il42xWMMptuWfKyGWu0/7J3wEFBt90rQot3x4samx2SV1iG
huTZWZRedTEVX9iYHZQnfA9sQljYO42Nc7P4gx6QpMHjhoTjXh11X/BiVhVUHIxq+PUxszKymruZ
U1Q21dwHvubOPJvhra9E+DHXCCfL4X1KtAafpFu3LCmD2R6i/Zh7HW7Wu4TAcQfoZzDJJEcwZesM
oVsaoRLHXYkxFrqW+NFbP5Lsq0OpK3e7qdAE27J65GirRxgtTo/0IISDx+IupTBvh9F9gw54nzvy
z90s/ffTn+8Ek3X+8oM60wWON9VQ88tgTLQHOdaFUpKwk5s06RcP23xu8eiBu/cBZzE6CDiNKfgu
RpQCKZ5IS1pcKNbYP62uPoTXbLm8yDWUiNpcjM1nmKLyXgq0MNdX6mnEAX2UWhf9HP1Ff2Bbrb37
y22Gdjt+coQ/4NIJt9dOCQRTKEcBn55G+9MfYcDTKtjBQUbtKYEK/jDqgbVaqEo053vhE80jJ/Eq
iperw7tM7Q7AGYJCWHTrzuDwb7SjI59quqgUyFkFUkXpBRgknzPh5WThsHmllfuKCxeeRLvBJlAE
ksrfT+uY0gy7abuMTK7Qk4ShYGe05QtJoqZi8fdnnhYRmpwdrufZIBEi3rlWADzMIx6xvryeHC0d
rkESTACXLxxYZluG2Pg2Y8iu3VGR+PdKuFX2M1IfFHhd9lORqzwaYr76wG49tDhmGtZZmUA8b9db
Mic/G8FX8H/LtWkYL3o9q7XCjB0JSLKdEmYiSnrYr4hg4RsaDCGs+JsRcEKu0H/fRQwtY6iQ033e
ZXUxF3axOGtisNEEXBIdS3dAlrGuiq9IbX6lNF1U/IsNM3h+1DnQJ9jtTwAk6YMchae9sdcpf7nk
JaTsv57cJLvhaZg5Rfp+2ZRmmmic4JNPaJ2Sya2GD+uGkiknSPoA26CxJ9+OF4JDucJR3S0civNV
OBANmkwRoO+qLnwYC/ebYrmgMVXEmCJ2gUJ+Y+hIZ8HrJr2kdep7bFu51DQRK2cxe6J6DO1uacOY
bSXZnxh16QHnCGVZFQAYW6gMizI8fp9M9M3Ljb8UERZJlJU1oCXom+9a6qTNiSHSHkNJqWAA7KGi
fL3fpeb23+oZN3fow/rkV4fdSbpO/meJ/NloXj4Wc9jV61TGZykvLvHHkXWG1Ldycc0qU5a5mRDX
Py3TMvJpYSxFaNjOBdk2Z9nxVeRDBt3t2ymWJwejEiKNEcNJBthlYIs5Skr5TBKL5zqHC/o9G0nm
F6LMmZGDMcUebXUyME8n6k+Ee9NI24din79IV/HFgjg5clsP0YHVuZ5JH1sB7i0aYmvSXEPukea+
l+zTT9J0jIp1G3pdxitMdyV6kiAQvT1H8Gf7uTQQhUD3Up2iFujnNXATXOUDqPueJ12WoWfb+xgM
rfu6K4Waz9ZGOZRukyKMS5eEhUegBzKEccbxymQe8UW6n2YhJeY12Ols/YDDveQFV63+g/CU+EqG
OPeLLFG7I1apATd/gdIhCm4KhwBO7AB6wCsDj4wT7q+VMD10EWQHh4qtMPkNBs8xc/WNMYc9poQs
54Mz8aMuf8sgNt7JA+8uoZfWjPJJhrcF1JN0zB5qi1n4s5QkFekpfeheNfBK7OJatnLtVAkNP0vf
8MP7Vbozgukohj/VrrE7y3bXwkfNWWXV1WnjnuONMqNG1AbDIChrQ/hgSKj167VzIUvnvPJTXKDP
/5mKVlM0eVbCrRfeInUbTzGKodNbhJV6rYyRD6l1OppuNtep2/jKX5FmhPlpzVxqW4UYDO/iCxOq
l3K8pfVgONZaPuFqsHfqnscbvE8Xu2tshoItrS4SkmqGwG58zLLXyFPXnsxIgUK5VZevZvkGy2N6
mH5TFimhTC76TUtB8Hp9WIwZHsEwqMsenAkzogackFag7HXKYPuNiX107yQJzBsEbmCLxlqJyVjj
Td/6MK9nkXla35FmZ0ul4wPQyGjaxwqrtslMtPCob4LxUGgGNRfp9jYeo8FGkCUdLjfd/yyEM//A
aoHZQ1bssLxDy4wM4tlmUBTTJfBCFQR1/VuDCvSfItaVJD8y1TfsigiVmc0iuZdZchVYaWEPvI6o
qXAV50l7GZ7aoHYa2VmD0DuyPdDfMtKUa2JHt67v/19pznPyl+CLYrW7w4NmHMkskuxEqI2F8MF+
xb8AeCSrhAFkf8DOvIgsDQLLlUPjW3Isxww7j9p7VjjPoyodc2Xw/g5WDJda71pKR3EKe9V2PK6K
O0lTDmAQ9Zcrrsr/xgWNp5c3/YIVUGX+YgCBHOw8BRNnG4Za0fZN1xjHHVl+6AZNIdTNEW+cnY/c
BnIMMY9qofycK7W9Y1ASKzL1eB0bj4PXFGZcoawXLXBYJkqI0BtCHsD5V3BNHcaZsBCDObxiFLY2
6cRu1YLrhbLLcZLrPfpNpJaTosx+mTzjYszA6Tk/jbum+kYPLOENRfGsHdFMoj/6c7Rk7wnie4GK
ZMtoIt1WIFW73I3Sw8Q9I4ZpfZXt1Mz+749awymsyilQwVHQNa0pKVyCr3NfdiVCrOamFaA+XPQF
2B/KWuqThG25EQmyXOeJ7WvzY2YDK0gVkPZSXOov0ha48W7N2VBYLWeoJ2LlErMo64izPXL/Dtqg
B4GZjvuIosjMpcGFYJvlym8ig0dzTEYrcnV+7Az32W/pZzucWOLGg+AujXJ0DSqqBcMQg+Qn8ehu
WkdbNNH+vKkZAd3fBxl4BjBVbGUhuuE/R0kfGAHpy8mOvaD2lPNz6B/qeRKL2EuBNpunpm+Pe2DY
gSzpWeWy3IM2AeHQV6ysGxGYTU6/2LwsnIIkZK+Oz0TdRBKr4/FaSzZwdkYlSLq/z8iCI9S4q69G
GGV814AymkhVeMPTwRTtGwg4bEJy7wYUi9fNptrKPV2DAY2HKDzihxVvbz8t/yBBfahK/32aypc6
ShPDkEm6E+9JN6Ce8wC+fZKI0F/aMwyh/r5qK/mDFulioYMvIhpEBhP4iuaw0Ado5jBKjecP7Jc1
anhI7l57lm0igRZRB41OfKq8WxKYmUjpe+MR8s0s5GvMzsXJCccJafmp/QtnM2Eid7jdrNU263Fd
DFZF+R/NEH8lxALffBhE1tGqKJzRcwybeEJgmRlIIlCFF3S56G/HYf2LlEChxG6b7YGm5eqWy3IU
yCvO+/Zd3DpfGPgQ6Fhk7UAw7tVyWqEOh+KxRTvJJrhyCrOdgTUij35Uvq9x4Vc3JsUItUqNSdsg
heBGWvwY6TFxwinxxpFyVFoKjO9burPeUUvpvCfKj0njSdWNgk7KxFq8ujwom6HTyTEi8yjnOVvy
DM5HK/8DIrHHUX1FkuEJIQa+e8x4FIBt3tsJpmfqSUzSFLI+wx9fTOcuR19w2O49JJ/qPVFh4ZAI
8sjYtqiaFx8Y4Ab92RUyYNgJYEXa7RekRv2tW/HmkpkurAUIIAMRBRWQY+DG2vnRPjpY9brVx7Zy
6LA3H0mn6BZYHe9SdlNk7uBrpe9gqyRJvDk+mjdvJ+2l1iECyAbyPPMMVAfe+va0rKNvDVJkV19P
GSJp0RazEskNkDGmIh+9qNWPtP+cwXsWf06upmbe+cV+BuRFm1I4uRsuQ5RxbGIkzlywyaFejtNH
IlqApjWzB40CJat0CDM4zRIl1myjuIhfzZtupS/K/UXGkwhLi0ZY1KUX8FrauLJQgo9HHNm0kMVt
huiisrzTgH4MICIW339UK0C2Dwnygm++nFPcpg3Wiy/x6J870FPx+IDFloBlddabYJXJIIQgMz7c
ukASv1vKzV3YfQ2un3fGiHGSQpHJpUR4vgMMREd1bXslR+Lac4d2c3aix1gd101w6rxTqrfFME8L
MKlcJ2pTPaCNJaDI8dwaJ0HpYU2wQVRRKVpi2UjXChQNNKbm/cwgzjQRl/jbjFeeWQcxz12eHLo2
QmK3gPV5ajvSFVrfFPdQVERJikSVqNEIja4wg0NvoJedRBtzjUGbnh/5xZ+LX6+U8dPdgirZipJ5
Rn2rmbQgkilj4QQtlof6rxXzW2HmCEPcrQy13sKtnGl3XM55K8InycKMpU0GaHvBo6U9pcTBHZ1d
eeveqpIru5+JmVrsjn5qdJBeAB71PQPqBoxt1CO0bKQOc4yk1yUzIe7MNJJ94eHahCIIWfpxInMf
G5k15OkziVlTcOx1bw+Xzbgu2+64mDLKl03bGXj1C3mII7ISVZmFkiIxg5lrquadfLuPsmnXASLV
PowDFaKrG1qXMOMd/mROTrr3ReZz2a6M20T1TBK46Vu1ke6+MVWFCtASydPOG9sKwWbfg2loJn2Y
l9sUfLKQXmVXECiuuHnsiJB9DPBjqyn+sRh6QYpmJfhn5tlP3QsxyourX12iH4xMfa30m51KNhki
rx0xM+kaPAlvcdgEgakHNiC3nwKjmIqiPp8N7Wdyd2MzbZWb0LbsuCjwi3NROADFTErJg+9N1won
4ZYODOhEtRutGVow954EZcRRYQe/+SsEJyCjKiXWa3esfxRyB7MGVE+9KH5c4kEbts7Kp+ZM9r3K
/fH2RX0IpPQ5Tl5Jll8fxWntw4wc8xnitaFQPp0eqfqRgCIjMrDtf+q1gpQbZdkewsO4YlLx+KV5
vIMXL3wSEs9Gk1G+XHGJ9NQj4jYq4rb39LDglSXFfM8Wm/7d/VBid/fG0S/lnUku/Den1KES3eyp
5P816zrBI1cuyT5De9A4HUIrLsVvwCLAVL+BTSvuoQDM4x/RAHIdDHgsMO2AlvAO0QwCPzubjqLD
DqoRsyRtCGkGZqxBJ4yDQ2DFtWQuitOVRnjOm6ugdlt325rbidKiNrPTAiET1PNtfGdPVOSVIrq+
jfUer9ViexAYAAhX2k+CYS5Hmz5iB9+aiI10aMuX1S7swxYKMNDvUTZZNcnPwFkIcHRfTfrtSLtC
ncL4RqeQ5/aH0y5TJVpK+Rxgdtixoh3dBFowKldV+vdqhyz2DONH1C8OXmfp2DV2QZuUjPKqrdR/
1R074Ec5TqTOaMvgj3yNVTrTLKlEkcBB2GHs1Q/ikuHYyq6chkorbhkGUJu+BWEVtDlfwV1Rz1uV
9u0UUMKu8LeHghC9c3oCPm3jTdjt7cr+9XHaxDhW+MMNQuk+uljnfVp6XmQOWqTYiyeDCrcKx/zA
m4BznYJBYHcyY584Fabk9oYjakXqniCkTalLMxco/8GyWVpTzDjecl7qjba3BG13Uf8BZk70N+jv
Bft7btLBjeYmH0hc/DJCb1ekUp1PVVR9T7wus1nUwNMiEapDzOgxgQ/06iamvoST3t3w07Ib5Ofi
7rD/OBKY3qbfQX65J3pXXV4p/C/1gXXQOteo49R/pGo8oHRr5dDuq0VGyaZt2AZaHAodPjtFz4aV
56l1xxKaUyXeFHw4DAWIZ+LKmHzkKPyfAcQ/yjlzAKOPcDhUatjvxGN1E0RwtNrNcjnDOjKmRD/D
YE/31aLLk5DSY7f56IoLZirASbpLHPyIG+KfPqKDXNS6h8iBwJCiTFTvdjYH1RkeFNJvwWwvqQnL
pyX6jHx1pAZH64KdfPjVQ9/coRM2iuemJRvBIFPziQfVeDjfBwVVAf/N55aVNdBkKx4IMRO+0/hX
lw8Hb8OOUDDkkrNyewiayUCmqcmmdWsRpCRThI2jR6wA9HapH04ZGBl7w2IMoiwWZlYdXpdbwNiL
ydO6QXDQ1MyOdYbA+TAhfzlMK9SdrZjFffkvAwmluDhTRxuxSKOnq9r6k/rtyKvqE39f24oocY0U
f6iMDefYX15c2YGVR2gkTZnCXBvdZqw8wBokc4OTeBRf2AgHtEbIA8A/hM4ZuBrWvCADcZorGqgc
bCiKc+tlx7bweLlokftDctD4MiwtW+azUhv0VgmZPXhtfQWbkRd6qPTHNzcH1Z8HvKyA3OQ8wAwe
PX0SwsZeBZdDFyC3X+aX5TnRMd8PaP1JjVeVOt1E7V422piyswU22uaKnkqedmtfbJSyHo5/3KQH
0yYSHOiQ+Ry0iDKH9ig+I7IIx+LyNvrX5PKgZ9IiM6eSEm9WJZRfAocVQXaUCevEQRspvs3WgYoH
JaGQ0GN0W783pEvnzJfGvncySD8doz7x+HHibjdnbmss1JsFPppSV8PAinHmsjVFOQZTdXlOvZ7f
DYYmyWPs48GK0qRbSkVJtBemujI/1XkcynpwrdP3o0yEcGnRccfGqRm18V8witVlIqiD7rpyon1t
RT0G9QdlLDMH7XryDXefaW11RNRhr5sfos40kU/ifE6p1g0af80E6f9mqzZI7gRmcUp71P5WCcfq
+vJPgZPr9waM/E+hnAWCleWdAO3qdSc7xsOgxx9GhXMLvOhFv+Q3mwwWED5G2UGvUsdmfOMsmice
ZqOzcqewsbySfT4okN+1XDvAR8bYNXoZ6AJqSuer8xKYxzRc95uq/SoaGwTKO9M8JTZn6ecQXGdl
7nPLwb7XPOfY0y03X8x/VX4v2dBvb/v2bN/32Kqm34454KMekpklWVAL/+Xem1T0MjZhEZMeC0Bh
D2uXNrzcEnP+8O8s3r51WGp8smD0oO5trAMz0Z2QuQ8FQMHtyKL3HaQvIPxDP7RQY6nCJ4R3ZRE4
W1ukBKJ/nTMkzkLiYXdIdlvJi2dyeuauLvzhQzB7Ct1tKnNG2Ic0Vfr8IG6hWidMFV/Nl+mcg9Yi
fOB7o+rl/5uCBYI8YTQLG9TEp4dgxTtGWE0VZd8LOAuMrNH41O1pl4hz8YlaYBC23n92jdvKT8lM
wL3Plki+Ri5QiD4FJTw2l3Jpr/FI27Ko0ezUXiPnip0W+OJ5YnfOAOURkMx76zAUK2d30/7+alKu
bk1AUzZtPNMyEOFK5PFUNKXTdVrOm38GB9vOAziJiRykJmf002xGtnq/LZ6KYeeNqENUNX7/8Rce
uC4clQuPdxxTZ8UZ4ae0mtotvpWANccOZsVjerPTJSGglyMWPcH1gZZHo6ZBld/beY0conhyMCUC
hfdnUKlosZcT9szyC550N4lJqRLWQ6AYAVaIsZayLAfKudhheuTrisFc1GSI3gPHKWdubVKh3coe
WzZpkJ5oqNGsseoSTbQ8zRGmcmfwtpy8s75n12Md3bEJp5+pzJO5o4yncFrkZnpWUNpNn8u/4Cw+
nGWa5Ffys+tL1lW0i5FP/XJKDDh+poca6NGVHmq/DjWgZDYKX+WKMlFhLhFxo8vaHtLimDtwCE6S
dki4LKkfWZKwNbxvU/gHFhgjx3HwXV7Ji84+5rRFTKp9NcUhc4IM5nkiOoeo9mFc25PRYaXZZ9lo
mPZfiGh9WSGRd3SEFPPkdBA3zJ1XW7RmMq/Ir9y8/G1T0g9x6jTTXyd+f5NOGGeVTnV2cQFU+v6e
5RSYAGZ7svXdldPOFWRSJtjWD5DJ0/SvosxKURe2OM4TCcXy8LN34//JJA1WK2r98Sk/nFbXQjYs
Zckmz9Ty6UkocofksU6eRfVNMHCBT5+QKIC69uMfIltCz8uR6queXAkQ9ehD2WSolnYs1PVV+0jB
j/dMQ30Z7lugOKiVIZnT1yb4Q2Q8d7Jnd0X8zHOiZB0GYdvneMcF4mnViXZCfD6TG8Cn4bZR/xaI
RAQ268sM8MA65U2tnZ8h2pIH167W7F5UI5x7R2SF5GTNtA1rgBDo8Vv/vVEKgzQsqszXprGWqqn5
rNekyjrK/ZuyZq7YJth3GE3DZE5fUjZkohRZ+w9pRe0NGPDn+6IKdMkZCcSmp1+zA0sZXpNNxmxE
fnXfJ5G58zYoEBnnjtchz2UwFW5RUDe1cs59GFNeAC+gQTfXIyx0ovIWMzQW+Hve0sXqXDldExGx
2/WlqrGrMrzEfer2gPlHd/HL7up1Uc0PJrPbyi3DE1wECx0CNn1sts8UqXH1K4bKUvpCTpYcDE5X
id50OcohQTciIJMvG97uxFSPm85Uahs2yWsimYe3izaWb3BoF0yaJzl7/JUIjZGC+uZPI8l2y2SW
OL9ssyP4GsMlgGuopZrKwI76eG+RDBQ+cSGL4Q3WRNzR4q16evacKcnOUdcChkqECS5wk5r4r9DQ
yjNTbfrO8RqnOzTS0Pi/ibbdslcrT7oA02pu9R4sJdYYikrPSdOlVKJ2u9slQU38cc6bWLo7rpz+
5OK204Ts2MO5bPAT/k6gvFguAT4M9QQkA+R/c8OA56U/Ehz0ez++I3B0tGuFk+CZaLnIz1CZwRCw
mpm3MCRVE915MI3jEj6K3WJAS/y2unOIf56xuFIOndOXAIUcu7Sr1moMVCDIXYI1vt3+10+FX6RZ
RgW9g/eJ4FFiB6e5D8RnVnVknX/EeaLmZ/3OM7Z1MuFybB6yt9zSxE20crGNwZOBtHloHQOhkieG
qf0h2dS6Gw92lMJGbaeGYSrRROvjrlhsbjErBcl3jGgyOV+SQIkSkFJp85WKQjuFPKvpsm1gnuZi
uoz0XhnsdPwRGtM3si7cGHz0pUhOw3cZxUVQqoBlM34v8fZqa6MDaK/CzxLpytX8kZU1x3sUcAIm
mvvsJGHVewPvKAwT6Zw0bXzaA3FCss8hdyLHOzG/xRCCEPrxVQuuEM5ruydGyAgym7bb359D/UQd
83cpBgURK9RkJVj/3xI4Cj3HwGE9M+AbjJUgrZ/dvBPvwpg5tIFSwDh/0xvBFv8OnPj25qLj3etO
9kqf0hfSwcXZ3Q/lSCgGrtlNR0kyOS+PzzfTzCJUj51unqVSxmhv+h5sY9mmdyz5kRMarralSryg
0OL37telEvFRjZ7QQ8KivG8st6ggOecnGQ/crbNUyoxIFJCp4m2QTpezrWOa/F6sCsvWjFAx79pZ
LNPEVIA+j5txQQedTBhlZeUmqI99z1jTrI0WmPk2niJmc49/WvcOmYv0v4Fzw9xovLgZ7eC6H0V0
yWA2UuI84QB6VkNzOlVaXoa4LyEu8LfUDLat5u+VjVX2VmZr60o1QzsNjl3Y5DTTKEzUkiv2SmG+
eQo95aHwtDU/TBNdmptswuMiRedf9Re2gBFIw89WPoqngYfMnaB2gN07XHq9k/z4i+JWyBf+sH2K
T+eOcYbyGp6Pxzr5ekH5+H7Cl4Axgl6stb0sc2MbLDfwdIZUb15O1X2OdC8Vsk8QldroaeZHEq07
Q8eizZ+ICUFiKKa6guyc9TmFhOKZSXmW3yWdKgBYJryrBJEYD92X+qL6d3bhPzLC0AqOvERIMhdQ
1hPc64eIAbiPjm9Ur9J3bXVEX17gB+qTbEtD0mfH/ep2/2p3g5cg1PscfYQxHSZTn9p30h4mbQ1Y
xdlJzEIomM4rfrHen0H2V7oEabMwbaJ5xVa9Jh1MXzh9aZMIlICC4owIbXzXPZTdZLNjQ6u1U8ey
RBT/sF1NODcHcGfuhuSav7so0/AkBeF1HPf7afGA+vLUBz7p/EJEQmYBYsTjFcTS/J8cY733qL1M
I8ztj1iI6OqcBTlMwnba6OnMj0AlDMq3FwF52zlrl2frhZ+L7diQ4iQYG+RVHBPJp+SGfLKXEm8m
vlIlUpfp3CQ5bRL5e2qN1/2SuK4BkjPzhe/JIRynq8diDy7Qnzf9AkAPnaym/gBoaY+pk62aIrML
Y3fBlRDB58k007kv5Ztvwi2jbFrJAfuCt6fTBTkqFhw7vp9cfGcb85GDlQn9KBr/bNUgUztRIX+B
tiSvScil9F6YjjBxk8AyAIEw3aie4Yyn5YPHtv6IQpJVQ8dlGvjdO4DQFxRaQ77Y2J4/7hb/g58O
9QTRsWHVkzHDZCYZLi06yDwQieKa1xNLLo/fHOIwuHekd+aGhBbd95EkBtyP7lhOwCQjXfsIdHoD
n0hhDngHDpEUbZsJfh8mXMfRLGSeIeWwsZrqhYeQi4oa/PH3UW7wzm2bCyVWtKIzoiR6MW4T9e1h
T6H/lqBMHq85dMV5WY+OhnKZw1rLvEkkTANKq27V7KcXw0JW4kEaz2zjkk0m3a47pq5W2PnmpVe8
8E+E++AI7a6CFQa7lE0gtVqqA0ssBfwJIKwlVFF1vedwZWBCOwOfJMmaf6ZU54ickKhhjVuGDMgy
pcQiJHxGt0ITDozfwtU8NtL78z4qnSF+UsM1YZgIbbhYk/aTlljVIBMzmlYsujmdIT2y9+9YSLR+
9RH31XVOxsFF/OpmcHXAcVTymzR8S6Ir2bO1OUloHRMtqiZs7lVElFzNuUjr11NPF8tR9ppCstXg
bF8hEq/Or/e1+WltccyPsbhu02DaTzaiBR42sSu7/XLvbRlqeYI/gzBsSaOcZW0gpHcFFxYXfUvd
r7ScDOrbFKgh6JDNS6PWuyPUDR+uMsVfdgo6Ana+7xt2dfIc6oPTwNJc0PHhd2PPiDePjc1NCecu
XYD0s4C7jM5eh4Z9KNecVfEPYb+mWRa5b1RI8L/cDfcMIJROcpZ/1h/l+Mez4yK6//4ZW4Ap1RO/
uXvKMrgRHKP1pHTO4FlMPk8fZvh4TTomtvkHqFal7FLzD+5O+M36Ov3F5iGE00DxuyuDZcFVI87c
q3ob/HckgFe9QB7SxIP6hMWi2Zb95+GBb8rZ/5105T+FDRTKagpOL+Es40rZFEzXlyPV9rO6tc2C
gt5MYI4SD/6BfrZuJ1o4/drCKnpC2HYBVBHEiSr3d9obukJhB/8xfNeZpIL3xO9ycg1CQ4/e1eQ+
aoej5NM3aNZ2v01r6A76K2AXVMsCjhp04FJcyH4duS6IvODlC0bEAQg2l0TNithDQGtPKq0enS1w
VYJxw+kkmQoru4TOqPT3c+jxQIFQyMQL5AlqmB96LJS6K6Gm0Dj/YxrP8ZVWY5pdPXSXqyO/Lk8r
f5jjR3jd2OFHO7p1AuNCdT4E7b4D6LxbiySnbYCKDseR8GtMhvjZ3PFX9ySJwAaR6ZoUDR5JDcjw
J9FqnbpLogFuFiOZ12QNM7obpn1Ic0gcIDcv2iatmZLLdZq6neBpqkJExibq90Jn5MOelG4vDION
dZUu+gwKjA+Kgcqs5wHjnpDY1ukYLVDRE/9vggEtz0EiLOHsZJW/jz5nYCLJEJuj+QRTIhJpMuIb
b9qRfu/rkT8vLvIir/xkjo88gq+lOMBiG8rlkUA7HQ9sHwBfNKntm7hClKvxjuhQrudWvhi05reK
v8dc/JwEcB3QRVKkj+GkaBcCvu+jr4cR0tChofzDCBVhjId2hQpoPb+1xmXA7wqoPTvkxXn1NJug
TgOESwIM0SqLqmsHtH6i1F3Ro4NM/0aRxp6dKOMVZyWlAlGk/gnax7YXEUSpDGcSITg/fbXWgz7i
guBY9LbPfFA1/HVgzbUojet36SiopMuLTmm3zcOZZMJuBFFyK10KfKINujUIbVKGTvZHulSJ3dWr
+FSJcf13Fwd4nvdAyi+8vzZv3tOJzHEekfUpfyetcO/3F3LH+g0UuaxyxH3OhgxXjwlvZJavV4ah
x55xSfMa0kE0FPvuLPenGkcf4neff/5RfB0kTTps46JmHwKvif5pwqHoWcmlzY3pecUCwTMBJRFv
hZ2lDWbGZ57xcOtejBmqDfT6FTCP1WfbHvBwDLXhHNYUI09cynkPCW0sF8w0vnwizWhaAzRyfoPa
eu+kKqxs0ZUR0Vb/GCcK91RGMbjbyjQQXE1o8eJXln7c8U+CikFDKc6ZZPA1I316KeDS8zpCbHXh
ul5imao7PtM6c1VDQck1JAtcgFrhLgraSe9As/CEk2u+YaqwL2iBZj6+slN9PoZfZP8+rNIgvkPR
HsGc7+ZAgb3MBnlCxU1EwmRC/mQtuw2jWeze7VvNrLE4SxegtF1bkXZQHOk7D289y5BcnXBLXySQ
s0qFLWS0Nz3s6hWp07r7mF87lrA4mqjRGD0PRhZCFbGTatJfgFGb2HhmrOUvbSRE/PRoNw7xmPkt
18poQ1QDL5Xln1eHTiIhcye0gHbBq2yDRX5tqMvsCARh+0n2FfnGTv65ULgLz14+BVNThuaK2FFw
lEHF5ieFumtwO0gbhERgatB7BlFQDtPg0KiO04V9NyUCd61D+KkALkvla6+PVIKNXWYOR5yO0S7n
rIq9OT6Dbp/5MUDFB4TaMokQhHMhjBWk5cot6HFpTq6NFo/tBu1V/Kw0U26kCbY24q1sPBqTeOEI
Ck4lUQXYk4xCD5vvR/8t3ToFzvMQFgGYMP6Sn8LP4Mg1rluT9DeRGYU4vM1X1OElXSnasba9Xx//
QagDW3uOUqsZf3zeKnYZqHPzRBVaJCH5y6jN9lwAp7P29QBLHxhZXPLCYYvTL9AwZvaew8LKRAzH
XGhIOBfOc4ze1xkZhUikp0jtmqGCGlYIWgq3R4KxdK09bugTq1aXlUXXAl11ddOBjkHrP2MiOFqH
HQ0Ddws5fElrL4QiTGzyqGPswve7yrQLTPwxtFzpDNviUnMo1drMQxketnwFWxnzgsQg7kO09bws
8DpaEdm1bEdezI21A+RFQubIqwA3iG8lYnuagdEl3h0GxK2vt4sSDlCReVBNIYML9H/Urh5Y2MZb
duZLqgxahMtGJe1IngMc50VfzjOr+6dTuuZfUFHTZ89Qa24cFybYio5RxUZSN6KY83zqk9lIET0g
L2ZJmudUG3ad3rVDEtKmXpfW/lAyr5LrZdA1aUy5IVRLOBicmKHg7jUrNZmsNYBn09jUNH41mm6j
YWp4JDHgOSym7xvbyzK/a8Hfg+bkvDAuGhNfhmhpeQakZ+aB2oBdMg31hwsD+6u9tKqmAjyv+s/g
nbb+vRdbzPw3vPlpm0+/iflWJuWLpNTgB0T8vT0Z2ZJh0pWzXcP2m4qR99Iz5/cXmBl0dmYUD95L
Goy0Yghdf9olwANPAR/PnesoRhERDk1Wpn3YpoSK2C71fLI+/9CSU/pldT6oLw9/K8CNQJ0+4dHK
eTXobBPNexT6//8apyOVM3ZhAu3dGbmSIvSg1pLtylmmjM6rPfvw87NVjIJ9+Rifbc0JtYMpR9h3
zwrXdwLUZ49iZCgoK7dW6/SYE/Jd2Y90IU18q5iv1MpPTxgjQ5wEATWLXwlrrh+Iu6kborC7pQzn
elXAJ/kLoX7p1UpNt71+ZVBHP32W62sKF36LCHA9tKYn/0R8P8XOBJr2reWN/YC+y/Z4oSYfDApx
VKg/bM/+2++1cxTE/5hdrvucPOY3jOhPaUCHBWQDPtcwpVU8I/jPJ3IUcDUVnd2dL6OhXV0wayhu
Kxyp6sgMvnG5eB8HKRgpwxTcLpUtBacsBQV57CAyM5F9pXUu5lcAFTv9B4B20sVa6i4FvscKPrEY
+o+VrEbErdYC178Q1V3zL89tEHRvSLjEWE2zEbgnso+9ylJGXrhkcD3V3q932wybzxbV7TKTR1xr
O0RPd0oXs3M1znsSj9nSQbeRl1oVpqkbfX35MLiL4DVZu1+tGxVf/UkF+9ZqnQQBOKzhZW0k0tzi
Mr+TY1/vuTpedZK6Jsoml3cr4gHoB1SVpjVLiZ6l241VQI9M82xL8ebhwl/RbySG1c6sHcIq0qRU
G3g1kGdPopZOcYCZICmYNNsQOsuUuHLHVpqJ4+UK7yjA5mCRH2WFAkCSZOYcKG7kMvZr0By4wyf9
aAdqctGMu1cfC2jdsT9TPErYVaCvHrtCI7ddhm/i4y3P9PPNbZ3Dcafn/71TBdzXznhwMweHAjh3
aYu1QvF1pNNXZgReQ7DEZ31IMI9Zpnez1xslC48rAkRuwQBIqo7siR3ZpklKmQyQzLeqFk8QeoNs
Dw/OEL9WbigHI8c+zbQanJBpdkjrPfB+oU3EfsCgKJ8Vpdri8VFmeqLUVMZhIJZ4lqdOFD5LDRjp
SpALNpwvZjfELk238I7HnPsK1s1hk5ONdRxV/mGN8ltmQrlWFofMWjXb4B/cfBuWDunUAZ3cNN7M
Huq82117TenBpPfNd4I7v21jkEtii18SMxI+4kWUTIUw8nScGVZGovEOGJSvfqer9HwgJavOlMS6
rm4+UZRavUEiONDEAYUMLSyyxaL4+XmpviWSPULSwgiu1L1Imb0PGFi5o1ukGegiVUbtdZa44f3F
PLY7nMuAYZGsR6vP7nQdX/3cMJh8z7SoHybk3vBAZIXH1xIXk5dJYzqYaUXxg4CZ2Dk3tIRMZuLx
Z2arV8+ds4CxGZ+QGDQIWfJdSWhf+mNKSbdv4FZuOBwytn9q8o9E9K91cplKvI16yqQAYWqBvWMp
zzMtoQ0MyWJKM61c+pdZwR8/4AgBo2yt8f4bH30fgB055kJDo4jHaiT88ruNkCahKoHNo572sIYi
ghKTWyblGkBeiAaMuZeivtXoFaTZfetJ5zwOB06F9eeH59R1dwkJo472TUyIZ3G6nXbFvSHfgOjl
i97s9fCzWRHH+E+heCqs4Hvj0qw6dG8b8sLw4ApA4Y/gW0HseAH0OLgF7uywK26xbM5iGQIkTGSX
Z4q/2TZpB5YodIkC0zbF5u9aNy+sT8j3kXP1hoGGU82DZdn+BULf3jcj2Eb7XDHknDotMqCUGmeX
5srbukPaXrn6HHkvx+dg4W60JBexi7rZYUAkkBEJ9qxSCVQLaElL4dkVmzVarHFPhNVoPyDbia8s
36O+T7r8DCDK9PADWLMBOPaSuzVh1f5sUdYyEsoxT5SfgirAEXgves9f0MxlRwr2JImJEHRFsxrv
dRMHfteL5oHnS8lDhWS8ZxOhypPApbYs7vrcmXzri/ZkTYpHZTZ2g9LNCN33NAtWjPKCUzELLdUp
jJ3i+GK1+DdFvhDxGQZe3nVsy1XyAI0grIfJ0mfebY7kG12RatKXoviaV+qXR3z1K0F3T01SFRb4
KwdDbI+1T1yK1H0gyrVL/o7VlF8jT0+E1oeb/4slam4GGXoX7fnk89aeSWujUnkB/pK7iTtpeodx
eFats6NzHipxtzqD85kQSRM8u1Ph3ZRG3hNMy5G7lbYiBvliYuP3gOQQbkLMU6HnTRO4UOARkgB3
BRyRVDDB3RVECMjxZS4Pw7hkJWORyI4+h61+VkNi9w5R0pL/QL4dfh49s8hsTESTr6Ibz4TEeIDq
iLiA1+OMMS3e7/Qj9LU+MqMml5thQKfyElT7sMOkLLDPbSB9Eqnr31yLLukrb5aOspBAzLqJL3o0
F7zww8to8qNVvG2act46b6K0iJ89leCZWYvebLNHUpz7E/BODWlovGQ0gIB3CJ1dNp+nbr/6nIec
rjpEyq65pynGRjqeUaVmGLFrHfr3dVTaCm0zl0wtb+SySOSsdhI0VIWYgaq39ePJsqcEWopVF392
TnJDfOCbQ2O4ud4QKd4a2jn0MN26GDZCHp0FWtYneDrsATHkMO/VuXngoEjInfPhqGPmoWYpi4mF
IMIjpkIEUq9BM2t2ZxZzMn1SfGWIEiksdztmOw9/h0sBpaExW6RtbmBQFeYHsGRv7P/PhwzoL3tV
5ac0q/w+pZz9Hoze4JiblAI1fA2bLuHppOlqv0akXC8fxwKs8KaPsv8G4Hy+QDneSkOKrAcT+RVT
EwDvFYZO5BQrdRcZZ4PjLKIojY6YE4OF0XyD8yOjjpLzehRUiFNndr/GknY4wuHFO6zsEnI1u2KX
ZguKyXpK7JDhwyTI7F5AYUPkWjjB7y/s1J8ve31DgYHQrMZZAY8BIucmp3u+1lLtmLVKpPi1i/W7
4YoccNfbRmVUwGYxy19LTjbIoaRcOVGYCMnRTGcOeYq11BgVif+Um0895xpzpZPBLLPHo+2ALY0z
uPwYlThFEBL4vCdw35x+aUC8vh0wgIr7/72BM6S8UkzBSucJacik3ZghfWJFAUBPyNksL/uV+/Z/
Ic9/YZGYEi1Aay8iyEHWG3sJIu0Dki6TV17xboceWqTlN9zi/SPAhXy2XPE1hMPqpDRgHKLS9P/2
l053mghrJtsbMkLI3tVg52y3+TldQAkqcNtHCeRFB4g/hp+2S72+WQ1b5hoRpXbQMcFo8ww+HhT5
UkYffwMtt91Fnevh4SrLl5eFxORTM8Ku1I4j+2OHcU9XK5eRVhuqt9mYGInMAXlzHl5WwNAMDC87
xh4d/i0yAOy5sibIzZdYp3Iy7ydp8Mo0pwAW+hNI1O2RNCCa4+E5NKkeGpMVIMW4Czp+jbkFq9ZC
+MYe35OMUIGW7flAJ4kfB9XGQpTuQi1RVqmUiTNrudUFgJ9St2NWL8BrRE/1uxFr7qLEhFAzy6Sd
cInhilhCJf8Sg/KyuDB7ZC5xDUvA3UzH9nE7IWHVKnUnQTiyhhKDaeRZj7VUcA+eFTi4sYQA/zQ1
tOQJcwZvuCkKmIRHG2jD8poO0GjbXpBceXbvwocbCLAsOoPfQadHihGug3rdkwKaicXqA3EXeyqc
khfJQgfJpDxfDnylAM1H2704Xeoc55OyAKImZw/RNMtEpassqlr7Iv5wvtD684vl9Bicgh7+xN7J
HxVtlN7aGbvkZp4Er/YzBC+MZHGnyErjMSEjI2ClwwBRbhqgs2Fv3a8XkJ+ejhDn6bcAUYOYkYKN
ttK3W0ICEaLA603CXOEI5ZsrA6zeDzMUdIjeIBq4kbfpAPTSkKX25xghVOTCxEvcubE/6wMY6VL4
8pCpZQbOjAYSIDCQbuT6KbwBUk9QPf/FBheUFn9pv5DTeWE1738vdPy2rdDsy8uiVJvFYB22yVWW
rBJsR6wKfscqeF1456HPbninvhs3EdvA8SkXVkHc8nv6DYPm8aCmI/WWUz9GBezdFnsbD5C+EfQq
QwG0MYoamAGwbLJpZOOtDKsi8IZUaIEIEP10gS3CGrJaCvuzqN+J3RG95I0psoBarXogEiUyclzo
ycfz9Ke3vNe+XOXNIFlMeuIysJKzNIOu11e9Otetmf8Phfvn5/haEZ+Bc7h3bR/EIvh5dBeh6ay7
t+ab40zywYdinWIuxR6/IoPcag1Reko2TooGCA4C7E9fDe6SwgmIol2r+P3Q3dCX864te18ikrEa
9lKFYQWBqONrid3jKxP/73OqSHToh4TF4xQ4rGM7E5DJYOEaPccFu+qeFTeD7vVmbwjklDTzIDAt
eSIOcgaLFjt43KzsXI1tjfOP92I98IEtMR1/wns6dmoO+kk0id9UgIPwnscKUanGja4UZ9pcmYTX
x/WGIFPLTmNqCPsc/yeP1wexFvbyDFwPIeyn+Qve/Zb06WZlXjIMy/+Lm31tY/nQEadoi6S51LtP
srpOfulP4U53jk9pGXatI7SPupWs83zRrb8uZnDRd+7iLlioq6dEdHlikpBQkep2IGGgryQu0Q3a
kO+JdCzYKrtmBOb6X/Y3kOIYmtpkV8Anhv/9vlWPp9A2tYih+5DXf+UYupn2xOWIDNwn8fxzip8z
zsOzXnDWjF9OcvF7wTMt6MRIuDCTKv5+XEIQ1xFEgR0i+ykuPWC7O8Tcv93yu1TwHWD6QmzDVRFA
Z4rmyvdY9lK/p9HkmB6ycACIan1AElluYVwoAqBnnMiP7qNw+2ngZhs/WkmCF1sTOEXokTB9WJjY
EDnP5Jtd3f5dySyDcp7jMTbZYyfTcG8jXchA5svAwXFSSqOrCMIHJZMUfSA1Ujw2McMPISBbNy6f
C5f4ST17ZiViObmPF3pRGghT7u4fGVoE/Jf6UNQAcStK3yPHykhXjErDXf9eKw/twGnJNzrEpNaG
pMnQsf3u6xtUOI2Ce6r9U5TW/fkQgITWmYDgfUET4EbHM1kPODJPCngq6WADDDNcBBhclVDrq2Is
JMJgJNTuEG1Xwk22eUfNm1gbo4XlzkiK10EKZ4cjFRD84MVnQp0Nd04Mai6S3je5zJ+o0P8xxPga
gu18CbU7qAjF9BrzLcAfyId9tvWs3gnBqJpLtrjvbCTNjIArt6si6KUaW7Y/h11BOw9scwLixQyJ
EdsOd3S4qgZ0lLQxHGvgurcUGjedmPF0DomGcflVcnWXCk4koyXZTRYbfYr0lD8M0SAGY6RcSmBA
GLzjr5JtNupcnwDJ9m9tZAmjUyBZ+O8/wD03c/fvGwS///Kjb8WuwZXE9mx4oGw/zVl37SQC+8aC
bVC0XJpOzriDQl7QfunxZqTdi9dVmkfTNZkMxaRnkGBP2lcO/4Z5UnDh8Kn9TEtXQq/9N+f0ZuMe
WWxOEU8Nfm+sNkcby7rNIcve8bnriZeZOWfG80a2DBrTwFB43xwnlKnSTZPGoKvxnfs59oJt2yfD
4gVaQrtzDBEFbUv2tDjfDT+vOwj0ckAeQJRI4kXvuT8MlyG2Ht5FZszNXMOWaicKwCAQnJ5kqYvU
FGkdx12XFGnokt7oLyoEjPq2p+R5cAUAFnUrS0K9bkVaUBCJcmrh/xQgypkpRU3Ovgu2UzLPbzMh
HPSt9MtZpIwDgApQm8yRDsPz5fgRq0g5dIQ9IDpbelsEh0usdq9rqjN4RO7z/CWqB/Wmvt/LLbWU
yjkZxsEChvnsqBszO4APhkl/NexsP/cl6aq38zgHgyHYObvwaQhW1oPNPwlbMyxjnhwVxluogbIP
DHBVjJ9d1yNgVRfdg/OyD+wxgvQH4M8T/3S3Paogm8YCgyp9KKFzRneRXv+Gedj7bG4A+g/RUPIZ
Iqp1Src3uW+2KkAlTGAre7xmcvYsgqexxgz5kMKmOogy7g1tsWHoZu6TYQV+3aYzoMu2qk0O7hxY
MyKvmQQuUa3bG8yqtPpwuiAn929VTYIjY5Chg+W14ky3oFdNlClW2WGQioAC2N3AsTyAlA1lk2GO
6ipe5Qo+ICcoJ1PSCStVd5BY/+o3oGNHkEVHQlWKCBLMeCNY2LtwNJuIG0DoNwzT/qL2KJJw9Dyy
QkqS2OcXZYnhkRgja81pOyHJ/FzwaXXvumLT1yGX72T0WRVa/i4Gs1PMRDOeskZ5p5LwYswpCJua
a/BbJpo9bRJCMdiy8xG+CLtXHp5ft/hhm042+tTSfcJr5TfExTpHRBMlv4uJuFlKsuxtpeHQfjLE
5gBRO5pyzm/hf2o9w5pG5jIApIzYJvw2lHH5kqBHtM4ZPvupV6d6DtSUt/guCVVpT8mIL1xyVt+S
ndG/44JZEigv8BJ7mFW63AF1TpfzQJrpE3/qN24PcdmvmaXlk3f4WTm9vouNzLBTlOQC/7hB5ukR
5YYG9NwVi+BHI1O0AfZ2xZ5Q3Zkgn0Qj2e7fw7hAe0t9E3HOvYJQQdwnrL8MxeLjHEHO6thsiyvB
emIhoU+UuQxUkuT5HN+xbBU6Exe0loH3pBApwPFe+ka9Vrsgw/gg90zon6l0emlbhY40MyMbcr9l
amOGcAcwGdYitzFkWxkmKsCB9K/ib4i+dWAOyKHzkE2d65lBZKwYt6Osp3WL59DVObPY54semsyx
vkXVacaIRrzRyUBKCiVfZTUUHI8e+axyaujOpqUvnonUQ6vseffPaUKKNFyKCAWpWpWs/OyMZca/
qhwwx058jWWWNzYs8FWhKnFXAZEIHFJhGln4/VgGnNVUoKM3mTloNRyj6CxRg7AyL5iGni0mNUrJ
FaV3ycNm3a3soX8lwHs++JF/pvRXMVNmaqOr/hXO17HY2uPg0hUN4HGVZRarW7TC+eUnPbX+2kBD
f6A9Ui2vU2TV0MFI2nntM6Wvr2y1jKworFSLHdQJ5W9pcyZLnxf6NML+aqoXAhX8XXw8vRX9CNQb
jqWxcUbp95Rpy4Gi9J3SNSGt78zeuI+IfthDWHHsTrTk6047HF5DXwY3SoxlHoiMS3GFFLEbW3An
fu3gP6xfmUoF/2bYi/EXccrbMTYQ0tMcToKp4DXsmlPpoT7e6IGhIlN+iHlELvyHf2CL6Gaktywp
H5vNgn8HpozXJ/LkEjE0LxglDBH4YeOSFwqqU6+Y4dOQKAHILjpBaHS/pc1mF9ebYbnabkRkOpwO
PxlWw5Cat1sdsiTA2Lq6VBrq6NgJ/8u07vL1MXZHCOPGht18Zzg5fEz34uy0XTWTIlRRwqAjLU4D
uooQkOH6cCnux66YcO2xmQ2FZE3zR1v46THJqi77iwlB6xHdJ9pRI4epqrIIwtbSBqepCgVotT99
YDmlyfASNKkkU5HwsZNvlC1vQZ1QtKZtxecMrUKqvsEIYfDdmSPmQ3MKOH7PGkYsgf0E/H7lhiM3
HPU49AZO1yJCSnM7v2XIt/FtEaQ2nyplFRzvugJzNhqjiBEjhznb0WP896Ug2KSGLkWamWTejWsZ
yB7QaGxsi8LecOCT1sPipWMi75br+KWg42h9g8Ds8JvOnHEuH2fvkVn+YZm6P1LGXRoJFGU/24D7
VY5xUp4xhkSWKa/bx9lXzCxk8KUAWMw4IRq28Vk3tcTQYRmwS5wTqYVDzR+nweApJvIjEr3OTeU6
HMgoh5Wl7zhKWiYGk4fFG4zbFRQ7F6t6aL48z6Dr8HvFRh1V+Nlpg5X5amsnrMCmALzK2+5kQ3xe
2rtsCMxnCI73k9b8exuPdkKH9K9Fjhs9r0eLJD45LHdzGHyfI2H9mMAKa3lNm0qew/br1ccyhNh3
IknCz7It9PCeLdYxyiZMWIILrnAhWAAO8FFMCvo8A3GDeOZbr/IQkH3NEJoLNjRDT94jxK5MZVGK
Me4y26EHfsio7XwgEhy5A8va1YXROMFWpjDIhcEQes3fk50jutT7AKT5xwfJCQIbKqDNXlFAb/yY
J9n1Y/jcq442OWNP8BxLymEQKf/1U58UCoXmG6hm+aTkTDJ4UbeENIY57/ugzV+KFFWgSd9Vl5tM
HittATf0aP//uKXUxqfwP9B59LPtGNqnCnMJDsaRkiL2Nu7+cyXamNVLcXte09iav7JzmC8TNtn1
IoQFNIUKwU7v9Ej8IkXHusiP/pKFU6lXVuZS9jNENnP436ye4RJoYiOBUXBixGuOM3bNJV3wvbGs
R5azHASRKm1SnjMUOz4DCRTWjgXJlrclvmfvUPnfTvaa0G80RMI5PHMyxeFI2Cn/uYEYL51ElMdK
5uZW3DTMM0W6FEkXBMLyMqWo//3DsG2XDqwfsau/DMENRhHS0V1EkWkOzspNe7/ex21Sfd5qE5Zj
lhWt4/kNp+QzTkU7j/XWWd3cEq8sXQyK3DL6vvuukLREoOw9k0oL8WnwCj6MfLcGlvJlzbpqpCIZ
DlopMf/y274+GIfoqOLXrzBxbLLSxjdpvlXRbFtp++LMZEi0Px5Tq+vHAW8UHotAPjZzuP5DPl4M
CsDZb1B3zxgnFFXij2fgG79mFhezULzIo1aJIV6RnAZ5jNRfDxskK4nawkWhyPvrAH/yqXD2V82g
fda1zgVk/FBpcFaqGn8RvYoeIjdiwjmartCr0hxu9NpoJokph6mPXBwjDjPXbQMPP4XqJKmZYq0D
ffz24zG2wApWHTXdNPBo/kco5a4t2eYI0vmjlj7c00GySO/4LOoqMPw2aVynIKiO1fZv4YSLMOdf
y9Qob1u4AWEKcdY+QenBCYEIn5C7KjvWxYJyH+Ivh8YZ6rk6WsC8SWmj0hTM7QOW3JxyposBQKCp
LAOGlU7iB6TZOQQcQ9DSECqpf+aYMZDXjk1NPX2v1OvKMeloQ//fydkc1sIqCKQzqcl+sCH0eLEd
NMVoFfCuETrz7MaUxfjdHnHNPmOBSyftfdQ+b6qAAqbesQkNf56ty9gNYfxBsKr02Hg9QeqNjwGh
i+F+wNBj7exN07gfybabAjIZGTPjYvKl4uM749Jh8XmTN0i9CHPmL0/mzi4R8+cp3G6A4V+QQvRe
nNZLfa588mIPAkZWw/Y4Ef7kbPr3g3t47SajiVQ00662n43wc7BmfsyC+Omv5EFIp4PwUPHM3LDx
Yilhf4j6GCQi76CwrZ7mT2KGf181WISZp7fmytxNbuCBqkHhkIGJvpEs5woNM+jl4ojFouG04V1U
mytCbqCkUYTsFa67fWTzfOTWxMGjZwcEVUKYUUpdLEKYwyt+T12SJ7rDJMXSjgf+qA4hL+himskz
eaR1ajG+DrtuTN9XS6XUL/dOEwPLt9t5C4BFKpJqsMcsEzo3myJtnjBmB4KBQkULi6IXsbXSBKmN
PpUONW2tRisUTSIeHzdGZLRK7lppNA/6IbBOXZq66IZxGZSODdA4AQwWtBpHTafgqOsWPc4nnZr1
/UPX9sTtwhuhP65DVPoJl/frimGbMt5ogtxya0+xDC2Jt/jFr32mNqYA9Sk7oCgsrqjg14gEkNV8
HOvVaszrv759mIYuT2P9+mRUzAINBWPY2do1GZMg+VW73ToZB+RIdcY8s7LXuOFmReNqQyHmcuJj
peZcS004oNsXnBgapWIMq3v5FKLR/32D7IJylEEFIQOd/0Kj3xdi4eWc2wFDacc5LwOLWdJskvg+
JyFK4rfVgQ2VbbKMjbil+MJTyzpW0HgPC19VkPD3sRFhN/Jtm8P9kV3wwfJpeZHdh5mp62OzG4ts
fbUiJZ62NbSy9QB6JwLJf30jWMxHAEH8Qx0uWPAp6MHYrYjLhBlzkFHDhkPOjJuGeozKT+2Gbvqe
1xu+BMi9B77/hO05BBK+qu8NIyX+O2a6Jt8E1pAePOkOugd46e9p/k37SiowSKefrbcIuZwfhifG
2bqlyYxG2w1nBsczXMKer/PXFoY2zcdmnej4VbaOusBiry9j9wAID3XGXbvsbqRvT3qYvzwaYSw1
Pj15QAogpPevALzKM5QZ71VDQPHby6uEcAPKSH9kCjy+pEAz+7qsBNMGJhWhA3X/bVVkSTWioTev
4O/rUoL5hl6FK14bOGAZvWOoS97mLFGH7Com2f5P7Ox39dstJtPsAWkpXvPPaWX5WviJ9DMyrTsx
naP6V7eKiFZfAc23EoyfCpNi/BjZ6IYvbzeq6hIUg7l/6wx875ABEdY99R1wtE1tE3QAbZs6+ZKH
MezSWC+ON81lDl3XK81wXeYjrARHYgVSxFF9vHeE9Y1IASwQgNca0zCXVn+Zm9CM1MuOhr9mjBsI
SQKKOuClnAjcm0SrFAOlWDP2iu4LqQ4CJv0u2Oqxnitk2kxEC+y4yA171wgheZgdEXHyJgBLz005
EgSWhJTkOd+OGrdfogI9zaF4qCigbORXU+JsNZIxM2ISIRc3FiQgMq98m9D6IzTWzoWNmdW3+l5k
VqyyGgffEuO6t/LNxGAOIpDn7amTOwnt9d2Nr1gVzIzotppvtoXtmnzo5Ls8jZAuY2FDwOqfcN7P
Z861JWFF7Ejm6mFKWmsfhqJk/Spd8ca9DuB1fhaRkEcHEtGbbWXDvQ/TcizyAVBXr9YCRglaNRi2
sLAyXTP/7N1mvCjYCSNnvexXPnnpV1+n7djliINR1mM/VyfivjDM8rkr3j4WOxM0jUUBlmXZhcaz
783l7EQqA1C8AJ2ny5dCDMZEMfKi+lhrUC5ctLsDizRBUbkDfT2464aNSa4lnCT+skKD+oyMSB28
K9GvF2io5p6niUt1XORfiEhJJ2ELViqNNPtq2I/NLfJDZffstesZCHThRLCqcm/hMa4ImOKs3+8x
NYv+qeVfs1RZQDdv3OVkpmgiu4X+8UaI6XExph/usj+L9jec53pUkdKDGYxlCARclMHOiHsZI2GL
ySTEXsIxayWTsgKlZGoRbMhcTpqFzd4c6U+RDtzzauLnFDaqdOIzmnlWtxNOEZKN0qXQXX90pWtd
jNer4Dh5of7EHwQq+tgKZ7pnX3xDH0fNoqNFHXVQFFX8KSw4NKBPzIMufcBJShLPpbJ/vjXjdJO4
A9Xqt3CsJbI+Kkcb9JFQGvw+yp9sG0vz0EXpo7Aufi7/0ZHt2TTSRKZZwRCzH48i0Rlc6B4thA5I
4o/d7wi0axLV4iFeIYWd7gRdac1G10pE17TV4mwHCTDLaa4wYMVxD8lt/GBiC0VhrhrOhpzR0+r0
v06lPzdVekp94F//+HfR0AsqpSs4u+GXoUPDdiAiG8tYGZmgRjlMHwhKlN5ddMQBTZZMoaIxc4PM
1QeVcjUnkGia2F82Nd8LwvO40iVeZtOEF70WU4arXnaMY+DOca2+3yAO5UaSYjVe+m7m4bSDs8In
ombOKlFKv/F6k5HI1Y2bsT1MVvCzlWK1rBsvsDMSYPaKg4htOJ70T88KHkzLiaN1WiJH02K2qtQW
zzXYULTLKh0TM1NGBOkMcXggt1tTaqsQnYfCUtuYriC5CQw/26S9xdLhlCsq1cnAN4Z6QwFPtHJk
Zp8F1/T3CZTFVRNv34Jv/Twp/QHecSIaq6iA29hup0QELG4lRhKSB+ZYKm94Jn7xwG3N33G75T5M
iYZJjs54QiksIj+Jgh4e1j8ay3V8/J5rLPjfI7yLmulx3nz3sl07du4OrFpy8HEbKCOGm9A57ITT
8Yqcmw8t427im5PWmurryYWobSAYCxD62Fo8BJ/2+T8tM8p7PWW16pbV03PEmP3Jbe9nBXgcRzed
6YJHrdI8+MhAJvMGwUiwCIT6/gNG1Xts5nqc1acTKEpNfGhE7DrqKcLuNzkK6CjPZ/197BWzwY/G
I3YT1dh2F3/XCszUirsLmVGMlpI/+LlYbmZmcP1jv+J4FY79n5ARcujT7GvcbR49Za544TGvuAYw
fBwPod92Oo010rA5qtP22LwiJFJmQZrYMfiQxmZ3LMUTCrecDs2vJsON+fWf8+YCk95nOWvH/Vdd
R7B1gyNW9ora5dvq+eamOb5iS7AxEtO4TqlOfihpktUr64Yp1edJMSpy2lp8I7GxthJ5mkrF46vA
UYakz5bWK97ffJ1twKm4IYO5iAB0LDZ1OL6LmU5xNPdBXJ9307uHWZdZAKElCbJez4MnSOISerYu
VgKStpalw5OkxCrdDtNXUMXKZ+USBg70+2kxYQc99cru4/e8Wtn8L61TsEEsYgYdzHqs0J0ftStQ
gxH6EyWXPq3HDa3gQ1/qsPnxGCySu1I6zHTdhzl7/P7olM6+7AS36y2QyGmyTEcSlaoxuda0hcry
98qRC8mQdMNrWesmzV2ITPOGxxVOgFcwMQY8TaPs2p0UsQWXg9DW0eIOr0lbYZcK+sdpZUTpeBwe
MjmRJcBUkRy3p0nw9n8At1vZyVEcXd7h/zWbRAPOo3VGc4hl0vgv3bVLzSF7B6EAFaZRhk8P/hfg
Jn17V5fpa6WxspF37Ojcq7Nb6RcEbWY91VjLYaHdvkS6pFU7H39yeSxKpZ+wkPiVFNMbVQHC+cUi
ZunyMA6xO6DujCzXA3+usWFBqWHj9/qBV6qssgXb6JwKx9/LI22bAvdiQdnkJV6s1CEN/oBsAjUC
ez+NytNRdEJJLL4MjTwlmU/iPjFTRZxs9NNC58ImOkX8n59qO7yLPxK3Y0dfyun3Q4MFoh+mdRBF
EX6fCVGqf8Y8CV7K+5HL44csuUdJTJDmX/CZlQ1sIsfq6J6kgj6Xau38mnHw6eDZPYdlx5JT33Nr
hsRc/GlQ4l036boseUpHsznqTLsJVzzjJxhEdLKS9waC7YTY1zngHrefil2vwpUxQECWe3CUR9xF
qyLAGKPK6flmgXoEBaxG4b8MLCkkvAUKhNl/PCE8bKlnDLc635HujSiMQ6dXtt35ZV5knpi8iOec
Jku8oHV+JAY2JLC0FG57cAzSc5TFt+xkadR8uoLkw7mbhnLkobL0ULpBT+jlMHh+XaSpmGyWLh1j
EWjRUZntSYpe2cdtGZa+P0uIEHiGnhI60hBfWiOy6PbgUTWpqYJJGXFH1ZKmf/Npk51Aa9SRoz3r
WIXUA60xE8YYPilQdhL9GG+toYCtMhsEQBZW78RUgjaJRXYfTKWDn2YX2/nqH06IOUII00Nu7u+A
BXNX/GIVoG7accm/yksDR69xuuWT+S46FfKg9pST+Z7AmvYMd1y7j+Vpik82cF8KNpiwYBwvKv7O
91ppDZkFk4uGHjUOhYTqc1h86/2/amMIi2LojTqCXBAhF2+370+w0wBSpsQosFngeP2KNZAHqVeU
Z5S3zqYgoa0NEX6nd9OrvstjxgnNvqH8ftjCIrvAewL1joW+vzXwAyj8AylBuf1kqwRDUwWnOGrE
L56ypN24Gaf8ERxInBbg9bqsyufahJ+DACdtSni9BLzEp4rpF6gXxkItRUtEa2SFQkam7/TQiW/E
oNmrG08fbvI009D7oFVU7Xg1PmaJeB5u4WcTZaYPYiVN7MU7XEe5gytxEYnevMb8DzZ3pfKPOEpX
wsCdELwCSjHFrkc606gXKwsgclK/hsWaRUuZFTU+D2ODeiDg4uC9FyCC0w+q38055SgYoi6yOK0Y
CVkEJh/JpfkQ8zG7wIebrsJyq2scy4+mzxGnXTyc+KhGf+6W6j49WzeQz0toTcxoodNaIyTf4hLI
U69hd0RXVsL6aI4pfqJ4IAIzRAjGk4gItOZCKZbU1bX4lo/uMylWEJa26mcTOJlorBjtADWdHtjF
mWnGX1Dq9jCTkgUtMdPCSJkDeFtrSHQaqRCzaXwSlISQiarQUK1JKFk2btoSludjneyUauYPwFen
OAuosSjpgqvWdmj36XwFpaEny1qQcsu/c+0jdbYHUAdlMMbqbT0lzUOIxFLz94RS6m7519r6lQIG
+oyyvSBPdA1OrmSvqwBBEkAtr3tYeNU0NRCIcHA9SpdaoLo1eMuezA5IQzTDBEhYYgKDGJ3cHi4m
AF9hnJMOZ7LlzJ2+CCN5Md7xxML3oLSieulZybmYmMqZxi+b0C/bjm+bdgaJSXF3+ZwYWS6FxSJL
AyAooFZ6ScaE0GXasAyNVb8GXpTQGm1fj2fWoajaib3CoGEwz0bfJQZtxbRZph0OfFuWKES4dT24
ABser3/tQCEyCM8snwoOq2odTKV9PZlPSmRJ2qGgUmscL0yloZE5SNaAiXNtxCNBL0a+Rw18mX6f
0uj4ESyNa4iWNx+BVjHLzAfoCtL6oj7oEOwz5UcqxNL6VKF8v4en/LHYkpltoXvpn99k5nxikCXS
tvDAFNSw8SzJs6X5MK+gPfvM0FA3tTMMROHnq2+y38kI2JPicVJw5vx1CLDguJKab4MX9KU3ELoN
LLKQLzfEViHoFJPPZX+Yz2H0R0ke23S/2Y6PalaP8YswlD0GovhXyzj553HjsregTCA9Rhuy8Xcz
L6YeMXredORocz1pW8+NpLV8sVkWVVm4+o+ORScVJoynEsjooxAX4f9Bg8j/PUEJl/CYkobX96Lw
X0F42StEiMULriR4Qy7uraiw4N5nZ95L9WQ8EAjT+M4aXpXNrR/fgEjjHRjFygtPWECSwrk5GkEQ
Z7DUFO9NDMbVeRNLLtSU1OL+gyQU8JEc5Mp0YZ5G+9hLaL4d1TAEoczEvfD5bMYkzh3CdD++1pI5
Ul63FPKx6/i4Wb0djG8DEoYx9F7vN2vRV6F1DkwpSrRvS9ffpiaiIscKaqIAyOe944hbJN7paGSo
iaWYt6x4p0VCfgBKSTOB85uM6MD1uzWddlAF0xqeWDUXIdqcPrN7elKNcRs/MFO/KIJAmtvkh7tJ
qEnimBx/xUXi99+THDY6asInxLd54uIKClDmwR5msTeJLbg0Hbv4Ls0a9wjFMQjwO/qhYZblShT8
6/lYZh06NMVePCVY/mvSqCO6m0/mJSQvn6qregjsH1PYaLkWxAzBra5F0h5eq98q2Evo3auafj5K
izE54Q1/0RBbsIcna15ac6w0yZrd/O3jm5cg80zqoIlkZOSlE61TdMGXc+dq1LB5XD8ipmPJmn86
3BOAK9BGAGFat3fh72O6UZ3845W2v0g2CtRY1CR+Oa1SOHVcPrPNCI+wkecze9tewzc08wx2Uskt
XrKhyWWSpZ6h2NNU3EDahksXbVMQkQjTDIOs3FGZeJpHuU0aSwMTq7FHEGQ7z3Z5PtVVWdHYiAOt
TiV8RylCf/mo3onHLHOwa90kkayEa72l67SnyBwGyM80U5ckDl5fZWtb1V6DpWaq0SGruGm4+0Vw
oNhXt4An5hY2WISBKVNbWlLUuF5boJ2pBcZmNQcCwa3AOPeRzKBQVcusLQvxl+hNZ1mSE8bOEKLr
AErHLWLY7H022y/NpgyXU/xHAq3NuSVM51vRjm06KfanqmlIe9wr5bgUdjrTfgn2MWtsp+SS2OXC
uvNDZrEIDmEJvXd8N9GvVkC1ZsIleRk/ygkg8/r0CBshRW3WeFrTbRXRKYLxil0NPiiq/m5JB6+8
xqDja8LPrZnC8RgXUBQ7OrvFW0pmqBCAW87rL41tv2T5FgOhiP2/NloFUnkt6XT4piXfejJp3tY5
4n0dRZaqyWpy5/zUDqwB3TXkhfBLypqD177HRfDdWHl1SrmggkfUiBKe8/rNJPYsbS13nuFC7bRg
abU2qXuxi/JxSwijVTrI11DFSI4YugdOfw+SAcwtEOMfFZdmdDAEwSvJSXeRHusD93rYhsJ4DTFc
XYwHJu28B7JtEIjUoyOv6mgGCIprKHGSz3J6HomQOXpthtpQ+gOuKf3uwWu8W38y2W8SRFU04m3F
dUvtfVP8Awm1yFn6qJtAg1cHodLJbUnqxpz+oczPH+g3fTMoMKUx6RGPszTvTTdNqlY1MfgCpRH0
hYNlWDx8EWKfIrZOWMLA+1nZllbZjxz/CfqULuKxJkRKiWgBA59MaalJAf4gaIJg1yfhrCCrBrcg
+djRzaoX1VOPVwD954SQ1qdJyw3cAFEcS2ny/2WvbyFrsYTb2ilbUh0b40ZhYws8kcCx7qxzevNp
1WpoklTXvsZG8WDGAtsGEqOesxr+HmB8+wPaGFoIUT0bOiXFDhBlEHY9ooSpk2zYhWLPoyeSkyOb
SsXBcyQeSeLne1zeaW8shUfrWCsIvtXbJ7Y3gH/iucy+0npDHBXfDN5pcd8ei/ZnG910JuPo4caV
lEUYS6+sjYJQu8btZcQ7yHSR8LsF6Md7zprQYdYwaQsA1BdJyQIjIHRLc6h/6Xn2rQrS+690wfGI
h5/eH+CmWwk7oeAFo8xCdyax2z9eeBi8HteNhBMvCOGdIol1WrpmuiZjihaF3g5FGZqDYSmwyzTc
bviq4HBtLQ84xRSfLT4nog4jM0SHndIbbc07aZvJWwyOfIi0dO3oPmKYTbssKiP25yahFrmkchMn
ZoQWYwNSclOy782WpF3QSSkSlaXgpHX16fpuuPQii3VCB0figlfXOSwdtu4LxNB6CSSzBLDwhHmQ
K/qqBbpHpk1plT+VMyPJZvi6ayk4RpUU7y122OpePjAu1bP49dXE4CxDP6K1np/mxAdPtpToAy2b
uRGjiKt74XAcv6z0qDQJF2GbySSjtG/sIymxyyB/Qdepf+ZE1Vtyj2Z/MC8HdVzKScBWiH/fi3QS
33o/0PQkvezn4fnJ32YvAzIFVTEF5uwWlwiHixrkObNx7/Nx514D+zv7QPlvQFhdQh+HJlM7DCi1
ARKyhJ0j8F6lGzGtLwDVUSSW/uXSIKEJHRn3/gxdTbo/Ca32n1MOLjizFbGjoXaHKjoJ7VOgwyDD
azx+12kPxAB8/W7IkBYEjCkdhtu4ghA9Fo8GnaZ9Qwl/+VRaq9sUsse4vCVURoNGsUr4oxfGyUXe
eywC38up0DtxJoC4aiaq3BC9DCe4FSSUaeH5h99/Ywra+fcaLT+dgN5PQwrVrim6R0+Z3FbCCbM+
RVJqBFVGrwntciwyY/bUOHo1Ya2S4hP0woG8sXHymzWx++SxMvl2YEZUAJHF79J0tM3NRHs/Nm/X
SVXJ/uPBPg3nQUGLZ/e1BFWhGhrZkmGKlRJkoH4b9JjkAT9k/IJdJcAzRjjpOtZ7I6d0VG3MyWnX
Zzo/wT0YRQyHi3KLbNC5dXUndISRQQA80UyHT75dEoPfqe7DfIsVhJODW+ZaqWUbULEWNb8Af0DV
nw3npJE1kCQJkaI07wvtTYL6IUaq+u9DqcWPhaS2f07aizfpaVgoPJKm+keB2uWHqvh5PLVVJi+3
dKkwRFEaEOROp3g5+L2tvBxPDTI/L2geUHDhW+UJHkQyFZmIw7zGxj8u0VoWqgFq52oCST+adMI9
U3jumb2RBRLVi5JN+davrX6VVy2W1CMedTT6l7VscX/w3qdY7zergo6YcTAIhc6pus/AaQehpmXN
j+rJ0uDd6hgSqtXm/fLG4CEtug1e9CKxADlCkLiX4t692fNOx0ee9lArFXi0RCp8oiwBRWEC7cUd
UxtIdhuOt9KAUfdgsM+gHzfwLU0PgQ1zEw7X4Jlk+UxowYbwAOeC9V78YHbMNIkiqCwafCkX7/1f
7/3TNBXy5jTZwYiJf243GQ1niZdYsHh1Fuo39dzNjCfrqsJTv5ReiEhn+zmPexT4N2brFSeTjzWV
llnMWqYXN445B+7DdZ96uh85iprmOcZv4txizNItP5cC/emQSZLVL6PLV63qKPmJMa+zI7qlVizd
F0zfpQW+pJ6bXTt99IbAhNvvbEPaUI7ELASSQemDbjwG5aaqjEMBfzip0N7ZZ26KPWurriRn4TSf
IsYuZlK0Jz6UNK0MeVX45a8hMjEqqYoIE8De8u6Stp3xKihClm4++RGKcpiJyXomprIgHNXLVmAr
/oHHqcipiFgGXC7kzkpyRM8lD6162KHL/90sOZvh2Ahv+zA5I/aP1B/BXecs8lqLWil3tKs+4EPp
R/SchNqB+dxYXQ8SJtBHjpYWr18zu4io5mHFW+XBdoWRQJaFU5z966k6AMd6MtdnGmQxJqsMOrMk
rSSLsnHM1CN7Xs5fA5pJRw2hhXcP117dC0IPNYWj1D/RSzoyL/B1fDgRr1nuGBrAxHYZiED31VTP
EICmgDrgprMLoWVWnQZV3OEFnwEKJIRIJs2yzfKn1EXty4Y9k90kAKUNOUlSQDB5zz5fpPykmXgs
kf3JN0LlDynk1GmTN7OvahscJPt8ct4xw240wSoA7Lbi87c1hfv12uKW5g/IgxKVlUyZLJJrK23w
4w/3HaXH5NMVyZnlU+8c84QGcBIJh/OcbmtqhDHPxajwuE7kPyrp4X0dtuPZGV4AEQtPk4gUiqeh
D+yoJ+g7oJBhcTQRDY9Kw9FYg+v2ioxfZk8skV/j0c1sERDbjN7KCSninLNoKFKkR8cmlOd6Uix+
Up+xnRp2sWPGuANBURKDn0OJVKp5tn9HiJidKw96dk267VjWibnNklDtOmSYx37wxatidmPkv6S1
FRrXVx+J8fC6LNhfHdoYsvGT1nisWCxwLCuDtOdMMonfoKOosoNoGjcW9YgEL59CF3jtmer9w09x
I5TDD04xp0MHeGFjkel2wm3XlIZDn7n0fCRm/jfD8T3D7dEDCSoiMgg5tYqI5raXlelM2Jw8fZVf
m6QJtFq9DRPdySveFtwS9rcOxqTPiq6QxL0HQQjXy04At+dJGwmJuEZr+lGnNa/eBENPVWU/uHRj
oLbbsSg0c+zLPF2gfOGpf2a9cZFTxqMOxuPz4FU3GQigDgFebpyNRR+MzWABVXisUVxMCpZtIVG/
SJcZm5qsjEvXXRMlNGmb1sjW+v6o4p1eVeC/HJh3Iv4cafJYWLetEiNgwVDMoKchrTI8kdub+rIP
QKlnHAyyC1tI5NTc3T6zGteDYhm629/AY2X0dwiDXA46jjr+WZN65l6ZdyO0D/TDzb9Psyzu/Tup
C+VFU5Ze8/xtmB+oqFF4RRT6AX7RkbzjstH8kPfPtPziPYvqiorNPScd9oDXfCcP2MImWOTObaa0
uWy6YdYEpaUdunmFyAivEKipGylkDsPZrMjyTqLmHSGPkqzGlgQy+YJ20kFDarTCLs2YkZ6pR+ZH
qYHhqbamVx/7S8hX/Cti7YoJ0n/gS92j42rC8LrccGoW6GxISNghG2NX08bEGsYJgcvjgLb8cG7i
lNrHmX73tPpPnQw7M7hehT/CZn4Rjkf+sJbY+PZ1C+oehtXfdsp4FbGq1unoDkeqw6HWCAqox1HP
hAb7BCT2kKHLTy11SSD5y1EDyp6KxKlI0ZEGLjx6p69hVX5Yt3DK5ODbPRE2YIO2lOuRoX2/5lae
2pGZGKE3WEPBTy0kuh7beS2ILbZunMCoKpzrCWeG8/uxmXcp0P+TsYiI0ldS7Uyi7ivgGmHJYvfH
rieIxbu8Trh5/farjzVN/0qWEWGWj5NNNws4nTaNhzuAc4Ppet0wTNjdvFvUlnYuiVdVQ5qhJGav
V4PUDpLpF/Vo3T02zBvPkXWlP6z4dhDcSatK1+H0RgBMHbFuzm3W6VArC7Uhy782N2DKNBccKmJX
bHSFktKH63KgnhFDOxbjKGERwZXIPn4wBXKKkzuLQ/+/m6dvUrTbtE9oNCmM28ClBNgG0dt1FfXh
LmunZcdSnc+YtvNEKsztOKgB5Ki+eojqP7BN/7rBNWUmDy9cWW3PqDquOjIMmOjiAOShuL4IEmh3
miPkJR+xEpJqtgGIFuWjVBWT+TMPBHk4hCK0OFCX9p/2siCp226bxEx4OkaRfRQvjt/vMstfYuat
9ojVwTiuMMUKJymnKs9Ogz82bJcW1gWFKejFt9lOTsLftq+mmfnBN7jyjdzW9hJZvqB9b6tBYodE
l4cjLPUABy2ouILvMhlkOnyqamdpqA1iY/F3uEzeiPqxeBltfFYJv0gUt0EnnWPbTiT1R+MaAaeG
oUsQyjZ4h7c4I1pPXpJXpye4X77AGrI5H6brRC3hxTq5u5AYxC8b1nsJaDzByC/ghmjPXXTIaTuO
JeG2nNDIjKYGFYhSY/SPyv8ahvk+8skSynFuBo3HnDTHuoCx1QAaofJkGchRx+YHfWY06OlO/cLZ
4XFYkI1qirUB5AZc89ldjtqccRkUx2uJDnXvyldloYFwkzkxQmXnI5QMPzKYELH0yfU6iyszP9ur
B0epUO/ypoe7pGPkmoIkXevIUWGETSYeXgwmYZt6sm1WDrx0SrogzpES6sOUOotv/JYFDl9bBB+i
UYFAyRK/FrH9t4eWcQo/xbPayvW89XWnqjHP9qxsHwfulPNSJKBCP8QeyxMH5jAQMcQzkXTwSPvp
BeveVCyGfViEpD671pmEVC/CgaCRgiCD2ygPRQRw+19GrKvEEpDrYF8EuZRaJKVF17amnsPGhko8
1HNk8WW47/ikkeJse82XQEYEH0Y66a6GkcE9b1Ji3rF732J+cAoTT5W+e2R9/UJgPje2iP8he3IM
m6sA32d8bkDRhbvCAlc6zmZe7D0jvUgoucQELQXHfuOyd7ZPqDIc7lgyzDFoLSbnifQ7XY8XD/01
Ss7oVTHcMiZ4KmJvN+LHB11VljPahsyhKHmjFS9apXxSpuYfVNg39MHlMetD0nReS8ewA1mNvOwO
1KfYbIDs8b4qW9JUM4GwHQPYuINshttmNnBEbrHOk8/k7HLaUULZrc5GYop6mIVQ37JNthkhn1O9
P6UfpqaaWqufU1hV3PBkXFU+HtTaDly9kX+rd6IxSazzT/NIt1fpJRpSJ3QadBlzu/4RkD35U6Vs
ZXAPR3t46woqWYvIACHC8PUM9EJysFKhMSL7R1h9S9XBrAk2D9sq5k/9huUCPnqu4TawPpsG5O9l
Tj8EQ//mFXWe+IzYGSO7tzLaPz1y0FuUsGY9TzjFCx8DuuHfOjTY/KXs9XAPzI/G8/5oMqPFeIde
RIogC+LP3duAh76RrKMJszMQvcTBqm1ERnLBhbxd8EXZXf/3rmzHvlPhBxL9OzOiQgD8Ku+PSikF
vSKFRUy+0nv0SjK2riBUsXamQiytDIg5ScJ6Y0xEJ1VJnlOusVdjvXFXXTBAh5Magjg/pnOxUIrG
0cPIthAJtUU67o9YJfkZk8uyFPn84UGFcQbF50MembgAtmuWzyujejRHwkvHW9uoBn52KELGiJYy
7nS2+DqsgCB8SrScP1WdOFiiNiEEeDXeR0qouuFlmmbwnrhr6rC1/zaqNZO7aj65cH9VlzrirXGT
AfFgvtMcwazh6ZBn7aKRWXavJJQneHUAU8B6vJ20za/Zm3yCIyZJLIJQCd44aKJ4g0ZJsAvLjv9m
NfWB3e6eeG2YQ9bzoU5MiRUG6DfJNksukmfm/QfgwiV/ZZKrWb3l0n93IyndjRMfAdD9rz3kZ34d
5RePT6wyOb5zpZnqkdKNSALZnESTHpunwWhijgATaNYqrszyr3BqONK7vJOKlhJo+rGr4Ftpk0YR
0vkoCkbimFrFYWLl7I1rUfmD8Ksngvi0NTgL/Bp0w7vATxhmPMcG109lZdOIGCv/vn5AjbFGGiQk
Ocx9glyPvZEuhufF6igsZ5eLI3Z92CMF2G3mYmkFlT/3fhU2x1U19goxyhjqc5gKSWLLsBHYKtkl
iBahYMmvGIsELmLIGolXeziXCsZJXXiVGyWgrud1VEhMcNaSlPvl7qbYp2QBwjjSwvgMFEMUOxFb
CAQkm30cWjUEfi5ByV39tITg2Syase6vW6gEYGuMkRwwWI7wJ+1krubBf5etdnEJurWmCEd/Mmhc
/3CJM6ZX0cVTllbzvkZ8PR7pJViWruYujMsJ7hTGzKI7wuqj3zW4aKAG7odLJXYRBoTOe70D4Sut
vM+MYvFCpMXECeeecYcSnarabhBU6MrKgSnOCZqNN9L91nAMDhPDHyNSY+qqjRWr8HNRBPTxcc6u
F1+e/RImyFxoUH8QMJRQX1L3eOQ7YW3++VDR3DxEpCMCHAEdFNit1mMFdUNXExHZIKKHZK2nTi+S
pFFUwlRDc2h0KLXoct/Z7SMeaQ25dhQz7B6MiU2N1Ns/lF95JDzp8y0+5Lsl69CwN6/Myho7oG1u
lONJoFysaUg/yGBvIUtbBmR05AU2Gs6qBwDdbZ3IiS22wQszC1BkBacAaaBgQA8BbjA32b5sEAQ7
mUefDlzhYE2n6qy17J2/0K+iSQHAr9hapPt2ABx693Tx4I0lpZj1eLnS2WnSOHulnWa7m6YCfFp8
UWRzJEJU1ynBk5uLQRf6vleVq9uAKGpMDtgXUMmXmo4mEap49Ipw/x1FSXwYpB8CWNKOQEG8Anoi
+aQPi39QoFgolQu/eSb65mMqfH7yHK35BsiGY8ME0ta0PPkv/ikr1cqj73nSd+q79f00/6BJrT8x
gYCos7w3EAcHxFbuwCbxIu/uuyB98WlseyrR1OCsLjcKPfl0d8tLpU15w8i7d/AjuEBWRQ8BPfG/
Hddga7UbnAPpBkwuXakADiTebBYAb7+BJ9MuTOfn8rVqWtFXcWXhO7klmETW8nQH55yi3IqYdAoV
OlEaamwsfurz6KfXG6i98hpoj6AeeTMyUmz3U+irmcPZArKA/JL3JkLO+Oru7M5mnb3XJQlu//uk
u/X+p4p84LE3SKABTICqv89kqgk5qEY74rYCxdKTaGOyJm1YXG97YcOZlOdZyREMlpcs7GKPUJXr
KmAhn8D/9ZM/mjusIK/xQy7dbXSutRecfzW/qMK/b0oIbtswwWx6IrLYf3PvR1FWhExKaKtgc4kW
qFVcntZdAEkQ/q/5+aLVJH6uLTO3MmUJh2hewq57ky+1QLvU8k2T7L7SkMZDqv7Y1XbMXWBRVXOO
RllgsPkpvFDlXEH4BTpImNzV4N5e5memAPzwSgHK5Qs93UiJr0FCRHIsvFqSmcCFNJLA4j+fZ002
Q9Y8q9UE7UNyPnGAS5m2ZuoQmGOKzf8es6cA4bA8kh53jdpdQOmxstdxAJrriyfx3T5oadmJJ9Ut
PekCHk2UB8izKnmhuvb916RR/oYjQQRRFHHJmegv0cRzzEGx/3ORQSWooMa5+MLs207QGDjjlfaA
rqHmVW9iDkRFXiPNIH5dBYW9NJp4e4ZGcrfXk+PkEleXd23rePk0rPEGB9Busdc/mGnNxRBXLH5G
P6cG4TXQIkMhgCqW8CNp3wrPkCHnIw8oNcxOXSsWAuA+ma8Wlu0A0Tui1ntQrxi7gzRdTeonPCZb
SR6jdK3HtgOXBJ21ENhfOSFls9ywHgX/gU8ZWyMFF5dtxFgIsB+9gKoRfFDt1TaHzYDJevR8PbL+
aRmTGAC0MUYSm6qcZ00CtBNw2nsjfjoGHTvqjSY0e5rrk2cUPq2obxplbJMvzTkF79oUCdfJHIZ6
JVM3rrRpJMRx/dREs5qE2iKX6URYINEUdGagy05w1mE0pFwOQQ6aU6QelawN6/toa0v15qiZN9tp
IZSNM0cWXWCbxc8x2QU+UKj4JcGHCmOGMu5j+VntxqluZGrjhMYqjSJEhk50jbuGys5o3slC22yE
OQ5w+uSW1SlXtaeFXhdasUhEHu6PAQyZV7DftELzBywHKMjfiPu5+Cwzu/LIpgYlF/LB+2D1gnDB
VoUnaxTVs+o3pcHueyUuwEobG6XvZZEMtzlco9tXED1jAfY5f+Jk9DtUhJIFpfF2zC4+CYRMnel0
7pqgLcY/a1EckXkec4e2pXmHaDfY8NJ8Rx05uq94BN9256OlDIZ0sPb+sDwyGyUWXeCswxYeguYK
nEhdFyZKkyKxMhiJxE+GlHzLkOY16CjpoLXA6P0QOnJMBF0NQO5MzVP0l67OfVhFBz+QLOtDQJ47
J5J0z1GFMfT7ZX/LBIEYxbwV1dm6qubN5DjUH60Ln8RAJfZa7jhQzuabS12H0iWR9EWWi7aIjhwH
+bXCBgHQDShz1EtMn4/TLmAfPyYQpQ3cRgL8fQ+LatHShZ4DECE8gDcS864q0OFuXNIzG9D98P6n
hzWpkhIziZTr820PmXQVGI0+2A43tU0aQblm4RR9hLj2bqTyxIyZ/gmhUb7+WD2HbcGtJQoWGM/I
dB7fh/1lS2AK2GrHA0irx/XbAFzvxQG+LOCVaE7XlzexAe2eMHAvWcbjhBK17KcM9P6SDP3kN7kl
qYe9FbiZKxJ2gRTCkEye91Y+0UN70n7tpgFsyWlforW+rya7Pamg2JDcefxgTshnyPhukufBpZpd
4ZFIQtwBL5jN7C0IiqNHXAtecTURTy4RCypGPMMqQ4wUh14jgjHtLZThkdtth8XR0RQlcbalPzbn
/P1xLryl/EZtyNsm6zo77lpzIun1MBw843oCin5tcMI0Uk+UBPr+ydqKysMb+vUHNYhDE57HVwW9
iOGu+LzQe1qttUvpZFLlIooAStGbUhTGHh1pLNQQv5m53YJLQMVp0YTFfPvBP2/vMMY0ABXBV49V
CMrs+gXqtqZrSl+9bdn6BD+J2LbOJD88Fu24X5RrSGGxdLzMjjiTiAyYrMhWM7xoDK5B0y+WrHvw
Nu3DaNaq3EK12Frfwe3gG5ogHosDcqxBmvOe25aIGgM8B7ossIjcNE/SQVmed7OT2Y0waLsg7Q1L
042SRUUyeOM/sEsuL0l2ypgUSxmaelm+jXM4HD4p5lJKaTzjutdIIGLDDXikS6cVWd7odFMLZo6v
wZq0DJyhMf6MNG0jnjNwyzFPd3A6H+CJROeXQHiCwbMc3TW0uJmJTpUs7cQY5ZKygPc+V4MNs0m4
6Om/lsk2zf1yi1IB5OYcQPX1gvLTPUIqU1C7POV/R629YUVN5LAgQX5DHdc9XmQPlqOxhjW4OcBX
C9ToRNVeBppgN9FbmjKlBgTLHJCNNsA/rX+Cp7XQYVNERPqHIdqq0SDYm/Z2nSJijJ4vopFY391T
VNMD803IrNelGp4iKnpfv1Xd8/JYAzCxh5V575waUnK/jWcO4EbLraHuSSQzr8fvnLcusbc4N9PA
HE6v5EjsU6yjOqZuYn+QH2xO/l2px/za+9jZ5JfVyNofVLD8Lk6Dk5l73mBZYdC9PXt5+AEhQxVb
5TrsKUs0BrtV5VWd3QbhXmzx8NUE0F66bPsXj+18AtpSGgL/uQahRp5ru6KhN1bynx6DNejHuh+u
2Z2CfjKEcuD6llNiGKAXYlDpZ70+019EslS3vaSMjUHnVZdM8L0wSOKs0YZG6Mw9e2xPjVYu/xHv
AiCdAVTzHMXSgP1OcJP1cu64euNiQWy15C+PVTtWzv5i4sIRq4OL3GEzR53aNq1ongH07mKE1VSp
Br/3ccXh4YVLhYNKIWxz+9ww1ydJadKtr/ozfyMkyWVWz+AS1MMECSWLSHrDmjQqTYxj7GLBlfJ+
TtMr77CY/Udt7F5BfIAS9D3jP79QNXAHXejk+Z0vYgj0fyemvhE3enRCqP6CDhgZb2kaQrX4X9/c
XajDUjJLZFc49JOxqQQgqA8djObh8ZYDXGrJ+GfeRA+aM1XjQ16A/my5tqorCLIiVoZDTUgjeEof
IGWeu20+mZUE9wtUmbNqJA8NO9lm9K1e3x9Pelj9y2Rw4AfC5Cj0dIkdag6uNn0cCCKKlWqgIBW/
CzgUIEYwFqavJtAa0aUmUVqWzlgCX7F/cAqw/dgHCRA0baqV5BWfjkBDoR6ZyCepyeoVLVaoATOG
zGbEYAtjKosygkSCexyryOuyavlhuk+SSv1BlaGHiByl6ULkdnbV9NnE3UKgadFfKKcGdb+oVviV
a+8EuhDS7qLAEoTZdzByHMmtV+kMeAFbS/8rT1wzK0bQbRt0r25QPl4SHjyPLoUUGiVUBBj1qEnl
FOp0cm6FG08I5+cx7+OnCNqnqjG+vxlAL96Ys/pWQ8mD4pTgM+WRfbhPEB2kOcEgRdgs3LsBlKzZ
P03bZXAFPVZFgPZbmLvGkt1zJ+PInp+rcFOVeYcGeAdlaSOEjqKe2x1RsD7aQPVKYw2/9Pp0dHV4
UjtY66nmy7FEFdQc3THR9Qipb4dfO1IeG+JsfxWM0/98kRMdg5VncNfMApwiC7CSGnbkkhx1fTh5
HoKJYbTORE076rBEgCG+yUbHKme0hO3j8mSW7ZGH/cbo64x1MurnPUztMvHymYl8xfXQWn08k7/R
g49NFR74F4c7j5GXI/CSwYEyLJIkdzUetULaeptP5M+FgTzSgPYGVaT6tf/GRbgEP55+Gd1h0lC4
OqzWffMYJS4ZenhBgsTzIZh4ZIi0ucgOEjLrNVcmWYCcHstcHXAX86e9QmNLLcjQjYmuOqTmSjuM
JUHwjguMAJ9qm6iCGaVZ810qSjlHvWpOletDpSvuOCa7A6BIY6krRDg/q5nvVPDOkmYJfPqalYh/
wxKFolx/1jZkZZdXWW/1uFmjpZ5/d8qYhdig/X8ApDRJhLYSmpxZovSrhZnHAHvXJfJFUVltxR52
9I4jkVUWbCm9ILSqTv7+/7+KkKoe/v5C3WrBzn5GINk31/X3KCAoy5yJhTP8SpIiKVVuW9q9xNDu
Y0Wq/WpAUeIVbxp/FUDL1dCPfTEO6uOnCbIPqDhV/D8wJtsYI/cbn4YZmyZdjZWlARZ8TCmeYK/3
ktmxn+zSho2OcUwAnpPvdnTP/zMhiiqfbmsVX4eRGXJqCV2/iEYnI+nnTf+i3KlEDrb5vKD1Ra6+
9R36xfJS1TWqeUdOClDqyZQX9zg0R83XRTjTzru3T9KQ/3+CyTFbgOMPkhEx9Y8v8dajB+cLCw1+
1cFk2OAXE88Q8AmrpHfxSmhV2DGPUqOfWHkvrMtsX7tF51jkyv6XLyLGjSZ8n0D0IssFRbSAUqIl
EREs9M3ou38DqyJ6TiJk4nFZZe7ZXEmHWjQgZk2AKEKOvrBrlxgZ71IJNNrwCSKYxiGhPBMTHi6Y
V1MdH37Y/mQhzlqlqh0+SWEC71WYneDnHea8Wyd1QYdrXcK6oZi24hQ/Aqsfh8TRf1ww6y/QTABH
w1NJZZXvF6WmDvBwGJ/EnX9El+NTvuK4wephSFEt/k7vSsSw2gO2pLjbLe6hCkw11KgnBXwHrRDx
GeT86jrNHwtNYkoMX01bfnbuaYxLIJEdKjZruIVD8WmwhBgydVBrIZOQfNbIcWcMF+F6+4znXDda
v1MssMNCeQ5iuSJBWnWhM/wsfNjGjcXC7++/iNKnh72GF6rPN0IOq7W/WBbmevQQF8m/hRHi3tDo
uZx8yEZwIh42bMoSKGdeeslEMwEIbnQGPSwzAh5eZzbu0JxMxt2PrPuhVNWy0aRjhmVwHAuJKv3D
1g/SJQcAmpJx/EWefDLbgAjnxekLjueHY4kE4PjYRxAw4BtRQ/hnVndAddInFMrdaVWMkZ5TrEIp
sbBYbF298y6/IReaIpHIQ5UGinU5wo8glKVyKnHL21+KSHQC8QSAhC0OJ2KfPwI34Vlufyb6JxX8
PhX8EQ/lcPz92486yxQdK5vyhSXgvj4A4yv/zKKcEA96Wc61ezqjK2/hTUbJRZsHKTCW9os6HLrk
vsN4QweLiORdATgU45/93Fn+MBmWMsIkGV6ywnUxphE2acTrFnbBfi4Fn7nkFaedZi14YWB8M13V
ph9/QiJatrZ4v7lMXpMXgql5Y7u4u2dX3EnnJDgHas4IrL8bKG4NNh5p1q3uDn9RzlgIkrR7Ygr2
q4wk1rb3Hvimsk+XFLxE+bUTAn3Kin5SUWKO+WvayL9ZO+4Buz+99oV2RaQXoQOc3AW2OIHRzQ0i
jTasabCY7+n15h/6hiJX3CV+eNqW3wvafBWfgecz3y9qFw0+BVZ+U0v1727msB8YWsu12KinYdFR
VO7rLX79ceTuqmf14slAnEDPyztDZB/LqKXQmAyGILWK32lLukJ+psItM6l+Ws0jNtW2khcHtPpN
fJS9x+/pQrUDSMy+8IE0KSx42CLg5Huezhg+8uEq6Uym8k/VbrUcX3fNpShrSE5Kn7/kThN1beFA
ILU+8FnBY8i74D1pAIgt8BkbNVFIfj0eoYJYzRaGlhYRefd1J1ieschoMBW2B2hPgmJmFj/SPl6+
g6YuxlQFeS72RlxWze1MBVW47KKKoFtepbTvVtkkwM2qGKtj/TvitytGRx8HZSYOHVVsYOUyOq+B
3fO2F9QY23N8In2bImmYVuDjuvswpPNWadEBd28iFMB6m57tgV3OU0XW7Ua0uq/gDSXeT8G8ziMh
mC96TGdxdtHXkJWHw0vyRgBanPG+HNLg1p43xHsJ5epz8AMCOmlhJepaIsP95W6Zl4PArf2SmnXF
Rg4xs/VlTEnZy4cXrW4itr+9MfOewrcmTR7lXO3tGS2v0J6StZCsclIfzo2s/7rEyyoEo3x1mcB8
9R68GBUigHIhHDYQwxuDCjPlrke7y6sMwPD0PGK0VHKU20TnwqqfH5GDjcJFmR1hgUq4cg0DcKPZ
Cu9l+fryNnt2//QaM2YULcQfAmD6Jhc/LpYpU1MSY+jlRjVs6z+yVCF2tBoSo32+NRUGYiB6QrQj
ls0VTFbCqx1d4YVEWr9x6rOajbaSpCM/Fp/i2JVC1PsMhkXlomamVXUa3EerdAv4KHdds2ceCzoO
zfHzMvkm5ckxxN4aOR2tvK0TtCHXjVArUnWTNcgQ+S1RdISNFVbSvO71jsQCyzLx8FtYIuVa0DhD
FB9poH9b8tgcVgBgderjkUQfiDZmkXHhw8x6exRKRwhKz/LHi4z07CbbdtlbIxRHvAQ2UhORvUvx
mHEAToZcC7rFrQ4hVCQkBSwPnipZaTHWDN6Ld0n6tMDgiZSpDsn62i3dbJdc4+ODne4+caAKg8Bc
7bmE/Ssq4s04T16uLO9x4f2CvUoU60LOsQvnU/RBKTaYp+xjCpjxa/4vBFTxBvghqXRpQKQbMQP+
MPrwQBApekizDmTXFTY+8nggvMjolqNzHfhnNFQuxzRJsuYE7egPY2Gl6bcMnN/hKhdwcvlSN1WX
gOK2fAFDVvuHNtY2MrMT73RtBAcn2gE0ftc10eEfgw5bk9QUA2y+PHModnkYvnghyXmf+Xe4B9OZ
dRG2bNAmgOUl22Go7WlKvH1Cptlyhak9NJI6aZZviBk2zoPbef+dl0vaxAi26+AUzNdI0c871lVn
xRtvYCpacQ/c14byoQYcReB1Q8R8tDjmn0KBDVLPUVlpS4DeyWb3qOrJorisN9XPwtEC88FqS8Y4
owuGrkZxN9ATiG4e4P0FpgnGQt+X/FH3XQMN03Knb3hK3dkQS68XdsPmgEJNreG0h29FZgIHj4J5
3GZ6eO2zNULg9MXEynxOsaRGzD7aUpMju2Npxnjq/4H7iw/urwCjjZHnKAzxG2tMnAhlwdAZCiRO
IFUt2RH/UZov+/b1LvsedYuVabyNRR072ZlWXh5yT/htJfgUIcs9BKvcD6apMFqAT3vW1Je2xB3F
KDJtaPO5xKuopomknBDKXGUBOPVet7ahxqjt4PiERzzJJb96xPtop6JH8UxhisUNsk/XmbehBZdi
FrpzeJrOrMTycR6tgQyXVLyJHPE/vr7JmNIsiNqMOU1+raJn1H1pT35hjiSVCbp5ZTJRcNGZHfHK
Ra2zo5fLV0goEDxREnBELLp+5IcZDUSqZcEyGaBnMZEQH0uS6dHxKjEALU6Km53tU+RnEWjWPvHQ
4PZ4iI/z7hMzk+PYwmSIIiswIwLdAEkaJSWrDwMyzfO69v6zZnpNdxJ5YM9+06RcqQW1uu2xuKTX
Y+EXiFfRfixp/RgbXNOPC+RjQSPRk+bz+DQQHsjXJibTVIt7Np1G9M1AB0uB+6Z2bxuncXVcaQi4
Fflqf+o+9oK0zJ6M6yhAPMH72ILLk80ZaE58bxIqGwlyWZh0Ltr9BgwpsqFbGglglkRscZiHD4c6
GuK+ZtML3V0GoL5Ib0DLBmbZI18GroHXC2mYzLGl8+B0wugKwqTUJsFP4b1hZjoaN9owvBn+eKBj
VBzbTLRqJ8MLXRgYBi1RNEW4cW7eZ8aS+TuEKOH4TvOGEEch0jvyhOsBLU20hLpmD/wkBSr9k4cX
WTwgojKaVyn6JkLEF5MPLYbunI0AbZ9sbE3YgGEAhUcrkBNvR3zPhSbSPqa+Ryjv4p/WcC7ZaqgJ
86xg5tqEH9oZr7g/TbKxX5neFKY7okEY1pGhsqGaeVfrjQEl1ZwWwuQEqHbEJbH/BV3fpJYVyJl8
TrfhDpQu5d7x2MBrHIZ71wkUjHX/EVF206LpcFlRzbEBgMy24Yv0cSiw9GP7mtZzbZyELU0X5EdQ
bvqrsmDYcYTUtFKL/LwjwnM77uiYyMT2RLxEM9a9adSV5vOuZK5oeacLwpXt4TIAFF0UhtE+gVyT
qic15AFYIb0AQAOwUFJ9lXKSYI26l/QUaTgbN2/SQvkYP+8ImtKrDlqpRQiI5mz8Jh6FfmzSBziZ
67Q0RrDKG4X0zif4lZ9KHVLbmX4xNpBGqu0nS5K/+OydZutHwXcjbEjHXYD9ZqdhWEAQAhlNuoOD
EThQ39rZcfM9rXc7PqhhBVpzqE9051XwVFycWSW1VAfKWANW3Je9xZfehWQOZr4gRLSw4A660D33
sFarE2U5aEysyKgPLzPXcxCDGEOXm80IpZuP7tcY5sF23J6c0wmCa7DznKdBB9lqE6BO2gsxyfE6
CfKDB9FCy64ZFwtCHuqgPX24/nAKtDnimZ8k5fdbisu9V14tViKp29IVPX9xXN3y1Zv4jj3fw2Pn
lXhafB2UNtJ7nVhQzJSBc7GdEmM6TvPWGJiyWpLSpNHrMURkD+VZyzJpLDngN2JxRwkkUGYhOH7r
ZBgnHhGDEiDaJ3RmRYrKDiVXLEKL9v/P76uuNuO6FXcnHpyABs8YoFLrB3mWKXThABxU+iFz+Df8
e0Cw25c84TurLJ/oJmMXKLN8BdiRC9qJVxK4CpGW8BFbPVtaHLLd55iLDko5zZWq4oFg96K4uPDf
Z932YC8eTeH4Bs8HgEDN3BDpN3/8v51WnzqgcHCJ2QYxisXc+Y32Gm6Xe0n0T3DhJ10bugVIj4J/
6B4eBsEeoHqFGG8b48n/O62TevCpLq2AjUj3JrWqTzajUUFY5aFURAF6OROt0h8Llb4+F7+pDc4M
fw5v2iHx8WBA/9rOOAsOfLz2SwKV3PA4gD6yn9WDQtDyPdMwuOo4285pOCzYvwFUA5jsnWXNVcWz
HbEBdWkawkheIgKNOs16wZEGDt5ikadeuA1rrPO8jo6/ercPk2OtpP6J6/UrGKtG/mfK7vA4L23z
SmRGssiH+q6sF15tACpFMx5ttyy6SGxvAeULg8M8vCRD1Qy8vpIWfnU+zhChV9yZiiAca7v8Apci
j7eqSkz0pXoZ/ZHYKoGHiz5aMm1txJhKx8arA4vyOg8HnIrAtXGqBDQWI8FgEiLWYGYzHQoXis67
9fIPbjRF8+b690JYZUnUJXvzDtIjfDuZxx4LZgnQIo8Juc3D1JuPzEGbdSxS19Kfvf0dcWLw+0EV
zZDdVd/GIxr/2lCxfhOwqs/UMbOqX7YQQ+RPJ3RcPIageZVtNFbnt614+MJxcpGBe40qzbB281Df
qsYu8XhNoOlZIpMma3wuaSyF4YDXbWc1DLcQ3Q1+PXy1RpnVFJ6VQQ1NlsLtrJxEcV7/1LRFld6P
twaZ8RfQmk6B5yRaDNDbjDsMSXtWGoxNNxsCfOFPXyLbUb7k1rPbo4OnmgXFgkFZiwL7AQLaB8pz
PzGVqxjN9e4fMFP4jt0syYPEvFRNVLRi7rNr0BgSx1mDszjbRQNNFrZwhzYGe6j5F2gqdRCwHRyK
bK8HDUJk1n/YYcB7jcUYAElHi9Wzk8Wnr+iUqz6bpamxGZ7m81HojCYSS5TQfFDzdcCopJ+4sLTX
NQZvUqaAbwU6GHfrqpKJoWuRZbbhwoW80niyjkFY1MQvMAVPbJrjHf3wUf1jukpR6cpbg0s/Cf+9
2F7ZAPkF+5tNU86/kf23GboIHkL9fDUP/XJoKSLNM3jH0zPkVls4sfZq5QF2mz3gjCLlqhbeFiCJ
8bPqwTwmlzzxfxxEccy7n3cTNYzSwZG2XuJ5btrkZkhPO2YhfWtFEjJekBvXTJ421qkqPY4ywr4V
lEPvghXniJNvz+FXy5kVIpBXP0sLHd+q4oNRzg7fHvSPYkFdr7ABtmshkfsL6QmIZ4H84kOTKv/0
mq2wOf0eqwrECegb02msIfXiodtQpevLtjnHyZZJVxFXUec4Z1cLrYWTuLUma8qHfUDK0vpcfvt+
TteiIW2e1c1wa7PsMqDU20Y+icXWh9yQ8ielirSNVRbsLa0joo8LTyW0uK85vBEejOg3ah6iy+IN
WztgCD+vuS+4C8cQOwI4r4fhtNGluR+IK2oVfR7I9oyQq3JBAO9IV9jUMiBkYGu+QrFCa352Cbzw
4kgoqXSj9LQas2uD5pta80tqZFrl4553HgAvT7WPPxGIVdq0dWAYVwuOCQLX6nyo3Wet56gtt0a+
WtH/wYOu4Exjd4/X5Av2u36hpzTr0GYenEtSmyjumF/xv/d6vgt+SLvtjHCrRjOOn9QL5JfsSueZ
IgUMrTqj6IHKJ2DBwjU3+jsET3hkmbSyn7UspRW06FmLFOeeCW+AMnQC3cqxNUaJ7ViyiIv3Y3VO
Jpm/6dA6BQLdb2BZXJK3hxnXVodTqDC8XTGVOepFCI6Q5V39bK3/BEBt1yUcD8FqnY9S9Y0esUvG
ybaBqddnPYpgso14qQLiyjBivMTF0FRQ7q5/YI762lQ66YpacGTZaqRe9JQUpHYsNnwAYCmovN78
kguuwWt1bDaYiZmTeR8WK4P3hBlIBfMSceP9GH+NE8duTwqXWP3Hpj/o7i90R7gGj8mFC5LHWXPW
uQwsrMkkNL5R5iVk8Q4QpVqyU4A2hMG/qAow4Z1pt9xYHT8uWfQzr/rd5L6hp2Ye4Tjkc4bEg1z1
06NZHl6VQ0HtJFiYGV23z8uTAT9piZ0KRzE+HDkJ7sCKRehVrYbJk8+7aEq2LvF+q532bV+Dn8yD
KopMRcY21DHjf1FM+j2yw3BUYv7WY/TcptB3YxBa2LbxUotc4GwyioXf7Yolgv4imfHvgEWK1Rmo
vss223ZQvXvR0kH/W3l8fGM7ZbIkh9ccr1jX+TIk4Y5+7/dtm5cV4h66dm08/EFvtM+9z+3JVSbV
pMX+Pxr0fJhi9E79vOty/v8y37UbIIWUvujLPfAGm5MP/abpxnuA9HI6jErMjRJd06fbAZoIXmZ/
EAuzCllfRe4DySShez8oWs9GGaQjNI+G4ycqaZm7pLZlcqgYBwBwGoXGfVLS2am8TjDT2DwwN5h7
Fhto/PSGxPmjYaau1aoeDPFyKJZzShTjHuRQWj+yacBhVKTzQvihyIZ1nQBTjRBRIRBxDn6qUKOr
OR27riHY0cr9Sv0v5yxdztvojULa0mcoQcDhRlLaOwRhGeyc/zXFSkPbtJycJlj6efl+YX9HAAzc
2J/C4NGuYg/665+msuOQAc4th468zZOXvAcVYFs7oTqC22szOF6VtUvMA7LiDt2/C5gAjC/rpUUK
6XVZpf99QQihZ2gp+hbGiFyvHnn+GRUIAmSQNDShvFr1uYRd896jz6KcNHsrvwet9tuQJGQH7lfE
+GscJoYGIYq2A/lLlQ3Gfxcvuaf8KahwWeUYb2III30r/7v/5o2wRHgcLS0/J8EPLDqW29/UK+Mz
GFJnz55zxrNK1hEXdpcnygNqQN5Jh1zFVoUHIVI+oDsN1NwqQQPF8AB0Fu3o20K1qsZAl0u3MOGd
wTMc1GpqPNjLJUIviWlew0uzgbfTyktgBY4H7PyNcKmT6t0pFWNCAYTP4NNHGDKobMV+xK2vuv4X
w5Szl98f33g+G6vnrWcG1c4j0yKPmMx53gk0PpOsJGt/S+jtdqohjPBosk8ElF27qGO+sirF6qld
SVxBWwqVZVTnK99B9+5A90/9mv+wkt/Xdw/a5BMmroFICLWtryPG4kuX3IVigx0nlIhuQEewhNhQ
r3FR+ad5L/w8kSzDh514w7QXJpQfkORK4W2QATMX3cxos5aWSky8QF/VERxdD5PVHmvwsH88FqRU
+YXkMZZnXiOyFUVaAh7OSIEKrrmCTDwG5RGGFuoF1Vad5I0pG9B2YvWG5zmaivLIZwqCeIzP5agF
YR2vvnEyYYEHbb7AFlBTFL23sl7tRg/2Me9InM2yXYJPjB1hWjY9xy2PuAhA1obIk7yD3caqN+Y4
qOgQpO3WDy6IkrT4/6hQuZFD17TgGHqgBsYx1flWt25Tb4uT9qR8YJN7v66nuEzsQjSf7YFQtL5G
4TMezvc8hKO6pTSKTX3bl9Z9vHcASBTN7qNhjk/e/2D5zp3d+2lCeQXzQVVummr/K54Xx/X/e0HT
D75r2tK2K0e6ODa0/i7cNz/JUmuke8WLPUrZP+nvrg/8HMxK3aUrZVyV3gKJBTPg5TQyADoTDcWm
NLP+leWH6IfM3XbybH2lqQW2qcyFadkhiwyQztB9iiE0cH123TZNWLlh6Owb968I4uTYj1oMImh3
LpZc43y7OWrx2TAYCdrT2Omh+TeaGg7RLcux9yb8nW8Vsyj54mzqY3r6pwZrK97eTP7iO3N74K8q
6S0vZ2wLWKsRhJTN8dsUgHZc9ceZ1VQSA0/Y2fJPyxfX4/q+2fooSjzSH+R+C2VHVVoLpkwcSHAJ
9Xd6fJMPMde9RawfXJl5vd4eL1pTyn0LccHtpMKWogV+bXz/PRHyIeEONKs4erjjqU8Yo2mKJhWG
0yhbUgNqRDA97AibhS8Sop1ZL0vlQGuC89zEKmDMU8IPY4eZiRoecMJQwY6r2JBP/+XJL2LBWBSv
IuLpfipcua9aQUOCfVHY2PQ25aivtxVbBBu7yvU1994GiNYTvQfNuNVBBOnTOKEQOv1F5JDVSmjo
FKGHL0/iPcLUVz6+m8zu1byjJFw/OX06rWs/3JosZWrk02FCmZQVBPI6jBiJ6svnnPPHhBd2OHBB
DjZAZ/yb5+Q9UUYEw+62RY03MFd6lprBI2LenJUfVhjA/QgeF5ey4SsY9mgvnB0O9zHHY6aiuchD
gByRBFqHRMINngbmze+wpNhIx04LYqS+TJPNdYNay/fHreF0tZw6PXh4yMREK8MVBRcJ+2UcGfdb
vPo5yof7GLWg2G5khoKLal0La9wuo8DjyFTJTGZUJ4n/hzdSutVv9S1D9fCxvDNSxjAaOeVqjq1L
bQSTujnBl0l0w6xZt0wGuVeJst1mJDVTOAj0upwRJ2dOb6E0dBeS2Afqv4r6fsw275C/KmYlyOUD
rJ7PaBQ1YzDWHAppmN+l7UPpHsCjTzQG6BdeotNMvOVqqrNbBfZa9pbyz32gySLpapVWTE896hMM
DxMtf/z9VKsHkGC05l6mVol2FVU9SE8ng22YNM97dnR6fAbkoqWoKiP1J/JeQSb778dFuhZb87YO
dQN5e/sXK1uBzZdP3Qp9bbaVQOZsc19hJmkSPTsFqpa11LtSniJtbSjpfa2FRdZQwkQqLBFQT6y+
wS6egXLax+CK2JM+6J/xIXayyRzJDuzk0S+uj0Ip3ozWhyOuaVdchRNHRKvgMRyvtWTDTizFxkoi
nKahp2dTSrrH8MIScJhBEu/AZ/wqvg4osYPgKBXbKHl1X7UvvbNTvDkcMUSHwfuuI7K0fH/Fxt2A
WhDXFOVT+LGSd+G2gNKci7HTniOCkqq+v8uMlMmMzP7PCSs4Oe4OGW5HSMx3tb06IeglFDS0U3jx
VNonBP03vPiEQpqDLymINFzDxbIj3J+v36wy9uzFkYHHZ/yU3efog+aPzPhLn9yTRA2ilxXzmjD/
OQZjA+Dr120i6zNBgXKRKd+1kNMjpsOdb39XKM0OxwiTjCQgYtdP7rntcvTPNxiHI84LhTlNo3j6
Br7dDARSUIzs6VZK03gfKwizKvhnV/dRTDoQXRF/2kDRSmG18CvPmJHzeYFZ+VMR960g+/FYo9Xt
MNRh6dWKldEcVQDlTOhdPjuu94PBUrHpgHK1TgmmKFTrIsUqrfL0ycP6nLwpw29UvLFAqaKANVMf
3v60Te2i8ZtsNotHgtJ45/2CHUzznBE6W1neoZSQuxtbobrAMM7xxOZIV3KgOGHHUVnT+k4jgnU1
lpN/RyPeXadlchILb55S+QweqAt62m5oDIt0yOf95vaA6SunJZWrUMslxrfP1l2OUBkGaafbqwJe
/cuKl/tbcZQqV8AdUVs583+XmL76o26DqWInBn7IFyMiDj6F4+KVuX25VH5j98Vln+aklg+KXfgQ
JCJ7pOUd3GeDU3TVG/8fRvDQvcQJcZUGmiXZmjNfDNcoeGd6YY8+VFr/18AskmegftejHieCyyfc
kySIxIAF8CFTowPfPiC4qA9M46Z1CpkF9xVrXiFY/+9Do3i7OgritBB/gPpwNLfrYGF5irgchfm/
sM0LXgjpiGRqlYNzq8vwSPpoZjsMx3kk/d6v8Y1NrAZrdM7IF4scxIa5973CYA9gx5FqndsPAAx5
nEN8uh/gVJ2r1b6fiJbLBf032DUAoZkIq4bwhA0ekMxGP7U4VFePQs4p13nvMYUnhTzs1APopelk
3ZtLFVrqaDJwg3GxdJfWA9/RMfl6+6HTgohtFf5sYwu37i8qc3M0xzwvEK7jjeiGbUEuZOKoVLZz
xltSnsVA4T+usJlH2hX8WCZe7O4axAAfnClXI/CaSe73dxnZ1xsJu2PX4reUEGsTgbCSoTa2dMm+
1MRQqH5eDRVWOpF/ah8wCIx/6/S7mGO5AnKt7rElark172LL2bo0CBUe52XCpl+hyVvUyyKw0ROw
DYd+5DoIzZNPZxCem6EB9PLd1RtKyPiwqM4EFWeJt4o0YEH6FMb4yY4fePLGuqpQqqvqtjjHmtBX
OTOspptgPzD8QlGx+zakgQ9TJbZoaChEZCFjHHRsY7bXtPck8wOU/c37/54ehIxR7M76Qdq95DL9
CDTCRGEWM+0Y9LdGssmeHUcshEXZ4Qf4r3xKhSO0ZmAkWCylOK5wLw+wseDg/t0FPDbwl5DrfIXM
9C79m1FuIkp5INyGx0Symt0ZfGb8LM2oYE3Lqwf5doFjorVvHLnjo4AwDpEgVAJM/vhi5/2+GgFf
lZ3Wzb8938tda60hUV0dLsdzqqMTZI/VLGhzSrTNYtYnmEE54t1RUj11XPWVCozmuJZ9sb9wN+B0
aR+v1qG1lYeY01Yn0+l3c5mxciJUGpkiDLeNuWvfVhjv0PXiy4pFw5NZ9+9U6MCQzlvaaaLbpvcF
Daf7K0iS1O7AB9JI83ZRmqxces6AQk5oRVd1V7cjZNARZNKD3Sq19hdKxj9tWS5GJhmp9LIPbJfR
e/TnA2AHyDzZaEBxKXBJH+xEQ/hEc8Yh9NPxoGxQfMDT2DNiGdArFnhYUD0AOh5ATaI3l9yK4kLJ
nFLDdvWRkvv8HDIQMF8SLRGie15piW6LPwPDWnAQTMJBnlcVkZucgtqvgrVezSFR0KUgFTKVO2b/
juC6dYJEli1pvbnQUHbaNna53mTQyOKWxWsRujq9kx6b0zGuiOfgZRHr+4r9xKqrEDMazIHw1Qrf
cVIDId0ASfoyZxq5oTqrRI6kPIlKMW8dewuktJLxGwPilPphEa1sv1v6zUpH2sjvn8tVslg6u2xk
UfQqqxGkp8/V9jPPiMAaucheTJS8mk4XJ5ffNBeMd6uB4gtTr/wX9H+4CRHJ6LsCojGlVbvTpZdk
hCf3YZPMG5GyQTXuIYIW1OgL2Jn1JnBkIU3moYRBKYLW0lGbBqtazK4mdjyFXlsrVa+5uhdThILE
MkimDSkePPQ6oJakyD01A7MW8U5u0/fMAqkjw4pxiXxOnrozWxNKi5h5LaHZzBO0q4/edmSBk/bJ
8ddlbFZetfs2FYXLDZazI3nk+CuVhaUQyUwxoQS7KbuTGz2e9B33RUprA+LfJ4IEqEoVARmjfcM8
g65MrRF9zlTQZIakmuPz7xIdOBpnv6k/l1yToFysxiXNUkfdQsRxCw/79uVKCmpUc17xK4u54frc
4OUVH5I+bULlcbyyN2n5G9WFUag1DraQWDtJ/E1O87Bem/CC8VrQK97BFyFca4EFFzsTRfo29gY5
xOY7z8fcjUfs0mblPwrB1wGYp8gQsvDZa6XvvcZcvaXhbGe7aWk3t7WZiml1qTn6FxZJplQlIh0i
A6wKty4+qWy5zjldkEuBALgGnsGf8biptgp/zfRxNI+I8dUwOwnQvR4QLhRE3tVIetXPd1xo8Oqa
1/n3yzvQu0yBkJPYaTdRvmnRtr4tRyVh7OXFVnOwHAG1CopO1nG44vI8qthrs5zucX6xkaxuiJJh
jH+cmbSutIBNaxR/NoYv2zAVfyyBU4w4Z0pQmsv7gonRAuliGLWqqW0xE7QxIhN+5uXATDst5Kmj
CBEqVe58Sg5c+cCPGcSSPr7AZeMUVqBQDAxaRXuSmuVjQNe5sWgCwouu+whBo4ibWeweJQ949NSK
io2oaNCnTAjPvtAKOZ6HqV37Oog0mTJ8WaGTa4Hj/sdAInyMM5HbDUtwe41wpJyNS6eiYhgoaQp4
oJ5OaHqN+zAsgfNcauT5KVyQ4NrZ0q1cOeAoSv8HlAUiQdrJOMDajhb6TYgZ4wScpCZATywJerx9
Ur8oC8euqryR7VWxIbypTo0p+zZmh5IwSiBi4JLmzpf0whA+35SUqNaFEsNDL8xAvpD+XcrIO08e
HGnIt/+lPRP8rlz1knnCcJjW4DSD3E8MEWfYNcuhOPRcOYZsXhmfa3z9irrEg7yV9TGJblO6jJ8O
4CNRQBjeKBZTt64idm7fITUDlfx6RYsm9j1tpdEsio5Ra4MgjAzfICIWwfHM7DvwcQFTywIYOd4g
YIcw19VilL4xqYvbcjHpjzlXzIQy+0TUkhKErsG+X3btPg8lxj5XvV3Q6DnBy6Q7fMsGFoFQU8sB
tmfasAPaS88H6goy0O/ZzBPGGR/42vFlZg9x80tXpU192SVeJYEXCvwcJf+Lhrg5M+jSobT4oGBd
awxhFQiYdaVqQi3yt5EM3z17TeZDSWHGkfcH3l0GxJW4V3TU7y+DxR7cas3Pa2l5BplGUk7yuZf7
jiwrwQo4VaFkX9+tuHu/HcYSwjPMrr58a0vx5T0X8ugjbj3S3Td9blxns7IcyKTp2uvDXOvZSWgB
wtFtDY39kQ8gpVG1sycbpv30BpvR6Iq1U6j4ytMoNu8qR+TpoqqztUn6DBfSxRAyvv/vgglXqkoS
1dCtcUGfOtjG11C3LGUkZ1mAxcKk+5DrVUgFg+PKrFBO4zJ7g/XW/pJwdu2630hpPd53WSZCk1sv
X2m17+eBdzrI3FE5zQao26pFYDM/VihUrlFqtpevVhm4rzxN7JMx4kmkfxzMedZm2j0dzJUTmIOM
gwwRl6Y7g3nhOHIRIIV7iqQSa+b+9em17/A7HIhUalVOJvhWYo1Y0pYvgZkbpwGNPANNR6YaxVnW
wItSJGMuPqN45dK/mazS3lW/0tO5jgTOAe1U243QUACDeyFKYtWTeIlKtvLNnXQwnIvV3/AKYSAQ
2gl1aETxNN7iWtc2+AwFP1ZcLHj4y3EKDsLaqCWaKsbF4c9mI9CcYonEOwpzywqnngiwuilGAcmy
vLkoBazAPhhyGs4pD0FYk3yB5VYz2JnBd3kgfP0poHBhn/se4ZX1KnvG+JvIsxYTzwbkCjMx+8Qr
BinjMGasivkzh2EEzi1KtRdLMQOosj+q+3oLTyPfTzervMYwIBE4QxYeORaMHdIZBbe7N++En0QY
bO8AIYvF0qdfuObF5E8iB5fUiutin0RQzFtJk+3fw6dhK6x5hSNOTClHJmkDflyShbXMaLKKcJ/5
feM5aQgn9CmX0VKWArPsjuZdyibaHcIalCJv4q6S9H5ShRi8PWDJ0/La1tlI+IzSTjZOemNO4S6l
kCBQDxg6LIpR30RHLVQQmmOza3gVLpPI8/5Bs/R8fXxPbxOQUrhbBpnPorlTCblW5SX2hn/YYBup
REe0JA5h2XRz796zFbAhgh8lLAIhsqCYo2PojPWMhCiLqa75An4JBBYKIwF9LEF+/zb+SVVZSlDS
Bum50P2OObjQQ1Q4On5uGs1Q95bVyGOY7r35TOpmvDirrEf8VvnpAgcS9D+A+hSLUbPko2xwusSC
7nU1TPOMeHH+zns2LQhU6MfLYPJ00IrSCX7v5S+ibdObpBFUqX/UBxzlBTd4rzjWcuhGfDXZPgI6
vC2zVXOvWKeh9dbPu6td+s3cXV2yTUDxherp0cy9HMHz1ruJg+VXl66QiU0atmDvgB+5sRyUSYcd
KSARXTAJYAGgYQHY9/DvhSou3N+XKDk33FfYl+LM45JqioecD+VZTeqybvNSuLZshI6NtJ6Dbz8C
a0qM5XDATt0oXENwoJlrpjZwo2xjNi4KAD28TrDSeCQO2Zef8HgGe4ZZQax8xnOrirogMX767rAb
aEZ/03PYU5G85TXUJw14L73EZak5RlcRffkfqN3fdf2/n1lTp4ZWJys+59dVuKk05fDALpGx9UDf
YmZvMRucBGttdq+2wp3rOPKafa+C3+xw9D+9bMpgWOAR/JT5xs5YAbJGD/yEYxE7X+BUjxKYRy/F
0g+wgG+qx2XuY+CLDBrdHjbLLMn7k2+lq5lYNXt5WycZ0g+wZJKRGRqHbLoeB0mhpyQxe5xmstci
EC6uEY76OkPCTrhJHdlCg4N1SIwXq/AiGc0X6OrlvFImdaTJD3qXAW2pAK3MMI+xa410kYFj/1QW
2thdIu37ktKn+jbws8e3By2OBxiMLYOt8LuyPTkwk20+FZtuZCYz8MeUKvnafsHQpb64LZI+0KGK
7GKmAZ58TBuLuS3u6V85Vjb+5lOyBXNCozbAaFsVGQCXTBZCAkfDaj4ZaS5fa3dOHLRCIBUHd4Y2
/b6LCsmx2oZVvHeqxxdj7YwiGAyXagsLk4g54YMZn6VSQY3Ww08hcazqh278SSNgmWlGnxBUNGDy
wzGHTbaZFlzmMetS6pjhZDMXjbrQH/1BuTjKlYRg0nLpNmY2r8i922yTGXUurrB7pHYg3hsdM2tb
HXqUJ6SYR2iZuHnJxRu+UqhEN75KL3trsBwjunuO/X3+M9E+tg0rrWgtdoy95scZjl/UNm8QWfea
Wav1LWLhALhEva4ymnjjBoY/pi4eMMmnFgDtgiHfbIUPPen5g2dFKuClxjVkUibgKord4Gk9lnma
igYkqHIxmwh1XL1Kjv49O5CcyXSHXkAAJ9582aKfjfj6lSFiyeVIVWekgvOkFRxUyvTuG64wlWoi
5jLa2No6W/Dh7F+XgNib9hO6JBepvruImMKUlsLu33J+Xy3NdKnGndU91pb9caJPjNUAN21ZFBfa
+yKq4SCzNdMIP0/Oa3Kq8Zqgg6+bLvGGuC4AHz3uEH9zAAfBEl5C/13262/Qdu80obQWJxoJvyTx
qTf0lEvut2XXr7JQ8YzLQ9KXXiw+9ytMfkCulkhm3KxtRxv0vS/qlCfKJUVsOIJP35AMEtsGGU3C
6XXhDSIitczEZhVFXyl/87vwBCSkP+9k6gJKHUSdTzGSNPLzEgIw055kcMYW/zGqj/xa154CjDtA
9zBeHT2M5QAJ8JZ/MZvIcAMNxUQ1SWcUT0R9nDC30CK+S+5VLkyVJw3AO/feD9UhhqtnMPHzryws
5+DbEecRFPDNog3rVwBXa2iRpUo5bNuU+lm9fSYOs+y5BfJoy8WjU+XIpk+LsxmJs4DBI8V7KFkk
I3mCBtaSMp4rTT7Bc3NrzwVDNpvYRJy2PpFEMPSJU6n7lS1xhkHHsaTxbq50r5bbwOETPrpz6ULy
2v3hM3PTvAMzIucHoqMdbRqoVtvskYosVLymICjaimyFbL8aliBDiXNKkTBkf0PBzhxZilRGAfLB
cRRBJHVasy2ElTMFC0/9YJgU1GBjJWFecLlvgcIYqdFmF5mHf/CicoukA/sLg9ljZQKh/28V29pI
rRDn/Wem/BDflE8myUjnfh3/X5/4+hgdmcOegonlWO+vYZLV4IqO4zNRDIKm2RH9VhdNw+mMWgdg
cQ8CHOESh5quLtGvGXsSsAv4QJy+j65XlWYsRaymFxWxO38TXVhwUqjzzyBmxfuH33OYFxaKZr8W
muiQttrvS70UTr8M7oEt6Pj3UE43Pb2erlgA4//1kDaK44WbnWVMDVLQF1I3a9axbO2GU8GQepO4
ItCk8xoY/TPrWGrPvEXcnnChQm/yG/URHC+1dA+tO8p1cwfEUoVqwR2QRrWsbsIFUVThIbhAwLx3
xdJ5AjfwFH3opOOleBKDUOHlnwtJxrBLibuiemDHZLh3W4Z76U9yojYc6efHQNeCIvxGzrDLdDMN
TmmnuzWGV7XukfkAGB4Ybpf2HRl9HdCVmXfrvd15QSDfrlsQIkQ2+Hbx9l+6U8bJCYI6yGE0GLnv
PtVDbMRatpbn595NtFuHhDSivNo0UvEujH5hghBhiVFLAfTji/MzJVRCIOgSDrOjMyqlAbkI6QIs
ZhxckN4/+p3jsk7Ur4G+t94/MnDYHDohmi/PmkRQ4btrEVtbZvd3NIQ6/pXyIxUm8JzwyziGoNI4
kwiJyiVyDtrSv5rjGm1XupD9rJv9R5xtpnMz/r53C+cz4PadnA2mTc88/ClAIBXbHUfDVZQviVdC
ZMbx/qazOk8F/Em1tWr8e5XfS46Xh1npNHEZ16QJAXBDAKe45w6H5dcaYUsd0fJpR/3RMQ3o/UEi
cEGdnLem70zBqz7RcaEuB280YR3mHSY+iARPq1ibSEdzVi+E/zI/2RSujtIQdcpkfiWDj/Sj2YXa
f8LHhFd/QqeTIOC90XN/Lq3sCtss0/gRb4EhV9TAUWVgLKsf1/BLtbGSchEhcbIxMcofkJjxO+0T
PtIugqpXqksPm9dq8Hiu30XHDvIn0E5jOT5WBMZfLaYTDO0pbYpweuPuXCUjW5vdaRxM9p2BHG37
Di+w4O8PS+AHmI5zwB1u+A/Ja1qqWxmQoo2aCw8FDFwnMASbnqyrFV7MRHv1CC6lzOdTNhW/GZr3
9RlQWCJHY3n8ZMMJvCRDoDO7dOvaAP/GUnaYRYgZs8mSb5Xa6lQC5mi6g0qdg/76gkVSCpQ6Ubp1
H8mN994qZ/C8edvHAgRUf2/g7I2I7PP6AXZj+yryYE/ZuXFeTj7OlQLdb4C4Fi9H6pMeOwcRjAdW
450NQJve8EAZKuRht4cxFbiK6Uk4NZOOKNvq8AqJlnLeX7XalmZ50tWqDbllMivPo4+dakZqYMrv
lY62HXkgwElhkvX/9IIvHBW7qge+Wa3HItBFtWG48Ib/pen1e+i0C6Wcx/ellpKXsMBUvZVeGFsp
BlHvQv3JEsT11ESqOIXfX8KATAAn4tAaChYrPsj3EInFh8ouV107IoUAu7YS9v6WOIHXhGyRGX6C
BZczong4jssO87vuoPgaSz9qpJdK/Hd4IA5SEzFCU8E+eHQ3v+Ya5K47TOoGvAPNIMwE4vyWTOZp
Cp0EHvVkUw4yWRqnxB8nj233J4v1TjfO+ItHBYmZDVAhdSAWbltRBxdE2EiUEPltc7W2Rlit4eU+
nyIOaeQpL8uY3aRuOgXdnzbw42H65yHYF+jeuCP2iVyvG8gGzqOfyeQCn/UZuNBXnIbe303BWWHS
Y7sOPBBsrMSsGz59SFDD7c6Nsr5uFJDGGrPhSrULngcWCjWLyyM9qflUmY3DxxPVtYheYtQuunan
JP8g1EPuvtDQJ/pO7RZayJRQP4p3aXB5xtveM6oRNY/GzWXrJ/mGJpIorH4F9Ff07tp0vIOC86e+
ZHIKaecQDyKxD6xEgePjJ3QwyImOljNFRSXWaJH43j7+GxRMO1+jTUVYtf502hl7lSsc9kS6Dh9a
xatSEyeM6HM88v/pJZVjxDMgHX+NuoaA1itlWpkXiA0o1Ng4mWDg/62z11ELc0EcKydbdg6mUX3l
gLxK5Od5/K9UzkyHnUJpZ+BaidSKuQNc1sngAl141zJjPUcR0n6v9Zi0CerQXU+bPQ9HjvhG+Y1j
jg3mCzWLePYQRkbAr3T9/6+hUJgcfdW828Abp+/gQvFuybGFTkTOVvctpvqOY9gvfW7bYFZa76SQ
oUoQQn8IxWVxlbwcrh9gAobBnheo3C+FQEA/FO48vBFljgd4f1Mma+4CDcIgVJa3sxBWP1IgCS5e
RJ4TBLkEwS5kd6XvKeCGCvV8cTYoUL6CCaUyEXnq5mE7vTjAzw7oW2xBYBgivlNWMzROe79wbqk3
D3CmW8zDAuSw9BoTiHYB69w39Bu8NymFpbTcVssqtXwoC3PWbkiwvgAHcYVW3Af/8AtuS0GeQuvO
uixsd33zvSIvX3FpN2SnRpbQXaRoH/5QFsxLNms30TxP3XW6FSTf4aDMqGltD/pacT+ESne0e5r+
iZA0FSOSEE21lo0JPL2Pndub8dmrjyBtiuLwEch02lZAJvgULRlX9fR22eZT6Eh1lPMksjRcXT8E
O2ysfVH+6N7vGNauN+hpLc857V9PJhWBNF6mWU+9iqm8GcquP0m2JNyQ7Zp6VNm77SHyXayhc/7Z
FRL6qIZ2q+som/hsw91BvUSGkEcRoN1eQwsSHqTi1nmm/aOyvbxW7asxkVX2EEw1Y2fE8Hfl1+Tb
vN6zOBkEF3hjAMT98jfW/cSQ3MF5G7aW7XKyemOlrNhGXJOfMU1bgX8FfOrFWtxEv1e0ZLNXHes/
NgPveNR1Z04g8CpAhTENLMfDsVsSIgv6kDDZM50dFjv0wjwSgUpAl665WVz24dQ8VSPxBBwJWo3L
NReFW1hnsbwL8T4fi8I5Ry3NqcHBbyXgZwGFQKrBoRytBhB1qpAvkAymKS5ZHtDEGgFfRuk1kWHy
d/OGNZNFxwLSb9kAkmQXg/6jAUbwqV6TZqPvtuguayZ1ER0uPUeTDMb/GTJ2MC/A2euAE9gR+rKn
kBYvj7biilRgWvOUJtfYCSwsLFYyMK/ueDVO8Rge1famaij6oUnPvasQi/Z5Hwp00NYZZMVPZPvu
/BkH9IzPlCo6HnSNTc5tY8slHNNj2cXO0i2xJZ3c5K7i3gcnlH7Tpqb1jUnAzUcRHCUI2g77kqVB
F7ZvdO+zeUgIha4sMAQp0yNkO2sPqy1Nmw+RQnhxdN1eSSKGBHFYb7//FC3HW73Tx4Q32CIJ9zR6
zUEPFqKFxSCNpre6VYZZp3bi0kcX/7np1iO7QHNMm6wsl/L9o7R6abLm1GFPkJoPUlfXkoRBOWKI
sxd4KLBb6JzYbjqI6Wgo/OnluLs/4rJYSHTwteKiIdZ3dAwLOZc7VqeXZLd72Zn3a9f3DT8YVS6w
mHX8O6+exH6qE5LNtYCzODS+E4rJmZLJA0p99RExn/CtYtCsvTvvbG+TiQkHtkyYj4h7B3amx/Sz
2r4slffwWFybNflcIfzH9iHek0qGCfw5JqBagaXv6ECBn3v8TJ3B5mCDEy/34NJufwN7kzPqM+7d
mFl2X7PboDw82KYnpDpfPAnjBWnq22UO0NfWbypp7kIjE5OEXTP6plvqKvTbK7Hgs1nE25Gx/Gu9
j8BXNI08+8cQtBkQOMJiw2haHI1aFWqO0DVL0daUaaJke8Pb36lrsryvvabh3MqGM3FFlbkGZKVw
lK4wCm/zDE0ld19BnUJWFqfZ5YhNyXDOHb/kO0VEichmQGLN9wqcfC/x9zi1G6Xx4GkEXFWDoPdr
HIlLWhWWe25eTl54XoC/Z0Xt4abc5BTvWW97W048ZBJWn1Z3Y7Cy0kF9Qi9MVPwvdx1svPEsHmcS
NjKAUBoa9Xi6DwpT3gZ9ZvfOjRkVP7bQ0u05pKtpHMpwR6NvqR8qYKAdNW4RzinIcD8F9wCfzVT5
Jg6MFDlA7fT8E/LdTpos/6qa2KXoXuxR/SYd4s9WsSpnIc0gCHvsPoAPUSRXU+AbOhqL2r5Af6wl
BPkNWHBFbNgvHN1SJE1ccJ0m5tTKgs3azey5W449XA0ZOnMSVIZf89+uue7gWMlk2eeZi1CpOYKP
0olMDStyztcnfw+tiIX+DpGXtuKZea+th9+rSEwguzhQRemIgFyGIT50khsJ9L9KYImkONQG+sT1
wjunrehIhY2g8x8yLStpw3OZEIeataIe98E39XsI/2LmOr/oagCT2weeVDeqynl/vZuquBxpv6gP
teFmAGxFD+WuusfLcGQLOaHQIewkF/lb9SYe1zw3itxGOGY+q3keM6YGQdpmuHo4w91hbZDZuJX9
4PPi+Qa2Ts6D9jFri8l5u3IuNoqFPVMpfzJ7PJjtWDYYdw3DK+hdCrub5Yl6WAIt5PxtMiHEpplS
vXFKmJFcwyykuGt5MJDUj9sXASlknacspBpzMLeHeUgNTryNgIlgUgIGmVT18EEUPqqMXQMb6vCC
2CDItMIv070AXq8zaGfMGL47+fQKNYRjIpIx8hGTZAqWS7BvER7wPzTcfxQ4KLOQ02INZWegnSi3
NczXkZ+Osh7drvqJL7zaPc/mF+505XaEc1GqGM1AwR1+1BrYG2ge1ccErl1vBsgw3/GIjMkq9Zda
ixbsKwtW+v+Pa0Pl/Ss65VK2+d3jBHKvt7yZy7wAFkkxyuH4V+UTG59QwJvTUALBAOtRJdK/zac7
ZTQH/VA0LbAkzE5ckJUl/K66BE9vIlGBeaM11B+xC8RTxbXKzxaDx2y5CIcBh9d1jkOy9KI2aIf1
7TPi3czomOroqY+xO9wpuQt7aItRhVhKbvmUAzZNcqZcFWgyjTvsQE6Kxpi71azBZEYrczpLFO7r
TIEZv26H3DozHYKBjyuVN3pb2fVOQnL/GquShszdvh6TcCv91NXWyQcAkyPu5Xg2uBQPxRJX1PPO
LanGOQa/rYrValxB0gN9Xf+D4Tb2t5AFGsng87lsLFv+lgKDAPV3FN/9kpbyKxdg6YFF9QQyO6MI
z8umPaURxdkE3Kd3IYBSoX4lLjnORTBpk5Ozpddhk0sv4XmZ3uUVT+mXIX9yrD4tesWBaGAbIEXs
yTr/QiFnGepUjiVdN+UzBUN7oEZBGu7l6s8e+psyIbAyg1EGU19+tXfMzRt5ENAcmfML7i6td9sY
6QvqImXFM/zHGFo/VwbdUMbz7ifj+CVzQ/4/W1odddjay3cq1hdSInpdiAEt78FWWmpr/h9Q/R9Z
ZAi+bhbBqWRFe/aV2CKdzwcqP5FTRgqFQeDY1WHod23V36UF0qWA+wBuxvBlqx0neN7UlUFE6kE0
zp/Ghyq1L6BS0zWFn+ZRW1ZdUhuw3NSf0o6NCHtKXa+jhp+X+FzeuY66M58DvVUk22oHCUW005HZ
Awl9daRaR3XLAnJsDQZdv4V2FyQWkj6xSQ9yC3UsRa+OilsJWz3LvwaJPDsdCV6vu7NMvP5grFto
GKldk9ylPxa3cnuGzK3/KrOcO7dLTgpFTAwSFCPsI+kJi/drXQGyG/A2W+q6WRSM/eSnYLVdFYJ/
QoOE3GddP5Q7ygx0HMG55A+4u6zYa1FFQWVFOSWun7r5+gWe4XzHuxPtQuPWGoqHIZqFC3gmHxqH
9V7zCDdo964V9lYE/q7aIGP/cThyjhd0nKavouR5XSgr5pg/897LKeoJBO/HT50Qd7nHAgsH9s8R
hvjABCf/UbCtVZRsCuicQH/QSAOIxoe5xFTeWN3xmHWyzGwFG6dRDNLhL96OSwYPT6buwYItHuG8
OVzFIdDb/vyGc4wR4aaVzWpnZTf06MeV5AbJ9czbqO4eT8/mCWkr+lLJhBqSr0+WLPUx19seJum3
sXIQgS3knG1kE2+7IxDGvaZ4AKfRt66k6mShO3PcAwq/t47mgeXERC3ND4aela1pu8DBCsEYQfcw
S792P6vRj5vqA3i4doQW95UzJG0+NaTIJxcqH2fONXcT/bMxi6ZywJTEI1yzxCI4K2NATDpAicpj
QxOSDJnD3e77jQzno96fLu0m8H+QydOdPuOESr0LWN8Rd5ZuPKqHNmnzdmH73u1rh7H5Yp9oDtC4
BPRGQWkQZvKkymN6SzL4sHjtbTjxjPbSByngTduvMJR9Z2nDNKw5phBYhxliFH8B8We8oy2IaAXH
Re+6NXkK8+Kq+UWfNkA9O2z6W7iuXUsFBgdU6eUcKkpXzA3wfOP1UOECE7S03M3vhFqx4J2ssjnX
D8CiqEao1nu07hRESoUPaY/ZqV6XAb0TAcUinZwtBE//fthedwCxSB/DEuxzbXbQ1AL7Q8eNDVwU
86tSsnQo/RwTh+XATDdTdBTHLpxvHkzFRvRXDTY1dZi71ZxepeOERRZDxW8mRx7b9/EFAp6zGpea
ET186KSO3wp2VugqvwfE36cFUgyXhsNb2UTSMrJvaqLqnRNV8Bu9f1kXOZSx5N2106aAxcwjOBgM
QnTsy3n1qSTm4/QTaDhjZHhwrwqMIXpSY05S6guOMtg4R5rJ1q/zO8NIhVkdG/TbIZTbtVJbxpro
gpFcXMyY6smpTqChyuz/c98PLvhQmIOJllSKkH/wcD5MYsj1GXdd4vMVFHcR9ea1Ilb3jx1r3V8G
w+vcjUsZ0cshQq43uKH08Tie+GPpKlUnCssfYzpf9kai38Uhtl/aULF6cNJggMONXIHeudobjGml
uGgNvSPpk6Jw8r1TIziUcCQo9+Zo5AafQvHgIrJhh73j4wsf81qmDljGo0GBZwt/jQKxERmMuo2i
00EYbr7PvPvNTsQFxGuYZKM04jiVfKwsB4lbDA0DjFiDR+tbjZAu3zN8Ag+Ua10L8KiDij2nic+P
xbfn08xaU9RjE7JsxB89pVRRDLP86+Ur6SGLGK4Tl5J3QWiIim6j1SNBmpzB2e/Qx9LRbE82FGp1
SkXe/KU0cPidJUGrzt12/oT9w6jW8/2vEkMOEhPUm6NXkZCKxFQ6rXYtVk8cgitmuvrzjnjG+lq9
0GCWPXm8gDw3gGTdNrKmL5XxE6D+9vutrk2Nb3o+EICTNBeH+iBxBAzjCzQmL5vRgtXvCZNAVo7v
kAYpA7LfnvZR6hfX4cNosoW2iRbrb2nllFDw+0td3FZGRUyVOI/pCXfdlfPC3GjmUZ6bco+M7r8D
mqUWvqyfF7uhmEgipEKd5WYhkIZUC5TmLvfeGYU+eOkDmWP2zh8olaEFpu85KFdyDNhy1+TtTbw8
6Q94uvNNBck3Wb9HCpZU6d/wrGA6e5MerrGsVIXZFkzsYuWsGMYri2MHAWPwuk26i3EveQWXcR03
D5rMFAcX+3blc0WEX5rgFqIp6sAfaeYtLrsnW0Tys0+JNw1TBFyS8unjUwPNC5035S893wdPwP2L
cTbfj6SrhZTv6egyLX9nFnG/9SfEzOs672hNJUAxwJEePwrc7o0KBQ8LxufUZXmlpreAgEfjcgJd
U6EMdakfmKCQLrc6ngZw8ZwIJjWB+XHLtDTfdWrZbNAHi76ux0VuEdiLB87QKnHae6mO2Aoy4ERx
sbD4QF81uudRlKkne6TIGHcrNKRx/IOcsontPIoXIVJt+swp0PnJj8xrAFdXYU0eA54yfQsms98+
gHbzSqO4UmjvbdPt4gyq646jgiw43ZWUUByEPTRF9gch8VFC2k9Cf6HO0c7Nw9Obc8fpcFveBEwT
Lg57HGus+GzFuXxVAa7xH1CRcZeWFIYHcq2jPB9Ijocl3RrCvWXV1OiF3JZ1OUnvwj6IaCiAen/C
moUtldqyMCuwS4IAycYCZFaF6Qr+sZJr/XznwjBqUpF/7flNyJgGgr6U8sIE4C14uuVGBRvjicbt
rJ/vUlSEHvXVKMdn+dd94/wIzekTvN2FlE/AVSJo/coymkPd9GXcAwfqBNyf2dRPHqFaI53mSPhx
sdo/MafcyTrq/B3MJ9QfUfE83qZdiU60jsaN9qjxfSH0GL2cU5sgIiuvSNhN0McXi72YwzBGV7Eh
9qn4+8bZaErR61vKxdT4RXNPeEUZQnooFA9+JZYMvGVfPnVTXWpdTxPTQAl6fXlKfPxQveMbIFjB
cnbFUjriQq14R75LkMY8r0GnQbMAR6hAo0WaV7BLAensUvANI9wFAutuZBB40qHlr7Phw46cfSUq
tv+GJrzKQ6bqRzk+UyQOkS5G0nlzfyRLp3xFPy+f/ZWsA0ER+ymljJmx/G65FLdmpcsG6ybZxo9l
x3B+Oy5FFUyqBhJ//g91M/ToVdGT/AY79UaLJPru0TcsUpmrkEWn2naoCgAAvUG1vbPvr0p7r9Tg
iDtggZCJMuAmJtJj9ooUnhPdCTLsKBaYSxwjhOY4ZmnB5sb3Hwlmm6p1tOixETzpshnunyxU26Ob
cRlzUuM11IxyF+aajtD3SE4SFMoa8zyTH6r5o0fy6cLtQyRpSMLzBFyIz7z68UPvZR6AJ6dtgtV+
M4fosKgjDgC8/9jGJey3WbOZeI7buxk/QFv2aXsW3hVG5EbR2biIsfSCeIl13hwAL9jlbgNX4iGr
OEXTPrKh5aOaCiyM/xPP4AdL7jCw4qBQxQ+5zi6b64SZF3Q8Moq2Ed+P5UP3zLAZnvIIxmzfI/NL
JS4HCF9RcRpKpn3ft/deytB8uLHSlH7SKq32X4+lijzAD+qbXWB6fbTmrLLEzLwfe0BMgtpODe9W
q8PZESJlO8v7thcr9MKfi9No/26X7r7hfzFjrIwtFWA+lZgcaFeEWx9i2oD3dVF/eeE1teDKkcwO
J+Db6FQQv9ZFAO0t3OSDRLcQFr4pouicQ+WrFLoYMN66S3ErR1HTjEvSYVNPSgCLRkzK9W36S0UI
VCMk6cKwBTtj55zsDw9wna33ObzjQJJwoFxCsJM41kijyUAuynDjGAFql0FY2uae/LId3xIXxTqe
GBQPL5rHYtFTaJrvXIcGqb0Q+/bPpbnwM4Qe6+dDoqy5MU1DxhNv+abhGppfNc1jPVRKHBruvmae
mDiUBdjWJo44noqHtvq/KdasdYkJr/8+2mCjB5fGV2YVIIZBtebjLMI+R6Sh2yPNLkl257l1dwai
qQJbZQsJgGk5SzOLHjZcRJ6uz4T0sT42G8nwZvf7h1Oa6R0lBgieD0bfB96jCcsHmV1vyMcARPUE
I++E1nh7rOuLFXG6zPQQzYnPlRip4AiBl59ylvf10O1EzbvZ6n98U//O3WsVegNbIWVSiQ8LwbZ3
aGkCnVi+GDhGa5e3PxEdBczajnjPStJ/QKADgVPxv1GdcNe6wmVU0UYLWY3eJyyUD3tEhB769WJ3
4h7xcfUkiPYTb2sUJjoi0brLdlwXUw7+TX05hLOk0b1MTa9RBpkJeY0C5B7VLfWhuGHL1kZxkO1e
vHIObtSIsgdQoyarmeGoHOmjRAYP+sHHHPT2nzJAWT+YTTPWoXto7ffnIc6Oc9CdE6D6ElcUeeIB
5gjmho5J1JHtDTmAXC9UDSZE9mv/u6tqMVvXNcs3w8b0rmqKroLiF8Tkv0BcKahN5O0C/tlv2OHH
mNUuBwSow+oOLq9XzwaBwA3pqDOi56yxORnM5vzJYfB25fOGZBNo+yXU1tb/bBJxUJ1uPzaw1xfo
QY5tscqU3SoPQfI8ipnGqQGrZyB2d8Czcv5WRZsVE8QA5Lrtb2bLlQUM+MGEEdBuBrbSotMlaUe0
792l6maS6fD75LFWtQMXI0TVToHHeV3wD1jVvBJnfqrZ+OQN+KBmqlCkkxRoXtZUyvb+j9Bdvv6w
nbMYSdzN6hb88y8bx8dIkBaqrPE+YN+a2SrxlAGLJo+b198zh90Ywc9veC67TN2TdACV+bJeE7dI
ynAZr5sy9ipFJgDnFqfYke1awzs0dXALoi+snMYBYuM4vfjr/13D8f3i8zOm2txBOe6F7w1qBysT
+JTyyfKUlGPstmhysQ6rVlmH66kTR4pCtw839JYB23Yh8c8YfznGHNvhVj7ch4jgyZm3ucJl9E/e
W1/h8o+x3RRvYA4wA5rZsrzKApeGximM7raub1bEDmUdEivkeKxK7fVt7qr+POCerH16UX9GWwG0
dVxmBHKS5e8UTXVKYdwxdrFp+VkLBS0Ef5RnRjBFUQd1fymfIB8aLWzln1iEa7Smnjqm5FeHMORD
Ez8ek2klfc8TOuCQRe54HKe1+5fG/5KY1Yx4OmMqWn2e6PRDvt985o0e3VfKyRmd/pCeKLDZsJhe
9+gA5OEEnLLIWpc3szFw4j3Tp389QtxqPefQYu58OgVd0gQ0b7cS2npTZa7pKyRjOPbvZtwEa75t
2niV9jxkLssr3qAoiGDUoiz9R3haRO92oSiyaZq4aezf57KcgjrOlUcIG/Iooac72a+bKaln2dic
rwdPKfv8BcrI4e7l1bO9DJxdr42GlE0eVZ5QFoJBY9Ak5FAb4plaDFtLbKK9X6eN7bMkgqbzOQ6G
hx++cO4q5i1EbY+Uafuzac5dkvjRkSFn4S52PMkIetqZfNGhQMQX5ZROLgh2P9TnKUalonvmcBa2
6WUmT3SmlLvV3K0gAUKcR8FqZfUva8tBrAc3TV1o+q3ObKCg97olj0X9SOroy2XG9Q3hR3daqaSa
cnGF4/bFAG7lJKegDOq0lSo371sT+5mzktzLTjgqQ9vOn43q8/pHLxwqjcpA2ug5jmmbFnZeULwQ
FvhiG2dzHFdYAMJxILVFvXdFdKezFnIHxaoCKvOS9tiWoNDbe7gn7BpQWU8CrMZ/FD4KTM/+MoEd
GyGWZa8SV7v9nm60burxEWtMtoJ/EOgo60OcYKyEOm23NrvGOw4PpHO1c41Y7krrf+hPIZ8SXD6W
W7eEn7rHhD5CZWIFqNXHJ7bi/86fOqLzSWSB5LGa76V0OceMDjaf63oD/Q1nucrVkdFTCM9uoVSL
l8xCGkAVdOy2E4t+qQTge/QWQORYkyaZTtcwrWge5w6B6aQISjvghp+cDW4/aS883CWZ8LThQi03
8C8cti5/j/oNtpK4V41mKNFQvVvpd5gnfUkio6pTY7NUjkqoxOjNfC0MDjSDtNiFvdpzeD5lyRvV
z/JzGAPeCXJ9I6/TIWJNgNyHRQes7gZ0rsCyzoEcv5PGJtx+USB2aROHHKFkS9KjIN5PWgW4VJwC
ku0TgxD40q4Ln+svbuDiuN0y5nRbLQl1h4yUGSDrg0UYpGSBj4qQCCQfBrcotBrC28Z+fFmu6Jn4
clhPeidU0CJWRb5CUl1HlpNXpl32R9FXNH6HYI6ap5jN2Tn5TOWslbBliUBue6ZUduwhICl1Fuga
VN0ONaiekw1c2gWOWAOFLGMTiip9prxdTanx8EV6agIb4HYbIAmbwfENYWNchyHRJL+sjbvKSL+v
1xvJkDpELUQsW5Mw9maDB43ql2FNahs6TMFhzbEqGAw/4CwDVZ0ZKGY78VaJrmjnP6S+/mWKKdKi
tKxRpPmH1cUvvcxlEVcIVxqx47cYom1bfyfqjbQMcQ+Xr8yZj+kfno5WjpZg4rDKfeAkEgCx8cN7
uUjeOd3NDxl0UDzJapfWuZXdki/+tBC292gSp05Iv7nHtiDRRR8TiOyzpmCQIDy6q0EMRRHioCbh
fY4X8akMKQZZilDLYf04146MHHky6w+e2KZohrFccuehg77IJJGlC1NOtIlWUQZaSFM2KNHy1k/u
IzGFoSdu691Nr5cPucnIq8QCmL0MrO8pTv5MnY2liE/9X3cvROxRhcgtOlgjvNKTOuV/Oyc1IQx5
P1txQWN35/TOfzPYFxAi53j8LB+pr9xA53Yf0lWK6vlY+WsbO2aJp3Vid/K6eCUuP9XziYsO/1uk
6P9Xyt3fup7Vi1pm/7FRxu3Xeob7N+iBdXTUc+6DhEFnjpmXF8yUVU3n0RCs5QjbH6SVeCHp8ECE
wiDuDQs68oKBtXaJ0lOFIfwMz3O2o3Hbkbq4HWIzxwqBRvKUASGS8zg3zythRWlQ/CC+0juK9LcG
BG4AAP7E3fM5YmK+XLoJFuKFzN8KR6gxUXWLmieOcscRK6mzVpPCLu6aC+wuUbsCGC0JUqrppmQd
i6RRTFzZh/9U90ol7uuYVdaJYD21tvKBqqlQcbFUACv2f9f4TYQYrVYOJXLgUZ0JRPfhxUkx1tXJ
dVoq3uWxt0xP0vOmVkQY/NcV094Eda0G9/oruKSK/Dc/saGi9IxI/54I1j1NWHXFtfgwcMnMDzb+
m8kFxSs8OuhvecnWpWNxTeweLsUvLcZiD7Xzt6oL/nKU8/fL6Md5jzETMg3npPaybojOMScMGAcx
TO20OhgVOFsE5ywAGzulecUDGWCq3OPdNTX037/9+sBjgZUbPRc9wJxTAoClP6LsvsOXstJIhf+U
gBZROEbdX/GpejBWMm+gaS+qpAauk3Oo6C0KP11W7uDjA6obIiy5YmJfLY27B7HxphX2Ni6z3QBk
1fbm3D2qRihK2m14xl+81mVJEfeHHbA9VMpY2lNJ09V8xK29J/SF4zqPEFbYQGFvz0LRT/0XRUXX
lC3evqU6CDzi9TS6binaVUaXGl1hbaIlRAY2kWJqngWrr7B/znm83P9iOiJkXErCB75jqCWU7+ec
Pg4IQ/NNp6v6mb45GfSuw7gtmJN2qLJYFmgGdlF/AlnYLZi6UxAmXS14wKZ0ot5q1NQIGH3641HB
AZYBJi32Is1dEZQjMdP9GxH4RRzZ2Yp+SUmvOpde3NX3uCGi8As8QgTFeHoPZbJOWRCbsMuPB070
WQPzpa3btNzq4WFUQG6Aq8ss/Npg0URg4UeY6Dob+RsTW1o57HhIRCqv2wT4Y5PWyNYl+rDSdkDA
muyJbRr7wCDCs+5zhP4UbxmSnzr+ntQqH0PT1lEhnztA3HZJGDpPtikoHfiZGl1V0GB2CzGzxjmp
ihqCkqCTaEZXe06Nx9lm0ROG0HxuOmfiMI5SUlxhsVT95zmrSsoRe38O60PzmPRlqu+8ZtBp1OOL
sAg4yyDbSIxhaxMYOI/Nw7Ya+O+QiTQx/msNZDpjxUbogvDG8dwGYaTOAzt9BK9vVyT6Qfbv+GvU
DDxMIwhoxebuRRRVjtfP1ZiwTPV9PDr2KcukG/Wlz6UV653q3vw/hN8WYmzVWb1XPiXOPOpYkIOD
WkTI8AExzWmtymNe1r3uRjh3MZ+oEiazEVi8xbzVvH0rhlCYd7V3KVglBkjscV5dAEs4cj5mPeUq
YbE6Zx2stXq5HUPdEJccptvAWENSku0Po/zEGzpXuKnhizpmTZ4y5iH3pPdWhzLWVWK165/6WYsP
JAvXN6tZT6flZSaP22/vqxA8mw1c1hxhRbqaE9QTz+94cjin4bC8O7x0kfWmrrfPlbTEg+Z0B4ML
05W5HiyJfInhMvFK36T/6mc3xAVXVNzxutmbGe5Ry2NgqQqbn+y23T7wof4CCUwAyunxfLO8cHYO
NmZR+z14gNMSCBY1XOoL0+FDp++pUVmkTIcRnLW8OTb7X5q9mnJPfkOq6BGQQu/k+j5S6epviOJs
BO/d4Y53HrxgAUDi3jJrZXtGQCz7jD2kvI1cA5nVg2LWsDCK7dIHIgtc3QvIQaD91cImhKLEHq8Z
jAYlj3duAcwWFOMM4n2P3NygmKiaPFAumLG8nVtE/Wxf583Y/DlsXgyFLAAfvgSs+IY5m+49z/7x
P6yFKsv2YS4uTzKIiGFCSkgPEA++wpVl/v8eoGC5uGAoNv6hjHhwixvkDNLyOJWsMPdO6fS+WSuA
bx4EXMR0uKwHeO03pc5x8HroPyAHGDWuY3qnHgsqX4hs6x/ZzI+r1jkvcovK2fRhbTEGX0xUaNAt
mjcEy1FOiIUzezy2Bd1kZZCJpzyZP4iF1Ve9PuUHdB8pxY3ouXwzNQtvnv1zz0/vMoRjtQR7SzVj
DVV4i4sLHMAemvf1VQNFOHT0xWCGCYJqKSQjrwWUEg+sii4R1tA2lBPwX7q6btxaCjfcxO6X/ibX
78F/1gqv283DBwakrjRuEAK6wG9tWMAsjEsd92t/+aZABEAiSDmMaQh65S586oXwDWx60AZBRi0I
/aWnWBa2D7drtVSK9U0BvlrfWA8dnskdRGx33YfyORUozwSbNEaC8flEV14sJjdh6eCkRy/oECix
oBHXGXM5wScIwkYrX86Fbbj33HwfB6JdHAmExcTTWa6k69qljdBOTn3MpyfIkzwJE24/TdLR2mH8
WBV++uOoa2/uAcevz8x3Ijb8IzoD0NYtRDrQPAyJeUqBKJqi6S/fcQ7CG4ZVIrLUv6KBme7gJYwX
PxolMjBLqC5md1sxamdMgl7wPNUk6x0bySuQUunchyhNHIYNrEkeMFDNXKSY+lis+eE+scG5gISl
8GlKBmjNlk+mZ40NjSyko78zYO+A5XGqXw75ReAQeCQ2Yvm1oBmtNDxoHBnLk7WyN3Z4H8VnX7DN
RwQkORcd7z9xwdrQsg/7kIBkdGZMEzO0kf4EYi74rKgjeRqLCxMVqrQsnFu3Nz6I4JNaUBBXUJ5a
K6FIYYW/Qr6JJ8W8Vb9meLQ4EWKR0aeA1ndOSwMeYLgIuKZRemdS7sXFtR8DsrMIzWFbqeTJY+qg
76OmRbPqMvMehON9li+3nDs3LmTsyNolLIhQt4I9NNkxhDO8k95fcZfs4rFN3CuYkeTYpfCn6dKC
rKoXaJv6u73wn7tT3fRAO9BNd7Vv5BJR7CFHBDpCnzDJmxOBG9zZtM5utwGZUg1QO/Db8eZ+fxPI
ywOQB4gSRlJdGPewlbxD3E6AdosBK6WNeHqHMJU6/GJuwYKUUZTtlcv8/KNLYjDtf1AuqRf9/YA6
cGhyFrEniHplz5Npb96qXxNcyRGl40r9Je+Ibg+XsLixCRaeS1FrQpzLQL6RXrUZn0mCojWCedEA
ueIy/dydav2L5nMBlFIaiHz5cTZD55r/Xeft/OfohEQMhnepeCoHaHzZis20toL8zyiWoScYuZFz
hnyrGm8eDthj9oy6JmKyDzV+ifcN0gVcLzMBFwca0tvlM52SSYv45Uw0jRJ67i5Ks0wIBNr6+zGs
ctCunU6g7DKV0qNkokj5ZMxyHn2Y02yxJ7KQIzdFJ+pqzkGvv7R3hFRt1WFuA85WAQ+c/k+wNuNg
jVJUBcE4qYTY0Gj6CyYVA6NMuLfiCW2kA66YUoN5xcev56I2sy1/asz/1pzH7aqK+V176ApI+LPU
Kf1lhbQLB2r4x1uicN79a5UeTEqmEAEp5H4W2uoI8rOsA/09+2P8aNXuFBEN7nO6fvR44Tz3bB6r
6VVscprehxyXKJrY2Jc33kbRSo2bfHR7k3j8+SaqrUoc07dkpmqm6ZRaXt4eYovzxtsOG9vgVFki
7ih2ZSAk+lZm46VmGWXYn+ksoLT5+TYpOk8etkhs8NYs0XUN5Pa68EvAvRYBD+3590qIn0ZinHV+
KAszNoyT92nz2aZNECY0mrlmRsUDR0LXeiXNoHXAXBChRtvm2zcVHXVKWN9bd3fQ+KdPFQFpkc2u
N3k9zgq1s+UB0q6R/fyT9qaXcG7i6H2DatEQj9E6P1sq2f+qx1aVVQchByLEAkt5Rjh41wf0ZAIr
mTw9Yxw/Ed6UI1eDk7+URdOpczldJx122MEWuQxWCxEMHwEIXdopLgT9lGyXtli25MohbHjKYiQP
qY9c33jQroWPVXQfEV+m7kqlGMlT28eLg1VSmGNJdg5piUIXNCFibQwBUT/Cy9hF0xXQSApOmwmR
6RHD5g6dFgQCs5sw291TvfdaHFuTRTADcbJ/xSsPezu5jXNXBljp/wEcGSl8uDHBmPR3m/mZQNOL
hRCdqVVHrZ8HifMHNnJsmQBlZY979ZzGef/9fdW1Q6qHwEyARtwAuBkrb/w5uLMqE1sHdGKd/1K1
2QhDosk2GgLUPBakc7m2ct5hApteTNEGstB1CVVfwz6BsN4VTe3cw4mYpvmnQIJk1EMQhOsYRUnB
tisGTQSqRlyBHGEpUmdBUPh7CvRES3iWuHIsCfF0+JOyHrCUgIOeAUQpyMWSN4HJiwSkz6zsouBG
68Npr9E8LvLGYuIYVtF/7eLEPahNMlEAnoFiqElT41AV9PG7VNwA2FfI/8oYc70OGKaOl9SivKvN
Do30PXsgLftVg88Xiv4POdMhnmqVLp/ZCAsF4f2+R7AmSuXAxnEj8JoYqHYtx3+itJq7z+6z2op3
jImN6Lr/JyWhl/VuJJPDcX3jZuUq7x/d5iChUR2WTFCf3ktTLljDiu4PiJvtwZUd2MquT+DSE9PO
t0oKlHKXPmsaSjMiVIRSuCiZZNE3JWAEGpnxde4SiOjjKBJg4Qt5AShYZHOxEJ6u8bTiYQbrMs0D
Nag89cDnAU1rEE/JwjkbmlwEYgdDYgbvAxY3xjN3nk0Eh3JqU3VqZXwXB1uLxId9z8C8yOkKeDqn
Z1VGjfcRzPtwxGOFzzQkk21TXKVV9oEKo+CQz/qTJ98tnq6+XsAdZzKub21CmCFE1xHTcyUFyIqI
EL8UdaiLPeYnrXWcqT0nSleGRUxvXi1uzKfqmz7sQmLRLP/o4ua3BF+DSHZgE2nkSYNSnvy2WMLP
CaMDQs2pytOZAr61T+5318O84Hmcf/pUNeo3/WlotXEjMtpEStozjOfQjgRxu+y90hAC7Guy3D5W
Ep+eOB7fVQ+2FkKo0xrDW0F3akmpkSrUlIhFbBKXhF21y8o9dUBKcf26a9TNnHdGKZwi9PYjnGXN
RKOMpSoPzyQOQv93UZIPFXzGuN1xiaQCOxRWQckCnNeiXX7QisBKI1mheLwrZukGXfigTnDE5mV0
HeELr9nelQc1SIfvjTMP+AwSi+wtbbMBzeDie4dJaSgw3duYJzWKcefe66xdT74gONzV5SzeuEWe
mglC4qLFIBaGUZxWys4cwtLZUqO/WpQpvEd3kXdC3+Gz2PDWViUVtJWmyQCtKIfq8cNxwWCoidRZ
qrZXN5GY3mGjLzEY+WglF9xHoNuwUiDNzng68jLgj/Ip0t3vF5uc5v3dX/9G+FJWVMtbB4bzXks7
07BH4XyfdoDQNQlkaPI8DHxXR8F6IwdcgDNARDt887p6wfaqhNImAVqd/FE6s4UIi46/xAth4Gu4
vu/Xu6XoEqKV6343PKCm7aunz19pn58lvIo5ItRu0BH66ndi/IYYz/CsHpxVDbuUrobLEI365xM1
7ujnVzbQYeznt4OEV903kwZZ7q7Q3ZC+4xhPTzhP0a3z1/wtFTrggBbl4inINYFjqzgwqLWj9Tmx
QDrh5q+GFp81cRBeSDOyZO3HXIezOnBK7inL95L6wEBMtwFrSgqYLzCJ1udegGSlJze22CGMaaJO
/Q9/8HfYRMvKX4qb4140ZvRldRsN+diGtewq00Sdy8rNIbrh/PVcCnC8a6Uw3HBJjZTiMSxMQj4/
iJ892hG9QuSvmLDTy5u4/lrKXwa/y7kX1l8IBgtC2ksNhDagm85FgpBeuP6wjU3j6cRNRBZpqnwF
nfUjgR95n7yiyPGo0ou7Va0c8oBz8zgEVlB+gPRvEXJcorS76O+w1HOqnAUO8Ji0Px2MZqQK41tq
7+jz6am6u4w5z7GoOABCH9AgfYuBDNzV6CWRS1pKilMpYRXNSziXdk19umFCNXPOEZqOqJTXEqle
Dm9z5nNP70RngH8MHgHoecVjbFpZtCvM7A+Simcmr4Kh+zFpa21/yzal34shhmdoHgS1x55BVdDC
EDtdfhN6DJy19UWLy5CnLqMSFrEmq38hAyJObQk2CuF9XiwHu0anREnxidyVpc7nkVc27uRuAifJ
hL95pAAfvxXXdFnGXwCLqbOA/f+GdOuYUyDKM8M4x50TuhnzwkcPDUskidFQLh2Krx1dVNSDX1C8
yO89rMQtMXJu4AuiQyub1FUiHznQbExjKLv4iB07ISu6xLP5cWPBPe5kAYVPo42eaRrpTtteOzl9
6Pf0B2eGDtiS3ZEAVWQKaI+L/ntDKaPqlP+kJd/bTV4mxUPtUPQ6YLu9hmytMVYn/wgQ206QnBc1
jEviPkVzK+uc9WEvuaOrnY0wcA7o4TJOFLmL6cFk8clDzoAX3eLXqV/RimwAEkyQl1rZCiw1mC2O
C2SxtY3+p3Uun2U8uclUUG5ePSItZJNKapNeiKfv7Ec4Aliv6K/sTVF/nq70a09bDH3r3jbkSRoM
L9jXPCoPZ5NMXsdeV55nZnjV13hgfii6L6WX3qky7W4PZfyzZKv0LCN3FumajB09CBx+/sL+SIME
mZ6IgMfyrHAvNYXXYrAl+OeHPjC0ajdSbPu6zKwih2ry0AfPY29tVxOZNMO0/zy9dpL+lt9GqSVr
ig5QUFZzdz5IASYB+g9BKXERms62SsDkRjPNyDIPUsufUqTbIUe5RU3t5SQd5XwNMsrPX7iLYPbk
us7Fuh+lC7eb/fgLPfT1HJEdXfXFFVybhAXm48huPG557fr/uewJlpKWqMdASyvlRbAqB8v3OZSu
I8VCEDzwYpRCyWk2nS5e4y8KsITuG1ty9ZRZsV4Ho7TDsA/3KUZmKyoYS+iUlfGwu+xD+J+lf6pj
bHamELDpQRBywMe2fYB6d6nZ0UQPod+jB+5pNww6JqQuYyEWL5uEwdL/HLBbjhAwS00zKVjmI3Zp
ORo+8k5LUkV2eaxLlrCmtAmfAGbBkyfYXI3w3I9FGu+M7g65+XdWCcZ+GNgq28qauGftFcvm18qX
NMhiwasgqaBCAdF8SHk4wOvWqjlVrWiGGT/owdspRV7RTjFLN1vpjUs0Sr+aMrWR+vue/TSxKbqv
/MWipOTgXj8xiAH6OFtTh4QYGOyjIZ6Pwc6IXNWopKP6Da3mXRhbl8+oVQNmLt74xpfXvMgxy2wc
TT8c5BvQW2E6iS7lDGGYSVpyXR6EZ88HrRRiz+CfyNiJlZwRKgrOHMxlJO+k93qYpC+1q3/TRBVw
V4tLJUQtGjKxfpcetaL/EA1PoEerkE6L40UsYIDrAGXZOPIEjqfpWM2lRtbwA4jaUZBLWbUqebn4
ZwJxdvt/bO6roIuumFQK6iumyik/Q5lct19ZtHKaAEhXhWRs2G62q/anXYDMHHOZfJsEID7J3GrF
Q/MeAK1l4lqZn6RMrqcHq2aj68bdgL2p8eiSiAgaeyOkEJx6dQhRyFSGkgGu1qiA6YJ7ud6lqtRS
dkhWS/Ffewq8jbVM3HvA84EJ34t/6MZr4zxVCninp6naaCR9Ta8j9PuCxXrunJvaIZ/8fMabP2RS
iOugFTSzNu7kfQPVMa8Ea7mpbAfOPRw0FhaLdIsw74d9u5GrySzS+J/p8RKAoIGef60eI7ASc0Y1
nLdr5okh/AMS6eEbCUSNtmGNWIaDlTBN7gPwNU42zFEPX1h1HB6mGR+zD1JnrRMMbuLBE3thj/Zw
ut+0JD3y3tvI0KsPYnyo8ShncKjQBabZM0kM1F7u5MVQfB/ZwRlUxssJh8yx7tZscywwKyvwxU5+
da4e/SPJ8XevI8K/4yRyDlYKqOfJsyc9SA5Zr+p3d9lYwgqCNQw+ttvF7BuXFaNVJAxfjasMISE6
oEdNIGISGf5pr4sLsdO/7xjn2U4/VYauh40dQjCTsMekon0z4dO75nCGn8EdOPOrXeQ06BgdtwcJ
YU4TIqpcPrMGjyZv3DB+ZAwqzfC6F/p7ARdVVBWiZ/2iWTJIQkk+PfR+azT+LuQBsiEsT2b/cXw2
Sro+WeTi1LsNnSGKDN8o1P2p9ikyowTkJynZdXzHpxJ8LS7tHxKuv+26dA4Ky9HRJeca3gvW0HDz
rsktMTDslkc5OD1Bggc6ydcaOmn3lSBVQinAW1B61bJ/HSdSOjFwSLNpNjQyeusRTHeW3YFAAA1L
31cWUSpOW0rDDs+nmw48miKYGJO45FHYZgTMq6U4ltL7+e4n3eAxZks9L4Ri8yWS0Y6zbO3x1YCV
13S6FipC0UyGXDhBwqNJVPS8O8FRK4R67RBc4szW769OvV+czm1O+3bmEBT/7UekKXJizU89/+QD
anG6GC4GL2UD8PQitrX1kjwHmswdqYIhCj8jRsn+A0zKEtxdJsRH9odvEhNiowSMnPUJmwnSlkH9
iY4Kl6k8K/mZnAvt3frxMuz4a6jKmK12vlssBso+gTL8jrZY0PXGeWCcdoEwuH0Uke6nJUiZSNHY
sHfpY955SiWELgcjBC4wtelu1P8aKoSUyAny71pTKuwbkpHQtiTLOUq4en+HKTZsEKklAAyP2gen
Z8vNoXSZVR71gjskdVF883yY5ShOg+haxwxoioYLBmz34ffxKOejiABq4TuC3/fxm0YnQ201de1l
8Vy3ei5PQPeBlqB2Ctbxut96lgK9LXFV8ZpTGczmUtCuiIvK6JyksFf4vxoPa87eWl6J96IWmGqr
f7Dik48QtiNGjemlLCYE5X7Y7Xi9GJ1KUtbdOJWCvlv082QSyVE/N+UpB6h0dS8lB5FjTBz7wDIe
C2sj2vPaeTIpIFYlumlUzrF88SL8o/+54f0W9lji4BP33aXwpAogiJKrZURMf1guQLNRagEtd5Fu
t4tS7RI804cvGB3APPdjBabfM3iQp8xFleZTVhgk39R1q+N99NOkZzLipYXG2WqZI6KDLXaOe8Jp
UrRy1WnEKDVonmAl6/N13NeoqSCeyuDRXbD2YC4KQaK2R48ukkOg0qJWqBMK9q2DAYNPG5L5bRd2
nBZ72ajt2dyMI6MeAFL2WTBxa0Ssgvi/pHnS0OvEQlKOjJHIJxltLP4Y45Y3LZVaB2ZdZIxuGBhx
MSSA8cHJHcje6lPu+6IH+9WaPdUS4jlB3h98ZYSumgfRVd3v90eseHiV2mosyVALAQflWmeLSo5l
ZHOkM7oUvXndAWaB2YTh1YvepTYmtQ/vZ2Co7NCaUwQ3ohfPExWf19+R9VDleFNg7Mn7Z7+ABdag
gn6v+SxBxCp8g5oA5Gneq3FR5xonZnQyMfQcsQa5q9H+X6Eeyv+ftsIbFYhQ/RhcAC9GrDMxhyoc
moJqfqkZPlkMsEmRroN7MRr37KxY/bf7VsTn3kE1favIEuRDTtKlDrzwshma67C0D7j/+Uw+jXX3
DbI/dIaxFrysU1d7LjC2kmqrBIyYWB2zeHjYnQck5Y8uUlY+DIhh8fuBLk5HyLxJiUx/RVatfnxI
X1ykjUM77b9KrkhvhOuivTU14kTX2DSojvTa91gGIxQP5bOGxuSpRjpxJ4Rm9FzV5vzM8bVi461g
0bIOAFiGt8d6AShTKP/Vrmvr6Ku/aM8bf6ZZiMthNR73dFwL1cTy9j1SQGIJlHU7NpwIrJD1yyvi
yLKt/Sxxk775H/N1tyH9iGqx62Eu653BUX+B96g+TyRo3Dn4/i5lts1gnE8IhBEicAlgh06d8GAh
TJMyJutn6ER8+ZUbtRZWxcuf7RpmcI0mUG/95xQTZOVs/21mVD3mWPVmQvpP/jVmQX9yDTuAvjpA
ru1C0O9tPOsIlhbxPo/75VW5topyIm5taPo58smMSJGxqA77757pArNrwP8KqyJrjwNz5AV2TcBu
bPt2qg5Y87+yGs3Brbh0MuVgJ+tJdTRihUnxlteN27FGb1vht70NnkTs09FXXZgufYSH+SWz+6i+
INwFth43Od7xUxcn7R0z3OvizP2ZP5a5wHkZB8ukU6wDU3bd+PMdlggyRGE9jk21HRfHfQax1jpp
GZgQK82GLDhDVbMaUV1MHOMf4obHozF6ZhbtkSHPuUDVeRx4obbt9CkGe7tja0Jj3rLYIbFaYPrX
zLxYPc/V7A6wa78spkRCmuRplMHtO+dhgGsoiPhVHvlhkpHofUjVqtX6bw8JgCOV+9ItZhFkt0iq
e2KY7b+FOUS+y+vu8bO9n5FlssIFSbHVVqFNb6KcyLdGY47Y/bLmwv99Z4Gehj4u6rjqkPZefww/
bzdKmlrDvzwrJMaM288yShZwzSh6w7hsOIu1XyOdzKNbWAs5B3cD6M2kjTQ7OYEb1EEvXunlEkwp
bf10ctSss1hMi9klb6SVJ0HBhz3+lloaEOlNNvQMOufV3LFu4U+dQrMACx9Vsk0HU877LqKzncBi
9z+8XHsuvYYtb8tQZQzx9dq9WBLjVsiyX4yZk2cO0X+mqsyrC3X5vmaUos5G+dMOazvFOjBSVCfi
bU8fNhwKKQtk5xxIngnqzmCFjWELEKDH3/5EcG6n0N+fJD0xLEbD49rwW+quJOxEPSA3BcOgH2ps
A4iKO1Bo9wRb6IFKg86l8yDKxkFadTv+tdFLWlNL77E7jOWkDZ0vEGG927EN+qqn1ubV/V/rXJi7
rvFoIpI9b+5qNa2O2f1xXgL5Sywk/V20mwbWznavDm7mVGj5LtVIXQIQfnxq1MymvtN7FtURv4jo
wfR2lQRgxeHeKg5qAiGRzZALGCgkWt6//Vvyskf3nt6E63oMWw9JiYqR/kYFJ74d77/8R7CCnoOa
Rd/q7Gxd0Qdbaw0/rO3tVq5yH2zdJVk0nJmh36s8YAzeVSF2TEQZ8niRBQri97mulrSY19yWjmOP
Kl4hEk7qpeaYUtMnka5jsKULknskFJFoTAKgz4wyXZrL8OD9928tT/bdD57/qWBK9jrzv+RDk2LN
fWL1RFwaBiM8C/mVc8Egu4BRu+YktqJxxAYhkxurHNMFR7VkHXyIc2uDfYPLRgJZgij4MKDc0bya
ctNDL3Ra/52TVk7klvERmu3x0RM1Gky0taoeMy5+OP5nvqbgsUFeXpEZt8EPtASXmUu1KQf/lKd4
P5Tx53Xb9vCqQl/C8ytgRZPC5wpURfeo15tcej1qAuR3VrFTRFSuBMH2jTafK69z32QIuy+cjTVw
oYI/75Lc17bIBJooSJh7MGAFX3WfDuj4kR5GHmzvt0YBz0MRAyPiHLWUmJUE2dt2x/AiTcG4STIJ
dyhtJsn/dnYsqJ2+5ysfky5pMdNGenzcuL6T1bL0BI8JfLt31HWbvmBn3T61j64tlqAcoohT6QOU
EG1yePFnsCGPnoxd+v8Eurz1u/loCLHqFwQB4ZFhxnwhjTAdPb4Hn0SIWxR0pM0/l+MwpREHBF/Z
unM+F/c0P9rCev2s64Aj0QTKImdJBo43zawQ6EB19NOdONcUdFV/ki5XovouX/M6qr0ED60+KwUi
14Ej/wu1HkLyuMObYRvH+Ao9YMCvyZW+1FyQtgqbbe6PnvzA+lKlp+Qai4YTz5miRaI8JT0AxC5o
b24tYGzI5w/2chFGe8eMhEzX0JizO0ueXGQc2GWuSn1WqKvTo060Iq8tlu9FIQxnkqTz1UPQXKjH
GIxntokSGSs2dOv/43Ap7vsJBSoGWlPKn0DJxiA8kOv4J7vl9LJsWIXcOP/4Uqgl8A7tc4U31PQ5
7wjskQu7VJhp2RQpYyGo/RSw7UNS64t5B9ec+Q38PQazSuA7TESjE5+T0bxqwCoq9rPzdH9AToh1
sD6M4TUuxQJkk4e3JYZhKwLkdFWv1SOMG5UsQcYOoKxfdIJze5XU6N3WwXgzMGAzfbz5IB4QFfp4
MTDTKzKZFrxGoos2weEmmxsEjaWuodzwsjNJkjxwtM4RNlMt6dY9/izYyTBshNpHeAd6SrzOWQ8n
veuZAj0n6XFzepvEalEpND6TX08Y6fWhK6614v/+Axj/73IJ373gGduu3AHAnwAJQ1vYpTzEtE/V
9mM+TpCqY5QPilxX+20UJ8sxrt1u3WG48TsJO4eUnaCGH5FkNsRFKG/ay7tE49DxKwGAR5tkVQLB
UZ1EYoqmBn1KX7PAaHkmbzGyTq4+WANLQO4HllSFV2r53vzN2e07LhJgKegCIvw8msFWl+tdAlcy
8/jF5PIAvykTKKV/vgC1sj4A5FyXhIaCvsfo7ibIF3A3T/5JOvtmQ2QsMWEHqTjqN6yzLOE1DZsQ
D4HJ6+/tK8+e+vL78DQWvNjxlCQGrxnK2D8/qFf76LfUz5VpDJZvVSVB7E4FofS7/BhKtPedB9qv
q6DnwFHVj0+62QHEQZZa/0v5pv3LthSTKzX6j+RHZ1UxzIxpSPheL5J87NUMvzkrV0hMyFaTtWaH
GRkAD1FsKl+j4ydurBrcSHomIsEKZx0Rca+SHTgJ4vufg5e+39TDXOS+ckHtrYFnGQi2gL0Z0yFa
4sonh5GXgvbqdBOniEHWpXSqgxU6gB99IrTFJCJsg1PI18XQ7iBsznxilyacL2jlOm/wwG/BYtUV
q7NfRjQQTXM8DxXiVWFyEVRcy9utV5qsE61AzDBsal1xfz0xTXMea0STLpFgcwSjYnR/YkSWfaxI
foiJ+H/+esDaYsMQx8E3Gm/4BCjQgnImkjSmLSPijNguwoggDaQdDfwCBdja9CqrlU3BfXuECSxB
f7T3YJExB9VVaxbUWw8nOhhTGcbdmdVhmmsHbaj+y0dwEcnzShzzjXb0CZ2XtRLQBrCg6qzT4R2t
aptdz5OGsJOpBdgVkf9q7XIAgO8OJrZrColCyAdXWaslviMvBL9Genc153dZNewgDtcIotl9qmdK
cataeC7GgMDike1H6QGJTsGg3EgR7bQdXPJVzovNr+OW7Wj8odbbV2oY9aMllWxa7HHTM/Cm1PQw
Sql+94DtBzCajcoLAK4qvI0LOGsPNCPEVyL6OCKhjbwiIXEjiELSKsOxUQnFZVCadIzC4edQnhWD
H7bS5IN3YOo59kRiM1XjYqPqLuJPQkEqq1DkbueSY9jmKHSn8VGtsMnsI/buwrfOaw0kRow7LJ4f
iWsLOKnpF1LntLfXtZyMVj8F0SZd1RyI34926pPs5kqJgds5FZhSfGM7lYLTrTyrpQb++JIVol5v
BdPviTk1XGyMd1/5KMRfnxlYYTFd4yPCYB7btGBenW/HPPn1HhJjD60/Up2CAQIH9xvtUiNu6sUV
xOfh8bEtX99+YnY9QD21ccBC/BdI0nfjkZD4XWv6hU6Jq/Y3MadTW5nT4G9silP9PaEFjW8gEH5r
hfCo8IUQKhEmDvb6yK2aGGTeWkNk9Jm4KVWU+75Jw5bAbOVAvs8ud+67jPWZvhZoERAzk3/2M655
1ixUZD/Q7xtZ8yZukf39dl8TxjDTjKl+Mnaa5vYDJzHTX8LtePxof0MBZo3YPOz+rF67F1mwaipm
XAkU61Udr2yNi+Xw+X9MEE6hKtDiOD7bMEoP7hKvEPozglxAdvFBM28z04G5mcJVciiaNcdYejpT
Z8jngblPCF+t1wn/deCvOMLXBIxnF4Va0aTvF09+5KDmMlanGh7fmQL5DCPf43Zuy9Ik2y+WU04U
aqHGZzGB7KZrWO/swcx+HegpUh3KfWjSuL6Y3DKzv31Q7l6z6YY6rarp72FKyRGJa4xMXIXhcaT0
/zVL4+ZzVrJQChzVPJxIH62TiSmNy9llaq6dQ3xIB/liTaPEAHVH1xXPKAB6DcRlUU1mcMklighd
9CKwkZMbB6by2GK0WCunjUepKggT1RKFIvKiVTBpTJOxDoyiVl5XMWl6xPbs3q6Cs14ZljLX2YwM
f1Rsq3hqdK+lYuZCDI4Nmd/uTjOcJ8mRrcfqhACeko0tkQfxQG3YXH9X4nobVdeJZT8vMIWZBS6T
aDItF++KbQGEtdgLjkVPtYjTS3yeEVew2cVE+eYqKsKhIJXjQDX3G7HBC38/6cYdOyoxSAjVBU99
Byh1dBYmv9IllFMpeE1ixfCY0Rkm7p+wdBpFiRxdZzPzcR+pK9lfIWlRWv3GNByb1YkEwcy61vEP
ATIdjPqQiyPz4/iwen+EFoqPUWN/pZnH6OfVv1v/Bhx688w1OOldDHipk0zJ3E4RzhDH6PLm7nm7
vAeYKu2U8OHj8jZiYVWY0WBuaN9HseKqXtscqAvYvgtC/3IdSIc0/IHRzt4TfDQVw8qxwt1XMS7y
HMjl4b+KpCVewQQWAr5FINGSTnrzZl9raevQv5280ObDAjlnkb/DBUE21RnXBNlpYiwHwRlPv7Sq
guZ+dUc+rNHcaxZu3VW7LWsKWhmAuVb4j4fKBQhVn2i43aq1aiughFTrzrU7HDOqzvsxCfGEwdKV
5afaoUjM6TLdnNUkvPCAzEjl6CXb+k89c+zENARQIX8EgILYtPrgNiotVaOoDFZ+0fvCoHT3inft
zyk6npVhH5BHSwwXLxEeN6nwT3z+HVg6HmHgqRHjuZMV6Joxf3MLcI8+ikPhd6fL2ZRJHoEqhNmC
9JCG9HQqnvrf2KrT5VeinOy5vdKZXLcbfstUIXQY9nsKd+FFPWNBZsK76NvL9msHgYS1+v7cFTC0
vY0rkHlcQXYK507yIR5tsfJUBfQW5hbajFJ+8UUqL7VXBSVoEdCNrdH44nEVobun8BVlfbmXn3Ms
te5kPjRPN58Ud9ZjhoYeTdhUv+C8u0sabj3xzOrmOE7HNuuJmSYcX4uxeKDoojwzcDR3YIf0TFQV
SFyV3ssXBWAHHOUQVbx7BUJzOt67MJ+Ba1mE1BqOPkEYhihZPPgrPqTmdnRca5rdsjjVAgFGBOW1
oQ958EW5b/UgltRjxymPC2yvuM5Z+tDoX3a/nhgS77HLwBB1wOMWkSzBYxlG1Q475EoOQy9bvpa8
/yG70UHzp5FKoDrgLzBWMks8FuUwA4gtxzAjW3Gg3QBBUbrYVz1HsvH7oVXOJcr4y9D6TzttMh9f
TXpNFG5KBw+PtFJqEyCE8z5o0UPM2D8EoodjgU1J4pLuAWJMDEwfnn8VFoiI0XNaNyNCfMHWrLgK
Dx3tfnWAN+rFz1hKzKpUyR8HpdAsVU5g7e5aYH3P44wbvMSZ2YwTxonnSLPQLn+a7lAdSR56wAkR
Ht36x09EF6CCX4Vip2r3MbEr9/rMlKFUcLb/kPGK76E3QXysSj5UBDuaHB/Tabr9oK/0hXDyZ9YX
QbMXYI94Mk0qmOysni5xgb0eUl/Pc6EAkJq4PCFxXrOBHRQQUviCqqyjf5KP3M2fIxIoqg00aHe6
0PaDmdsOsJJJTKXgpwn7GagjrULCmbqGmWsMX3Ywlfwy4p4TC7A5GWRfizjzl0Pf46Ec01+wHKSO
RDL+IsJcEUDktpWKxAXSH9LLifLahg5ZxfRJUutAz0FA9YKmLh6tkjee51uTyA8f9+uZjg1l+lzs
t80vmdROEDfKc+iPBN6ziVIkUvr0XeQEJQw17BBkl/G/WAp+G0YRQP9FuVrx+z+dkmgSATdsuNOy
hG+lH7yceOixlikcHPGyGetFfT1nDZ0UkNqeA5cih9oRtVgXtfYsHhqRcpeiK0+LRph4ByIxV3hp
lfO/qO9cA9kes46am8Wicyb2dQ30sckyHxzL+IJAk5rmOd09K9Q+yRqXVJPG6jMk2K/XhgJpDAPd
bfb0/uIOUwdMAl3HxIqNX/Udn6TBo8PcCaRm66yMplrLtUGeY0/LYXzy2q+PMnvfKYuQq7HFip31
irMgoHO3+te85F4jiW4jYkf0xbVsbsiTxzUG4/QWND5D2IOBrGWr6BjrrilSpzxiRrIqDVEWgSP5
wrNuENM/qD3OYZ+DQU+5fVhd9jZFrfuYyGOx/cWIiB8F/BoFuPefcjZLw3mtA2jH5umx9nAT4Zdn
S8Ynd2JkrJO7cwwJsScCsMWRrVgdYRP9IQuLIGAl7BrxxjTk2xEvA3CtiVXS7KrOSajzcW7N3lbB
+YOUoFYPfodisvVD8giSrBm+Db1u/hq9Xf6JjidUBQUMZbuQZBGxJp8p7SudA+EiMPUrBTFggN7W
4E0lcn4UiX+p71aWM8wq1bviBhAUU222Q4gGDGP1W9K8hD9W/vb27BL/KgoBsuxn9PL0wV85yveT
2J3VkYrkRleH0fVhZpzRuprLQq+AsE/Vc3RSndoZ0Lajhv4yO+ZqFWvN6AI0HG/I+6YT0HcLFH0A
RkyJjBcmYlJfi7UgQpEdlMYegcn+gwbnS38sYBGbxS1SGRuJksaK6FX+L8b4C2Qe3deNLhK58ZVn
xS5+F2E73oERbt/bdsOdTxCRK0IlX66Dd3e3VgHTm0+xGV2pkiXJ6F3raEl/Gpc2Da1OXgHjbSae
+rOaQDdAWC5JZkWhEfseSdrs1afv8TCDzLQF6lFw545r2fqN6XPO1V+Wja2QRuEqiDdyd/IemC6d
Fx0jESLjse6wFy/Aew0u+40myJRBpHGu1lp0/04D/T89lqRTDFmlAV2g+U+LIxTZX9oyr3EjMKKA
O36MwlTzwMk9kxOS01O8unUgtwLnoJBlW22uIWgahlxDVN2LUsmxsgK01zfMssG6AJE4XEkjLGzO
nuynJixm+0Z/1zey7Fa2s5U9uDKAa7Fw7T1H14zfgjE/t+oEDg1gDc291zwsiFQPG5jnMRhWgYKW
JFTPfIW3Fxwfxrab8Q0OqTRQUIe2Wl4WRgV68HnYzqDnq30UCC73oGA5gCn0A/qCTOeb8iD+Cbbt
tHkt+ej6HcmZlYHLyztI6rrbkJTXdxSaBVWXWbPADZjjx26bZ/4faEg71jEWPjyocwcXI9dT8U1x
VpKWUWwdl3zqYZVQT2BKGjTC2gWPwIuiCGpVmKe1G+KN23ID1JLRteCuioWsI0aZfgLRgu0H/KbD
INYbpgCrCBE1Hsar66ApSdHmcQmWhqPO3B5Xh2lXE2P2Xxd49WzqTuSv7fjs0wguLsMJM/veSfD4
R4sQATWFInLLDwcx/bkKe9lpHPc9TENuYl5YCvrUXuuV1/FoJqD6x3m48fHulGnOZ3l3q6QbVzzi
WWSgiFfpikWi6wzPo71iKXD8FuJ+jFur0CP/yvsOKpIC7pAa38lS15oYvphBb87sugSPhgbyaFEt
KB1HV/S4r5tdV6QYm0abSwF6rW7/llH8t2gOZR8ROZFl9E+6FisgiAVrOY4T6U8kisvEf9klQ9oS
/PvEq4gKVWD4p/mysTG5NjtTSaAF/9Z5GlXZnN84lD2PmHZ7cIiP9U49vxUOzLrMDNl1r2M7fA9x
iKYwZYCocoox4myVZC9RFMWddvt4ePhdeP+rOW8wDJhfnpqdWgAvGBUKPrm8Mbx9Vvr5KrKrzRb0
GiADMxGEDEuVslvtsydSQU0Tc4ksVO8PLE9zD0GlC3A2pYPGpgPicSDzhTbML8UAM96QYsc1WVmf
M5SslwLLIH05cFhPUxi81n9MxCqR6JrVCVbzhTU1Pb8vlrForZFVbJo3shSbkJQq5twCKlqNk7sS
qV3JIHHw1h47LP3uvV6MNxDvs4JLaIE1Lz3GMmWB/93flHVhmaLn99MEC/EkCkRO/yUTLLdAQaBV
aYt8BsmRGNY6yX/S0KoOScy3tKA0DJm1tS0vg+FryTWRlzBRdWxlKOQlQhKPZb7g/5VWA1AqS2fC
VMAWDEUQyUVxiWLiFIG6KBTKrXL0+hQU2lwPwR5l1BjmXTKUYRHIccCK1FGWKCrk8rMsMP+ljft/
eobIk4zGWzNV5b1YzXxSHEDJD4zYgpGuVPGUrYvW2uT21bTo/RD3GGHz3DGwTXUwdsJr1+/efbFf
1aETrgSc1jJ5wjfkr2p3XHcrwxK7GvsP/oxMF65+jqGXsPP+peBhIaGzIrGeJF49y5RM9YCaI+xR
GCmObnvfS8NOgdOKLXHJrWeeO1Af+RiDZo21qZbzypjf3LneeRMTpqzu5BQ/D5bKRs4PdXHEKvlz
q73ktHJtdgb99Cr4WV5TJfRN3Vuuh0zyMGP9mst+FB/UtoeN4AKa+41dquS2AAsE5d9dV0Je1+9f
aw+yG3wU/QlnIxhKhvQsJXhUQ6AUE7C+h4QmAvSBTHOSSlU39Vc/clPg7HHu8nLgi9wnAz4r1K/I
RVF7WhNlACav/g9OcF60nEtoKo+qsZAQG6z1IGZ7iPOfW4RR4QrtVR9BY5NoKBJoYXFVxJNeTog/
v11hG9Z1zjgz2NCOVKutid81Rm7mYIuGPPdvTh4AhD0CuufP7vDp/q8132mLKHDMrrUEnXba9erM
c1c+5OQd0bFTh+NWdVTW85X5L3KbfX0mVtsz6wWFVBVfyPK12NGAMJ+dvFhafixhpyIFrBnPwCSX
QBI8exVs6aLvWW2WkN90Lqgr9v8ZfzaBIifHzFYglqmMFpNTn1L7Ml45Ts80W29S17jI2PceZG1k
x57AIoTk6nF+bgjQIkrri0pBD82eo0lAmhn5wahffhS84c7YCgNjyIgq49qbdgZRj3R1ikF8wZvX
PE1Grg9WrB+HA/yDBQ+QV6j6P41isEB5OkXG07b9fcGivcqVFjh728vNX1D8h3z3ioENKubDibsT
m0qLlNjF7Awlmd72LIySGKIgGtfQiV4WB4gIr+qC/cuKqF98Wrq+rPy0T7HWYIwF+vdaa+G0szgx
hMAsw6wxSsrapgH8b4+BnaNHyd6cyCPO9ETgtKv2Zt4nLgL9+5NJiNoTNuUlClRifhbM+GLqUU8m
+Lp3ADBE2fCj1Y/oP8l2+0y2bswcpUdWNOdTedBTsZuGTs4q25tomULebZz3bWArT9O8mBezS0Oh
krRoUQAyBS1LmqvdPXJmZyRlUcP3DHoQ9JANwH3Ne1f0HyFGWZ1wOHcg/eNl9olxUPEpfR+fW3vw
6BGqCSvIRYi4LbghVM8uOkjCvvgz35sC1oZVd6OulV8h3ZXCWjwzcUeKC7gWTYC9l1wW4ZVE7WwM
jhS0HGLnoosz9BDQBWmCIWrFlJLycpsRtC5OND/1y3/ZXIqNWgTqn8oHsrxn4j7ERTITH1A1ff/O
TnxQa8NuH349d4jybq5iCmBnxIYH+LY1s+rWqvEum+W2PxoeljFWxdwAdJSp4OeAW6PizNlae4WP
6U2pNL/RJCPCiPCGPmQ8oPcYAA/wqC9WsfxronesWg8RJ1JmCPHuInjSi6njU1BYR8a4ug4uSK4T
4aOg+M8tl2PbRygkV35qHHMgNZ3fPHezbD8Z1dN3z/mwhDl4SxEzfUGu3m4FOV6Vn2ezRmw/OiCs
U68NpocwKfZ7x1WFLxHM23nX835nhUD9nB7c6DRlV6lSo6/UibN7kzm7pFYrwi+A4hKWhtpDfvCY
7mwNMiFhlA0wcyjGclawdJrTcj30P4lWI6tHUGUlar/GnISL4FtVohcTuLqk/hJPcsCcK+gtCiV9
ExT0qHDbaL1SOHT7CvbT+B+r0rkx4fcKDZHZkSAes9PP94t8I30NX1lkVIsNPw0SGn+czbfzxdZv
OlbokE9nt43dedkOtlF85oPGsOgLvT/2Eq8B8U+KlQ3i6yaZiM0OwXmOJGTg5BuszGNwyB3gNVEQ
niMRr6TkkPeXeEhd71A8odqB9gmrBEpENaPKLb6Vsa3UMqNv2W3VsGvJ4uPDZ1Q945y8/FEHFNYo
5SljFn+NpoPbtMDzNzSvRSuD5LzCtprtzkcVFUxXG74mOtO91IStwcyidi7RpYtzNEcjPktLHeLO
mbx7XafSg7L9c4eVMuol5zLrPsGVktGDfa3pg15mLBJxVdoJKvq1h8+AgAPDax7KzduAejYk+hRF
PFTh71ulHdQlSjXRsx/KjCsnZZEThF5o6GAkYCOnPa1LHRAVCf/UFUZBklSfcUEW01vkUq15kJa3
gglt+3uJax6PkGN7Q9UeyYGxVt90mR/rLyOXUt+AivHBqLeynJi33LTPeIt+qt9699f+cWdhTpM0
BmH5Wwxi7FIXnezXDAGsKHZ6hPlVO30IwxxayDg8kHsBDpMM3B30OlZ9HZ1XQWRn3ZJuTVRoOI92
EgVNL9N7eZieBvFZu44EeBSr9NdjcDj7uBV8N5bIbzYTDy/gH3vbenmzhYcd9qM2Uhk+M27TafD5
ZuZP0V9iTiR3LZIFn/ZQSnH1xK8eVZcqN+fLcxybEFgFQGhIXjSM+nk2HjUO0b4FUbchIvZcGOm6
5XL0L06CSUcEDzaBtvz61ZSmYXNglswSvH4Xt8uw9Q5o+3+llIh59GZQaMvQNjgUpFGHUz+nbVDQ
AmRRGTbUBSGqChvJeWJBpqVTgpA41kbw26cF+rqU76ogwCWtIZR0HWqx4Lqs0+btcKZDYPQm3Gy2
nsMNuNAvR8BUmWwHHVrz4kZbkkS8Gh4LDopaUtkVb0FRdyfh2dA3LZf8pxS6EKZ35MJ6p5TfzPp9
w4e5jfvCcOUnUiRY9sdTahJV5WF1eXAikhl8qQTy80ICDqJ7jrFEBV8sYistwnIksezj/kOOX6o9
1VUiweCoxKpV9tb4bjS/7b3Wd/1Y/qPIiu27UxZJz3WbVp6bIHSBUEC1wuTL32/jCxw8bRPHRlpU
3AcVE7Ko3pT+c/+ySWeW0QYRwCYH8vsG6AEWYRwtB5Fj6+/cWIpSsGb5aw7F7rD31GyetqXUfZjw
OawDC1ashnTkoOJzT3KgJfx6rwIzaaiNuZVYrx+gfRTkENbITPDKUC4npQi4eQpX5Yj2pKPr5hTm
sNtvfSvrPgccLXbotG/t1ugBARAbFBeYFzswsqmBwrgknYeUTvxPdar0cH1QEN61c/l4HceS8mar
DYme1v90n4fpelPg/eP3SuhiVghMxamUNI64DyTbYJU+Yx9q6BY795gLJuFa87xp/zCDrDFIfWzE
Y3vlHlt3P7BiS3hrxS9sCrnZMkJQ6dzbNRQ7qt2pR8V/2Zx7tQd1Rj55iAMiBCSCAoQ+i+ADo1fW
tN+kMkVc/LQaNDYJRY5rI3FSp/4DFV0F6tpmy97E/kG4XFKTjW0+2x+C7RG+yg/t9/XlkYz/njXw
9xxd4xn/PfuLUb6audn/GES5WXnuAsbDSkdcg/WJjxBIW4O6WRlUt4fNlNu7A6zs8Fw6sQ7Go3iC
dQD8SbIEkTGqdr4JJaZZgQuKeBXeWO2jn8eoHsPfzk2o01zE05tQOgl03XJ2zaRnn6hk/ufZpjKp
+eJoZGLmRkdPBex+cjbGglD1gMbZvBLTe/gCCfOfOh7OfMfzMxR38Mp9ag7lmdlzYa2bPTD83R56
a9eENA+nmLPn9TOhQwn+NILEXK7cmfQ74+25lBDZL9PiQcyzLo3SNGRsjWjEr/hbcg8fCs9cC7l0
HK9ZwMDricDGiu2BItQW14y/iTxLqvAUZNbCYeL+TJc9L9z4pbjiewxjI+GzvCGpWnbANCoE+yo5
0Z9eOJao8FTz2vzt+B65YlLpVMe0OyQ2i/S/h670rI+YobaFpdTtkr5anzpHAFmn4O9HkY0YRY0o
VWM9LbLYgz7hanvj0RD7XNydY2E7JrCGZnNHZUmGumplMSa4ywgnO3eKl6VFdovAEH8aS0A5dq97
GGF9xmohISrsh+vvofkJp6JpdBAtgI9o93Nj6VHcR5PR3wAZA4MgAv25rSyuTxr0XKHMhw7lhEaT
9idsvzp31rx7+FXdSDaLq9aC3xffrUFTak5uhpwVKg68Bz4G/L6kCUq+Rbtp29q8NWsVo+0h4NVl
gweWfq2I1wQROdRdVPNWBLRFmRQmnbOegyRSDdMJ4Ytltv0S4C3z+jqzUDVYKXZKeUNYrEFy1eeI
Ye3L4abQrl2ZtUY9nPQnE6vKFdwgCKx8FtYxcQSg2HGpVZX6sVM0vMnM+kUh0sji9MNkxGTJfO+6
OnD58jri7zu7jfwaAZtxRoTaqCnPJ1FiEtLbQ+Rf8M6HBf3Yl9p4U3No3kHo6N0nqeFsXM8x5X6w
Q0yh7tdKDw2F32SG/zBZ4eFxxzRjLoMCb4Y7YLFAMsdj56Ao/MGUvyQDHB3TkR7khmnvwI9VdGLH
shDqHSVuzDOs3/rCfvDEnxA3yzmF2G/pzfcoqVz4n5S8cnlki4jkQX1o5IWxmARf7I4yyBHbuPxe
hIITLC+PduDk10uFI4idqM4dWK/zNyF89pBahqw00UBeNjhG40C17VL2HfZLJUq7KBXMiU9qWJ0m
kVJTpSVSCIeN/unzXzXfH8M+HM0mcs6QCwUE3tPyi/rT4GURB+uKo60wzbJjdsCCC/0LCdjK8OIx
pyOCNqsbThhqv2Z451VZxETGi0Jhx90LBuxqJ4JMLy1SkjCvs1TCHr9yqGRwC5opm/23cXKC+WmL
7Z/yDX4bwTXOWR55G+luSUSA6IvVfD/X6GWIPlbfF3p5yXDwi039uSU4eDk8gofew3gG5RwYEN8M
BclklzYP006PO1jC7lIZHMOoNr2VhyTmPeG05wm4ABfC4AWlODutbrvU/GVHa8cJwQ+E+uA14rAI
5QYOa5NoZyCnhQZRNYdaKUYIlAjoBnj/FUyKbhQLoaSoUBBwZ4MBuhqwhFZh44iXmX+7FZP7JvBJ
OG7XXE47PgBFbaODjmx1wDnZcdwVHGMliKsAkWv3921DPKLS9ljeHYJNWQpG86XsMc/ZJtqADCVQ
HwMM9ZIBSxTz5RAJLBFbJcWo2yJX17hFlqBflRhOV5Wu7xOVIxhH73tG7geXFzN3a0lbF185Rwwa
U/fd/4LQZscu0cf+jK9YmG+wbGJCA5OWR8BUQhlspf1eDDnarTnbn3pRjaq2jyl0bCy6/hpLVqyD
ZdtCWFjd+vt/yF4qjryOJpKw1mYKethdV+CHHFhm4bL2siuUJZI+cCvKyqgsZJepmcYy7NsuPhuC
k3Emb6vX3Xrt/5jNKDfWV4kfdxIH4LfZ/iGVDhfCCv1a1oRHAtg5oqTIZi5wBtnO1oZsYmzEcFvM
LnF9Lcxx2tlxRZirKbMBGlB1dB+JdzKApbj7ByYRlIynXVgi4MYR9coCAE0dkg/oHlg7pO0gtftA
Od9lhOzQOgBRcZY76X5h3fbecfJ4K8tqufIL+tMbXC2RTcRg840zAoZhBYXp1euDm7cMFxdqlHKb
sor4XEZPrTIBB9bOoloyfsReWXgW2EjY2NU4ex0JX7bx1Dl0PGLh2m/SJTtmsWGXQV4lAoQYIYO2
mWUA06rHo3KMzxkfobU+m3MRrQhMF9UdvT0YuaSkiuUJ7mXN20wWQlOiZGQZ9rsycmoQyrTwKZp9
13iaT8TzuzCST7iAD/8Q/RBVSvc/FqdNaXMEoWuX2TTDofdGkdP8Qi94b3A5mLHZSP6v2PzFfeL8
QdHqpeMpnk13DxsacQWuaNAqiAFCp5btQBWzw40lUWcPkoS6HqyzYAu/sGdBjRvk3ld7iwMuU72w
NpjrNWizgIMiD/u0kP/QAJaUEdqOtdIvMckKWOPzUSu1smV03XZWWF2gBBqLmZAkPsFUYmcxYyR/
bBeT72A1jI79idr3MmZhcmuylV7Fos76pAOofnVPAzcKRHwYZzODbPatBvFJPexc9VfFTLftU1HR
KITJ4kZjh52ZpjtUEU7vi2QB6K6rXLzONhZQ4+9HAJKxY9eRJgo51LSoWgN3lgbmBvWvSKXjKwaq
avl4bgpyEOBbEkHU3BUT/RA57oZIvStpdYTMSMHBzAo6m7GD5kNCvGM5aCRfHKQx9HNQ+xbvftkm
uhmvS2KxmenEyRvewrUmp9I7Lq9RubNXay7QTcQZlSNYXmd5/ddGuCGNh/l8EAahpGCJ2iW28nRE
il0MiezGm8R9gj/ChcLu9jVxbsiVwvruGH8Fe7dYAJEn2JSkefQgXRr02rZaXBvLn+ObXtI0sm2b
8gc8FV4qungN07fFYdtAdjyZHRds9AqgfdQ7UefNsRC2NE+58dvAxdjqmZl9k160qQSIdhf8p305
GNJxwKWDGH/xRzAUk8s6aQrQPiYFeQ4tcMK8WVa0OvPmW74sreRlVrqD2kpj3UqcarSUUli6rlth
lql5eqkBdLHjapm4z9tO4KGoBIrsjlMe1WHX7bPCwNKWTk2Al0n6L6nSfC6hKVXHolMAD9ajjhIi
/gQmLlTG7K0WLt/a2D/wMqKgEbiuRR8ZZ/cVpFf0nqxpEVhAsS4r6tncP7Ev1w2ySC++5JovEqRX
rRNXc9Ui13L1TQtdhQPL7Z5btUi8BC+ale0lvOKYyLYNd7dpXN+w0NP0O/IqGcpoqPrfVguQxrl1
wE7o7Uz94lHQGj9YWCLcsYDldQYXLiIDmnuwxVi8KjB/nOdbdi1FP797irG2HuXGQRonUoM36k1o
ikS89/m2F93HWx8VQwOJp6wHUg1Hhcx23xHNJMcHt1MT5FUbuAmTwh6qvIbYV6BSfuFu9qrjGOmX
1eTUsNf2Zi7o3h6fBf2wJlnvRGu5FE34kBt23Hft1K/skUOxtfKgpUnj2WcYVrkPXGYPma+2ltAh
Mcy8zHduAlu9nYF+K6zVC13p1X2Xv0D4yrfS0kYXgohpx3X/QvwoKG641lz5IDVsNqiVfF5/K+RM
cC76OYUh2jMZO85NSXnNIb9ANYb+/XDJeEa4oGzsaOaushM6dpY6XZEHVTO+QV0nc7KNELv2fuvA
8jv08KJLD34mFEmwH1fZkOD9cJyi0sQtt7q3CHhZgTQ7lEwUJewHhhmIAd7WWwcZ+5sUCg9Tu/Yh
1HWyXGGZuDP90pRl1dCk86z6Fls2SWNGZTzOBv7Sp6uYpIDhBSzfK5oJ2m7c1xx0F2GJqfs9A/L4
EwErC1X75BNhDJPrluEYkYw4GLpUWZI5OY3DmXvrAdbc3JdL1joqt4Quyhat1iEVayVJ+oHRuVko
Hnq8Pi8mw/DsKGbPi0MsFiVY4XPzH5XBeB3MiXPDmdRBWRitzCTpZjbDuvEj3yyhcrZnlhUATgzB
DS8x5gX+3d9R9zU+fBSSwX2CGtE7gDpFcqgCIIw1GkfxhRrpG8wemSKsFYXWUfFB5b1OAu+cQjL/
RZ265cjHavGTxFA2r8th70qbwfzXG1AoJIcBRU07YJaqqduv8BYhATVSCJxZdBDhD0uX0J3FKDHn
4l+xSOfFxjiqRVmpgNAdSLA6IpIRn8PWaX0a2Q1pwFwy+446n3Rtt7aXAb5+QFeXE6SazgOtYhqj
enytpFozx/CWnbfIaAc2dBsRKA1wR5Hz//oQcnBuDMawHWBwa5CUdLqqytsk+7wZcxDN1gCkOR1A
pfzxvaMPSxxg+I0ecUWsBoHlKaevx+U68hepvKLg+agK3CC/i7P/+Vq6nTHC3TT3hOdn89Mr4FAg
EO4U/WdEVAdRqB9SA71nn/LrcDjDB8S0T+KWp5zmgKpAi+2TWN1krUxg1qOqVweXsBy6z+eTDFpp
Gvubvo5oce9nSTtJf84w+u5mBdNHOM4MRvOEmV4xESH9lHNtJDIDLbiXOR9u92nc7PszEK3gl2Js
K2fg7d9kbgw1eULYD/8BcuulzegpaOIG0bA1mRVrYta6EXV4lMpV5ZOjUEv5+X0w+DNetE6vAFB+
UP0VijT+mAdvxdIHzBvku7tKlc9n4lM8r2mrToPCdwJCPu8wpwVZJbmtPZBB9dJ3VdsCM4B3TYD/
Mxh0kFk+ro8uJMUs5351LBQfm5rVVmAjHkzVjXHICVHuVg84TIzAAAdEibbKUhhaY5EQ8Dh90QvS
VymXShN2LHNFpf7f4VSvzY/wc/i8wOjWEEvE3bcjHApfvl9a7cM2HYiGPFNnKZ695TzrVoKLR9Zv
c6psbrOPPrkC02AnobdDVA0PVIOkg6tDufmoCtE/AgPzWxmmgWCDsHCtFWJ2U52goeJaNF/xmvSc
GodX971gjBfqtf4zX7ZVpAWRk6rotWd2i166ouRHfszPftfRR+gpYB+/SjxTGuaIykjq0CFuhlVV
DZeggiBGdgJ4+2i7IeLCGoaXw6VD2c5WMo6tL9Tk6T9OFXeqmZk/FgyFkLZYVhH1tTl3o0c6fzYt
6nyYERKOKfGDL8e19nZvxIp+PIsNBuHrVAvGdmLUBNTcjmDJoymMHiXdjw3X1MgoICtJ+wUeATiu
OlwsYC+C7/C6VLJeYFA31eNmEIR7siwVw1ct+CWOvtbdIa5dWiuVy9mZS91UvFbkylGv1O5o7jcw
3PqBfqcr8LC/Eh5594OB1TweZSzlol5cAStIsYyVW0N3iUQM2WdTaOZOQDzQCQz2dpnL+VglgQKw
9U9X5WNCPQaxbhtc92Bg5i+u6zHb7C1PpSCUc0K01IWP/5WlF3czjTJdQjb96hF2hsik+ubA2eBC
e0VAV0sxDSsqVWLvzBPePzwEsclS6WMv2m8A9LpI1rUUxRUkxECGkaaauYEmNVkOesnZjG24lNbM
31Kto6R7MsiqwtRyYEpHK2E/mUzwcoHTx56E8AeW/V5TBGsRDLOXhstaTRWyNDzfltsM5sy8FIwO
DZ/7Kuo6YzkQVAtB+3ACpU836jUQQ5bC8qZL1gvxRjiT64BBEZM/c0nf/NZg9pgv2os8sfc/1amo
1sU6wwyHXIZokthD0shYb5rCLZYbNM8lIZsmCYOr//bsjJNi4dekNx+vlwJlc225Q878yqkEDNYF
DF6WJj+9cOYk++tlcyUXveQOr3qq4jZoIkK5QnTI+Va6OyLXO/pcKEkgJMY7tPpfMdJkgA/mqkCG
qKHPtkGIIPQZJFQG/WF0XDNRBsZ5SJJaD8UK8wM2gSnxyAwzY+gSig8I3Ya92CvpdZSeBEP3m4wA
mveheYRH09DZqHEBqoYBppHIQ3eVIReWMTjP5o7xKEOXm/mNvlPPE9Rp1s1vTJpQZ8BgC5TuVc+x
bgmwLnIHKeUGlD/qxSdAvFdgE/+5jzpg6JlJHferhI2MlGFr+cAtFx3HdZR+zqOVFH781mqSqjCg
yBzni7X9hVIQVVZpIeheoHQAC8DJcOF5sKHCsjvglCZfH+NAkxPAXmujrdHnVZXuTS1femUqNw8q
H1DgCvryi49MOr/rIardgUrVtqDsaRmd+Jbvrv24F+V3SKPiJabxb9e9fNMKAskPEAI47TOMAYaK
C3gNXy6kKYOBWYlUR9/Xilkg9+0QNL2xceiCzpeNp8We9sOvrK8lrCtyxs8iEFnHd0Kxya5y0lvO
a4uKB/huq4QA2KXLO6PuexdxdRiivl9uHRq0LWlRFX57cnYIruVIaotJmisXglTSR122hVJEEUYD
phs7P+ljclL89sqLzdlXVSPu1Q97cv04zbGHX/kDh17b6HqgTyEeCx7V3b1Rn2GrDBTjAXm93/sr
mcDKFYC5zfk4y7tO4/gtMI4L/8FZ/MQOtdqzMyMO3pvNOKW2msc2j13EJJMBCkQM12ebHZxXDQ/X
2XEuSW1Oq72Bm2AGsJ5IuGpAEhYv4GTMg1exCeDXRRS1f5G41jzm7dSXinqTdS/sB2wrGFGgIVYu
cz2lFz/hpjzclqk8CIkTUhxU0fUtvfYvA5Nssx9ff3CYWtr9po6xx6wgwA3t7hoXL/TKZi9WqbRq
VEFr2V3+orGNQDKDxOg5ZfnHT477hmWNjkgjnsXVUKzN/w+WGjUjUuLnZqUubWGss5Gj6y9NJtwA
4xgKKHlOButwWSwKWuwsth8kdRQb2BifzL3lxEbAFBWiu6Lvn1OolECijntinx12udUB9q0DaBTG
EVp6uFGZZR5r0K5dztGoaviJhwB2NGUt95RKugs590MyaT+WjLmKNtzJvvPfepfh1+LARK8+SRZb
FLnjhtWfs7MgdDS2Rlso4epMwhMNaduY8agwWmzKGntDOG13MZ5iasUSTqxmryP9OO1Csc6tYZi4
Jfxh+uCUak3uvkUPFWsg2KmZwfVCPYHAijGfj7/S+e8nlQssDYm3XVdLzslZC3GbT+u8FDIKWOrd
BeYapLTBcs0szxgbGvgLTqlh1TDmS8kj2nbI5MEmoLus5uJHYqX+9vwCIDGrxJzjR//AZlpP/XNU
8wAY8aMt19wjuai4ypHFxVZ2wLZjhsd/Ax+XxXKwUNcSKAfxXzS8b2Q00UQN3PjVHvLH6AIQY5P3
NFZKO83NNUYB5n3ZLlAchEGpg/z25ee6h3y2MwEnhhxNWwi3KP987Q/LCvxEKIKI6Zf6glf02Bbb
yFNb7Pq7Ns0qxF1Atw7fXXdqxrWuoGMCd51h7FFyP9TwJODN3TUeoDNFBGkVbw9lSHPbElJrFIc6
DF8bU5JKJySXTGbROiInX/TTQ12O02Nhh3V9OqqrdCv4j0g9LFMbl4kGGpkkUAEda0Ds9rzx2iNi
m8Ilp+toFY45ozPpaBQRadBuDW4Mq7c3GEuZY12NJAFlX0SrYtAexOXa8sCPvQ0sfaBhTA1sscHx
qPVFuV/pozUHnqlrITz1ybK/Szlhz3PNhJOoKi2/Tmaq3QAlkbUpffmVz8rXsg+d0AENtFUPqHhS
6ncXz9C5FIGjMZqj+lrTxS04n5MIoTsDKdGqX6gBZASP7b0Skvzzb9Uc10P/benk64LysYDgsA7G
vo7unsi5RuxH+HHPh5vk8B2Kh5Xf4FLuh2RS64JgGfHBtWBcmQXlPAdQXcYYZeZzaG78WrkN78yP
Z0DAx3GMNAoVQX08AY5lesTeWPXl0d99Kb1XPP9xwgVby4SSNbuHkouA9HR8MCNCti4lBxbPOUAA
eg/f88aKra+Tk3U241zi5w0EPjR3WgUxz+2ltgo5VlNXLT9GGZ9nuF6fSlUadY4lKegQeIduxZYv
Hoi8riuIQe5nZW4rlUfAwwzVadC07pzbJeYirbUBgsZkYr8Ah5kovRJm+HJFvfOq5ehGXW3g766D
5CM5eHpqNZhT9K+Y8/Gq015h/AmNl2Uo4B007fRUzgx369u1hl1bwrPnQuymSJ1kLng8MWa5EcNe
zQKWVbBWfK/nbfn65WjIdq+9Y3L69rkwHO+R5PQRsp7KsFIIpoC+XvLBJj2yDl9wTfRsGqm+E3iH
fscomcSOBWFoVO+0Vt7JooLRMbLC5Seoj5ujDBU9mCP5ZBlihA0s96+vdLyo719lI4duxlk/oD7L
GFt1CX5ncrxEZo6SVObLlAdfVNNwaG+RUK7/3zbfFNg6/4rXFxaFD3jz+hbOA9NKFuGZOwT0ZKsO
TW0F2jJb6mhnITyCP29e0EJvJ3DcBNkYD5gl6H6OIkjhqlCb7uJG2UAW/yiCxklk2IvCtqv3mfll
hm2FEYbMl2JpT9Tbf82zg9CUgDnok6A4Wv6ClouaKNRajQ5gfIcU/dnqK+4VbqD6WpFQoWOtLAJs
Y6yXuGwDrrnefpIew5UD7b3tq2oru9cfDGswnrdGRb+NOL13NkfDfA85eJWgpOPBSyCur7vnDbbg
8CcsVx3cP002HDLOcNaWNyvZ96xP43mWOmyFO5RncSJnHD4JhqoHFne+BidF28HeUjihCCaOAvxc
XId2lLLb0j6pnVG8jQiP+7u1t7m4pyfRjA8wgrUnxkaYkvsq3Af5sY7INywA2YXDl0son/Nswzx7
jwdqFStPuGgfYKdsPFHqnTtZGRt+sJp/y/DVOtqiOdYxPAAPWnJh+JD6KCRDQ/Ghtbub0HS+IsMJ
ntTUP31tprTLZ1oEj0vTXLi3r2UuB6jfPyIjU8PO3jrqD5JZjY3bjHEanqsfa5zK+eQA3GmNTjZs
uODs3zA9WjIiUD2GKH2bVbAsxq0Ns0y8iyPFlsYuerlg6GxcQJhrN68Z49UosbP56cq+0ZRBhdh6
Q8abuV/4Dr4kQnpXkqHa3fG3kdaSn4qmhPQ3pq5K2ynagNlkbP3TpyghWOYcESNxTd9loyBwN58p
7iX86Q25jJyctwj/9b/kZ+SSKXbYSubyPe6W2SVv+EeBviD4Ule+MEiW2CTqZdY5pTEJe+u+1Bfp
JwfvSzouDorh89U6SqqSXURDh885uMQVMRf7841+Jy9DYikO9IZXEZnTkweZNSBoPYijKeZxoC0w
worPlERTknf1SrBfJcU1CAct/Jp7bHF1P1LsNi9FW1sv1YxJ2SCgzvmhOEtBiCB2i0xZCqJVk4aR
+KOeG3TS4BRI/gGUPj6RVGjD1oDQ5DCcnffNJsMdKJw5dGnNAt39udq5j0qhC/A4vRq0yZbRB3o7
Br6Mxnr4JehzCf6TSBFrFomVKzfgLpL4cqb1c0NoDuTWX8n10WYV29OTkpTlO8guo9N06UETzbvb
qC6kig6jRvibpRzXzG99wU8HfliQQpy3L+IrJtFZVkTEnMUY0tVJMNP3qwoILNdaDviaLGF8otad
LPdJfMUjlBE71NtxJxLEx/XDlXN9r/Q0OoA4O+nRMLTtaNknt5NUV9RYv2Vmxp1UjwLOnNex26RV
qlDPw67Tr4qS+fbLS12WHUI/g3A5/gIhufRHiy0m+pJb4n7NODn9dzT0sE2OsSd4U9EFqd+rpCgL
zzh3xlbiibI8gIb6X77SaU480YN2pBn0ePyKQ3fNMTWtO+By2DIXv0+pnDbotggBR6nEUy+5YMxW
RWHpGWk5IuUJk5mP3/nHfNgxuH+ksM5pLC+beezi1TxwOFfOOjWmyg8IZCnMJJlARSb71OZIRfE/
foM3AFRXKqtNFscC+CuguQGr7rWQN68V3Os6zr8JknK5c0KfVoaQWQy+kQ0uVPQAEdE36g1trDi8
RQSrH9X8Ay2mF3NFMek9JTeRAAb0+OY7cHHRGhXgKLRGwpeFJcSeQJbkbCAPi7IKxQ5kvlkKU+EK
BED78lxL6lDir8FquThhKIiGJm2pgFs/jzDGpGe8hc9fUc9McH6x1R+uxQsNXG+GZFw2kuByAdkc
Yhe+Gecxgu1cKrbDjbnSzr1f6t9YUf2p4tEWUrY4UMCtCO7V9whI0/mn+S4LHtFmtogUscjJfYUv
MbBUki4sp8l4fFLUr6oZBJ1kk3iteeIiqobqOIt7ItxgV77GAZI/5kTijReZeJ7aKIyHRWmA5fh9
7VO12p5WvrHsq3+2zJY4Re6TfM/pWjR+E6SsocTyLSMUCw/xA5UdiqDJYT+XSC8V3nrveKCyGDBY
KhXo7oH3ZzDGHvuLwBFPkUuOiCGB6F83B59a6Thb8OB+P2tBMGMnMl0Zzj2MfmyjpsCh3FRiTM9u
BkXW4rH/WpQXiHDxsPj7YrWP7mnV8zNMvxBCAbnzE0WGTpzMGmJuKYKfAN5KkG4aqb+bE2Mz8Aof
Pon+El1tnLvsaw5tb5TEFan8WYGG0pCWQAgwn2c3FziEF9DToWZnp/urwbwEX/z5IhkCtaT1DeKo
yTLUrxIo8mo03LjW9/BuVQz86BwZj8H7PZmumLwmOOIz6WIVBsRbmUvj3MIHnYjKZhBEjIxKe4E7
lip2RDcRaGCDcPNqeI/fP/wRbzOlZKHUDLIDo+cWUo/f1QjfEOoI6wcu43Hu1EYp1UE0QvPwHWat
V7X3AXlu1oFni9hi6AmcqLbawM9qGvUnSxJR8pBy92EeMFoaakptacDwVQNhGLyRJjXS9vrv71ur
Tvf1EUgIgh3wnWG86vvGN8TS4eHqnRNOnxscNQ94h/t5Rn8nSiVFgzRzZwcpkobC5TFGaB/ZeQr6
OLtYfBOSifg4JfgyFyWD2XA/ra57vFlBOgdH+ytpv746pDdDLaInMQa0oYNKc9Vp+ZKXQARrHITu
oRTx41/x+s+e9ZCYjcMCiruuKvIMbiLUcSfqREBQW1jsrM+QnOXd1RXp8snyiAhQ+YOARokqX/5b
XJyOEDBy6oul+06uaiKL82taKgpMDsgFjBElmVi/8HmL/S2deyH2nuov25ha8W41Si4oI2DaZvQ5
B7a22brCZ+fj9WlUY6MvFUP1lD0mNqzTI06zE9YwA+EA/blSwpwuiUwNG4zl9dj/qKuD6sJ8HL08
ZRRN6gSf/kRcU8lZKqemDh8Q6hn/ur3QI/hrHUPVkopMpLzsKA59yMvEhcWcuHVfzNfL0PKXotOD
nbH9sxQMPx/McNf4XVc9ZBMXk7eiHiHoTMH7Qn/EyKUrVMoIy9VKoW2+nP1W2noa9Izk5uIivuHT
h1dPHmOEvCbIUw1fTmKx61FTRDXM75jk8s/D7KTtkqcCyUEcZUj+IpM+B+zXiX4SloOxGwIEoK+6
YB7yUKhh4+fn9Cm7mzcfY9f8WFDXTDots9YxsYGX6QnOErCuDC3s6K6yy6KBbAlOITX6bQWz0GKI
ew76pV8BpYHs1xAMJUBOYRnYqTk5WHixsiIzxSPnTF/TexPlKs4PIEGQ+8Q4l/GJzckLHUT+2uFd
SuZf2NTm8tBQKYA0E3w+4pG+hhF8uYubnkPPzy04VnHzNK9lOZRfovnSxgxq+Q/yN7aMySbZrGfT
ViqKDy3QKwbBPW2C7gpRtfU3sf3jp1nDF4yXeOdzDedHokan6iQKTEn4W2O3mCvZr3vOtV0OX4Po
UbTO6YZX8262jU+Rqb3UAusLSmwHj/InPvGRjmgqS0JBTd2G7smakkOO94B00FX7FkdXaGvYrlgq
9OgTNGWcA7/kItHdjUGgyOeMgUHQCPHfcwxux3DJT8Fc0fx2DNapK0kCUJhvYyXAldd0xqIbJ9ot
GiBjs+KAE7iZSbhmBr2GUsRNnMpzZk9cufOIPZ9ypkwoJNfbHrcaV1mhxrgdk2Y4F7eoZKm7hx6U
eqrRYI1+XcxZCwlgLPqdVwNshdfsFHhFKWSoXY/Y+RemVvhW16nPcL+eWa6KbzqetwldadS4ZOBW
c5xHB36cHQvPmF51f9irFyg2gBtWiOOozwNsikhnpHnMaxbKOT6ZM1huNyfGdqAFfFS4yi+ojqBp
EFbcnJFcnlWS7l0kmduPyxrSnz8x7SE11Mn1rHGglS1B1OAlhDZ3qfX+ZseWoRI+oTwJSG3dkl79
YM3503brZaVXm6rLk6JVQty8WMRh1xtzsoY2JL/dSiGj/1Wb3kl/CaTF1axz59MMII1kAx4WpDKU
j5uPlvfR10kxGbPttx0/XPcfkPe0irRscw9Z+UbELfpa35Of99Y/5QqR1Vkdbmx4HD6cA/KCAjEy
cCkn9cLABCf1YNJgPrNsbeZPNbN9jU4np8bj4c2IjiPuWGgWjSehwgn6T2c4XRnN7M0GRcZDBUTH
XNljcGYsP3zWCqIhBhlWNjl/zoh/u2eZxoK70VW4mNghh9YqGcBMZ4ke17rV1sOc3075e0iXzCzB
XfbzdQx6KaLlZqfTSpRipzO+yAkReEeZsl6PcL0BvWD7vfNRyQfdOfKLWHpsM2OV3lkV3wS8qJDo
/VzsLGZLD4OrS9VO0BT6FipP31MFpBfmvJjUJcTMcaAJ0qMFbu88LfEvNlWDWjOu9Ldv1ls3sXxU
fd+3mW8Eah+tMtijA4xx21PETsPlC9bOShuAfmWAJltQcJnP44i8+f8Esmb5U1mDz7bzT1p1Pcc9
az5yO3QxIwS0uY1JRUuTtChTkNrS5xGQnNPqvMbspzfo22blFnfUnZHL0HCYOCt/QORIcFG81ZQC
TqlSZPEnmeHXWpAM7qq94IZlFX5z7JC9oGQo03iQWrxgTpLzAG02WJRl9MrvfyeAVSAqr1kiyQ7J
gMQNSuQAtGKMq3Dfl+Pfm8S8Jc2EbBsWUZ9l1vdJqTFN+sP1u7llLstve3pNRc4pU7Ng/8JKXOpM
P2XL3H6PjClrndfhi+aauAz9GkOutcuW7uf4oOBzdZs+bNBnCMRv/vKHVJL7iIjAvn8dFfsoHDfB
hSa1FtzRapqrcPwZ7GmbVBFuUJa+oMUVd/HJwMji9g42JHPbVKhe0RQdGu3Vcifyts6+awJ34x6u
+dIexWAhcE2xfsyjdGc47dav/1Hui8e2aoPmaoNAVJrXi6FZ17SwOjJH//ZLeCz+V4HHs7HFYfxR
+fRFmQEhpDLiLt9D3BfrFR3VIdcd8bO/2/2faKg+LPYAb5BBOVZ2sGtY48NcNJr0X3dexxvtvPzu
im/jnQ44YJ27Y7pIPHQ7GXDE7whZgc8pasg/hTtkJPIVj9SBf6nw2Ti902idYSM/ZPvoQ8cWLomy
jkF/G5nGnDm4wtk1A/nncWuTajEgl65kkyovTIENTRxY8b+7/98H7NJBE99YlQflOFYr9qFpnxnx
14Lm1A3kQlzVBnDLZG+nGP+3Yz9av1A82xcroINH+6geORoo4HQ57NbmIThc/wrnDDsAy6ty3O4/
wY2SqxtJI+jQTUxWK1gYuguIAQcwNegEwzqf1vNBN5nITiUIF0aLk8jUq6QKTtK1/AaMIOSXNKPP
tUCEhLv6ZXNNy380owsrQhGgCrvv8ZwG3k1znrb5Nx9kpsg9DBq8AYOyWyaSKCw9AoVafqIF6PlM
+AakD24gxyvRyCJHLXnX3ZJHB8BGW2CS5OqKar7/S7EZHODKLAmTeVI3vpSzO0Wfv7mpE1jmdulp
FkAMMfx2sTWzicUgs/zvJlogzN4Zs10xnYimH3mL9TNH/i9qx/mpOYe1oLD95xdMwJtntAb4ls9a
3aIqs1PGUgqooFvz7cy2kTU2UrGk3dQmyjPPiXGJMvKirj2Qk94UafCCl/ARJUunyBldg4VYtF8k
o+rUkOtJ9V235VClD4ofFu/3BTBZn0TJVA+Be76osgR7VmCm/zFvnsOOXMS/c+oGIZBIEESRXSxy
ScH/JWRVb0TfAJWtGAg3xZIuell33u0EdwB1kFBcqyBHPTh1LTdwT8fIXBwYlccFCA7dPP9QRnQc
cvcXJelJKsDXtuFI625r0JCvSjVDd7n3ju8hN36s6RFDiyHGjx8sunlbO/MBomBGyZs2gRdMtJUb
NP7M2bJQf2vx1f7SQmIAHYplZZH427esxITm/zPq5dULMFCbGxzlQ5so1o+HgHnDDnNUASO1FFh3
VBdlDF/5XocH5phDPHpnnldHfz+uONp9uvZ52lYVuoEFdwb74lk91qOJ15RmszHkhyoWJ5GjOvGE
kg5ZrKN+s+nG1g2aE3qO4dFQuxsgLo23z1TgY2gKtsTcXSRKEa8/zW5EbaWIY0uovp1u/DFSsIS2
Wt37ZTi0TgiQ0tYHktDEyzyR3XJnuTihuezDMgbE3kPDO5BGmhcBfwxXBvsFVr2+KCr5waN3Tgm+
QCJ/SVMf/wsDPgJZq+9t+fq1lCCkoJGW9mIx5ja+lu+haRumA9asaTArSDqQNu7G5MEy1BPVp4Fl
OJaQWtN8u9+gRXAdwSUMP9bVWHGK95VmlsXOkS53FdJAadt8xYJsxMmoQT4m9+hnyEmveXX8AhFX
GFC1MF3HyEeDpC3D0JIt09+9IuDv2dPJE2bfRYT8egydVcS46HXkRBj1Mm9uHfZUTUgvDphkXrTQ
J7aQ249+MpzHJW0HhKndesoygLY63aRTD3g7g4DK8ViibvWG1WN0HlyYWlmCOc8sbMn8C1nJYUT0
HzetQNhJu8bpi3u8vBwhpjLQ9CyrQZ3txl3WroB7S9Ue+embe5Xs/YL47PlcQhZqCXPG6BX5ZYRv
gbqQZeqGoxXxoBHPAo7f+qDl/7/3mNI/QNIact7nR/uQuz0qS8YdrYEpA5A6iVFNuXYYu5+QcZlY
iOqhoJBbjrbiI57uIaH1KBkcfQjj+V/CscB/XSjUiSxa/0XmVqCVhFBj9ldpzg0Rey85uMo3S/Hu
yjtEttDRt5G9SYYQNf6BnDfKrPfrS/bLEHhBKLSKQgDSR0XvzpDhq1kzlq/I7f+wzggAsK+dQgrR
WwqLiQcIpJK5GHmp1a3q+7pE+gVCfYrRCS+UsFrGhPnYJ5S5YifAIoFisqWkU3RCsLT4HiIGyp9y
+k84xSXgKhKGLPvnMy25kq4EWU4vuZkiK3u35UBUXLn3Tiz+avalcho78WdmNUFWZ1aV0e0A8yhA
VI7AhfSsIVMN0VuMLvJfeq5sxzW4v8AvPCphfj5VQrdF6AG0UVdiinoopstBHU4YgKm4ZaNoMP/a
ZK8nQVb2OkPa3QRPjkteecnND+eTmJcWDd/vDu4Caor6jE2RAKfmYt91yPRrQIqBPTlE40wQ7Teh
Ix0tEKyh8dlwM6xw2F+bng75BU3GEDkIC21jTUt2kuuQB1uCYC5ooiEV0Vzh2Bovd6HFgzKrELFP
K2LFRYpVKRSCmJ+v210d0sMWvMkj1AWGmwojshD44DhdwCm8R4Q7jVk2LkMDu+CjjRxGKFrpEYSc
eaZsbJEfj0gnHZ7tM46qzU8ZJJdMCTEglFjyFxZnxSraG50GARmicR1iw6mxtMQJMxbB877d06+u
YZI3Zb4TFRWWBfcI+wD6egCu1gpyWuw0SXrbvhuxHFNCnXPv3REvcGXWyLNUOl8FpTR7l3ozm4Wx
MgNHH3K5ttEi4vFNPtQBW8p9OFGoVaOEyZ5E7FjIdmd7kHwhT6dUciFwN9AWLLKpmR01p5hbrgxA
+PduzqaX6jdDTogwULRsJS8383kyFk1Q+uB/Bz7tvAwiqt3tMSod0xyoYzi1hatOvmL+bhaN60NC
66SMHVLLxv4YFcDLzDB5kFsaVy6DOvHBVMeP+n7U56kHqi8QCMl3JhVonbMEEM1kSXVhuJOd0zRV
gNtEEdG+T/3RqCE94HrTIkqE0oKirbve2dl6iCNiZOcdSOh4PPW/6RDHrM5Nd1JYt9tq3KMT/hSB
0lAGMpIL3N9On7UsHhNlL3qV4WehgRgvWeJR13kxOXc1oC82EF53A4lOxdQsgKW7Ub3zXTxKZsaD
s0/S2ltwEMo3/fIkamPNtW0oVSMoqUiVYVlNDhjVuky6AUH6MXD9C5tX/J0/63TMHwgPWNOXW5Av
khx8ieptaC9ltpgqEQPD5k8ORi7wtNW0ZcNoFuIfT6IY+BWMxzbhde6wWG/okfWAz5QidlUDz4m4
tzfRq80j/0Qg+dd4VYrX/Yhm69g/T5NBlR4QzsXpaNreEckw+hGUX0mfyvUzVvpqMg8drlSRo6Vl
qp58Ma4BwrePkRA/k1LkE8HdatPmOyVJU6iY0qQU1q8vRirZ8ULiTykOw7/SI2YZojbWk7R7N1pg
VbV9IWXKmHmtUCzcw7IgM8Zb77I4ZXY/x0XG1h1w3ZSHZorjCXdZxmuAOK/dUl6pRoZI+/H6OfvC
IGqMCxz7vByppY6od6k7fomLtArTMvr3JgILqIqAsZ4XbKaTw7Wff3mLIIDtzo0ChwbLXCrUwZ7f
3HKkbsgpT+ilvpU0IPUgDbl+VO/ZM32qv7fr7MLZsL4R9wrxjrMIyx8091UHPm1YZBLGL8OP6QJY
pcpfAcOVIDRfICJ6+ZXFthg1R0AUVQYJHpAZMsxdlaLZ0ak1sZfDNXN3HaCtk0SaU6aanSvkvMii
xJN7ZVy3rjpTZNSD5XmBBIQhYe5r2DmKeB4HnRDa6tMXCczC4P3tnXhRX7btUB06A9q6jVY06Bvt
CjPbCC5sQS3MI86o14aZL9sxb276SyspGuHqdh3e8pMNlgP/XRGww2v1vtJjegeppTQkjkQWumn0
1p8S8ix+NGDo2ZVhGPc4qRjOe5PdyTrxRtKnPRuzupS3EaxgDHRpuOVjyl3uHDesAx8nONYpU+4h
Q5Qo0zTZ7bw7wFRkAmd8mBZwYpYVKQpeBRYLNSzpVQfUGZXwodzarcx/4LKF+443j4Dw+bFULxOJ
YCIi9Tg3YJAqQMrOIcMyA8m92+hwNDl1s9CyRt95Q2b2Px7s5iUEbQ6wCqAlefT1mdLKKbAhrXj6
Cw5UisGeRo+1sBHaQqmLtflkf8w3XejW6hYD+Vk0njNwAwvxwES/NiHaMueti6TWe8To6yNdeM7W
0LiPlG8wHFUEWATicaE7jEXsEx2+a5549az2b009KPx40bGi3OC4CWr5u3gtG07Apd/SUO9/d/ta
KfzBP5X7SLqZ3wGIyZ4ZaJsv3KO/BO7NRr+JohkjuA5FXAo/sJZFfLKhQft51d+k/RCwMAESE6sS
5Tt1LmrsgK3iQZ4eaj09xXRE8SBshOnjEZqtLRrRa5Rw6H2UtW1kX/QQ/v9pCn8DFQ08+qAxaaeG
7cIW2TcOjsPGEEo8kOh20Hsr6+zLQgaiHxyxMv5npAFOy1Gn64YE1ZqHjbtIa6tQi8vA5uJU5wVu
kWquPNkWOg/dy5vAbLQPPGM3htPFsGi7Zs+iWQP/SVU6nD85dcbEfKgMPtqJ6sQyrVAhvn69f6rv
tnZ+JhUYvSvHugP0D6c6lw8Zr3fGVJZ6epmYWRWzo5/CS1TM0ttXRL4+b1wkeB0Tsa9HZci4JBYG
cVly5suMIum+lcUY0ZavxYq8ndf7Xemf2XMHOExxGuNXlXuDFSU0FjOZ+jVET35ysGjodeQA1HTT
de7J018XgpRtbBkW4BLGc242/NgpzsGQtxQ56himgy8IZirAr2Xjq1Q1aCneYM1NBGgygxm9I0A3
nmL839zwhuMG/oiU+5ZrNlfPE41GnBMsfEszMzGufk95pVnDTgmP1A/dvFXuAbm1p+hhTHhLIMzs
UhRbIM4nBDnSRg9u7bVJK/bzJ0qxKJx3+FeW+dLiuR0SswqZoqwGCNIBdVrQX1uwqfDPx29647Zi
8R35FB6+m52zf7ljeTrSRA1aLIc4YvqWmRrUL7WjG1p/DGO5p7fXYGV6yTBwMEtb0rZjE1gkpP4i
S//Vt7Ul2Mlp0WQuY7pEPGfedc1jcaDVh6DM0oG6ImYbBeuczcAyBCewTujq/G4k4B+aJu99ym8U
k1eCbbo9//oW4hsE3wbLpZ+gSqE5Cur/LFNNhwPKj91GPLXNWBYYEeyEUho2Sw39u9ptVzcQNfti
uhtmmbNgnRnsp/QUcbVNWsoB0plxH2Uy3vfF+AmeBjACc4Q9hbaoTN6bvYQ3qBffNxKBl3Bj9OQv
qg4jmShIXsHDRmmOSOf/VjGZXDNc08segg3e5EhMKyk2XlF7+Mr/p4YeIZv69xYseJUzlZv9clCU
cTzMlHxIYSDqPlok0IsO3mFy0WEA8KLnVYXXy15J158PR2fwaLUvE9+93OGzF/2lUuXuF009ecyE
NhnmvCqoISzMKRNdeCPE+fsAkzzS/x7AuE38Bk3+IVTi6wbgYUA+EXFcKsRBFDFM7j1rYBHTVI4y
ZyBRduyzoYZpXY8QFOLPFBQ7pVSVOuXNdO2m7FogJqgbxiPkXB+nLGqVflg1WobC7xXkrPS6MfSx
oZfX2nJPscuSzeUnJOsSrpoarlKtkhC2ACQ8fyieQzu8YaLJi7u+15HK66vcnzWERnBBHrOkM2KO
5ymjt41gDUoWTOJAl6htuZTLJ0D9xQwEbX0mum8kuh2asCUX1179RELjGK7kV8LNlMlL+atGyD8i
jZiskMaohBVKUuCeA28/pSYqB5E6+3XPTXMu1i7MvuDfQQ7tKh2KZjRiTVn5F9yAd5WS4mqhnMws
TTAZpq4rLbL3S92v8/5TTc6WsZZJoU0eUxtkjKVj4s1VAneAn/PxMeWcQwGQGU+7MuUrNqMdLVM0
rjoHpoKhB71FjtAk/9+LBfBYjEru63Zpdj0Rde7MKrBEs1+hj/F1oTaU7yGyGj7loMPn/BhYXlKD
JmQGiufN5XJTXG2DVODwt+ocfxDVCNzxaEc5feiw1b/iJrHQINuCHP9Y7zULAwmWrO6mzpdQPKGp
w+yVAvB0zzs6e69JWOZVA7k8D2YP/Yg4grIdtzg+F1wpaOLyylrp+0G1dWLe6zKUPwGAckt/8gOV
SSI+/p1O4t11JVfvHa35D328ajekDAp0mEvMtSamYPypJALuI0qagThWwKmUUkH1nltUYsxfmJZB
7jsXIBMZm8AG+sv1MvKjyb28wURenew9jIz+HMZYtK+QFeij+WKyKpL18HuPRkRnC/bc77vL+nN8
fd+3cg5DBc9y1NPvp2E4RaTPdf4hppDsoBROZ/MdvojQhWg+1zqmpZUXqz7gEiZ+ZsWseXzSwlkZ
0e3Lf65lD2pQSIhpnK6vxYVrRVwN7MIUW9jzpXmAKvRGnwRkv34B+J3gTXaqLnofe7ydfn/KzBUm
OXxczg09cDqugVAJp8bkd4IwtoDITnA9udn9LHu0pdZE7bSfGPljOb7Y3LUtTsjlpzo2aauke5Do
GqP4R9R99wWb+1xrn1yk8Am2ea68xdMWbv7fMY5f15EU/LaZcSzApSFvomR6MFEsdmaK8dJ/hrQh
75XX/W7b1V4ZZJwzGfvRKiEwuZqiO5hV3/ldh3FwNAHO6JL6qexom2fiRRqfLwgadhRVFRT0pl8w
swlVOj+BzoRDvYc+zR8EwgufE9pngaROxFTtBkHDtjJPBtmzci7SErAbTcqhPg4HSYf8cXh6FF0I
WBSXqacrp6hI7hHJnjDEQrtkJ0E6ss2I+DnIuQaqT3f9E5I4xR/0jLVgcviM0IeKyd9N7DV7SszZ
ZNkN07KmkBUDBowUtNKQJ8sBG02Tb+1IgDq50ey4uhLJ1hdBtq59VU+NTWeGHPupkVnWalf+tpjU
L20Ft8eaic7iB9rzMi5YcXSz1WJaJySiGzIFrYyIwVVONFiwefv6MwSAY2HTemAC3uHOvRa0oQ7L
xPJ+BVobtiunbF1vs/53611H6n1gL7x+PbROI+h11ZJVmV+01KZM/nPSm16Yr1JWDv4HbChuuo9i
0i6Xp4FU7GcU0XtwN7o0+5/grq/vf4B0RhF/Li+qlma/NmALP/xcCMgaA+VZ23K3K9Ne3ufV0kff
MRAXZyCi1GpUsq8QblNPEpI7ilhhkInp7wkqq0IodpCnLgxDvC9RBdhFKc3esV3eewoO6s4iUdsN
tkKZG4zC7qyEvGgKz11TswrZ35tHF9XzSuoNST7HtIQ6ptyB7ZOdlpJuDg3muHXCaLenQOPCdjpu
6ZasDf3ACRrtfzSto9wN0rMph1Ixb6f7+A+N1HPYcW6M7WnQIUdV6of0Uv4FvixhGk8nXiHW6ZKG
jrhYV5t2QV/g+VaOUbblTvhU8A1vYQVS0baxCKTsJpeaRaOOLSuIcDVKRdIZ/tv0eoB1uef+p+mE
Q6EdnMb94A3GahFtyqLCdE2Z+p2EhclhuMKVtwvx9UsKvaLqxYsZYQIqyQ5mk3kaAZYw47Db0BgI
i+5lyIUc/MB7UYDnPJs5Ivs4Sph5xYyf8QR6REXQoeBKA0VcjxJClOU2Y/fP/thb1iawtYfIgekE
eyQw9g1XUnKsER38nwGzhfDyO9DkzBpgpdV4QXKuncpIzC+ABUWHhFBzn3d4D8I5rJxIkSj9HYzq
iqutaKxw4W9VEV21DL0hksyUTYDzlqkIeUq0+/otxQzprdYyPAYNwNv+PNsr1dId+bXnZqoa4Ah9
GJg9sBIhEfYJCeRDx690qBV5eZCBpCjT3kObzGSMSXHW6OkJ/O+pGD2QfMkTcdjK6LAagqfUDBA7
HTqPFPVD7M1QPAa5x3jnBLTSFcLQ+SuoHiXr6cGLSHMICikUv21EMcVM695jIPoTRRd4xIGqMQZc
c0sox6qI1A54e3ZlMbjbnzsBTr8RRvumm73dV2luoWMli95HZOO4B3b1V1negXamqN46137mMdkl
pKlotrJH4vxEbELaNRqhTU7ve173zAOe1ufRGjcBFLxTxQT8fE6vZeU2TCC/bL4DOSmMOX8aRwC7
zRIAfM0qg1GQhDUVBzpdacxFXFx3KjkKpsKgJJpJY3OiuZ/HaoSC5EXeh2hSo7EbLzcnP+ZiiOTR
kqs3l3lyYgI/tWkV94aeTjLEPWUROe/gl3+MIw5aZlkh4FXn1qU7leDySQUXJxYsGNx9LYG5mZhs
4jy8xEdhqnn5vI4p7xtpYjtS/BRcgMpG7V4zFIVlW2AkTvpu9cUIgDbiAaWJa+9iph3DodwvL+Q4
X9If9NTGMclM7KO5HWolsWBHLd+vjb+n0EcSuzLq8ukR4MktDewfvY84X7PESVkjrk/5fMyPNcxV
9yWc1A/DQbkPhfnuOEpq+PAdiggnM8BsGyrWL21SJFxjDHJaUqGVZOceW3zlkqN4gG63mzKUDekG
pm4KnvAil0eCBLl7dLhtuGnsy9rhPKX88qjAOwYcSGMxxcDlOEgDQznp0zx4TzTEuxX6GuwpyU1n
vCZZbZrHUHAEYrGGnfr0Rc/9JO9y89bg4n/Io1VllyBhIT6XvKDQ6sN5+CYEGWn2aEWlOvFnTAJU
M7mGtkvTX0THJVP8fGeotFmdY4KI1WuUQGLjdE3Jw6U7ESWwtM7KFDW1YQmY4a6p8axxsGxDJRgK
+9mZVMSGsOxUoyaI6970i5SdJFs21waG+SlMeefanX0xe/HHjaqLuSY4nPaEBRcEw1OBpNH0jfYH
gFG/p3HZ/3/C8QKBQ3Qoh1hEp7rK/RHCDhUxYERyZqghDUhcVaDuCEIy2CoFH9dMiZu34u25BH0p
+wD9dRFX9ogyTThaomuGEE8EXMptwb6p7hFInzjEllP5P8pVr1hRP7VV8KBMNY4jNMO77Hn6G4hf
yQHv0MBmuymSmx/Maig4paHMOdTbYjyn7QxIP6Rq2hb5Myvwdq348OJjWL1odAcOuK/5LuoAZwUC
sTpJC+L7tw5wKVStwV8cxSPNkdps4M16/YzoJEYpKWWIfnfI8a4aWQyViqPSETVHhfmuc1U/ZAJf
ilojzdjrkhAIYY/f/hLoI2M5hyBRwJpeonVpbZt5fOkV68YllE7VUEZpKZjAkYlWQWL0EZY34z5u
RWRkueleWx8aVhVlz78yNGLfrbfbbwl+VmK9m1YADeCTscLK9vo4coioOW01T9nE+zJNz6l9gVm9
s8mM2MlyuJRdmk0fLgqqnY0q0CR3Fn1+nhbhYGJgj8lWzndu/wD6o2WGM6zftaJPh2LHIKVaOrS0
kjrcUBd54bvYbdjjMLrg0503YFvKT9WTIJa45Xn2n8R5IByei3o0JKMlOkSAUh5PzVRfruthM5YG
O2IF9PwlBpRKqnQpkOw25xnssl4WX8kIpADqnOXEqUFa1mbO7CPse7T2KZY39/ssB2dW8DtEUap0
kY7k+AvV+ZigqYf4SouyYxFJo4OdYp1yMwTSde/93Lq1HNfmVFwkaH5gPfz90yp4T9OzWwS1uTZC
ueYscEnmYReQhvliqGiCOHUpqFxQVdEJl9XoWbJQU9u2J2JD1kIDedf4fGYY9jnT+Bkw0uCFYyRM
vFN/uBGmflGBfuLYWga6OG+jufFqB3QyYbxjem+PN4Uz0A/oiNk3U45IlQkJSlhSSubAwXVplnGP
rxrYjiH2bBi+f7TMP7KBpuLJCfQdNfxnZzPca+/7hcqATwrsPKWHuyhOeDkJuu4yxPAi0WaRX8Sq
N7VgcrBzNajjf5qPP/8GhYtpSb5vtAWrb0QWeCyhFM37VygAlU/PZn/c0MNhGlbO8Zdc529qm1JH
lxpFs3i4o/D3uNM3kXnsrM5lT2tIZCUv5cNcSTQWlQWNFYB7FDds1/NJr27nzqnYsLf64dljUVft
u0gGzxkIp40tlTDXzDR629AYkpWWYXP6JaMh8rDLT52530BHFwGKTbolQVcz0Ci6r84d5JQL8Vb4
dX08vbjhEcBXBH/oJEKzUA/AKMdz/Uz81HXUohqHSv4GSq5stFENueL61G2ysf4RDgrI3cyHgFEW
dJR8zwLaTnW8I+Tw3Ur+BmboSa0PIFpevklF+c857dHjm9JyJLzr0/ofCK2bO7Fs+QKCtbBc1YY1
x3U6vTeBUC5eEAwAB7lWwoJ75wSaFxdnlGxIMibTUgCPCY4gtVRQ5/mDAQUugyezNhmpmlayo3R5
t+C06jnE72WFBHssKju44IXHjfk9YgkTD8J48Mmhbx94HpNN01QgpRAChlQ10CUSY/CtAKxlNAYJ
SIV/XaJZrmUVzDVQTMxf0JSvqkTZ4XlC4SYq5oSYQNFiaEG9V2R1W82x42LKePxpyzgRaRtsjEuN
9Ar8byPMCJ1FrqqTb5IqWqtPISKGDXWYoV0e8qQDzr2Gt/G0xGiJV5PgJs4FnKJFP8XsMeS402wM
E4DdVbx4F0KQX6xufjC+XEB6vCETHmpdgPAKmNQbJmhUZEipWGh33mTDX9i4/MYPIxvT1aP1H+oR
mk9xpf/G2XXk/R3fc/d4oBFCpZYdizsk9mnEtrN/q8fhpq3/MKtPsAM1JM+VxA1Au/gXMKypPq/T
6HYLQ8TmjtQxUXwvj7djWGZNZe8sRj0oigbAhAISZG//fP/Rgolb7N63Se4pWIAiZB4bOpm7D/MD
kPvHu6mSRpwxK0psCXPScLkTGNXdqDK688QOLgTbOaPsLHqwJNPkcAPSpsfI/QVCRjZk5zxIqFGK
uwivtwafqFkcoSR3OP068B+DTBgbEFPKLMMz43jhKlX5YCneOh/UkBvKRV/VGti3chpvuixvcMao
J2332AZy/zEPWoBvOyoiPojeq2FDe5w65VBND9LJdXBRHJdKy6pvdu2Dv5SwKSz7HZT08qScBvso
Qvn5sDbaKPZDbAlkBt/wFV+DcsmtiwoRAUggR6EIr7/KDVzeC5LgxRUzgOBcpk6O3hHGCDMSFs/Q
swSfhz+XUV84u36xFmoh44u848MEEJd4dU0mTNuvSRYrfskZlIFmBD50W/jtf2n+6Jku9qlJosvd
q/EwMtCaa/hr3L0wiqcXW4AxQCn9VXxFrJCtPUqTpBK1Kj0IygNdQtVtxR81a6tIvLsPWjB6pj2a
2TVCmVt3svZE739u9rbqabRJqA3q/MEGN2PGB8Iaj9QjCpBKY9tDHYOrdfHR5Q/i/lV5oUu10jmU
Z8CxJG5hTxmFecyxdPgnxaRlmX8i06p/ce9qhhNZNfXMHtOeCFY4j2HeewdUvFDLOaWtgUJ11Qcf
DdQyKDhzzRksfypCnpZVLhNadMgL5hL+mEfERZf7KtfBQeXAapPQ8Xa8CzG5PvmHkDG5LJVjBDIp
gc8iORRF7TYaxIEd3D73q/+hMWsrIkSVieSsbMcYsiFxLp+cGS51HIzTQlE/gkfgV6whjV1WmZLc
2Up4h+tta4YPm+d2yQZbF78ETAMJeQqMHWcNc3UyUZ/jyRdfc0wjliP1PIgborLqSMVqYQu74Tvk
fEX8Hv3e5X8Z8BV6SyHnBCIMz7iuoAq8jRdSgMv2VCCCqIGyGMOTPd8DLp+CTeWQvcv6Zxp6oDIM
G+nDK31mMlHbqaM+l0AvNKreaw4CBZg7G1d230b+AlqMK2Wnu2cXxPdTJ9AX5n4tJ9iqx9KNpPts
Tmj2wnhFSXNfQq+xoyyl8gl0B2TNgpTQJJcVGjpKPBsWQJzTwEmK3KKOcxdWZwH93RzyW1kqR/Gi
2yzuiusguyw/sS9IInUvGkRLK2GEAc2qtIRV4nztnjKZjenR8RlRsozPjloD5uDFFrG7ftgtogq8
oDpvp3QXKgBH0dyiCU4Q5ySEML4b1w+bL0xjrXA8uklan0JgHwbVvj3ez3vR9g3WpBOPaZVFhzxX
A+iG66K0itF7c0Wvon1td8PPrnW55vQFTUs6FHmosbKAKo7aIxu1RrF72UW5peAAmwn95GegjiZ0
ETAjxSRVjgWbF2c3Iq6EtkwEKVfL819Gz0iKjJuNaAiugg9mF2t1Zc/z6Npspgu05aJKUZ5+xCoK
FxMG2vfFJVqj70SaoRGgFiTBTPwD7AFbaN20XcIawte7Gdn7jSjiKgWEJKJbUJ0sIYiKi7dXdHbJ
PWcyTjeinp9oAZT+w3uwv7i2rWYHKNwS436bS5THEXv0FgUwbqOE8fUxNPkfO7mOe+NcuPW1AeKI
YDkm+KiGc96GO8NcSmHVQR7E5EhUyE1AdOozk9BsDPw4bfFprV/Su2y9iF6T777F14ARtW+9TpNz
P9astzlqYTSztXfwA0j89hdrRqrLRkjov3rRHX+9tX1bcVyY0zZU5Nt/7v06m3P6s5u0wEVTUP4W
J2wB1pMyDcMGI2Sq0pfHsvuwEapHCagLf6wgk0/HEaE1X1G19YNaWJDJuTi3OE9qnSjk8eqJv4Uh
7VpfQZ49WlP/MjHq7v3ZaMQTpe0f+fonVqo15+BUASAv+sGKALPRX2NnbNTQ/2OAlcZ4BIYzSNy6
MfV0nvklIwLzinbOq1WxnC3MM9dJZOqaN7UzIh4qvMUltGJbJWPR+js6ZxM9+7kJtQbnj6MkYOBa
sGFPihHP1ri299+cZKI135VgLJWbacUyElqprZQkC4g/FMRKXd5SJ5iseONXTnex4ndSR6JoDTBJ
bFq8MZr9SuVBFiMCmvk/jAYLWTWxcy1uip9nQzAH8KfdKNhcRLgWVEyxJwTDs4SdXLoqkisY3In+
l+sngyZyCl/DafdZayHCdMy40gAIsN2I8bGjjMSsiAgafC8gDYQZwCqFl4ggU1Sha8FmJFFMLgtk
oEnrmDm2mMwfMDWW9CuBOOXucuPHQ0VyEjxUg20ZeHQwcg/IycwMB7+h5IFbWIA3feTAbDfcwlC2
If+4eKvWMSmoR+4PY4oXxpGbmzaGgxC5N+hkcBXlcbu1aJonoEyayVjqDxH8yvq8OB8nZEnJh6Tu
tAYAOhAR/X13bIk7Owlo9HCYHZapMQ/G8XXqaJEUGHv2DXkWSMYSo7uQk1Wf1JHYW9kM7f9ZlEE3
5d6vnjpbgeHiHOPXPCE3Dgz6hBxUEqqw2osraQafkh2YBDslWwD1bO/SLGw8vzq0LM9GBLaMB1MY
zkV9srumYlFIHlXjNBGSIstvUnl8m3FgErlYnKK99GdCGvg2uKD/22TQtPneiULxetXZcB8Dy6G3
yhoeZ/inZrMbgcCmsthAZ+GYKUQ0p5cPIipkvSWDIZZBfE9Hrzj9Zc7CEgQ3QgKjUwjprjnRPUnI
80aaqAmQqLIDLWQZ7y/rNL8RjMFsdFgOa75yHa01MgLsVjb2/R/+qwnc3gpBz+jvMey/NZG8kbuS
dt34prFViDbncJ2vD5uIyjwh8lqyBUS5v35Cl2FVMioC0UqJ4IdiYxbs4nCFVBf3rCHRpMDdOCQH
/AkWCP6iD1EoX+fZ63YDlQl/DxRePp+yBsv//pUzSifDx3m10pyPLkiHjA4grggU80QMRkFb0A+x
QfRoadgmxugTZ9vRZg3Z2fX3w3zroawCSTo9Q798b4zTlwHnM6gYX5KsS71zixpz6a3uh7QDN07d
QxFrdQhBVG3UhSkZvPzYQQ3tZoV1TXV3HQmd2Yp1GB9KF8bpmQo3xqJqNMjTVMYhWRjzkulvrLxP
rVSl/JGsYvfCg+p7BzT2fF9IcnhQKcEu3/x2QztnEsn+uvxc79m71+YRUEyFVaPQcsvg58ygSaLD
yiP2hyfa6Q5lMnlNaBGaC2IMdx9VXEA2fhxnZBhajeNyhd/ic6WrORgrp+D2ZKRYD+74Ky0kxuNl
7lrpmTLeaYw/drAAFmUMSPrzb/pouEI+7AMBC58s+jhDFVXRiEO2GfXgj9rIRgkX5YLXW2YQp2uJ
8SGo4wDFrEvZ5VoIfzfGFJslVQydHt+hFsxM/XW1toWmV255XZfeBH5oWm2Mzgud1GusClRlj+v0
EI594HHYQav+fNz4hCDpGnJFbw3xi93JGBcjV8asXj4S1MpC8Jv26sOXbsl38RVlraFQh+4zmVzM
cAOJrtvSQyRhdeacU8x6MzsW05OF0+txLYN5IfgcbLjHAZuyH9chHPM+em7m0Vz/VgSF+JHH8v4m
4N5htd4/wYAjfXJPtBsiNf250WEWRbkA/Dmuhk54Qjb1hj+Y0h41izgCOJP55CbbIvmy/3G2T2qx
5Jzb8m4Vn3QL9ZBuOeC3F/KYsenfAA0S9eoKrCI2sE+YMQlvCA7TKkm1n7MdFI+HsYbE5P8GgmXV
mhGLHl3nchGhUO2X03Jr395QtmAc5kYycW4VHeCDrkRpP31qTS82upQPGzpvcABTGDiQjUZJbhLp
vx5UXn33N6rkGeB6GJe1vK8UL2Z1Na4Ty/12jQuK8fGfNwfD8YNpwz7Oqp4F9fMtNH82pZ7lswcJ
o3elEXRe0HrktKbyY9DbxIqVpIeRAu8XVcfDcEPdNMpFkWEKPrqtomEdy87BW9AA5NKToEXlzRzI
qSdU4waVHi6H53SFCtFjDZBNAIN9IyvTirMOVW+3VNi8hW4bqDSP4w6TPBOHbVe/Z404ZJ2SLo4C
RdfIGFzZSgXkY+8oYK9YhI6yFh2KkTnxsmL7KP+jXbgNkpf+SvijAGD+UNDZLHSY9a3N8uUxZD6v
Hiz7RAN9eHIVMknME4Qu6n16jCQ9nfxJiawOrs09TLFzdj1MoTuH7p4OClR69egVdGXxxv7Uktoa
QWduYwKvbwRb3VYfoq3zUDW2KEzrPxV/hjVuZ+H9lOZ8N/4MfTGkbYNIlmT21mvQzJjycRTrNuAd
UUninwcwY7pBExGJ69YS8p4PwNbH9yAmK5qQlWsAOyhsK/bNGC5++2+N3UcTu+BlX6ERH+YV8Ehy
wqLhBdr2BlvRU1Q2dfwzjM8vKf2Ug9AsRE9d/Fm3oVhhUkg6uLjh7nB99zRjvIfxkR/Kkxy22a9G
CHwgaa9jow6XZu08UDpkV69+/pVMeVk+yOFalcJqQmiDgOiPyN5n/Aa8G+KsmL2F/vw0AwB8pJ9n
hP2X7ihux0JiG91kkHEGvMTKh2u0/+wGijQZdf9HmWpl+OqhCysI+OBPmWT1Gy0MZOu63go0XwKY
0qq3aVSYbVuPOesYOb6eG3kgVblGuzmz1Y32EXAmubw+HqlCWUAnY0Rn+PhzscQMekx9Gb3E915c
onIUVOmhh5Bco++nUDdPzlu1hWaUDGDTF53zlBWpMCmj0dPOzJrHmkRV3UGKK4vn+PaZglDk2NxI
IOfMl/bZVDlPqVjZMspY3a9xXv6qneO4i4RJmDIcrLBhSDIkEpOoogQKRao7RWMoAu1E8AHW88PL
D4R2JzxVNNht3VvsLHK+pOZI+M7EzYg/oEH3COP1hROV+WBJcSMp25XWW0ctMa3q5sWSE7x8zD8q
9OI2EjjIB7CATDpq3HQl1RUF/J0ZoB/FKU1QOt79Ve/98dOzXO1xkg9ketlDvu8A/QyYgRTASs/3
VKjOpnXNFS1yYGpsRACBvFbbiLz5i4S00EpgwmTLXRYHgCH2ESNQUj51rEQVrEE7DnBCv1xhTSV4
KyVG86H3SraVMXY21va96G7AV7Grm+1I3tN1OEuWa8qVPjnYC4bIUgHjDSghlqX77gFYEh7Cr1F2
X+pFj7hnUUxI18ck/Ft8mtGz537VobPmQTwQJDXjk4wRCJ2f0x3eLLI6mXuclvmgSqkgDt37yI6s
xymUOfYLV5dcVdObH2MkK8mRxkt6dFUYJQ8wtyyodYUv0AAZyAX52fvX8yUInWJTzBCbDVXCAwiV
SgD/T/4ic1trpC+MfiAr/z5HNrbwHBJurrcYVW1QaNtbaN3yvk6O0B+Z0tqPANnLx4wWGM4kzdLU
PLqH5mogubA2PekDO/FiklesR93KgGU+7NN75DMhw+3j5hEkLR7SyR2nud+OyKMBPCtTdNdxt84b
EwwN7YfoA7i4gyn8gMxEp6TmLanE4Fystydo73NCAi40nR+q2fVsY1Gau/l/U26GQjllDvwOHeUB
kr7p3/u8rf8rpEGxcMD3xm5SDoUwMY5NeuKecLpfrg3M97QTYflBXZCT2/vasqOQY+xCTYw0ejDV
mLPN79fEHcrPwSRvuneuZMJEIu2/cZgqGTWqGKIy40BjByCXWrV+uipimYVZEO3pV6NAyWnm9fHm
30zlkatzjx0f2cvlEv6VtOdfjdO4ENCrnoPkL78J3oAWHXRNGg+gHKtH7P4hM8BWx2Opca8iXOtL
AIE6RxPh7Tm5/s7ZODTUrZ4vRDyS2+T7cGfO5tiEr9UM0E9kI0IKWYdV8NWe9dadRgNaDfpFWxeV
/JgOA9eYCG+0JTuGF9HhHH4Mj/Qf2rC5JxnE7Ots36g+aK59/oTdQWvpFZdi7dgMBuzYniminWSs
bw24EqE/Uf/FTA/Vum9vW2RmFeUtaHpCLq57QSeR/d8AiD0wBiw8ON/p/HY6AW9MtI76ij7dsRBq
A0hqHBot+1rXsKRZpSjjPc+IwN7WBVjItwNwBo1uyg8LL68qMKMvnlRm3nZDJSeh6SLWLqPiRzew
ejEwtD4KE9cIklD1xnXFrCwk+XFS92L57S9M3s5xYc3CBQD5zlVzruXsCAb10z3bEcGylwMvBeSI
QBA/z3Ft1uirg1eGCRG0UHTXUSiS2VLuDSxOlkQ+8WNsGf+a/RixD211WIrVoonhyUKe8ygu1flA
nG3p886qin3I4f344RCRiKO0+gkJa+XVnVoYYt03sAPkXtOyQEdgbFe0O+6zKoSj2sBTKnJbw7Cj
l2IAXCbfuIKq/2PcWjQitKlge93uf9mOfwrfoCYKrgxRFoJPPDheUJtqVvOa99cGqwKn/MdaqBp6
aFjH+bPLCi+7kNr0k0Und8h969ip6IN0+0DtEnLWhIEwpzQ3qHtDYO67gUWG2DORT3iqBJ7b9IEG
6Z/X7BF8NcQ4XUBULHnYoaq44+MLHsowpIajrdJN/v/zOWwkP6TMJuj1QWafLSpegChwv23EgcDq
+ELJinduL36sH3KieEDdcBKCIckIA+lOjzqcJcoaZI2wrRYjhgksJSV8lHtPKcK+Gt6kPou5ROal
37EtP7W13YdkHqIRXyD3kJnuPQj0FAkiz4140XltvTbhnxFvUW1k9hb1DzrjHvsA0m3qIuGWWAaB
paRG2XO6/AZn8mT0GFozqXKnEe1oBf2zUyeuuuR7H7xgOVfUQjF2dOjhOPm7abF5OVagcXm6utU3
qslsDmuK7ctzVq0lSVPUL3LB5DD7mymGKsGM6A+DXyruhATUcH7kvsa3cETpN/Rgta3hg623gvOi
1qQUdxhyYu5HVr1+Te/nuJWGnAbh0v+85lW+qy2/AXC24FKHGrEMw+Nuj69E1cNI76XZYFYpr5dJ
8VbL5BM2DupdnqRkQ2S6BK4R/Zcz2RkWlTFVwvx0zfVt8d8ig/e0cyETXWwg2P+iquK8mNQzN53O
D0RcD1ARK8ock6ddBV/XUZIIHysao6goLPu1nwbsM0guMnhwmyuzHLMlUS9DtEspLfb/qdOW8EqM
p2Cqy+O5/53yDz90UoZOm7K5SePDy4lcrAuHf8N4Pv/T+upm3NUSMCCfd/DX4vaDO88wywLnGBkj
InDhFgsb34ZHRwVMJ6L1g8XxJixFQ9td+vzZOinIcmUnLCRuB0nZiaVjVhshFErbQCRDrvUXGouB
1c//md7UBYdKtQqCHgxl1CE1SzmsWl+a1b02TSiQxbWI0dBhfvDTCD/udLKHet89GC7deIouIPmi
1Yel4imVycNY74QlRfzuhhN7ATJeshvtPJ2d7cSA9RXzHn3Rwc9vCriNDEICaOURDVXAtBpdz6XX
KwTuTjtPOhmMuTF1Yo8ImqdJlwhc63w2jM5Lh6iOBlJWFZIr+AQ7P8FpDW9BCxbN9puXOMhXsL7w
eDGBoIKSsuK0JsUiF6+HHrMy8lVxUh3wyRq58jESUURI9WG1TjT8ObvRN8gYArIpAo7zx1qxGpsf
mP9A/u6+IY2Kbkp5318G3c5WWIbiFeTX2dlQMpUIGkCsw7x0hbI56L164HaJhJho8NSTtHpNc8tS
UPpao56KACA7X0ebCpKXxLAG1gK/h3Qa1x7oqsQT7h8Wsp/YNw18PBpWbiRcIAzadPtUGLe42Usw
VcXuIVENUgEdVsMUspE/Mof94vg+jqq0CHeryBB/DhFETEAaKE0lRKigGQdJ27V8AcWZqqOtbEio
ZOmEgaiqCl2DfVGkQ+vZcLl9RVIWp0B+10KKWvUVp9sRut3oTylSzy2QviZi02GKiuIFO+1D1p0T
DR5ePmC7Zx3Le3MVfeT4RQpEj4ssc+MH6LrqNvL1IybBU/j+mId0kgLvqq2rtsYVAJiqPBVsZwPX
fdwRt13+OQteYuH60d6oZLF3oXg2JnzVSP0M8PyWpu45uB19sQSUQM3hEDPEXbRvJb2PQaGhHaQH
W9qXjdqvy8HJErFnMIxviaXZ0GPaJEYrVKsVGXFbe6QAcaQUa8gRGhH5faulo6LniWO1ne8xhfOt
TmKlcRwYR9+0KVl7meSEhOU38x3LNOGgx7mt64aPN5HRDmvnscuFans9aXIwEgKCRp//cTN3HwIC
ZZHxGA0vJ8azdHKp8BXt8OAyoBIHiiv7UcRDaGJf4w3L5+MfOfkrmYBuAeauEFHBADv2nrGSe/A8
WCREnkbURcCStBO9B+kPHDGVDx/VHreLXZsI+L3u2OBYMK0DqThqtNKguNTo/xIo9KvhyA9/FHza
rTwBUhqDO/2g4Zb6xtWCdFKTdrhVZNfozbuO4VftG0a0BjRUvyQd2QhZZeU2SAuJKOAuDYemj4Vq
DegL25jwCgbqMhvJaro/y22xN5qccYreE6sXk9E2fBD0AeqrrJPpvoENEd9bGNIHKzueC3uiLtX/
gdd+EBysBj15OKK/cMIWcNIMvAB5HaNFIKs8R3wDqEUHwzTcKzeLDkX59HKZU3FBj6hnDpfEXWoh
DAuHw9/tuehQcpo/HsExxsgmEoM4FnUXXiSnnFKzAJvuq3XvFiYOywZUcWnORmraHXCeNMU+DqbD
22oKhJeDKTtbzFAzATpS6bDVAxQQiRQWxbJu8kHv1XIvZGIYxdcIJ/OkIn/gB/zj2YrArBuYcXGF
smGNNFeqRBeDnjHTPIK8ZYFjiS9yVvcDM0pVqD74/e80Kr8OPAmXKk/Vn1Iu1gW19QQPP4NmlB2f
Xzh+SpvHqdKMUOgR7LFd6DDV+iY7e78Jv04hLgPlK3brU7pZC6rlk6VUMBfIvfCVHPEmpV6qy3/F
9bloat8dR34AoDil/4gQIoXTRcVxsk6A/2PDwQkquvoOFLBL8oXb1zahviCuZ8sLfeA6aE3VEK9L
xu4Ll4HRjOi1dOG6IWvWwhOcrWeU+H5EFb4e1jdZX27ElhNOvjgq/FsdAcfBPezRHMDVblD8U4ws
trSydXAXu9YyoaDWnt0fkAoDpwMNrqdm3VlLsy8uEq17kst9Ve+ND7nxgCO65Glm92+yyJeeVqGg
ZPtqJxhNV487el2nUIwtm79p6A0NGC7w0GzjfCdvZU8xkiBF8Xc6KFVjStGPYwCr5XdI8XuHFeoY
ulyMyDhL97pkKqiHWGVAck76uAVdFvmy6jdh+hM5r6AOWPzhEc5DXAEncyOetqpLxYAV1IsqVOWg
YPCV/a0y9EvEssl7xN5RidkCt4g+D9GRuWnQF3pr1boOv+GBdn2ytgE0jXt3LPwhdZarTOjbP6Oy
54f7AygQmkWq062ZRclJifYagfSRW8xzjgQfKBNWzqjJ0QvwOuDmJ2CV/JS+e3sqdlcRBp3fIi0W
FkwhG7cQ68KUIjfYm1tTEKWa3egE38DHs/DoJk2N+xwNoaf4b58aRSWuUzZ1vrvUag3TcNjOmgDc
cnGlOPHNQmTMyuS4S6of0WNYAKzbpeWAPl6SeVh+Vm/1EL087wnAUDdkLsZ4cTa+VkJ3lA2/v+Id
ek2WacvgIv4gfqSqvMQsG3/XYea3aklccvwa1lGsbah58MVen4vfhCH6yHiW29fY6qPbQnFzbZ8p
3WDTsrhdqgHaPlWOomsn7zREAsX9BV+Wk7oKMjvhIirtSNxeUdRKmdcfiBumGd0tHCPXeTbsQk0w
eMQEfi8KFzN6h1pp9XdY0jS1OKFuB21a/e5rWgrW4bx5BEYkFKwRPeBQYJWSjeD3t/oKU565yodV
xB8ZrNn/ab+Y/VzX69Ds6y3EQbW2X+i4rXaGlpP34C2hc4rTdJI7Z4+Aeb5coUhF5QpTkkV3i5Fl
iJ2s5kQY8fzGZAuoRIqkIOABj9/esjmUOf4AEBNYWNcKYDto6FAAyLbb+mKiKaJdThZgQ5CfS0yw
VyBvv2s1TFuTyXUrl/6HbcGgNAm3tsyNiKipcobbNN2i05Y0Qtu6i/pm6vM1RS99uaBLnPZvaX8K
k57WoLWpKVIIVvfd7g9tQ6tkEtDiD3xixAQhQXqsg+5IpBnK4e5+PysCEfIMsrfdUd07ERT2tRkf
03se9RmCDMcBhknXaQ1XvaQiVcgDc7IWfmrWK+lCCsLpx8RkSNOg6DYq1YJNAPuFfYAdis1z6N/f
47EJHwvEarf3TRRbJnztmwZB0l0icMmI3Vxjhyojgze8Jkiq7vSAqtzNJhAyFBviQSnD6g3YUR6B
h6n9ziYCI3/WA6LfvL63Kee1nip9Yh74tJMfWKiX2+3Ef8IhE33920uvnAXREZVY8s6AXFqqBEfI
nX0A927FIoPfPA6AOj6sd1reEnYqFpe0E3FvDftkrh8G5FTozPIAGRY3VxCsgTwiPV2u5xl+pZtF
q0385AAJ8jSWpO4Xx1PghkCwrg/yUTF9LU6Sp18XcHEptKuP4msGfl13ImcXopbUQQh3kqJAFffW
aEbFgKqVxSrldNlnkVvMCjtk36Tze6NS5MYunqbnL0PkptgciN/DGkBNRFm4ikANT0Xfeev7ziGO
ER4sNHfyh584pQLnKtI5R/oGgOeEcMnkq/5QSL4yxnoW9gwukQ1GWrm2xcWJU/NMzdy/DYBSt7EP
jnUZ6U9ZHLk1sW9Pwcug0yYDrNnQIAdSHpR00UkBiHL1c2jn6OjV6VEwKQFZkuV4nUyZApsgvBEg
fC3qitaWCPFHSDuohLPxFXNw7NrzFIIoyylRezkUBajBH5EFU0uDfIK+dT/lL+drq9FNc6lJyelK
37uLT/vDWOPiGweZgaOejY7HaaxfnIHNxZNW8YzSYSdTgnF6N+UB8M/Ehz3JA1NATzgGcDlrYNwK
PNnAkjJomGW/VnmjkUc66BR23sZ8+wU13YbzpptzVbN8uL2wtTCv5bRHokwMH/AMdmjZYlmE3b9O
Ovz8IH8y+1nptMqoGLrjndLNTZXs7WZ6OcxQ5kOsQltsAum5dNLppFeqEJOgJmmNjzrYokWMHKv9
jmrOKxQpLeCrPGJtmYyD9YM6qrnr4SF7/Lzrd629iHhxmZ/brzH+XH1hMxR1bPD/aKZtRwGlmbK8
V0/TScv5ODtIq5SvI5GrseAJpkbIOvcZw4vLOAzNa/fPYrW3ttB2QmWnQyreAiRuUVZoi4CXDVib
kfzJu45Z5H3gdAseCGJ8uJunZFoWErUlx20fdfceu2tDqQzTWHCua1QiIK0t60RhNedq+a6H+qVr
6WHGkc38byOT/YxVUOyaDJy6oTD/7HWVlB3kG9F9ymKcZIjvivjAeAzoBZvnx0twDhRM0a/awERP
eg0Y+yMdGq/kjOhtMoblV4WqtRSsYxm6MW+924fr6iYuWP7V/A4mhq+x9Zue/fkxqgr98oFtQqwF
bWv/i9JrvZnVqY/LYohJI8lmabBfwHfnk9rv+dAWLHjZY6bNM+xbh8VcHbsosNeS2UCZUSof10fA
Sv4G18zlRvGut9eeiWJxnaZAP8TVAGQwuXz8Ul7LinzVwqIG+Z8xDJIvAZ4IUgPEjn0lo3xGoFf2
CfXY0JtEoo4VJBPSgpEktR1thJkXVsS9yUMvF2NSCA+Gp0I0tW/QM3973a8f7LTDyFA97CSi46Wb
JIjr2TSaMMbNvd2Q6J33aytp6QVGCiNKlUs63YXUljwBRtLpY3orKaZ+XrZyU6LGEmp8y3kDw7DR
dkMd9H5hixkrmYkgHPzPu5j4stAIE8FDfFGKSg6HgfRiMYiEkMi3KnnQ6aJtdEHW/TRioAyThT/g
6+NbVF+9vKzghgkEc9GybA1J96WE4vc0OD0ICCzQ8gzG8KrKVSep0XPysb3LKx9qjvJ+ALn0NpLF
mI3fJvqYDVo5jS5CJ3lfL9VrVPmV3tRio5D5jCLPcYO6m3wp6QwIgDgt/3/fHLHcuF4IJq+in4TP
SUaCRW4vDV0i0nlxmhp3A3QQRa4+7WSxgZ+mJWcN3RkAfTTTAPsyj6jo4SwPzsu199hRTDrERj5v
PNogIZyBE+meM5DOOtJ7MIyhi1JaeBp+zQniPGbn2Q+bQYoFJgP3XHaZoQQQjbbyz4W7hhdzRbyV
Fr/kQlN0xgv+fuFcmK8rHw6xpBuOOMSj/oFzIxvCRo01k1T97WPdu9CdpCL1xu71pU+hpY8hK49g
tbnl7LVupRH0Wom2xymgrii1pgOAT/E7xZBGzDC5MPS53Hdy0cuoE7CZmcqVEMd6tBgGpRBnw5GD
3Wv5x3uN+r3Owg/ycTfRiRzUGIn9Os2OVY1WuCPvvGyK753YQ7c92su4l4J4s7HM7clT+zssyq8j
yLTMJ5IGP3McUxm6lR7bO1lCcS75GM1JnwxPRXzWpLK6PPdV5QuwxdP+Bh25QwV/7bkaYsYoOs4l
qnZ5YWptqsTFBG86IHyzGywdmunCK9+6cCkPjIzq9/AVp3TynDXXa6JhAUeuyq39+1Vww9aXj90D
4H4FfzQAq88vYYni97lP/MISmj54L7CjvpnaQHk+YLxd0SdwOcPnacEBb/8rVHbu9M8ksWY2UpQV
ZEPt2vDbuZEVDG0+4aPwdGG4b1ZxvQJzl/67TKE0mEn4NumcuyAEu8i36/4hFTM1JXOSygleR4MP
sRyLcpqr03HBR4Y0EnLmSjlmm6vdrvmZoDHMTZMw9tdTE+9EcSK+BPe/pZ+d9q08Sb2E5/JpS0HN
6Qh/BpdOjdfnEmOkTqiaaf1jqMGSsecOecnlv0ZpbSxditMgUrHThQhGGCIdv7eGmeeu/MXYLqMn
q+OJJHuDb25eXSvux9tFe7X22rDFlRVu9SWYAx8I1Qr7zwOW2FFHyTV1o8BK6T7esTXO5grf38+V
Es2y+/IaIxpx/H5SnG7kL7avBgDsmzuqmKLY8cZCP4nPj2q88UxzhgNNSAQCU3m7wisc6n7TK2T5
6f15pLEtPt7bZrTbkt+RXtXhpeWyRFJibhboqHuFX0uJmaslI48DqRDS2RHUNDOoMVvyf8Othu9Y
a384XhrAZ4QqnQg/CwAKdamqLqIZNOE9GziXf9zaqhdtIla9NjaCmFuuxa/mvAaAKmU3kcuRHfbC
3zKYPJYpSj3LXf98WT46lMkLd8r4yX8vkn1FUPEq5ts3wkCmBMS2ftby2Ev0RuQLNwlMyLe/+lnZ
okVy5CTEav1NKom4iM3LImSAI85QxjxkQL6uHNpUsvBgrB2soiSnueCd6q81UavhX/+TYLLx6J03
/wrKJL2i4WnGqmKgLFmJre+FO8u0RHrvGfGuzun0xIl2T/wX0fMAxEnNSTBNgrlR3qCz4I7d8c4G
maOb7mI9ds0OkfpzcTllF9102uc35zGkdqGT7441iNqnDTeEU1FBt50PtSJpbgw/O+a2YGQ7jXBp
58N0UvuXDBKIWY5bmuYdYO0CKcYj9EC1tLOLsc225jiz8Rhfgkv7TsWEe/KrJ/gzw7mc//oTuJ5A
qKWf30QYjcBLxocRe6ujOj9o360qpL/2uni/dyAKlACNKNwwrNNCCw0+alndNOwQlBuBEmh8QmbP
6Ine7W9zbdIpNtmku7hvpHY/4rKnAqxrhGcL8JHj/5uGfXYVKqlSFtxgAh/mie0oWKhPsUJU8xcT
lMvKxzcChfaKga0kIx2FgNVmGYHo2S2AkgLN5V3KoJWeU2sqTGnQWdbyBelmzRDIczRxHURCTXqc
f576EFW2A6V1bgcsG6jHOQRlJ2J/37AsS1FEhPPUcevif5ol+PFVpUsDkdbA7604vKtD3ijP5OWU
OEcaQAP7dfUQm+j0cfnzeKpqEGDI/yY2io/4NQSta8XS1DZAsn4GEjZTCo0CiHweMevyAjQaC+G/
GLrTsRGY4lJHg8HOk5YxF1ikMXEDo8M0ZE2k4sqDdtIK2TXNLzjPair4qzJD8Pwck8EJY9r/6HW5
2jJ3e5jPPwP+LyQe6dEaIYumzUYxC84hCTqFJrZrYV2/R++Bigi1EBCqzKu+ypYUJGU9mPe6HsT0
2+7miQaXaqyfrzuJtkO4DnNTPoYp6gVW9UX922lTs5LaUGg5U/+lNlKTfMnXoyCJUvzAx0BW+b4T
KL8z9V2lHgsQb+Xbv0trDYj6HyEfViqBT1Y5MMLSvMLE3HpfYfS2dIrScpkdKHBFMSKCavlAW4Nk
EkS+6HTwfr9iZXOgNcvWQwFVc1oWNjv/DPhEv84MbXiEi3GCKMEA+SrATjXZXh+YsZsr0oW6SrbI
i4NdUQhkb0wjBkp1HxUhMJwJwdb4/bhsorVlhuatwmYFnQfJDk2OOtVA+BEAksdmC6fjhdnx6XiH
5sJRUeoIxxtMl402mokLREYqqmaTWFwIkcffzqyRFhvPv1uVxgLXzzhHXqrUHrVaUI0nbqQ7JwrF
pURZyUg+yGmzjfD1GZf9Md2siChTB2XY/laJ6hqOONY9e/bWLF2KwcwL0WXCdCy1wIrtonwMC9c7
3V/qf9l+pL8tm4EXh0SaJEgxSjNcuXDxIOa8+e+C6sIOEh9ydicu6gzdxD+vZ4tMYd1iSFUFpF4O
roZeN2Yi5P4zTfFQgieMT9fkw330R3OTwmRON5oWxx4wz8UTfRdtJOD4vsy96UqsPVV+WULVMxyU
gn615NZDqAAnh9Q2itDvgkz2OIyDfc2Gli30zf3imPlvrn6JU8e/QgrNGq7jRFSoajxTASB8a8iH
LP+EWTwxC2PYGoWtWS7iVGDdtLSLkG4E8aS6OpUxILKPrIxnMNLyIgD4maoFBhfQ3srowpSLykLX
Kl270CL+VY7DswHXvdzO6IwdT/3xgnTUjMl40tm3tncmcboIT5VGKSnFxBTUowFbk+vkEc5zaTdc
8K/WnRH6B6UOE2C1FRh48l4fX4hjo0E98wZptuYys3LILhV2E++wQI0ofsAhH+tjq7PWkeLlrIQI
7TqJlMLqUXnv13z3cESjcWLgDcMnSnThjh3l1ATKfsHpq+W6WCvw4RW3Q8xEnVS0dmbkXTmdDadk
qWAeNIfSOJ6cJAUHAyUqMkiFIOK9/Q+eKkEMlibLff/TUxZUo4qR1ISHg00JS5dsEJ8R18JWWOUW
Xh2MR0F5RWiyKpaQfjroPqv54748HXW/4GkWW4GBEIBhtG0P5wMMme9Ty4Uv6BApbMwzODeCxa5z
S1+3VXdI0ki3Wz8LGBa3FoinqeHJ8md+o9oY8s8F4PCirpHzTqkd1HrJ86bKPU4iMHF9FNipfY5B
yPS2Xuz5Wyo6wU6Bq85r6BL93evgmSa6YpyuqAXxE5XWwncgSNujNFSukr56GVuQxUGur6cM22iV
xAYvuEVoiK9UQ+0O66v3Oe356lOtbrUusEMOEIltCo2uuPmVfx/cr+MrFjczlSaKmJRHwovmj4LI
5cQpDTJhy5pqcb6whra2M2A4hLHCQJnbGl+sCJryeUpH78in1+QScm/i71BBitA+iMDkKMWYtMA2
7Jon3IS4VUd2Kkm6pzhRHCUITKXqkN9MSMuB/C9qhMZhvfDps3istbWWrcw/YqHt+ItS6xwN/tRJ
q7p9lB/1wY2FKbLXxXOufOl3kc/LnFe4om7elkucYpHipn3Ed1mqFRrJcdphNGMp1/EZWP6ud8Cl
NpHZK09m7p6iqRtpMVMCvAXCiviuCX9Uosxwchlj11J4esf7xDkn2JKCjpuqfNevwREr4A3OCu3L
KlxhBIpMwKbbQ7Sijr4csbigB3UTrfV2is6sw2CibzEEkehEDqTcbKrVWxJFJ2On/jychNbyOjh1
keI1KUBKRgr3NyrD26GvoZ+gszDtx8DpucC0Pnk78le1+WQS3GrOQv1s6u9/GzEqgl3EkMpt6Vv1
ypIMsJTp4bSmkN+mnG4y+MCGXm4TNbJWr1+FkoyFwaaby/YTUSH1dZcdboQ/89FbQcMci6EYts9B
ORPDwSo4IfokmDuaD7j9xo4ffB0Er8zyhhJDGHJtdj9D/QlLlplTkb1VJqIc2Nx4fyQqQ6wj4CQW
gRPXc3LhTXPSN2p1m67lc3f/eln+amBrkpZblyF1oLh0/FX5amh4YFNVYQCLAn/U+q1gdBn2dM4e
N86/CpjTVi/Qa/yz1XJVlKODqJQEcoQ4tGPr5nkNaHdCj6iWmEsddV04CZURQvivJ45sCi1aU0G6
7BAJ0XatT5Fzn1gAFJtD0vUS2PngdhVBnV4k3YkYdk5lQ/bZ0kH6zI5ysWbw+TwUb57F1QNpYvB3
RoyaIDA39Z2GishtOG/gh/JzAXQY7WsGryJhbXKGxnbC3QTWxWlYU51k01R7Cy9YrPEkBbce6LnZ
gOAFqLhOvUYd0dnNMzoQNTEOFwU6l5FYK3dXMiGYVfpUgZ6YOJeaMFMxTtP+eQI3FLZEk6KR0W+e
vZFYhVhZvUD0iSN9KhWo0wkgKyNtiA3EPt2yZEgYCs85QVP017xxSO3wKPMmTaZfJKjr2AnVzhJ2
d3FL6e3BLe0rfYeInql4MX6zU8DVKntFR7mYsmoLwqcblHM6YHnjxEKwYlohXNHQP50n5hLdIkmY
HAuZUpLC/sNCtbbQTZr1QpmqeaqIEKaOt3BYYSyUZrQ+LcjtANZVSv/nFjHP+BUPKB6qBDRR8aKN
VCU6cwpJ9oJXbkkFAO0F/r/QgXVkJipuR/mLw8TxJHeiGx7jlzhNrpjvD4LDlRebTCRh6lZJqSq2
L4/NwTct842QuRulp5gdQtVV/g92k9eNBaX3KQZhhIRtReOU6FsDaOJRA7peClgYZ1G2D2gr5QUE
QOIPGlVPDDKmnQRaTioeNg5snStA3fdTGaMBG/31n4gK81X/hiDBZVD3cQQCn8a2CkqDr7JAv1xt
j1Qk3fx61Ll5UQOUzA7SSQYe8nUl4rxqjoaub+rq2CCOU4iRS7FCeC02HNQhtjPlZnL+AXzEP2Zo
rUFJv81+H1ISMu0TsT6RbENeNo/d5DFvgX3eTkveWOSxnll67hvH9zkRGPRomiMQyZbw6Wtjjfm5
mxgBHQmQtvO4yu3yIVNp5Q0rHiNV7isSq1PfrKrahYA/49OMzRxE7+PVPgA/Qrdpmwtm7gqZ57io
oJV1w0rlKTdW2omZU9XtKS4U1qDElsKb1Cw6d7fjSPRfgUBTNkUp1q9KfJ6xBjhUamJLjFkpc936
Z+OfNtS4Km9oPHJgnZ3yrFEH59po1tCPzu9SuB7ouljHi7lmX/jdLC0eBiZ9ENli6eaRRErgJEvx
mGTbY5AsR+mtwmliStE4dhtS+I7P+2zQ2mChDNLZqkP3PeGCNp8CurpWJYO8eAHtZ/iJOjxNtjEU
Kwzs+iKqOT2B9hZTMjalBt8IFLvmELP01f9jiyh5z2csWO1gMHmsASQzhYDiR3iyqIHng6hUnKbZ
mHxcNRteJpCx7H/HJDCXpWIDDZbQcJ5PqpeqUpswATWy9dv/hAa37Rhb7HERTnjEdXN35VxXpG60
UTyoNTiV2dCQc93DkjLPBlmjnOY7PZFeZjf+YH17w0Sg9GfyzR2QQQKfuPcvfV/4SQjFUzYdG4rm
9CzeNnMuDVhJZ0CjX/c0j+m2kswlkqewwg1WKTu/BNSUB9YkGZlfCxLZf1fB5AABdkeaVpbfhkOx
qWuQSS2Z2UgJ1cDEkCaXO9l/1s0nszFTERCSQI8Bg9XZwhBm0ScLR08mycZy4bI/HlLD5sjM7mcH
0ch7xwcuGY2RTH4GCqp6K7HGCuBJonMKrjcazkMDHpf5vZVOIT/m+higgILuosp2Gz55e7loAbKQ
pbKn2VS6gewRfRcANCUEauodmzF1h+FPYl5eUvZBbt9w20cUuIV1pnG8GujZKrn77T1Uu8gtf+yK
ylge8/OLzKxZ/ZJU/Ke6rQwUKuurrc6+UvVxE9ooA2Q6qzA+psl05ADVy5chuJwVccIrFPPj9jvv
XR0RmkSDFA7vHetFgyyufBlyPDhR7tRMxVurEiUE80elBCT1N2hYH5AKvCMenB9eN2e39Oxge1IE
3z0CyW6VKEfyv3FOOby41OmE61SU9uNQa9kOMo0PDjw/8EkTWLta0qaT88YtMs44RKrZYxkesbqY
1jMKYbWVzI56D2KZIhcNfaJWN57Wz2kDWL3sBZ+D9ONcVgcaodR4gGWpDM2qmqusTyNku7Kw4cgW
vkt8p+nQZGh4xBfnT2H+H1r6mnMnWN8czQjHdDqi0+44r4+c8/fvuqyXtWnEcalawQ1aUSBRHvW6
8znKimjLo+ZXdlmDejPpqK9T911NNMuPuVQYPXN1i3iqOz7wPlWPSedT213awkWpW0BCDHk3krCx
YSixVxBOpueIVCWO8pTHT3rXOJBCl27VL0TDeU1f4WLJcDcoYbV0i+NcazQRiX+YeSX8h+USXkTn
qDXM1yStmRBF0VgwKU4+/AOxIZs92yiwnx6+sjsurmUBOT2gGewxI8Pp1abA5u74HX04BMbWw/BF
WQWgYeQycuU7Wg88h2LhmM29QOjUvPw+GnO89Rod6zJ5LtpzTmbsz3v/DLvd/ozX27Ko97MgK6Qe
wLYtlhqadKg1Qy1KjDbl4t2ys9sGAp1I7RO2f1pCYMVD+VsoGhovmtOveF2Iy7LJdb6fWwW1HNcZ
SpVd1yjDKPxRifQ7o8tNUdDy6+Qtxu8T0zcMd0dfA05Kym9ukLm8MP1hjW7JdvHGlQCSq2lrHsN4
q7ZRJl1/HGxPEW3b6kO2KFkv6+eT4hNNokYs2yba2jCzlcdhUcWsMbNWM3ecMrHhdLHVxs4PqE4m
gxAHtuTMddyWXjS2UlPAyVJaWK1UJdTOnAnnkmT81WlwDkNLDOfRa541HAN6sAyHSt4aFnkJDdB7
aUWPQGUjXPCvdL1QgrUWHiWyryfH2NUwXIB4Z8xKUsY01gXp/en9gOCO6wdAk6viErnJT2BnYSe+
dYV3NLVXpWDnVWoZaBQgpjbu1XHMsE3uKK1eRISfVipk2hdjWZsbKqYU7BM9XWESjM9f3OCaPCfb
j7sNkJOFxyuYgNjUkzxH2h/Zf0+QZ6disIB77i3IHxjAq1AovNmZtndvR8KkzZWcbjlZ0W+R56zl
ViHEDzrWuxlnXsxStvqBOEht9NupSGDej4G3VcE+dSWSIMAjSGou6PME4OOtm8GCJ9e++WwzmDFp
4iDl1aQkL74LARI1eSREpXUyokNtcBcTh2OiJb0150Hecz/tQ2jVWlEZBtA0GWtLktVGh+sK9Le8
ayZ8OlgPSdXt633AmylbmhPdAEBpjpJ8Yy3oNbntuIF2fMUJx3dEKr33faKHhicVYxG/DkW+GEOS
ydxbbdFJoxrZSJCFKDd1mAJMT/RZLe2ZMQCYur1BWQDUVljbWvTfsvHqWLk1TnzjGor2dsRiRu8Y
D6FhPff1NYf7w8/BTCQ2JiLCG7RRi60UXUymY/2FbidgUQraOUHns+XMajs20AqVnRPSV7EIfdlh
AOEflOqAbeDt0hFvM1WnCYixOckYsodjh8oASbaGLT5JrdlTonexeHPArkW6lZpa+CJgvRfNFBxp
E9xPgZFspjWksaL5PrjlT0mtvMJibEuXa4BW4yh6GXblL23ROdjOcRPZ6poj5KvGUTnX/ho3toqf
XYc7jSe+bCju9saMs1Ov/CxQxoetMnNm1D9/QIT/uJraHPfOl0ykBGta6YzRGfPfZZLGMaTakQWE
C1fG6SiJosZd
`pragma protect end_protected
