// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:53 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
R6/WZjIrPj2/X2qYSxH6BXPH1D85fwg2BjBs1HyO5Zldp5BqVx4Ps/MtcyBZfK1T
68b/uPUKSR6c0J4y2TxpGqDtGPbRR4IQXbmq/eVXBoM+Uvi/py2FhjiomPnoeZzS
ITgY9aATCf4r8oj2Dn9Cro9zX8i5z3UoHTnugymbm44=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58368)
5blwKCFS5cVMAk/dOHaYEW0iZcUWiydR8sM5/wNVsqgNzNLp/ExY8AwQS0/hzt3Y
Uk/S8BaajTD/d7pNiM1GxOabmM+B/zF4GqwCjUWkgW/zBP9WpFeYcvMJxxMYotaw
zFj02OywgS9UUQZPKZHk6YwC3+Q2gapHdgn2HyiBjIB7fi+K13Ne4QIhmPxOhoSp
AeqPUILVYRsrFo4pWYuSQNxGrxLLaP4xAUjOF4B8nTFyEVlJCPcXE2NDzbiHnvy+
gIwZRxXeYx0oUlHQIrDYPzkAjxXzkPKzmm0pBor6Nq+O5C0bA7DC0yKSVJZQQ8oE
+yr1OaaEXwOEfjq8XnelLZtltnC5WXkXIGumZYNcSorpD9x3YZR79hC2lHpjsaa8
1+l2SU5AwjvszoVJx5GbzNZF8PNMhMBpphy0Cp4243VWFWyucMDrzHRfEZIz5cO0
jWw2FmTZO+PjUw7yBAY10c3Jh5n+BWz99jMXXJqTvI3vWORtkGWqEu1dEQvGwnj9
xuVUF6tXMxYl1GQX36G2lL0TiWsfeUr5JjjAVN/jWqOVDF9smy/9quyxWzDUehwe
dMzM8WGPiyMJTbfGJqoxG8bdk4xsxcYlalgdclT1cdG3D2+4SvKE+uo3kcijMGan
0O+mq+q5M+TLi04tty22JRzBTLPExYHIUY0j1QzHQleQF7zytxqux+Sueeyr4AeS
Omqt4tUnVQSkHv9LBASPMEjig1PSKRqcGPbn7gmeBn4BFcYUo/ECLiZ73PDvmX/I
EtG6kR6xQ7nf4aLd2pW/DSUI4yzS4DdCVfpqkJNoF1i8z/oQYeIDzgSW3EL4vqBe
VdP2WVGheXZUcEyURwHNci6nVlRoHlIcq1afbQGRyDQZ5eCSj+6TDm9/ZY513vf5
Iz1uT8m7JFf9DXpQr4U5WUZuExeCMoGjxVrO6wBGU6AlyiciqAhcqgvwSXPPJLkB
ivpg2XTEkdut9NUzyvshbIinEVk0iCCs2+yRU8RmzsSpd0Imt8jMBS+XOzmVpibK
Hu0Cuxja0Lxb0GLCAuqMTCdsB+tN0j75kap7nKLqtvsikdHjCKyHfHHwP4i5wFPX
43rvelceJmErQjrM4xcRRqzUJHihOh8hrjxHWCCkGiMOtNqLPGrq5RuqO/g3C1J+
HnttJr7+amv0jbHV4WvgD/BJwo/6+M9q+N5JrUarEYyHpBFHzDm+mPY4x2dTAZ5d
tH97BiDA6FUjWDYUy8noTlwE0bjyr1caGW/jqx58MnImdm/JFhm8v5QWLELkOYW3
K5MDpv0cLDelwUT0nOH0Eii4hVw1AHcyZfTq/ri5SdLQzVtRDRYvW9rJGofaZKkM
AW8n+JzBK0zHMLuXTGjMw6fhtt1Svx4PCA/JNDCnl8INqS+rZx4QiktVti1Q0d7S
zZRyWdTy41fvXMnSQJ6DjwC/Q73xintfQOzfZWRzIaiRxlQtFmxZtGmA4cEm/9Ny
kFrpM8knWwmM/jUWmj2HhJ5cAOGqJZ6x/eYm70yp7oy8+9s5/mFVWeJp2XUzSPii
73UCfXTu/kSFBkgXXUm1HW7w8/o9kGwpjCBhLRFbJbaD2Vpg7/2aE+oxLOcdbf1q
Yu4ILA1pDjxAF+y+J1tyyf6TtJ7wz0ZyMHfSVKCU6s9DvSNuDBUKXxCNPC3seUeR
xPujaFeZ6CyuwxApqVhlYsGg2G3xfLtnNEA1YstIbDHYoiQYghNeYyqWzOUkqwKl
EdlBwJBr8y6ImtovGYzWnHB+KhdsDVDo99CZD7lf+zEY5xEHHEHxFvtmaLyM4GJt
x0E3Px508EJrv3XD9I9Clh4mOsOC28fkANBLESXU71dY1cjEtncfsbKY4xKpk1of
nfkETxpM9L2LFT4rTGIUMy1Qe36xoRCKIwEl4V+Zkla9LcSx0MNBuEu/skMe1wB1
u3FQzlzcYlrKwIaObSJyY1HNANXcVrCEZk9QK8TxL1Q12T7U29lJK7hzHKJQh/41
wCRLWpYMJtoKFT3mh+ixS0cTlnlgT8KSP6oB3yTtWYjzly4thMzBU2E+gX1xbNVQ
VGcKWuz1ixJU0q0KbaaNBXBUARX9rQFlZ+ZCenjUDzuGCPugMZxqFrmkYhHH1M8l
4+X3Fr38SipEH20s2gIVYlsvqtHYKXJKdV8/ls8FX6AVO47+hIffu+bFbJ3z+DSE
gH1M5/a245OZhIVRxtaQ+MvKT4oDm5snSLMUV0hS6l2wkJeS+EpA0AWz99QqyScO
IBEFwtVAeFaMXDO9GmcMCRTXyfNdQs8NEmcaEZkocnlXXKW+3V9Hcera0gpi5E6G
sa1SsbG000hUixn0zdFJLTeD0tFT2WpuuBi9NGnriwKQxYBX2vmpeTnjKUbUUiyI
tR3csED+3p3dkL/GqAdHhD3xsRnz334rQlEGCJUUa9y+TUNRFij8iW4p5vl/qsxO
SwY3oExdKHkRSMueCrIxwANPyUkLD/G1PdyoQQXOzBl55pn3ACMmYfV3YSeanyDb
rqbm9/Mc5v4GriOUF7N46ifeg6omMuaCIrnG9M6feTRs/WtSDB5pSytw0OJB7bQw
GLh1v14pOWQc0ZHWDTKHASbc2X/G4fu0xnNIoyGpnizlTv81CBVk+D/IRE18XG+P
2Mhn94oRj+Qjpv/MBUkn09dsHx8GwMYT72cwlkiSIiPUeAhoJwx5YK4cWHCBumDI
6glEyOIo/GZB82gMX5CsxZq0Al9UJQp1brWnVtLAbAquZxdkU3IYzSzFHLYSe6TG
ZOB9jeZa9MomPZ0r1izuK//ExGqKd5ieN+14+PLtEkl4/MjjFcAl+7pjx0x4ykK0
N7341dMRuhLhvnYxqFJp2eC4J5B7OqWm0NF+fQcP5P1CMvJn+rMZwTvqdmFwdXqy
IDm+9r04Htj7ZiIO428i0cDN/Ok0WWZ3eQ6gkqy96Atkp6nxB45MqgMm2j8anmsg
ZTCm6wTsQJ8gZk3WXgR5ds0OEwerrSzUgfnV0YABkIWUEEEeoOb9jhG5/RAndoyu
wW3K76JE/kcVU0k4Cogx5oNdSH3DV73HewKG5xlOI55mAr/0BK2MajRq968179rr
Q6FaN+fFVvcBvwtq916CD67wVqIthEo5FQDxx2cBx+P7c119zlK8Y2hu1a0Xg0IN
Q1JvMa4qsXYsrxym8yePWoNr6cRnj4os+rM29nh6okKg2hvcs2rtUwj/KwnbNY7L
+8iOgOFKE52Oh8N4fqlInTyoTdcwGRqzN28ui2dKSeAlkJDD1PyFofuHsOhE50Hv
y3m32B4YsJ5ODAiyF9jxt615NQTEqAEttBujOIoRRQLs5OdhsqOmcVd1VsZ8U0rt
cjjEoAOxu2QhcqSHui6QgWYlAQaOchH0bK19CTpZsT5ltiw9mT2jChGGsLq7XYLr
5/uT6l2FDnu3F5G3Sg8v701yMTnJttvbo/LonYlWlT8aycrq63+QS7RfOHZkKTJd
vBkNqHDVQ/x/jyizGDN7RSUs2r3L3Z9hJiBk0mXTQiMGM9TrFz04pOk+H4G82NZA
9DNoCEGgcL/yNxnVuaznjaQTouooCvt/oeynvDN5miJY0HPH95fK/K0LGgN+sR5i
yrY+sldaisQgiEhiwNhzTb+7axd7sxqcG9lCHpTIc5mD2WhXi9C3DmswK245vh7J
5RLjoPe6e3Xj75IgpfT46Di0AztOS6F9KGXy0A0/sAecs1ORuIfF1cEFOfm2s/nJ
oVrjX4H2yWPXB48nL089dOIKTrXbnyWLMcEYcOy9lm2E89QbuxLCA/Yfsvbo6iTl
36XX4HnmDxLXMjIUHq2FjUo1CLf5NSnlk5A2XdOIJhdrMY/Hhs3s90WSAWso1B4q
DFA8KHuhT0MqLK9wx94TmgbLoJU1VOzEMPEGZAHO89XmVUKDmX927vV14d+eiugm
RQ+qIofI9Arx89pbuFyKO10LiZL3Y85McdXOUjZaJ0e+Efyqlf79/S6Boh2Nwe+0
I3cClfkvSAPIVdEck23UVs0D4GFucoD3lUNno028CHQGt3PDv41SEedoZl1HgZNO
Z/BH+l62XBhCilApmzRHIxJWMpNI56gaVsXnnFKqNLEkgbmbRaoD472vSJIZWVrt
37biHlfqOauxQLKWC+jmdvx1NwoYJRVdntXiuzzECjVf/Ag39tjdGZz+2Dzjc13V
5zsIQx/WmuaDhs6cHCKzC6flGFu+FsyZUOyxCKC0jzsF52S2sRf6BizQVLI5TG4E
63NOeXdgyQ+NPG7gLUr34zBnZ4ZyS8VmZU9RWXRGior9iqsRsVOTH+y6j2ka7dhV
AbRD2WkNaxV3Nh+v2yWuFA3cZiz/DpE96ONUmuA+/SQ6BukRR/x2kbd0HtrFYsL/
CO8SQ/Rer/E/Ec3HuofWkXlhqc4kqIH7FR/ltNLczQH6lHe6yFKzvJDU+UDabjFt
yj5C6mwgOfus5IkEOjdLZWPUqzAJcBOAEJS2pBen78FXTkkYpvW3LSft1SCroUfd
XuyADaPwnl31bYVhE3PGLz+ioi/+Ltc/1DI7YPLjnuK2aLAHN6DIR2eQO23Xqbiy
oDg/CxYknNQqIVPjJ9Rw1oLcFJVykuql2DxeE4uEIYPMCfpoiU/M/zNuecZg49/2
bRxosixt0DTr2uuGIvEucb9v9Dj/zM/hERQzPhxwtHpqHCGIavJwTYiyO0sKpVhk
MnU9afl/NvSzUjllVI8KfmAM9pvRl4PaFZpJe2cJVAV9LgYz5ltCsR6LZHR4c5jO
B3sU9PonE1LDNfYEdGxT7DlOq8KH7SsCZmaQ5Dn1pJMDz3yEYYnRQKj6nujZRUvg
432KEHyuwKfkTfOYWe0tDZLBwSue05F8MpOQ0RKO3RAak+k/V4e4tf7FsBCMPIkS
/CgBXNhpBcbIsv11BnZN4zSrek1DoVMCNrvc7wpk8juEHUQbL6r8q1KuHU1Sgvr9
U8x8infQUETnh+rukiUUfiuWexz/1ATBSNVLaF7Auc+UalGXfzYnwstVJKxISdr9
E3buk3ZvivExEmEWsiHq7flqa3dJH++JqR1WyHTQRBteYSf10YOia7yQxqzPNuxf
TxnRyEm0AAgePux3zDD4NJ6gbw/z+l0xbIGlDc1XPP4OkcaSFbl6hIR23YGJnmRI
ddbWUtGWZGVP79oiPV4+wmhLWK87/RZRvNRATRfKAFmCgL2ufCtctNxrc38FoCgH
XKOc2QYWM2QeRlnlD89WHU0q6dxAPiStU7Uj0yl9FfNs35IvbHCCvpkGBEtaEWOp
0dL58A1aiRCUzztbOU8EjSv2UKnagyn5rsqH2iLF20SGa8LJQd6fEui2OejE4AsM
lIug5xU4gbGdCRnWXf5LpLV+dXD1UWZB0oSO3EnaMlIiAPBcTOmf2NN+jCXL8vQ/
+mQX4++nOa4waexABeIYI8ljlJiww40/y/CGjhjRK3e6KKV2qF2tXjJcNDBHN3eQ
lvpfW4kI1JVbfkTTr8CnzUtCrq9EkogXKJRGxUV7BDk3SrQJMXb91SE7ePKe28fV
yf0fifKUyXjG8wwQYEhxqkARXFyzhFQ5bjQU3uI2RV7ZtHqr25I/ZOnkS5YMbIoX
NsSrjKnmUUlMHe8XC10YnsoUmLELyt3zVPhYSINJDonNgit6qnx2v+1nslaR/C6V
Os2lq/js67gzyotVkRkN+PtW/l6x3XcwOpNwnugcZq0HGqerEobGvu8WFjAtoDJE
PiD/pdnBdqIxZ7rszmpimk+ZoEothBnbkQP9kRU4xWiUN2fiYROauBO6xZEI0yYd
CvNRyTIjLpSbJ3AF+/UEFJNhI8qXIfr4AtGON5PnLP/BPiUf4/qdIBlAV6wmOsAb
UFtQoPs3Xr2Btp8/CKAcuvcd0+w312gVcW/R43EeX1LCdvXBeKOqthNmAYqPkRof
Lb0pHh9QfmzxB3ZOSf3kiEGo/sbTtV68NVWIBTKdiPHCgEVU6+AYAxtW09tqHves
GLWRrM11qmKig2BMVoPTu430TxxtFYxjjkXhWAcNRwATpMbXN4bD9Kk2Z3dyPEn0
DpM4t/ZhOLKAeQRm6wtSsyVHvO5E4RsTqLnOcuZCxm6zz8vKAFVzOjF/+4pr3kn4
T9/kR7xz3nj+P8Au71vRKxjduK9FFoRt/eo1XCZLnZxYJ5jSI9VTzt6x4Nswq3Rs
VTxiCwuuVo9UfDSfY0jIq0mIkHYGtJ1QhtqYJPiT9mVe0dCSYk284moNX4b+YzVt
yCi69orzhWmu1UjeUz6LXcLB7EOeHp3/Ie6tdB7j8jXcCjHt6BOhEH3urRRnAZGV
t4sUpEyaZqMOJynw1NBwGVOWXOVi+MYcVW56HjaxMjBOzr7OWU+fy9n5MDk+JaMl
lrT0D/21OAmTi2CWfy6JhA6350MfxKbajwwjiRhexPI3tdJ3HOY3izJiCaPneAAg
V2hAdxT+BqXeAHfM8cPfC1+wXjeI6gb/R2CqXNVI76Kqkd4AwDlZHs1W3TJm6hfY
eSPKeoKEXv039undBAjEll7ddXl9o7k/7UK2w+CGX0npEDTmg+qc5wcJwujI4pbg
+fbK+lW8exVxqjYaESJ8OFI/9lt0zr8oe+SCsFa5M2590rWUw2WiNm5vYT0x4ofV
QoQxyl6ZPii7rNk3QG8vVB3RKqWYdzuwaGWUGQaP7F4ERdt9WJLX2LkNc1cxAm/a
Y0qZVwABCjhUE11Bw+MOJQ3oofKlIpsgUebx44cVDE//PHtfJ7zDCpk60OmDSMsV
tKOH8+/1xT5lZrCUzq1LhEzSLMGg2tJu3aq/3VkWWFeTXsE821QXvK5dqP/lQU9Q
fFAhTKLZD8MVf7lZ88JkGftgVg3nyVVZGnZf6xdY87JElIWzRJxQdOr0Nt+pbcw2
znlyPVkyXMoPkyx35zQvPUGnGnOeyUL6WG3j3SDH3CpI6H5f0mMv2HR630oRB2va
g0kF284h5yQ8lXm7ogpdBd5MwAItFGJbc0O+CnDjrnYlHp9DA2d8z2iMevYlQ6c8
LdS+c29ypXpclD9yVHXIIv9Wv1srsbXwa5vJ1+IbQWbPWdj0QZWArZPt/M3pIcWh
8QGja0dPl3pdqTSDbxTZNKMPiAL6TLGBZqvp6yvubuTpzNk/f+DgwqGiyu+pEBD7
XtWdQ7V9a9USywQDvVhIBT5u59IS4scz2D+uHxdKrOWJ2ELCKI6UynwbuLB+C2PU
vU/DTrjtvvHaSWleVbbAAcNFMPAPzGplMu+x7w08hNW1zu5M15tiez/84LOu14L3
2dD6OroCyPmgAUZwlRqlbWRZn5TSGeIw3VnV5zSDvwd2DUdcsU90+mk/Z8WbSFLs
joRaI+n6OSKjKFLNYWCv/QIWRunznSiVyWDlQ2w9aBNchSX3hXlAteu+LlQKTgZS
4QmRuXWYyyZEaWaLqKJ9w4kp7C+Vf5b09SzznJ+Zc0vJK7PfHYbNR67neU5Ff2lw
UDYwt7LSBxCaoyTOBb6P15jeS1J1cS99MtNbdz0SQki+n99VZ6ywoQgVAmNY9MVr
3XDTKl0mIcVnmWq8F7MdEFEJAgA09Og+Q8BDac8bKA3mVeZkXEbtau1bHIxwuErx
5LmG33/Ig1ZiH2R7awJthcnJ5KCev9l6OJfW2TmjHSpmwqZuopCTUQsQurfXSkgo
L7BBQRiL9daE3eqY9+CRsUjG5lkFrlF4zrFoaU9IZ7Gqm9W2Cv2aCLAwctND73YH
QOnz/UGP/McY2MZcOaaXqQkj/dQNc+TtMfPeqfvVp0s+xS1wAbIZjQqudtbOvgMh
UfJh9fiSomPPzxC6rgbO4TK3VpyPgUuIgoGs9fBksCutYDLvjxwiN+4tGRYnyoTm
liWGi+9LnC36OnR6CZ7KK5nz17BiuASZ3MysJYIYh4FqfQI2mma0790Xo9qv6PTP
WMexLr8gRnl6hv9wkOOH4K8sFtvHYZp/8Y+Ss+y/6SLYt+9CzNapboBaZ2asWFTy
IoF/d8Hy93/3nqfHE33/sKP+TnLReqNaCPc+QCvhaAiWNi+ZV+XNaw6r4i7uQp52
IQzYbx4m0ke61mlVrjU9SdiWIfZmkTdgFsIIai6d8ZLW6QdLlReaKProzHdStniR
oyTS7kSgsHgOcS5n705OXOeqyRfenKrHNnOEEu8QDNuBCmH8BIUlcxqBCusOjmvy
/wcHePpTk3/emVR75mwKHvsC8YhafKoxbFOyzyNwXcYhom2E4ngcPnyNR2CzaQ7V
kap2+8/Wyye8SLVF+LLsNwT6mx6hhyx0mKOvNTN0HWWxV3o9IDvstvcQnjrrkus5
iCk5LKT3aRKOHStB3vojmm99wP0NVBypHggSzH24b7HMx73TBTNY9TuQMJ0hDMTk
XQ0IZdY5tEwpvGgvq38Os6MGr3hCO1WEtFpOwKezgRKxsMRcVTu1CkSnzKx1cEfG
nAEOYFy6k5g/C6rr8Igqg0bf3TiJb31k48NPZ7y3gVdwTcSr57NaW5VjakG3Niko
e66BQ1SPyrYz1oVMvL6UGECyf5sOy6dKg/C36+wLMb6pb3HJYdmGGMSqItGHUK/V
dbmMG4+Bv0k6Tb+a94I5Mc+ov/zZ3H7BaBnIe6NcIubQQ1wErsukMeDFaB484WB7
oEepbQi7Ifd38tx5U1pNMjIKUxeqr+bqqEenOKAhHdjvg6uH+MPhheW99Yh70D7H
5x1JhdQlBlvgDlkjIUhQpBlD3s5LrDNI4f2U5Q2XLsCpwdlovEvmjn2CMoVba8Ld
hqI3AblxtFlFkseHXmFd1USnJh6qWUdItUF9PFSvVZb1g4EcxbggCRFa6iC10WoO
wuKdJtxpuoxUJKDohm0qN9OspDkkh+XuJ0QpzRwfckrmHP17kYO5aixWBa1GvRzJ
8DCJuctDA/90of8dcditKsL/qU60MxN/SUrMzt00vVc7E/qAB3FkLBCOMBxfNUKg
oDiNlzLpueq92QK8CIYar0pxrJlESW5X0p3zvwJ8aWFbe/LvmlkEzTSj/j7dJN4V
tXLWAGOopfUPWWDSUwX83xxV68WYnG2tZQyWEpp+dgBAIJMHKCkx4TzL6IpcpdVA
OdQp+XCNBRPJXv2xbsdL/UVr45gG70DSFvz0zj8Iu13QLJsYkhYSx+TzYllBUhZ9
3/5P+DsANmXGaY6laM5Rxcl3HZ/C4Dvjf57PZlMfQyA5GAWuQkGmVPanqzfeZMua
IqvrkXqzLMOD3x1q/ygZUPQHEwacP1Js+v5Ys392/oYfwURiXJQz4Jc8DlLX7wWN
3pSLC62Ez4hd+dPeksR0Z80YplyHOJutqmbWDJ7NrkuneutulYi6mgesOh6DFIjq
ZMln+LPdemTKQ+vEMuGvWEyqiVB3zBb2vtwCPRCsuzw7LgxpC+ycCZ5aYZN4Tvpa
dvDVpXl5PKuhuQ3yFKkVvXdGIwMRFBMuoYkfvgqVMMZ5I55U0iAEjqSDt7fd9Udc
b0/Wxr/J0r4ECVeVkc6NUP61o2DXlw4TNwYjFBfhF6Bk1/C/9rqzm9utYylJav4E
iDejc3GPCHsH4CwtMny30ygAjyKPgZEvuDWpUgImwvKOJMHwVBiijvXHdl6GPhDg
RoKVitkaY/WCAwgAQX8xMJ0/ccbqWJfkXGigLFYszi/M6RMuYyD7dlqLcw0cUhJV
gLzktZw6ubSn1ypM/W7BU9hcUWzA21I0jgLv7bltYya8WALX5QXY42uqY0X4ErYg
em/g3exqr/S07Xh1rm/xu/6/v9aGlR8rtr9je/J7BGDmtrfGXZtgFny5LZAMYCsn
tOjY95sJ46UYjJ3FkuuFBgsKCy2KsKqXBvqIGiCcgqZEiUQ0ahDiGe+vhpGiSs79
s+g2v3HEtN+8P/woa2cnz8fadr/+gbGbz7TLgEy7wGfjjH+MHq6AYfIXleBFdEd1
tu3Bkh4PXjytBArh9azJJU8pb9B/79eZG0/OM5D4UfsC7GesHS0yVAqOYZIuzvKk
sg1E2WZEkQJ//tmis/DAAvP+dI/5L62FwR5i25VJIldwOZTbI1DRAQnS472WHlpX
6E5a7zToNwKJkrb/Is1ipdzugGAQ0Dec+P0cjLGBFoY6K57wUHzksQLqeA0vFG8E
UXQ/xFL84NmMbJlfaYqsJMgkkP+QsP3xLZwwyMc8sLyKExttLArbOpiF1mbsM0Rr
BnCQ/1/ymRXipnBASROmg8Z8UOvtsPUZFYqN1FMz3qT8YHGpqc154pyY/K3xp5Iw
h1085K2doLM8mDtoUri04p/YJPfFkVE4yP6BbnPvVnnsSzfTzGdLqRnZhi7Siv1D
vLVW6LaayUY1i5tevLsiFX8BuVbSz4LpHvfb3OVoTp+kbDhOmgU19dGvWVRb3Ur/
5lXRfvTLRAxXeWrQY3MSJ1qoo3H3WHvhZMUPsXSsMnz8TrU7i76tB6fQQx2qCMy1
C5oGkph05cKKDf/s03gZoJNzrmQqG/wsxP00V/b/PvB1AIwnane9f1uaZRYLbqdE
YcEPG4TyHhW82+8s/yJ/wOYIgtyMzu3USJ42yPt9lA0AUpA6mL0WPbGYzkcPNFUd
ognUHEwYv2S9YY1BCnC+HMx0nrmpAhqCf9rxJ5uVspo6tb4BIdL/PYDFugwUJZtW
16RjzoSsgJjbtKV6YB6mricdPLUH20wB1K9Y5w+9YD4jQxdcPj6erK4+2bFu63Md
qBVH29ZyZ68RzxlD3NtEiQAuxdD4zXpLLb7wuo0c3tW5JRjhBrhGRtvFeTyizADk
QdeXrdscPd0GwwEppecthHAwhP10nE/GCuavsNcm9vRRoQFqy2b9/IyUBfqRU2JX
XvhEcqqlXjKE+ONMdQecF+dvVQPxJXfQmtX0b0s0Udvl/8gZTGPbARwXbFY0Wsqj
OjEJkTxIR2bbAuoHvUlTK6DK4QQh4dNSWtj96ZSkctz8V/hykG9wpy3WpEJBbUdg
IN9AJ+twOWiJqN6JuvAbmIjojxCn2iCdSexqf90R+vgSXGbOBSngy3PuDytM94Wx
XV0cxr45g7gY7vM8ltZOXvgkpNxC/bwGZ+2IpNpX1MnEsAu8PaM+Xn6/ii9MLUqm
YZnvDpBPkcJ2sku2eIEeCUzay1qisbsyyUIjpA/xd+g5iJiwMTMO/RMCKBN110/d
XzNyiRqqkb2d/XRT9e2SJtoUn3bxFXrIwAKeidz3YuBfJOGt+bpXi30oZkz+8G1M
je0oaqZSS92FMBNnGMQg7NVHg6ScD91Dah6uIZsd4pXVTLiGcUXVl7JU54OBCJ6V
B/BTgim6e5wwSd2fpwnHMfUhmCb+pz4QIkbaCNleIEKakHz0Cd/+tsHibgfqdnZt
2CzKxLBhKsJFW0BDwoMmG8hN0tZ2WSDwNtzK573Lhm1njbcLi7RB3m+mttPCYHOF
oIT5c4AMVTM91kHDgMx+gEKLgMaGy7qs76mvims6TMMKla9JVxqCbLFyA6/xFmuM
o2Pa2KNE3DsiMtrn/fn8luEWN84rEmmP8QgO3lh18yXxLOC73w6w1TuFPbjXmyte
LXBNCpk0mzNWsFV4+vO1XV7WIL/27hdezjXz44W6TMXFd8Sq55NcvGWGTbL6rrIK
gKnTz0CGTg9206ZRvs87NycSLD7vR0+KaNnLc0exvwWPSPs2rq6SVqbX5r1JCy2w
JKVh2Z/dWvYOVXdTRMm1gvxLF/Kmw48Ee1/229RQKVUp2BPiwp0jMxivZkyaEvSA
VvQ2BMzSFdV74VTRfBfOlzv4Y/NKuIcR3gvfMo12qCpQmCAF31GS8RgPuNSK1ZDc
IV6kGfFlJp8JuYyA6DwT8LCkctvv1NzBzd31Dvbm3In0WEA5wZAxsz1J6HTkzOty
A20do4gL8d79go3W18LUm7K+5jrVHOVubR8GX1RmqN5lb7+aUAo7rD3ztxOSz2hz
2M7txL8DBss27gMnwfFMDEvK43Peju8JeuAGwu1tZCZ6LV4Nek7fJJhpTbIIKxjV
WqXkBeQv9+kYoIXtjJu+M0CdrxEkJ6jwvUrAlWRlFN/pXS6c7DfRfWltrHBBlCZm
SxIQIxszaPT+51CYDzS3qBdRuDevDp3BVlHov3HcY44W7IdZ0x75LFD/dc7YY654
7/3OQcc+585/M7qDnZiXyaVioxJeXbefFIYqusPq/r82cMTHklYfpN2syESfBUzF
UfaDIU2hUYkQdk942VcgwrTVsDizABt/N81rMyxMc/2WLjkGXuxZuz+WqrR1/TIV
Dvh8xDj/hnGC/QSkzgGFphIRxJakiOvEjEG1wh+Ggts3mIEbfjfPiKlLFi/087O/
860w+13HKAl59J4oYPXTWuMjOQp4q3cfV8BAo7T6HU04EVrqUFMThLfQmbhKQzBN
oGkpJFzs83JKnTGLoHCconcfjWUj1cxygPaXACnOlic82K76RWQokOk0+xIzimdO
h5Rlb5v80tCGPypnC9+jfigckymA8la6VVgysSV3djfWTLKzNMrlcs46c8VBmSKt
tUWHsYPA18kcRghWbRjFZ8R36Pqv+dkKlmval4eZZsqgM2+xClqLNwVXyf1s7NPK
NU6VA6RdpB6C9vpl3KsTdAPk7bKqAkreNEtk4sekRrNgkb1i/WOi3o27gGqURQck
g1fdpeuxp1CVuVjnT8NslgPL8dDgIVc5KJONzfM8H+ojrNtaMVjEYKhheY+yvfTT
XRI6FO04/Z3QehYJ3F9zYijyNxCQCgvS4hhZ9OUaftlsjE9PkOHiuWE+tUR5xKlF
IpMWRC3WsSgew8yR6mRGA/kYUyFjIq4S5Y55PHXMuorPI9I5UUJpcYF5MZj4wf6k
mVPFYTJGs27iMhWR6lc/0iYJIqM9Rr5A2sfnmyMHYPxJD3A9lEfDpMBImzXpPWV2
4rMcooxsdGSLJAHY4fFs0gDf5Ed48SARWaa1LA9omBKWP+NjMoS5gPxPCSYxuluk
PnLgdwpgU5p+Os92UXQgFU1YuEFiyvzi3GTlcaWU0Eqm+04jRVnpBHFZ2sYvk0qv
bSDTl1t44DUgQNDHLjx914nLscP8a1GD0yxfGlqsv3+oMxYNQ/mGtSxSRgzVxAN4
Mx9/TR8KNJBNbWim0dCI8aN5OANL2TJtectgANrUBSMHs0sx89ZPS0pOHucuH+sq
V7C9Q2Ch5JEqhC0IVPk24B7fvk37RT4g01uvCtMu8qoo+merHx+3os+9oyJ7sHVM
32ZO6HOfQ8ypM7yuDno25gr66FWBE1FQWrm3aYulhCujUcctGsTELKRb9CRUx9Lf
dAX7ovMLopHURZg5C+l+qAdHSIuVYIkUeG6uiOsNKonOy2twFoV0CNQUY0+Jm9mu
TI2sWssKHHi30EwOKqgGwPJEfry6RkiPs7f6+cJt9gXJcyuHyz1wmNZdXCcWtWGU
cx8IXmuJbehohuG9w5C2r+Sh0w8uEZ/4XRXFcer81yvfBJsmuwbeMNJCQNos2U5z
BM9CPZIxXviZjELz2zJ3TjQAyVUDgMc9P2m+BE5zZVaqN5mUQrGVqXtm7QnUipuF
GXnMFcSxnI3WcScc1Q7fJr1roRqQ1fPpYj8hT4NjbXSr2M0XxJbzwzQJae2xHOGM
Kpq8zGK0AgjtO6I8OljG3UXGQei44HbHC1YQb/rLcgc4XdeNpRlfnNIJ5LnPX2+P
v0e5pQOdFl4Qq1l0Ik9neU8Iz6Ye+NWw0xUMKNek5mqHJtpdlFD2r4guwqlziWzd
r40PDQeEvl/QLBnn9KxDVWs1nxOgEBfxfhU/kvg4+iB7FcL4LcTrDSESlQzjUX32
Sx9GI82ZYHGvqWZMwDmvVRGCqLXGDE9AJHN6fqvpVu+2sAZOwfkXlbHta0BPYbZd
Sh7gIxr+YiNqB38klaLz+jjFoZskjNiA0de0HmKl8K3MGB5fC/GbGQUuQ9h5Ktav
1tBH9jvZlUcSkm4Y4QH+38X2YgxOrMCIFVZzYAL4nxllu7gfHZuAZtIOQcb+eWdm
ehlnSIvmsvwgPXYadnBQILhHn47H5p9wxeeBJYFnjnA1/QA/LYAwlgCd6A/WnMoe
gSIrb/SmYCucUZX3IFq01/qc05+XhA1D6VzTp94gnT2i8VsMFl5KGgY12xRWk/+B
s2CfcVLyEKl5OL6zswgCJhJZlPtB/uR2ds+vDBCbPHSfcfyDtRebdfudKWAT7lXW
H46pAVczcs9eUOiSJIhUf7vxIWuQboc72I678zWvMQIfZQrqzMwSQ73tAIn5keeP
O4joyPVMDI2VgQ8UqvIG+0YcFgF5NHhQ03smTypRCqE01DQ4QK3FCERXYnYcZO/3
bc+7Txladr/rt8jNo9BdRlUDC8HHvOSmdML0VAOfozZoeOXldm7sJ3JdfRsSsI4o
XvHVOcZco2EYeXVLswnIrs3/eo9nHpJOuhUVeLduo3DCdb8m7WzcguLXPez0YviV
ObwjlPOb2FgMWwpbSTRdXYix/ZezIIb++Fq9pmxz9J1CkwaNyX+FjwdrrUhMvylP
kbR4eh0qu5eyzjfKeCuPASrdfiIsP6Sbx/3lt5blGjSIZ/j/0D1Ev81TTRklH1Hw
gemN6dP+Ddm0GBsQW1WqrzzmrTsnMNNPiiHfTG0IIlYVR+tLgYoiDiF5ZG5x3WeA
pdP4cDLdYgsXifLW8nFDyOvZm51MNRNJ8UbREKou/ctZ7hSYdD//GrBgHLwEFLtp
socJjSnRbhZDTc0Gxz+lXorKGzPnFS1yddiNXvksY91d1Qx9eCx5iV5RsAVhaRF4
URu8kiz+uXLmgO8nZa6PEdNti0dNFvmszqgYRQ/Tb6acr3BIsDv9a+lV+mg4hDsf
5/vWux9EEZDyd6wr11XjIpIQ+BLU3j2+U0/KfF+YAKhSCPBKeMlN7oQrRbw9qbNz
gW4vWdZxm8gT1jSo1mLNFJ/58mUcDZJugvialOKtDneTnmMpqy3tlJ6bWpEgb9DI
a5i94cmEYt54vIg5BFy7nZJ+Lay3mTMzCfh6zI9mUqEFsA48Y2Su5/neFFpp72UB
owkfccT9/Y3sW+QIHHJ2kHum4qJNUt+GZq5znDoCHPa3lO0zGdr9q+u2cQoVnKn6
VwNxEwPHcfPg2VeJg9hFZs4oRG33utpCw8+wo72K0ivG2WSmeylCSVAhvEMY3DFJ
owbO5JS17wTJFmp7WGaRTydubS11DqIVx765kmH7vf1qkM812hvZ7Vyt4xEmPCY8
ruh6uugoEgRAIrQz6noTZXyeq+nZE3UjKnUojBIDZWYv5kq2USlPXm2XNQfZDZhS
X9kH5KlFxNyezbjl1kJqu34clDRjyRkQp21RAzb2ItPewcJG0JPHQqG42lj9sPt4
QhIBFv+HzxgqWgi8SK3bOLyL8LwjEwDPYeS0j7yXIbOLqSU0qu+jaU5Q4MaHv5Fg
l01Ilken6lwBt2Pz4Y1vH2VUH4Ii/QRZzJo4p0CK0uPTLBAUeji7bCTXRXMf1Kre
7spgCZqYhk+/z0iGLY9I/Q5p/iSTk1M15Z5V+u4sUh0rhirPLHGZ51RUWbs+8JYM
u47fYOTAlJlO6CXwmyFJjqIHuHnfh5uD2vyesYCMSdD8ySwkBfPcYTrMM34j91hB
D5k8CM3gpHcvmpNICWOhHEIZJqLctQPjoAwMBWwrWInJIvsEnXcmkFopaOrHqarO
OPLqkxmn6g0oGwzRLB5opVIR8DbmwG5ecgBYGhW6Ws0BP6CEpBoeRHMCWRoMmUQN
n964o54rkfxfmmGRM08avy32/lDK+b2ALoyoOI1YI+tYYhygBB7YX8uTzbOhRFoR
YlJEtRthSBwD1XQu0iYwxmpaEJ7GXSL8/T4Vip93XooVZNl8EkNUBfIPp1UMl/E6
g1aQTkggZt55XpbWjG3IOWDvrZGDy7+TdHQnI9sAh5WtuLHsHqYMf0bkQbue/TEX
V/Kt5hDoQlPj+rizF8TQC2DtvCcJj3woVKphJDZGLb47rVW/TbfSMzRs0x0RpNX7
YQwMquugu5TDU2x10gJahF/qEcFBCjRGT967P0zbu2zQt6xCSUfIhiJwBsmTZtmD
0biwk/RXLnio//KVQt4fXC6h672ECvW/68+hPEMWOKHfpO35uDD+2PX0QjlbC9v1
3rE5TUFQJnaRMdBIokudK13bWsiLIF1VXT/mf/XHuZ62BFtSyriZBNqWG2+l+pNN
9wIeqzBdMIiK1cnfN4bJpzB0ghaQCOTb0o9m5PaRxY/oyN5c1hn6Up+G7XdOBYlf
4MSIEw0u28SyDV7iBwCBkZED+kO5eeWenezvITtHVNfDksnJHdeG7dsbUWUqzn3j
mpuSwXbhBv8pED1Hrhkmfb3nHSp51rTvwywl7PUN6iDGsQxPcK2kqdCMNZRSK8QJ
Bjtes3B8IAl1aZWSNr/dFia38EJnZP8ajP2PGkwfNE4uCiPdubhxGsF95AzZCB5Z
uIb3/8vqF0TBtdX2CoqXrwzwkAatFw9cZwKgq+Gh1ldSwzTOvASopUyA0WM5sx3V
Xjb/nbhwZ2rrM6jCa7yJtxSxJiiocWwsDKaw4DHAvoEgrvf74cI4p5DuNa2A3l3Z
8YR8prEW+4GvPVTi4UMGtoV+PnF2TBHUHdZbRaqdRSJxaFaj2efpUz+tcfVzkay/
CdQ8HRXLC8TfVM9rpMud3wCIWQWkLAwcO8mH0kOuZkI1mW6oCqoiNI8qiu/RJNnI
AFlr+qkCZoc37VRFFO6A2UTtJYJ5vgp/bBLv9wWtS0z0pjHh/70f64DHzsEKSFfY
tomyME65fdGqIZlk7I9rtXIVDaz9S3uJJJPsBTvBgcEMEwaXNwVPwV1WDwR6pzIY
accmQYS3F5Oo0IHKyFDMSR1V/wen+6x1vkd5hXxXK4mC4bd9NT2r94xtdFokBHIq
kNyUAQT8FIo/bwoXBwZAqsh7s6U0Kew9zYEI17Ikc2GHCWfXngbCOOdH/mikTxMH
lmCUrRaHKe1inu6YVRmFH+BMnnAb5FvV/AtbvEjN9cU+l5trN25gDlTcHATXsK13
XR6IvLlZ9iusngkY98L8m/I8b+HbhDYa2FlZesrXgLGTwbEFQKnmu8Wj052KV38j
0grYTlgwRH3CrFrmyoMVD4/s9HB1GBJbyBrkrIw6FmkvmwziwSK/yXBpuB2eY9AZ
C4U+o07puPrW0y+kMUoiLKXCXmEToDKEIAU/Cl5TyOqzHU7rN7buyTSZ/L1iDNsC
zslAUrzvjR0XiULZ+l6OvoAfrTnQeh3CWSY/7ZVbM1tyxoDDQMXmxX8SXE7PbUsC
qgVMwni3RaoVxgnM0yacxfyK1T0taOq08yBwBBBW5Aaa5X30wCiiHWiqE4351W63
1jQCkd7IqGVgHmzoAMZE39vkPBO7tYgUGIlOqON4uTc8g0VH92KKZ62R1PXNZsno
cDtJ9e24K4DnqzGkzK6FjeOHTnv7eH9w2M7wcxuRREUewIMdQw0LKR+N9jcZQDpe
UeBKna8OunSflW+475pPCyG2S07O9qxK+uFxAYyNOzS0WPW3lyHBYo2IV4ZYxwEo
5zAZqUc5M/kSazoT+tdycC+uj0i7sAAW8IJHNuPkGZ1hFimsCca1p7OxXrbsduQR
NlH5EzARIheK41kG1QSwWqyTV8Y4u7s0ESxt505LgFA6nFw0myax165jeP25/DYz
tf0ZbtSX2V1xA8N5IsPzDonDppj3ZZbR3vzhD+TCSlD2wsZZJiBgp2D6iLrrVfuT
bwXhRO5JclvC1kUuuy8+ueShCqvSz1YE9xBMgbbyf/4iMzQdCaRTutWUXsASA/P9
STjoNIX9jmluRC/NvQ8OsyiH5gqriR0beF2mflG++C8XJOvJvMsje5KMhxjMdnom
AcVooQSH0Sin4qLvKA4aRjIH7RWKrsGwtj5pwHZEhEIUh0YCy5Ikx6Yl6t+wg3mA
b0zY0oFaYN2qba8Xv/f0Vl61K1al+5HT800ETOT3a0hGYEQOlvIBt72KjI0WG+lJ
a2z4rhZzl2SLIwJsRn38sgK0rtdYB8ubohf72NsPwUaUaB5IHQLsBFFDg8DVH0hb
IVEMKd0ZT79Er18+hfptT8Odt4eHxioEEdWYM8j9NURrIqeUDj8P6ea9xroxzJ4F
NaNmap/n4ec71kdWgp7fE6UI7p1ki0J7Z61rExmqnyC6Ms7VK6S2l2jChPDz3iUm
rMcaLsE499FT4SJ9Vb4NZc71oRzg7NYnfEMSL1Th5+rKcmt9Syl7pBcjRFF3rcny
d3M7/euMYeT5a9AHjnEsad0YG2wkXsTvZQ7PaT79OKTHm5xO/7Rm49PsgI4O8O69
gyI3xVcIwsYep152HP2sfaqwgrwpqH7PQa0lfRvIQ1GqCJ7r/TjjpvbpPEzOsl0m
E91tpiZefA6SpRuc6SJoCJKC1OjV/0T/uvy2Qnc5wC5jQk7JJGn7yEn4co/XIBUh
5+dtlBSKAp0NzQVoAjjVXbZS3o6qQEpfFXRkWKek4cWb5EiM/PXivialdUCOGDix
0VKhwjEDkFEY3LhZimLCakV5JgSTwYPKfp7AXuBcgOhmXAAxJ17v6wp1MUFqjU9C
G/ffG+1x0Ns/iUQEYbKNKEZssH0yKoVDosq7yY+zDvOBoRo0FwUc3mGV8WAOM1TV
EbD2CoRwowwVHNvPn1JjM5R53x6sd/V+XVjyBW7jrWptPC9vWMOYd7oq57AW2V3u
nzTTWPelHg9UZToyDhslL5Jf/hdYKhkS8KmGiOkk8pUMqygGdCfICB5BNKjfdiBj
CzmWpAB/d5hf8Me5t+WtTSs6LTNck+eLZe9ZI5+WioOiIxB2Q49awL4zP+pbGlbD
Aj36jjPdt1s5++hOQrkASD1tcc5zPo/fMwQaPJpUUuKaw6bvT2cr3O3+UydvI5uh
hvMgRnFxw1TrI3jk+zwMWSLfjRYDbMcoWCVWSok6kDXLlMz3EmqbLdQDLwvFnQnV
wcqmFybfD4glBXBz+RlAsnq68qmJ9itiiTsArllMVHZ+aOxmJ/LXu6E1dnJXkTU2
wVQIrixMd0XFVs7gX3eQJIof2h6IRiz4C7YBGpjOn4kr4styTiVImj7/D5ULvx40
3sTTymzaxutYRYh9Cx/dhZMIdamVuO9Rd0C9QkENodk+xkSKiLhjrTlx5f0mrhjP
1XWuyPX0EFXBLCChsKzwaruwAu3HX9nECd+H6i2k7Y1PCVyVBdQCFvPHLMg4vzpy
ozNzWJFuPirEdvoGNMCz/BSEZfyqPCVWe/Co+DXOKesZB3CeyxLA1BUHCGnCu0RZ
EqS50lTOKn34ZppYJlJRUPHQFdtJtRhHf54ZXp36+STv3aCAOdxZOe0G/HmCc2Sr
wmfYtS4gacdbge6cY9zfrv2RrlmdfIlyUI3UUplsncOPAF0sr6ID1W814BcfHccZ
ZDBWuPKl+XrIwfVSPtTV+J1/G6QlcHPNackbjLw44vGgUxU1sABIjac5jVnFpMbw
azTk9k5WFe/zQntdigKQN2LpA+IsoPR6Vq90SzeA8BxQKv1ApSIGGhW2W9s2KAFY
DvDbgBXJTQVibYvIbm2mhXzbgf5XEGU/2q9hpsl+SgcuBWb5/V+1B+Z/BEKAu26N
in36qKRciMQMu9nSKfSqgWiLa2nAH+bATKNqBkQPuSzVAcyCoxpFkq2Jz5JqZbrj
YUC2gZFDXna5J/qWjeRQr11e3M+MTCVf9e8RTCQbYe+MAg6Ea6aQyRTQxxk1Bid4
uTlQjFSrNWaYsvNDmbGPunG0Nbu+d+ecn4OZGZCHQI14ltLV/fXm4d6PoGDC7IpL
No9j7TvqnHYJ9b5CMIRaMt4t/8dwH0eXLz1RxJ8uvRjp4eDWhZGrh6rIfcFH17K8
LDeuxWFtFNaIMDTqo4C8c1/efTi6eYKobPDCFUZro7G7t5tNf2NXLRXIKIiM4hb1
z1eRD0y2i9KsKKu3Pv3tXt+3IJU7tmF7D19+BNZc+CbXzpXxV55xuSd1JGiJViOm
lDcZlkF+WMPGfySUNQsKwizm4xi/YG9DpKPgBS7AUmcV2wAVWVEdugXDgeD6+Kzt
MmQ8GxjPdE8xtU+y8UliaEZsd+pzJWskG3NOTVzlVIHJE07rmiTHLOueBHu/N/Qt
GLKKt5Rw5KqwwMpLfg+v3onxVmfMsIkcvLYm/6gk50+ohpHOOkth1CWVgCJ2uIBk
17NcEaTGhtlgDABK0wFqqOPr9Mr13QyY0bnkaihZnUvGRntJEttL5Cm+f8dm9K6X
lIsYbDZUwo+C+DkKMtgaXuVamtmeX/rJskkH4ycSsOYToLHr3WUaVtCPSWuQjZWr
UH5ZvbQ3qm/cOHFd5swj6LvukNFC5ebiNOlrbON5i3XCQmD15I752ApfnN6ProW4
pEjsW0PC0XPH/9nnwlk47UVSYSJ3F43+j6puxz7f2MJa/FPE9LUhreF8lULv+5Eg
GZ6v7PMyMVLQSt0Bin1n+os+4Z4NsPSMZha0zcur3+JAP8B8xHyFhTXn41lKt+Px
yUwYXG1W0dBBbSfWr5mFlgxr514ZrIQ4+xhxpVQqqYtVt0DTqMeSzd+1EBniecfY
AVc8EX/gCCeFRn8X4dahILofJdozBsAiCPCI4Bsr9yase7Sihw/9zVWYU3sxN/5R
b6OLylIcQH0+8M9ICFZBFzhT8a9DULMXZ2FpkiDny9WMnhdERvWdVDgtT0XheqtM
WkuKDT/umnrLtWkd8fjsCb4B7x4QtgE0n/p+Q7ZkDFAkpEmPavh5Q6VmYfxBUQn1
szByEodbtN9+9z8uXNYfzbdLpLhyr4bOWx8VaBmebNQ5F2h2LJBhHc2fFY+yLDx8
YtMwAaTgdCggDW6jff6WIGv6EF+ELWRrHhggKsw+VFHOcgvGVXgTsTmNm18yIs43
uolY3HgTrIbCzTbUD0yDht3T+H2T/mJsWxWZ2KLJhulioPpwGvKuycNvPv/2YF4d
/JWpYrIOmO+Qe+SIjE5QsXf+OsEu6k4I6Kn2yu72l+QuYIY2ybdNTo4ioJp/rO+c
LMC6QTzlCEE5aY75ZDtBmuXaS29vmwshKNgalzM9/zIKWtZ1/0VX8klXgM0rHjuU
UAkVV4Yq3Rcblem+7LFSzYYTCMlFyK8ebi2WScG7kSIQANLIw/+BtTYenHhqJU1f
901+YQ9RPzTbIXHCPEvlC1LziSKS+7aFVAVc5Uqj71c+4lXQIpIZHAzfNzPyzAe9
O03URnK46adnexZERpCnEl5pREUKztPqUn2zBaR2QaCEVyhczzN518Yo+gJteRCh
/0YMZBBpypJcT7HGy6KYD6ooSMxGL8SKBlmdGNlCrQpG8zhKDdZY3FeMNxxowkJD
UOmzG3biVfrneZEUw1IU27AMJZujzwTPqZXjSUKIjqiU97ZwMXPu4thPMJ1aq3Q+
COacUd9e/OCEYG1fWJJzeG+ljRoSyECac5dJ83rzDNKH/MOww1yi4/Ou7RDu9efw
yxeCQoiubpB9vEmolI2iugouUvQ8d6S6oIzQqGOVLqhRx2rt6kJjLeims96E2OzV
/Vyx7fksDXOHIzP+roMoxSf6FWVj/Uw2z6xW2tXslhwhmhaH5Gri/mAfpYeYrLLU
w7dXfcsqowlDv5A79TR1Vo38nylw1qHk9nNWOnwl9/x0LypNEBJYkkFgenf6bU+3
pP8Un8CjT1ywzGJJ+MT7SrCplFZyX9U8+Xbrn4bL5hCuHHo45H7JiUAfY2kp/oN3
qp1pfICxM1maONYwknpapdsNXQXHlcfDBT73GnMQqU4j0zQ3U2XQtPMn0E10Snwk
nHsfjNXuusEneEGFLjodrlH55UJN36PsVJ8xjFN6aHUQ+I3GJWhWDPGUnag24+qO
wAKC6T3iKppy+FINf+PSl7GCClth+kXSbxSX8RR/uuK114+Hi8P7owdON2UjnGi1
ZM/YSHy6WS+Z01wV2u3vDPCJZQv76pKtA0jLB5amnzyuI3AEHwYLQBljZTtCc1h5
kyStMsaegF9+QnLNeicaO4whvO8nEW6mpu+o3ubjtsIHW+WyQ4V8XFZMRLQgBg6G
eockqXAnWADsIXyEa94u8nVxgCVhd5qWu70MyPvy4AL0pp3fboxZeG13Im5QOEHi
rwWqKDnP0vfoQs2ZclFNKpvrq3LkjcGiOJnJoY/PiP55y9wXwwZ1eU2ZBgblEA+g
DmA4oRPEbPyMVT3dArS/KLvpL7YcAFQTnqonY/zAX+3jyb1pZvlTZgQjfNUi7Cgr
UqHZz+mhw/rGHP/UTRMO8gZotxRLyAtIDoMvMjM1ogP4hb7ZKtIf/PedmCucT0F9
69GegSxde2ajRNDbM1NG2Rdz+UeLYNc/aNBHJNmWjqgljsuqb/qbn0hA7Jy/euwa
r6HF1190oEDyscj1sXUcVEjg4QvgztSGcJ+DJqGoBjKHnKqjqnXQjwESUC+wcMzk
MKEXXeLw8mKf5nS9UvDGWV1Idnmthsg6ec9kn3qH0/GFTcGxScPbVL+0Wf6Ipq2i
NBpTUOSycr/+oy6JvKjhL1ryhfsfdkWOBGbA12yR0tbyoYg+3wEhYuUpLc0EJPlC
nvLsZo30Kei591M2RD3jyBBRXJdMA8nSnFVUS9RUv+/TXlEKVNUfvocnF60QPAIJ
CDYA1/KauXxTj/ylxMhOfIAutJXOBVG3OMoXGaFhdYkxIJBc3h4bI7k8kI1UKBa+
60mcWOKYW/MZonF03zQC5sgeu/3j8PzDql0dYSz+PYIPCNfoCXCdFiAu89vGr5Gu
gyAjP6Teg21E6Bq2fl/rN3PsyJwv5918ewfgPfMJjnRgI/6VaVqiZ2VJy7vNL6b4
2uHBGiS6E6OIWrrUjdVcrHpawgRq3AcSgAFRTee7j7b5ajzqjRlexT+hxeb/AiEV
L8tKMSPfr3NL76ubW7pcATRxNaGumD6pl2gyM6DseEP+v1Xp2y/FUg9B9nHlWuuq
rlRb+F/ZywFBm8jGbMWGcOer85NRR+FIkHDXxP5AkS/oBSeG+vdznTLAb3ioqvgE
CKQNi6idE6SbCGwo1Wak20ZIcBqJSQtH9XECBa+jxzrt13jTNmw1+uOEvFECon/S
nDbv6EA0WGGV6GR/prGH1/LHKFmynC0KyCQXnZ+I/yKfbLTsn/zWe8OybxfBfC4B
E1DZTJKI6Oj4o7JdryItBuOokKyvFBnus/iuzhAaOnwsAwM1pVixzk5+0J3qJyfr
CsTaWSdG1nc/Ja4oo7uy2Dx+YLzQVpuBBwa5Mh17tf2dOX8qdxmtNbNtFdQFqbc/
gGqCGKBPYwwKgYyGcysVGfwVXpNhQMZ7Qwr/IyISca+JgyO1x1ytpmpeNvCvJPYL
x0v/0QZ2A+LH8mSXTLhzwe3S+S86fj7hh8exYEmAghyVV+WKIeOIhBCHzX9xBVAU
2dpVp0vLO91C+4lO6KHP4B+pmOUerXV+BEHSHU4tO1Gi44n663J9V+bgH+hh7j1H
l9eqJ7sh4u0wxE/8XvnrNZiGinY9IuwxW/Wg/Gc7ZfB1GYS7nXR1negnGXmWT68b
5xBfeBmLVLYJp3aHnTTvLhhi4v0WQ5Qp0ACL4xsL8HJznJG/pTaoPSrU78vjJfDF
ZfQYuNVzbMZvrEn85RbBjxCx9iQoGlJDCP410d7gUHqT3FrdRiHE8ItrJrQfsSko
TTU3LgSb3MrKV1kDx4C7UeWpYA0p5IhK41AnNVtAxnNdzPGlE2mE/BmHAiSvbE3W
D04wNdEHkXGIY4YcbNEEI4kX3ONGram6+vOJXXvYt/hPWS7rs3S5ZX0nF//0Znzf
Lv2OoQx52uL3eppp6moXV9qAaXcE1ma/0KT+klfYwswr+RTqjz2HsiEujTnlywvx
LdkDjQZyImvlmF82KRZYlGI+chT7nLqnS7yJo4iM5vdqj8j0M3lEwfrUtHEGvf2S
buqW0u/0QPrzb6TiA9j0TmoXiWN6CZgOJSX6hMetmCdXk4KWw912W4p5ANROK+09
GQP9JiwQuIMRltWb5EjoFTHyrVmCfYIQZwuiv9qy+jbfwStyefujiGoJduBJGiAD
RJpy1ct5WkHubbokUMCn3DmRErwr6zx1vh2JzVepwazDHjPIR8Ux7ZmGojDGx510
lYK5w74jPfr1vUrCtqgFs/AIgg9XJJdrFAQDWjQkzV8uPajDyRTQ5Lszpg5DMLMd
NfRDFIfUgT1Ro1GoR7dMdqoPxKmpo1jkeAnRlDQjkVKZL4mWiXWZPcWyyqXH0nVP
fP8T6MenK+1w61HjC91V/Xgu68ONTL+07SW+2vdL+YhUxwkZLvhRCxfMn0g44aPN
qchSE81jPi25pRIwH9mUfCmfIDmdCZbJKM/iYukaG+TqIpTeis9MFDuArgkIS/qv
nLnXPDJ2PGQUR7xcnbnL9JIUZKLw0GhYb/JCvwPaTYzGBdo/ZXKEPVIqf9SG5kdc
FBMulxVd0xCnuN0X8tssJ+AjTQUGZ79W0Oy3Mmk4NWDAO9SdaWoRhF1lnvFBB88J
42CtaNRCeLWiph7IxeURvvOKpw1nLjELsLSaf78KYTIdbgkRM+yZkXWxjjPEnBFf
u3uc8YgQzDMBoVsuLI5j1m5HR9E0sYoDuClCxEhszHUJMjy/Tz71AdEJpOTPD3Dr
CIMXQfAipbwuPraFJBCz/Pmao08LoWR/mxGt6S+72GSsOIURSxWcrzaAhsTjPVsu
Cmqmra7BX3fQDcBNPhk8KcKJ9LM85U32/ORW6QM9zX6peQwQthOb3D5pWcmInqtZ
2bQ2B/Jz4wlcm7kTevvsKO2dAajJjlqWHnl1Jj7qDQk94F3cFyZpXxPIepiJiQak
rZZSabnykIqnoDTRaiz5mR1fUSJmxnKOIYOWteH008jOqk012Orb8w1QkG7ELbBt
t+Mek7OhxLg2pDT0c27r+OiGGOPbgxFP+Q+dO6FCdCIF6s9hXeLQvjho6n+D2rgV
TiOCfUmnGkreOCrXtZFcG8wc1U8AjnHpfy7NMzY3ivGqJEb/ngbdwHFFnpw2ol8d
OQrp+KazbWQiYxiZUi+lLmZPGHk2DRK4o3oZ5ukNpZmpPtsMEbD/K/XeTEeiSGr2
Zf9C7guXvJlzSg4tUdIAZyytfHKyZVVe3QjQxo/mJXBhAmCr51JKkwvmLfVdAf/r
+JwHtu7t/KgRKbkF5VTKCnloYj/dsKRT6gxPnXcgeoOBT3cIdbyXqd40EeIm7j0x
BPHvmORVAqmSZo64oyV/derG0ngN4ZMAssbSHNn3uaDYMCBMnwSyBS7hDkImYbj6
MQnYB6JndyYqk+IhsFxBrBIOAeK4wYiJF8XG5v5CqF14OR/6dK0KMLrcyDmtkC/o
U9VjQ6Rzj0E6ZTfbagCidubIcMi6bwPR1ih/BpN4aYVpOUigFdEjdNIKLoutQbFS
AHHYYWEWk8dZRq/YSanW/i26V3DrrWxE2yZC1Ud17m0xmKYrMisWrwM9GBxyTRwd
L0MkOIPkNhwL87ytkGAfWX/gT7iCZyzdy5lr4ecnphwXPqqM93rX/b8svtOLIoQa
6mqiLehhLI5ecFxWFF1msH3bMPJsX/cG43WvIonv2CAisL+g1DWcAYu49UT+VWLk
THpL0Gppw0Y67lO5evepfe5D+KdBh9nbCMMXY8B96aKQMcn5SSjKK2QEWKpQSiOw
/bTOdSoXa1pqRDrO76sCKtNb/ItGFXU2mdWFJkG9zbsNoRtAuEKxCbnJmV17WLeS
YOl0GOc7LrLx3OrF1h0A6yxtY/6dLRYYrqI4xKAMhWL7zadQbDkM/k4vsfUQcMdI
gr6+t7jk4As8njjCBDo1NK+Et3MyCq591mFF4uJzmWgxv59nsIH3EfM8c/7G7ka5
7hgclGNyfVu/F6nH8ExYbBysPb7hjQhJX6B+z9B2/ttmc/8xV2+2gZWDv2rqfpKl
fiPHjevb9TaldnJEMu6Lo+An/6xo64tdm3EU47ZTsNcqoGOYj927WRPX2JigH/R9
dwsLkwF001L5c6qDkSWQJI/mTzFRLe5MEcxqAONjtC2tAuNZxHGtHYmbiSEZwa+1
JveOssE/WPWXDd7KaAR9ciN0cYYx94xnR9gXgST6BFGP8Hci1beawGDKeJYzPEBa
AU/fEEEPdcNc4oHAlozXUNP6KCqTE/66mU2z8QAJvdb7t4G5jEttBzbpOlkiiTTW
DgGS1enq7AJEba8zuUzxnyhdD1AVXIcre5K48cAO9YbXIp2F9DUf/B16efo1XfFu
rAuOdDB9h1c/ZoTzIN1HgD7risEWvD1jPRoPwQ5RtqyKH2Be3OZ2Nf5/AtnsK6g4
tcGN0PlPyOppTs3ApKN9uS3F+jzsyFibBi/JvXBwZ9TEKdarAJNh6rvthXr4joQ6
8UUwXPCmHHXxtVyqds1L9p0Dx1HnqHA++1XSSJbNmEXrFVhbPQCjJB3Zqf3l4ZCn
bE3dH/dNOUUrtlxGY/LJ2Jg5j7LPfIimK7Is8FNHGXXvJbmdlu87ucxFAMmn2h6M
/Z9RcH7IsiYeK8BJJkj41LcNY6JQf9x8InFdsYlmENfVAjw4cOV2Ez5t6EcZqT7P
wr0BDiDg2f3vucG1xKa8imyTY6yrZK2GnljtqTa3gds2FrgBG6064l8am6chMDX7
Cwo1q6DhhLPoKFUdWQ1AQkGS5D5VOn+ZmTDi5gUd5RieVkxPvk3gq+8Pq4A8QLhS
d/tBNZ/Lec5nokcV7ziQ5dHHYwDCsnqMUS7BFGuaMpi9aAUFyArwbXfCerrFR1QE
EXd+xjPnTlIMc9K/2tSN2Np8hV5jZzQbioGINvQxOuintTbRTWmttvQgB7ZQp8kG
lzjD2OUIHvzyNTR39VSeH1SfVOtalhuM/vJWLWWDoq/eG/WjnWle9VOpybGWHdfX
Mip8tO9IP9Zvpkmo3lcBtmBJuNfOLQmPko/IioR//+l04WGb+KekfyZQ7D2wTswU
kqcvVhyD26gsAsLs408aiDxaw3176UrswPuMWMD8sxapLq0T/ACRQtGh5BTmm9Kz
4wv3adVbMntmEypk2mAiLMbbAgXAFYbLBhJyfKC4Mlq/PQ0tbErY4nV5jfrQL8MB
dbfkv+mrFRBl5v2nhAw8zJJJ54JMffhRtXhG3KdQWk7VZukzip1X1Ex8yp7b8uzs
GfmyXMLz5+RuCZ4tAc/3eNZNQVQUlKBQKuVqnPork0r74d1c9qEXSIxCESRkze5t
wZYRn2wha7J2dYO4Vtrz5c0AqnFy8uHt6RKKjosxyJW2FcsYh3bFnHwNiglZRNbq
kw+r7AUrNvAEwpz1V8DPra11/iEVEndMPmuo2XMzaq7jv3py8MLGXStK3W9Z/lYi
m1AERe9WUvNqKXZsIxrKLEKcUGjKOW2UvtRRHwRYsCGh4jumW/RAuztu222UghVV
QmzrdmE0omEwyiw487gDVMRguUQzSrWO7zDV0a735ebegyQ574f7S+ocI8PZweOm
9Un2qG28aleEMR6zxCdilD/b3ir+jkKowUr1/CqUcVQ5hUw/Mx22u7S4IPLf8KtD
CmbMTw9BHgp6TVAI3jo0A1Vp9Wfoz3nsNU+dKZ3iwioKgguW+yV18nK/NOWZ3zII
HwDCv0e6KAbUE4sWUZcdWX1Q9+gqET1+Nm2IluLGOnfCVdFLm+qQNfjtN7U5Zl2T
I+s2LRebLnmKY4PIvPoUj4MC6e5cpCh9iXduCwGOHlnD6HpeTVNQcaMSXcCvKher
+sIlJ6dNwLKmKU5QrPNYBsxPZQmQ2WyiNq9y3vCE8sx4D6935Ro1dPi4Zu38iQCM
iQZuFuLRmVAcmyOs5dTxbBVPIkAqPm5ibWhptdl0WZtlcAVsEEWI8obwJmn0DFwC
CdVEXlHAbjyvvA84S8rI+8gyykjYM+QGTiz7xgaGTprjUEOW8YA7H32tkl8WPglC
whJDiDIBgGPWZJAYYYLt6Nm9glpEA+ATli3Soz2GBytFrcNI77j+PcKT0TLTGLZm
cnFLiqxhtErgQ83r7pXDW4f23V7l+5s1pZekbfYGZzCGZRd61qhk2Y42HAL5nfcm
HpjzJWqJKCwSRBXGXofDvqkeXivuzpvoW1ws+HIlcAQiGq16Ok3/UERen/aM7Zy6
3Zg+i53J0pigaF7aRS667JcY/0aYEO2EmX6lwCsZcXrQsKOzl9suNyx1MQHBTS6I
GOflBkXsaO11B/cxNHtikj/0bmjN/CUpf0kC+K4+YaxmthRo7kZ7HnDjS2NvdSD5
MdzY33z3IRV2RCW7W7sfzpCnnQfSe7o7IuZG+pmJOQa9DBtCyouD0fnPMW9oCLyQ
yY143k6DP9RgobNbHFrND5Q/85yKqBJ5Yzp9MjwU8VQt2GZwn7Z4TD1Em+LaMM7A
hSLnsz6JGwG9Et9FVca/8GKLAr1RAiyj/yCTjyY/XERfMhw8ix6ngJH9c8k/arDH
TKbjfDSAeBLTJeGvVcEiILoNGHTBlr0mteZFYT0FNGO0WmyQF/ymp3osiiLhjAao
6Dlssiut6lLMcPw9bUIcsUOxYbLEeVwiq6x8C1c/CNhr+rrm5Z9ATATZ+iIVtb6U
Wsy0sFzNup+wlcBoY1FmjsBzHzc9TjaIBVoX23HAhIB1Lkb/3ZL9mkRkFq/jPfgY
CHVeD2h2vKU6l0uW5rDp3Qip4jVzWTidffrl5TwdFHFb3IRz1MqANz7pKoJg6gHh
fv16ufmSzFtGKLcr9Jjw61CXmIbl1NkAy10VwGnnM04oDNuP6T3+dX0F50BiW/Mp
viGVAIGCw+xdHeiAygzHIc9IJwCX21NfByvoMXq9I6cXpUumcvyk4/jHjBlr2hDD
TYpdSyf2Yy3+CSvQVmSMvkQnfNuoIe8DIDCFJCFGuSIMYhFC+9oIJ3hVv9Z5cMgx
TpknobGfiU50XzOb2AL+daU4lJ4rX763YmwAxn6EhSz//jH8c8KNdWVblbjVFPOx
6hS/Q6NOLRDw2WzX4H8XFh+wL6OFAanR3GADXVyIXZ9AGOhSEhS3GHEtub19rW9k
KcFG9odXTqIMLv4NKTaqUemcu6+iz0SRSXyt0nNhLAvQyOZfHcfaGgLsUGkvhpKv
F/Gi9TsLmc3p16mXm4hkGazfqsNmE4fqVH9juP82YEpLY1CoY/ZMvJAFiwFHoGJ5
H0tyFT6qE0kckR9TfCv1JDnWSoB9Ot2lm+kA4+8H1UjKgW1mtaFVHKY4QXkjG1we
nGo2i2azXVqx0/4nF9f0WXH8dDyPrk2QLDK69gFxBd595X6TfiYGyIcJrSJ7+u63
HrG3Tv9oGLmhLNIRjNTk375ZudHYnCBaoo2DBFKXb3pxtD2BI86cgb32BDZBF4C9
66YY8ZE0wJbZd1aLAP4v5W5QImts4AaVa81Jn4DR9eg5mfX7UY/URp57C3iVrFM+
hMWVM4sQj+DmykpGil4pl1DV2ZXFWecOiZp7/eEirqhJOP2XyYelB490k1S/reBk
+fe+XmVDr1528vWf6nYrq5tjLBCtAtEunMHmNAfaIGqzKS/TVUDpU2x+hS6UWf1x
tTav4PPyv5R2WAxX5RfT3OmpVAa9Iuafnu/U/EK0gtjE2y3IT+eLV7gWpxYbmWxs
lvX94ISmkLOdJWa+OPkUvcBSo5nnNMcJ2xUv0o2IcNt178kaZsDG9vWY2HYpQ91o
fxBAxI6SbKB0dfGe5jOoa4YPr/CwovMh0ha6Nq57eeHmaWyyGXiZ25DyXbNon+Vx
htnsmPucLHE94g9hS233DjWEvJ9WLNQJRF1W6LlcGfy/84i74ybPi3QRFWQSi5VL
8fwUeYDQCi2fHAO0h5qYWosERm7ItfBOZ/lIV8v3xaC+HayK0Binu5MaJZxVZCFj
wZPpIBS/9Y7/1FBQKFIha3GgKywiZ3ntiup3zt+gCXpthEYjb8SShPxDFGwoPJa9
oZur6hAPyNGECxEZSZwNiCb55CR60tRFMvCZ/Yb1VNlIsNHeqsiIRFvjJGT6o8qV
3D/0kRqts3ngS+rhhnsiO9LkGGlr7TFAU/IDX1fcxiXqF7E6rD2qCQiQkFElPnkR
R7xTXrzV0SNte0jla6KdqKimF470CGlXh639DvBnPkkgVTQYgZzw3k6IV+S92pPz
oQ9E+mtCQ0oUkmHy51IWEmjP3Tjj7r5cjQwyWGMqI032C71evox+x5Senhc7G4fA
XG1ngrnmw/Q1dJNXfa+UblSl8NtuLBNMopDFLb+Q2iU2gh1uXNdZcIZmdqnY9PTP
rwfVtkINuDmiFn1J3RBVE9xCsF4x74KPksVSzGy9IbuTd2o30/6Ha/oR9INgBa01
JY42WYL+GGRBAkUEZ81zKETBLvrxmMUzIe6RASvlnhEjQhEfVwRVnela+zZcc17N
GXtTCiPap88y7btBeGjsIPzGv967luSL4AT3Yf1ENwYv5K59m2BRVb0osBTiebWr
captwu11g6lXKcLHH/J8InVsMO2Q1U2CLptdHi342A7OvWzcR9ThHG3suM1OezPX
iaJYIoOdVfy6fP5mvU9ai07ccT9CMNLDeeOfXwAOk22Yz+IzcoMS4wo0nGE5Bb1i
pUam/4By2ell6HWjctF+cAC/k95T2dqZWgh/s8np7Sr6l+owd59X1hWJPZJEwawp
Vh/A8SDQ/VGKjy7h8nD508g8qRW6xHpZ9VbihcickjHXImTXFtJNibnRRLyjH5lR
dZJapArnVhLppa0QB7rxJAU2qRg3Z4rnJHeeXC/KtXNWl3ZZdn/z/+eJF6BWDeWG
s+bLergZR0CaU/H5EPpyrQzTMBqlm5uMVucWE8zTaW+1cmhAnaq+nNHMppQYp/C2
pR3xRI7YQRJN9ffW9vAs4qcrUsmj/7owtNxU1J5CjmdQoZsnRPqH7G2AqkybpK3f
LFmpgM0+Htg+IUE5V/R2X6arwu5Ztgp+Gchryl0Yy5yWsGRD2y+3GLQfzNo/q+Re
7vwBVH8vpF9uhpsQv1SbStIbVfOzgiSS3sIAqx6eSvH6HIKpEk2Mg7hvZDyebG96
/BwM+hlq93STp4FIk9zLfJwlqMLnwkoW90jLFkLx1eDHY2XqYZJX9CeN5SF+3lve
8TyJdiFh+0ZxnDgUqmbcot6meIaaPIpE2Xk3Uw4FUzUpvvkU1o9ZbS/6jwACbKNZ
jcA/lhqHBB43/7Kcx6gGOlcXc4vgx5OU9oO2DBaBm+LpCf4tU/G2LQg8Dc5Vumy2
1C0RFG5J92E+W/eMhaRA5B1n2u3ikaFEZXrX0qFXtHyFMT+L9YEmj/PLS6XPWxjl
wvFkz7WTOZloRC4EXhQOHwTY89KqcbdQBDyYBzNiC169pLc5XNows7ZQoXHgPn2W
sJEGMR7v7sH3zHQT3W6okDfSB3t3pypqgnSCTueLlRFr2ejgMF+ub0LYs8xpD++p
tJ28w+dFKF3aWGlTOTLJirdLClVJywB8vrkPbTGiGPtth6Z3F5EqGcC7fr7kqJew
BfvuNWgTf46LTmW3gXzi8qmyxehC66WXgeYA7SGVHOqWGWhwYHrOx3RXI3NMoofj
Su+MeBwxi+B7kAgeYfCUoqh7Mb9XGTjlMgUTIkI0yFtydtUQxZtfFk7bsM/OAev2
bm12HM7PmJWvjrkN+ieLjEmwQcEj7IVQBOVgMhYJow+Jf5RjE14aMrScmr6NP44F
ECZM8ytkKq+v9Bm5hXeShzx0Yu9fSaM2WEVMR/36tErQtKoTGpREZA/k3Fx8FlLR
jJdLn6Ki3aYp7L8rm3vA7rSq/hcwh/iwpH358FdxQEEWb+Cs3V5YNW0RiX11gwUQ
9TTpSbz7NbFJBWbvrFjfe//6CdoZHK74N5oLgGLiPCe/Bt/Y2H/ueIEIvh/WNB8t
0gVpBdKbo/38Dqn4fezehjkPiQfdmOt50LHPIQaLmNaT91KdtYvObEqRndOtDNCw
xmS2v+LpJxkC7P8ZQL+M/w+Xw79WPYTNJvII7LpiWVkiOYzpbUxAjoXQIFj8bQ7V
9mVvvKIWGELlNievgXYFfQcwgGYW2C5VEdL8+wExtUuUQNwnyZb4PplxVMs1tzfg
FKlQsFSuxZ2ORphUZgsXnnEwIDQwWGZizft0SKrBinEuAI4j4btFVEHPdivk/5JE
hhRZzYdecsaB0aDEf5he8uEACJZjjhg5UDGxCkvmW/QuVutdmiI93nPBxxf8grV4
2qKUe76J+L7rQS+lrRcI+lRW94+gP19QFTqTsDSGzkkNanxMJiiIbXgrXLKt7cye
BWX37+EjuY+5FhESN0jrULIxCF8oRZLaFk35PmUQSuKpumY9bk55vjx5KgGs0wvt
QfAQ03/fc1+sLn86A2WcLGmcAQiiI5WCZyZ82lZFdMX5uElJTLr+EuhnYYANyu2Y
KJUazvTUQvIc9bN/8sGIYIdI4ZQ5ZSo2cUAGYIa49c433cLLZlkr2Y5aiHK1vKq2
MGUIJgK8cGHRT5srYd8KEZkqZTZcODCZMJbAi9zpaGHLfj2Z4FdFBuvQJgXuVI6K
KsguxKczj3MUI0pn7vKMx4vvnIT6STdHZbCboCtaSQOiFG6Xn7qvQAPOc53Pt6U7
eIxCYnQ/rDu70Gjj5lBci8pJvj34/2igusGdmPPmsmptMzeVkZ1kCSzDG6BRnBgV
AZryAd//8+r9mvdrd3o/j1twAFNFQVyyITA2EG//c9mTYhlEODiXvWZthoCU/U3Z
8OIfchX2Wbe2EGnYIRI2RAxWpoeX9GV2aLQGAN5x7Wp9Op7ykhL2rRaJJq69YG64
dtoeKMmym6v7TVjaOnpaA0s88Ak1s2nNGEwde1Sn4rr/0sSaBIjAP/D1r7AKFKHO
qoP/M9Kll5RMXkrrLqjYTqp94/O+8GXqkNssR84HzP78DetKqZ0V5xxw+YoR9bmw
gizAhxE0B++uJBV8yrS0sN9npS4HIxxIN8KCBiFWowysmYQAkF0Db0cHXrlhraXR
ajiZvfDee2BupdnG7ExzY42YH8tNXs4pT2cZBf5/JP/sdad92xZghNE/GWe/mlec
/0jTgqKgmUNDO1lOZDcWml4P9V0J8fBRqA1zLTak0K52wjdzYtZQOLdbf+UA+cyJ
Q3dTXXyiGpTLvKLj28ap/esQKR90XSsa7NxB1vlTNRzSNTTIOQpY5jihnOGlTLvk
uZSKddZBYrIW2pCCxpPHY5Od005trIadR+Z+xZKzYMnOiNt1XxU6k5skExsmP0ws
NxaUv1L9v3Lwbkz1Ozs2/PhCjHs2Aq9a68IGff8PcvUWXDH6Tc64g+I2RDsOwgPL
6Ow9yhmXr6EAt7bQbLgX98lJVALoAgBnxB/0cdU+ndjBR8+AznUoVXNOwTgytQO/
Oj7fl5Z8thJFcGx5UO1vulOZM3vaLvzgtArUaKhcdv+/Q/4rJHgPWcc+Yv4IzWoA
SY884ah/J07X1AmaXXFLzl+nKd4E2PnpjOQgBRGDVCIJ7RmE7x2Aedyl5dTKpV32
+335f0DW27xdxgfuPEwAgeKgCTsrVgZ45hwOCxzfeuq6SDcPUdnYw/Is2G9US6Zp
RfOggdIYCkx+nsx9485hIblP1z937WpxxeSXii/fGDt0FD8gKb0p4Dd/RTNnGhc8
NC/SOitJFULcsmI/XqUrchitYzXhvpy1lTjAxZ9Llh5be83SJ/91azBbV9BBua+D
ncN/2+IOHtmrgONifU1QfFoprQHMjVjA7by83xQ81smK9AAVfIAU7hQq9uKcJJfT
Cp4LkIvJ3JsUgNhqNBmXAIp0O2IHfwOXmkLw8B5yM/gecWZoYsnYOqIFdgk5Znge
bKSxRmNn+eAzeZzAsv4lfV7e7O5QUBx4wBiqiJnvE+miP06eotgO9lVx5/wLaApQ
seez7OXVMNGubBVgAOM8/Om2Hxxr/zrMft2zmv93IEoWTR2+ywZg+SY51lz0Z8lm
C9FAqiVkpCh5VO/Wlb7rB2TQaiVTBUNeDFjlKCwYBhfxbvbShtAYeTnX6NJNTHOA
kpa2GY7lQvvlXLmSDlHU6cj08ODuT8uFQWFqILT7E1nq93aObRN9FlKZ3gmSnm11
E3f8exuBCuHelKV3kHTxBslqX89zarHpr1UhkxxqwmH1geooKzNbDhgYV8DRrcBr
Z1tJw5x8z8VDAfSIxOX10fWKqcoIHex8GE87NalUsH373VxBHBEauBxC28AfNqg8
gEMryt4p7sK6pnXBZHZDy0v9PJD8Gviz8KnqCVf0JPyfau0BByEZyru6CxUNWD+l
UpHA3n+0GAMW9PkAfK9CfzQflp+3F5zgjco7Fh2CWfH0Y4VwIOEE3hEzn9zHzUnZ
4LtkswdB3oPvd8fW2/e/8NpHgmvWm4iGpgnLkaQUCqLIb37LGaPDEd1u2Z1N5cLf
4qndBTV9M3PP7/6+0DxuIRWxDXbEzs15SjVKeJFtjTJWJ02MEYKsNybb5By/ygk9
GqqKjFyih4j6upTKw74LxfbC4htYQPt/ShXNFSiLCXE+JzmEwwmI0fXAgCCbuJxn
7P/0ORvQuv0lNyzx3MrJkTDM9VlmMetKhF55/XsNHx792B1728utx+mRtY7aBtnu
iFgFEtxIkOtZW0NO9G4iS04kXdZVpEr69ouZnRkOTsZZEmO0/0M0HjIpEVCr7K46
9fFhfndv8WT0Qd0FD4qQKBP4GB+B6tmjkZ/2WnnIWpWY46koq/EV97M0SwigNmmc
USfgS71OXFC3o93czfQwWRE5KXOcQDJLLQq7TwXsx/NsMamWwEHMzt+NSMFlDVDH
CCaJi0nOY/btYqnuXP0cJpU5Qp8vZqfpNed1HlZQ9l8ZvRGWs7Il/KBSJ//W8Uxp
3p7iEpK7GT6O+PSmz68uuPu6As9dYQQyVUiD48Mjus+JMkhhE326485giMrbTSQ4
ZmVnAdbr3pa9X2ANogiPO8wJBsjlz9e3QcMDYgUiRdsUxB83zQ75Rywy4193SSc/
OJUY0PbEw0xC1LZQIkahUp30RZugBtZZFQxdrIivXZr4ZaRpmzrxtAiGBPmHPlXc
yDwvwPyC8CNSxSlhxbDkSu8kIRGNg2J/Nu6DBKkvoaFabrV2Zuw7Mv5HhtFpRJdw
GrKxsMqKjni5ap0hu6jRCwQzpGsFrRcXBXhkDG9TlIFJSiF8GwIy+Griangqu0fg
7ePEXjLYKXwaY6O++3p1178H1smT4AAy9Wi2ybx5PtpML0QHtZcHEkx/Xs/VSR2j
vymTMwo+nMrLRkZRrxfZ8+15maDLHCWQLFY71Eq+MsB0uZj5Odd3hws2dsmyLZX1
qlQnc4bW5r09onEvR8BM8WjKiIsN0bsLJDoCwstWs86yObCUIzY8Q8eArYH4zuf4
GO7rmU+P5Pnl5uXMxiHVdK7RbsunVuRUswX/Aq4MvS+jSpAyanXWdE+SRBB1+J1w
wPWld+Vu2xK8tv+3cT0N2qr20GMXPl3WTgnIiuAU9pJx3/2Deogqufc4vjOg5BOI
axR+tydL9q0UKYcwxS5rd69525h2+AwTxwZMxWZ+kiQgukV1q7692/SpfZG+FvTD
1HFpMQrfjCiYnrVTVbSMoMY5UeziYw3fpgfVtqFBr//KZ6ATfbQUHfwlrE9lNUS4
zxr+pyExFvHE7ph4Z8o+0ddWu7dIdtcOjOXMbM80bF65Zk/RFK9yaMMXqJ4G6VxX
kIriTVwKSh3Kw+ULNY8voRmma7zfriwezKSpQjYdpUWqRGkYOx8r9ddKaFiKjBfX
Hq1DCF7tHjmHmLONeppCJulkQWe+ND5n4o1Vnlgk577rV3jV3K9pAKlqng7t4tx/
5kyg2D7ZZuI+O0soJoy88HvOJDtOPFgIIfzuU+KGWmvaxjIGxCymLwm/mAHclT5p
K76Dw/cyyMBVpMkfU95iQYv4MCOY2V9YBdhBDdh/tLM3rzcNBqasGLZdLCTOSOXc
CU2rfanBJIACMe8RjcE6jakYg8jpORZRherWCrXX/Tmc38juSHp1PpT4FDBirvQR
bhPAwiHOGC5Uq9I6ChZ+NTbVwmY0N+4GH92kXvvxFyMPM/RtDHq8CilXXoIzngfd
sDYlB54KAqIhH9KB8pw2pOL6UYBeqVx0FSMjb5MEBbfay8V9CYKQx7gY1xBGZhSc
hrmMGIVdTMsiamZKVJYC573KC/38JNdXT5NfLHv/hQVczr6wJ4Tr4binhoGxU/mW
aoryj99sgqyoAoJih/ENXTCX2jplekDlKqHNUG0PpIVy0OoyIXwNxG3+dgNn0TCM
tGIajPNljgryBtPqnDpz/cbCfEY7p1ob5q+pFfGFtL9NGt/Mi+cj0FRylDepjl7p
5UEkb16L6sj1ies9/TNiRuSyL0zHMX5eHi7C6bK9GAI/Ui9ttkNL2wxO8bYlqbaw
nn4bxWYidJjjv3IcJo/UEgCxjRLWK+av40VB6i8r8r9aJHbDjLw4GXJMVKap1OYa
TluQn8b+RNnlkklrGsgzqhJcoqx/MvsoVmSvbmshty5Xqs9tVlYm8diRpFwhN11N
LEoLGt1F4Sr5GJxJOGlAP08hL1Y7JMNXwb4M3NhNlS3d/YVOXydAEUhHKmi7CKYB
I6v+YsCHqHW5ZplDKVh33kR+5A0+lLnFuCUo10HP8/JLz0MTH0+GL7CZRD9KVyzp
g3M7f/iTGrMqxKAH/5M0+yfaksW4YfymcWlhplOUp8f8UfojLAh3EzZzeeW1IaZa
elnLc1KWPGmocDXCi8fYL5qROp9XxOgfgqLaX92gwgrw/8ryYCS6lm6QyeMk3nB1
Dh1BVIyuCwtG6DitvicRfrkUcz/1W5mupGHyVS2nF/hDI/mm/48Mv7zMzrVqeKof
h+O4Y3ssOmqs2skjZxbt5sRz/uHOfcm06KIU6TJYPAk3NUhWw4zD2lulzhc1pr6s
88XFVnwYgn6/dWtqgH2WkHzy4KRGvxTcoriya8K3ONtNwuVGSDhU4VimrkQ6Dk89
uZwWhuaclh1odhCnfaz3ODvtvwIT9cFGN85dS90l0st1xhB8Bqz9RzAugwq5a4ZR
76veg5LffHSPZCbKD3H9Rq3qWNCtHIgboIMwXFR00UbU3rc/DIUP/rq88o0GykAM
TDVYeXJGfckFrsvRVIq+7iLsg9s3eq65r4478yBO7Pmlfz+H0WLel80dZsCuygKj
76wWqFSH7S4CDNgl+G+LCoQHsrQoahpjj04QnwiVIjQhMR7DofPkEcqwED0K6DYD
m6c4o9udDZ6PqAQ28s8rV8Twjn+sT1QQenUXPChF+NbXlBMo7L/otA+VrexNTsPd
lVUCm9CbK4cU8E5CIQVOiABpELjXhq0fhFszcmv0V5qFT0aXC38T2rl+i8OfilH6
SVhKXWOfykQmPT88DsO7Q4nghQYTuRzXunv15r1iKUeKFx5NF5Zs5I7mDmG+hWzY
IstsH1aoF/d4+DQJMR5aS3N+h+pC6udZI9oQ7tMvoOzB4iPbDGCsUAvQUFV1WP1W
TSawEHQbsX9qN/AfPlKuBMeq+vRl3WgR6uaPWWHcrDcf10wlosg3Z+ejW62KbdGQ
xVA+cBKIdjOX9oa5X9qambM9yISyR/yqv8lummolSPQhjqkCk37X9JrIKDK8BF7h
LFXr3kvVQUfd+Nx5x8G6XrYTc3VM/5ZXjFA9dc69J7CPOO3wVyfAB99rMboW/oLv
gIozO3JeubUPn9yqMQZR3yD9b5x73l6VDySAgXcGl24F3ppcsJ5E2ggjwzR7sLiM
AneRDt/9FoMPoE6I4bY7dVfjvSEpCFOCkrJqn3LiV6WkgKYMhv5YznLs/SGZ9P43
ekxbqeZ7X0stDhhHjhvBboJtY8xIZAK6iBUHm5qU6AqU6VAQhO9udABYmB1LlJdI
vci5wxECaUJpq72NVI3oTmqpl3ImgMKUnaIMZBILDp/wY2Lm5NayFPD0L0KakaeZ
44rDNcd3PNhViA80zIadowWcYdrRF4M+Qht8K3P71Gr0WbMKp+BLo5dnhT4I6LEo
j+t2GTEMWktIL2Xw3a8T0ay5cFR16LfSVYADe+y5uXLLPTtGPCO73uFfkR3MiSWf
kRkBoyWytmi89CACT9Mb7n3jzNVMvERKpkeX/Wk7ZmoNYO7K12QQpklPms3L9D7A
DOHWHcJ4opkbB8uWapYcWoF89yfRuLcaHfUXLl6+mis5pVRQehhAZ9LU9yQddruz
bKF7iOf2OaY6Z9DF38BiLI4EzgzH5PJZCahJZIKYgMaEgsFTXuICKqZIQa016TaG
IL3hmVJE6SftbcbdzawsrfrDsRiKH9TDmuRApfuAE6C140CmPNH97o5BUjkHHww8
YK+bjfZaiC4vXCrirnjMv1klLxVo/isZhI/3yPSGJ3D/xZTmHvMSlDW1m+tPeS1H
6SM9imKlCbIRH5x+FYRzIulJtuLawLmnNIomAzi8SZZg4YK3fr+3AQCtWU0Us+Wn
zReaZYM3JcmOrVbA2M5fYgD9gCaWfrGx16TQSGP6J6s269fyvAQPp23s+ZfRjjOW
Zjoz8Hr8vdjIZBp+7drdX5zzUD9vc28lAz3+klKVhTwpEfHqzJObAa4ePoHfNfaS
IWNEtIlnFuuvvLVDaM+MV8239bDeRQSh8uWcoB9Vf+2hsGfdPV6SAeKczF7N5/6c
bT51RVkSZwO9QoT7Sf79QFhPaPeXmixivpohiM9Af04Q5fi5/Z9nCG7kTjplfuLg
cmTyChxLqmyOSNqbUpuUyqeRd/ps4AisMocqvMX+AoXNV1ruqRYSqbP0oTbAiZZN
b3Z394eZv/JizRK1Rliatpu8652Ptg1PVab0ru8EgRW1HoC0m5TaLEM9DbPVWRld
Eo+kY9+r9oHRfSwIWWZCFWDcwBkAi18XL3QI3S2g4VDrvl9l6tnLuJNxlpBaWEKZ
d9Pgb6Gg68gs71QjhOFBbVvszvSgZ1OEAzczWsYd28WE4l11Of0ihMQeuQt18/jx
QouoXltXIOMbUTYeZcF1bK4AiQKJHNzgmwhf+sGrCjrC/jU0tjAATuWyuD0H+DyV
l+1QVLnl0jcyHqAn6FiF9o785twLgfTI5p36LBbVS5lG+SodFjOEnFCZxlUwljIs
B5qvfVCYzdi28mEdDq6Hzs7qPwHz1W7uq+HxsupZgVAD1bWQ/qORd2p4iqPS0v3d
k2x+8CJQVVCwtJmzwvga64mRfraNYXQHO08/I0NJ1cZpcW9GzQBdSLPpNM1NqWvz
2o/zOa42W9DQSr38HH2knDyKPK3HJvGttX/xAbpsx6RYvXE6v9brgkjl7R1YwcBx
XM+ITHrl90LozT9yyGIy83wvR7Bhe94d8TeqZ8G9G8bmjZ7sw2v/uH+C5aeXbhNS
vWoQg0ek5TOmZvVYJQoc4WKG9cNv7ATKiYuXWpc8V80vZLimlQ8+V3MIqrYtotVi
QOYcUX1YQFGUpDV4iyeCrXTZfa+egAnesGJjrnQzwgl9T2RyJr95yTK7xlxqlQ1M
kf/rqCc+y2liQx0gEoM+EAR31QmnuXnYdwGMAEuO+FxuWKsoPwgTpEP7hnY3KVyc
yktmTJ9iiPKYomU17ScQX6zNyclTsbq4tBq/fKoGz8HiDWVMlhaAUn+P7GLU6KAs
HfObPJA4pB8adxyPSbNM9ncKZcfDaynIw6TW2UC2mN117G32u24JFvJVtwrn+xyY
r21EY7OvjXm5eL/ILZKf+l+pO0N/Z7QTPJb5Ftxmdm5+3sDYjcmv6xpD/907JvgT
oKI2KwPSJUs400lk2Cn2xXujwiJjurzzIbSHOtSQeUOaVy+fdxJguV99mdCSI5+n
jS1iiJiM/HL+e2qTx0WBtd/8oiZUCcWXn4EfWquR8eqHybdOccsxaKZMaiTcUtAV
sdJdpd0aG1vaMaDcRMpKtP3XY9EdX6gauZ9ODy7NfrbauKBvIUTvsxp+q+GGd+oN
FQRYf+t/iIBzNOZS1OaVQCmOxUu01hN+njmhmilWfEgtb5eIKCt3a8UFnvyVzmjg
bCGStAGSSTx1Tip48K6W+XkCPQJ5EnT5UkxLrJl9I16FkLvVS12DOHEwIHdCaKV7
VnUFDXRc1xUjMiJOyJ+mILVmwUFE1VMNU07DBQEhM3Um9JWa/dKM7hzn/WKy9KLB
KofRq8VQWOsPNleHcP/TmOg1ZbCmSwVZ1BTAnJ2P4QInp2jm23/IvB892qMHmDN2
QWiNauF691tfPg/t9IbAYcAyv7JsaItFoFdG8eI3KiULBNVFM5AUzqAaS5vA3BF8
temvt2Wbrj7YUyp4U+laPwyr5YY55lPcxHrKkHLrn/lJBvh/oJcYNNNPZOZ50Ikb
CaKZIoxMAtdkeiQYKZ0QBpD+0Ai4FYmgL4kcsZXCY6ZKB4gvmYlII97o/33uKgt6
R/7Iv9Z487PdvZGBJJtuEcArBb+e3S9q6HzVUMTy1/Ow5+TkANxFWFsYNX+gCg83
w5hLq5l/xASQquJFBOztwyH6WaYpiccuhc8sgBidgTa72YiW0IdYq2YPjd9lO8Id
qgIQ7K3C2yHxMspPyPcp3e77S0XiiiC1+w81yp1SqESnuLcmh0ymUd7Tp3nrUYvj
kQQAjmKg30Yf7nkh/YXJtDA4TnaNUxbF+cCS+OnvY/oYlOU4Tj1w8CpRt9DZ5NSE
5cAd+70WE8zY+r58SAjvIZERwR4Rxl7upEn8sv6oocUYW3Vbs1b9uX/FBYw1h7lP
dtfIVjr89Sf3zs0oOJFjegqBdtVQ88K+VvYiKMTlSVBv5OgTs193ZAYgZZc5oBHA
wIhVutDvQijFpDlZqBfg6kC722AomQyzdea2eNFn+P/vWHBFfCZDa9//Xy2epK+c
LEL3IEpB9njH2cofIdZso2M1gYoj1Tyf5KG3adM/0foNrR/ijWKwxuF7Qs15v/Ca
kQSMekmDGHUw5LjszMBqvbbEubrlOdMIcbhaV/g8WkjAmqolpXOl0Ja8xq2O5LOo
/y6Rwx9/r14ohhvzTth/PQ0dp1jJWeBW+o2EQFVMwyi3ZKTfO1QWCLLJ+gzdmCN8
LFc0EvgrnPUsHlfLeBFX0wd4V60MhcLM4Clz+EODtnhn66/2b4tBNj5MI3BOeHaq
IkkBl8zMZz9kdBRV8SQpsdop5oL97R/jLS+HzO1v6jDDGeVCU57AkJOSWtXukOse
GQuV/oV51EqFiDZMJsTFlViajdgk+DVfgPkO4YVdBy8cRugJtz2Pfb2e2aNxml+q
Q7tb3e00iZIphiEDTPnZBYqikDC6MPom+YQKMygglqacPyxThYoBPa7ldMmLYgxI
nPWV7gLnouoxGoZUxf9LaXQbpLNEnT2Q51JDBEx1OoJY5pItkj2pofOuCodq/jAl
Ty2R7T3PAvupY0ZrsLmxYRvHpXFS+XISjNwxT5OSY03zJh1JX0PQnMPVFRgEVFFf
sAmv1DFHOA51q56XbwBRdREwtrQLwHEW7fNrFZNOdDfdphiP27b/G7zi5iu+2vVW
yxYv6OISVZ1+UMEKguHXWYjEO0AKnAFVlIA4NGMF1jG0JzXZiDim1p6lluhIOjMn
99Gr37Xc3BPLCw+PO9e4mXHehB5ZVffnbcGD8GtJgznEN75LxiLKw0rUH6Tno5iw
iv4Gmfj6ur7DkXSN9XAfh4bC/yT3vSLINavSQtPpPvogKryPPBp0BvV/kNQ0yEG6
WkgWgdmHkSjrEAApaYf7VyRk39Mi/Bq4xvqfBLEFO/1nvrDyvxsYCwwkG/Ajl0UP
5kQa0DwFxhH7zpJPyxircef0zLno39WGKMoj3CrIkfelRuhercygeBVJX65j5mju
gkBvfwyMeNI16958w5FLmg9U1gIm0Qr7mcawQy4uw50fG6i+g8WqSU4UhVz8+TRr
Vsajl83Hb/B+NU5iiEQ+HATzV9bk6K6l9M4Ox9pWpUub4BblmlgzMJbX8gvfyA05
7HRIBYknQhRLvlVm9+dk2YPrrVLLr/4EmVSUAH/iztoPJWw2YfixSJcS5vNP6SEK
xObYTc1w5/oSxB8s8J6kS5jr5izb4NmHHUeSXIjr3zIeH+b4j23Inj9eUd0ZNnMN
ZtegrIg9WxHV+UBk8vFmQAUjrAEnyZbYlt+F89nXAceMHmVtoPXZ47UZltZo500P
JOI5U4kN22ZK7/muPteZ/E/TOUAMeyooNrUDcE35OBKg2RoMpuhIC68OnwNG6hs9
/FTGz/ZqN9Uga94romJyrS0temvGaNs2uJOH57D4Tv7e5GywOp1HiuFXBLc9xa+R
b6uzfBWQkfmDn07w1YMxd/Q4mhjrsJfoW+bX7VGnRXLiheSbInAbykROOesufZS6
2b/IH1EC5TZRvf1iswlFHhkoNleVkUmyVIRrzaLiCkSPOatAsZ1fDxh4CFjmfKFp
Jzezu/qa/XIGafvni01Hj8Gq1XmopMZcx2NL6cwFOinZP/zlGLPt0NfEsMY5ddQN
CV7BavSY4m6UnVpEEro1eKY8WSWS20S7rKxwlunllz7u0CwPurQKX0J9spIUVcEa
UfMJnnVlrSIau4ZaRf0QxdEsErCYuk7ZNLeJcfHaaIZTZ+8+kDJkQ/05ET6XDPGS
JGFFgofsrZlN5eWl8k5JR5AXkJLCx/M/1v7RwzlE5sSmiBE/et8iRF35MNl8dl1+
06vmhfxatjLnuQE3gNkrMCBVkTI3ArFUEEKtLaNr42EhJdWtZ1fC9bBi05xWFzXJ
TdU/lsh7PJvEwoISFaWKjycNdCItgCKjro1Gr5Y9Bkgp0OTnPHgbgy31JXid16E5
5ASOFOHm8ZV8aE1u5Wc36smdj6B+l55O2yi0dyV0hbw9ys79b41m54AC//W0i35I
FNKHb7hVAxKiesGHtys21HJnfsorL3W6oSkapLwCAFk8PzPhs9PZZTo1h1ySF5bz
nOJHNTAe4agXlwuN/dX9ekd/hWVYfIgDFocXGOjFzHLvWOee5gHQFXCbS4hr+lQw
5+0Upb2TsBt/2TvkO+VrmmzvY2UMjTuFMsMDLBLNZm1iw/pe0bG908fCRnVIsTLL
AhFDGqQWbE3S1i7AYeYn3MI5GtXWkSlo3F6xyrOl06GbU4STrrse7ddC36gT1Cqq
jAAYAAEKB22HzvgA9Ckjeb1PE0iD4Iwx+zPiq6PKWL+z6BhL5nfgCXIe3AikFagf
w0y3Anux1p1y9nL/nTmmqXTXRxp8COGAMRHZoIQdJz1jsucxhJJsRo5w9Nmgee70
QL9j7RKRjAZGP9OSwM8ZVius64ITNzOoDzRgUfD1Kkq+6FpqzWwMO4nUVIIMtbjJ
g43WBJQm9sQgiI0S7V0kh0pMQq5RmD7RRidIA7W6RRANPvZhtaYHfASkBBVdmcl1
kX5jypZBs33GhkQwPZxlRUBaVNWHv0GTFm8sCk+kQxBKcigI66aWVm/iUaC4K1Va
vIUKMkMBk9mhQRQi/Ca2QmgvxrD6J6+k4ZHOXsnCzVXGghE4404ADBecdNCqXYKe
sFF/AY/1+VUTj/vAML62jqcZ5P5mhuzZN5ahaG/IUQTIGY7qjCBAuciAyLnRPUMw
4ZFi5rI3c0xv8K0Z+Eu25PofdCSqRw5QFcaIu7nEW3O7nxAiAPCAWjN5eBXP4xuT
niiNxBhOZuftDGyiIR6+dqUYJhw7TLWv07aeS38LfRVkZWRWbIxY6urC3RXejbcq
OBDjaKXDOONBzLFahzb+Dq2vULHMrNMBbw26guiXZfBFzA647GyH+f8ZlNQqb7Wj
lv8sL0XY8NLDoPVA+y6FKgwxs35G5ryiyszfjgVWxRP+AlyTBJZu6est1zHqQHc2
ezIpEwWM6cihhp1inN15NbH+yD5EbSpq7ZKNiP4CjRuaxJluWGtfFx+1rxJVtNcp
AkkLRq6DjwNCodIXdPXFuYAaB4DBYh2tcqcLihu5AdONHvW+mPC1/H13oXVL5j4B
iyzerGBlCZlf1jMBFMfuzqsouWwFI18lOMULcjPdkCZEntZ3M3FAC6TMB4PjE+Te
gfF1HY4yAEhWVL9G7M3FrwiAIczCLMurizkKWVyTGp1bdnfE+qX7JLvpLo8xPE8w
AMAUz3lLB/mKCCFJZsnKUAv2KYqQb6pQjWcSnNqO11VZuc5bW3gqC80q9aZBToVL
0PICtq+TeMHnQ4yWMaTxAk+n/XDnfTJNfsZrF1mXAWcTEi6I8CridFclpKCVW6lr
khI2KAtKBMXKEtr40bge1isS8/96m8jY92a+p3JKB3tFcxDWbd/nF+3lciWgIWTG
iOvggIPOsfUz5Jk3OfyaunUDmgS84W3DNgTYplKHYRafNrJSy5iZiHleE3m0GKDw
m5AmCs7RjhxWcm1TUL47QbtUBR19zoe+lU+M3YCDJJkUd3ewKpFvHiW+whAjb49t
eEsk5moYZUyVh98WTuZFuJ003dAfAtVElMUJA0iwIv9fNoNoikAevx8OquvmDHq4
K4J3sGO1N2GBl17QI9Qg5OztG+Q+ZDwxO695xXYMpNDTdwAXEgw9WPSboOODVvdc
oOueslRkart8LaSrmQYZ5ZMZ7Z2sXYcXsZ8eQsne2537MgQ33cwXS86Cn+9I445b
gHSiaJE9LlUCiZwwrgGKEQyUb4JOZU4C7DsRyFGYzQF2jCHZUDUGr4XWMmiVgzLv
iBJp7qAe9LQ+gR9vjo8lP2IojXE0MTc68cxEjMixB7tdsSzDqF9V9T0IiovPJTce
TKI3DeEWNyH2af0l52yVFq8ZXlhSXiUe2sMZ8nKvnBSl32//xMqWin4OLYRhl5ZI
Ef0SAiu55p+umAhruAaJk5/utP+J0IKlKFT2n6LCzphT1DAMjxkal8JtIc0lIAUN
ZTaFBXpYs7FumZRIDGnwoNwfC8gxlw22CCWYG1tz+6Y1qe6lUdHCwAvKTP57hrGU
NkiAPVVyFPvYkmHm4B9wLm/KzJAtw8xbSPdIa8WAFJOqXYrf6gclTiiVt5h8VOrI
JQS6Po8OrlivHmkWMd6fngkYAC2ke182LcY+0Nfv8/+3/gPcMTgyy0GBehtn7oPm
PV9EqM13sbST2mI0vX/7xptk9nr2POUUvuO0jeKNkDf9onQMr0QlJM4uTXu/TuPN
qPxKKcVqq0/AWWP0EH1EEu25PmQT9NAny5CwItstnhbzaLRIULiB4ttw0pu+sRgN
mjJxPPFHqeTNZlNrk7BQPdti9t5up7B/8Jyamw5RSpveHJd+z7vWU7cnHwEdVfw+
AE0Qqa+98f1umhc7SF1HfsnumgXPuBpV0WnjWmIomVtfMQocVYMqvxtu6zbTmzDo
A9oMfzG8ZdH6+Wmd0JAgucnbVv0C6qkxDfq3tXX0HnpEFpCvaeh+aTgpIpOmkF4j
zvC2HVT08jg/wG96DrsxBNAsPFwVHI6vJa+VXl/AXuefGSMMs1pmCtU5fVshwUoE
SEgntClpWBEaJYSZoIH9n7WPKO27rvbPZ7E43q0g2Ja2r6NCiC/mzuz+v5mRTlQg
wSsuTmpXi8yIl3dwbncavyUXd2ppHkYowFWk3QTvIy99lp9+QpqGDaWK6NPvc4Z5
H5VYMAs81UhYMjxQaCjBmlegjaBIIiF4kSO3iN5wHBfcUnnVOKNA/MeGW/z67sn5
Y/i20LLJLZBrL2BmkPUr4QrUszT+68YJWPJUUazKUUrLKcc2icP4/Sfq4BPDtGwd
X/xc/SFB1j1SLQ27JM80Dk/XLt5wUyiBtDxh3d3zoqg2GmDB8s5IbmPwu8uB9xff
yUr2CHZODF95qonNU4HrvmX46/XpJTS05Z//DdzDgV5bNJ1h/W4cXUSiOLKN6fho
qJBrYeo7xdBbd8rUNTVQTGt353+soWRQRWYUAjaQCzvro7wPMM/yqpU9Rdo7W3RA
lAhqjcQfDbhlRbqKg8MzI5SKhr6i2fyQsIHwE0N+5t06W/+rhlL3o8S+PuTKrqsI
4c62Tlkg6VrkD2oNDEJzvgWczoARya3bFIYohKMPMqVs9zZEjA4L9iiAt2DhaZht
nsuCz/DfFf3ID3+0dE6S9o7BGsGmCxLNQspWIh9TjL++7wG+u6ayv/C8HuZJz2dz
gK2rytpdEIWaBdp3tc9QqN7Nv999FpBM52o/zx4oSjlvIWViM5ur4xg+on+XofJw
v9rHGQwXBFmmdbwvoN/uoquphxpMLfrkpkTILIgWgwdds5HJFOb3rvXlbX8OCMmf
duaE2rGrNWZQFFecjGjc/hZhDDqJ5hwxZS8Qh6FCZTtkkA4NrwVHCmRaCV2bDS7R
owBlsWxwUhCTcojzvgKvWD2+rNhVz9v7QNGwSKG+9SIhzsE/UtTx3e0eiLKsdwvY
9sEo/uS0ytlY0KXtGbcDd1wk06/6X11SDh02Pocbk8TiZ3amfEsLkCiqgt14BaAh
VgbWZvlVGUtfJZHX0DyA1eZyOJXX4NgnNtONOmyvK6ZkbY+aGTDQSVtXdb1BF/I3
vuyegrkpq2vOjc8Uyw5pWy8mFMeF5rzLQ4BM/NUA2ZTMJoBM+B4o2DE5P10Qxntl
/HUuS6Z9d2IgfPJ1+5Hu3VxvI5NrXTdlCf+SLflkVjHdqPgQqIGJ2QReqXKeNtu6
cUomO53xZdbDXY6U1MrcwmoU3uIhtrD6tzDa1kcOgS+DtvXAvjb6ksfyYQOV73wh
BvcGbjba+dx8J2/kUt/Abu9DoiymYoGPWImlK3bu0dJAZ7eHlJpGS4oZotvYhq8G
JG9xNJ8rdfPArGvCzCh8unBs5j8xG5SKqKyLR6r/u+El1UmUkjVCR21pbjmk4tDg
ellI+GIz4I0GHLEXwam9s8I1/x/NDDh2xSIxMo68/r1msf25TSoOwhA5NQmNZLT3
v51YXptUznmmDvYy/4z5Z8FZpXI/+gJo7SNi007zv+DfsQhxWNRH6HM/7SkV+K+e
9Unt6f0lzjdhzLgpM3R4/LwH55puY/81Vf+Zusn2eXUeKxTov4uH9ou04rtDOH9f
OMgMf+PPHT2s+pPJ1MPIeLy8nt6q2H4ukoR3k+dFPRkaF42EGMuSGQrNMXGKzMQA
t/oRoxEg8oA3tnVKUZxaCHJmDjV2N7UQ71dYegaB8hcQ6o0BFgtUiQIN3X5Xphr+
AA2ZTIYO7PfkQ+YLql4KTGRShTApIbTqDse7TaGeTMWJKUaSKN9RCBuXHc5rlxtV
ik2HidomQbij7NVT5kdHkqKMxJYHgjfzCtfDOpHyqAibVNJRu4fcY33FguuWbrNB
kQpN91Q/XJvEXEqxNaiI47ymafuaUExuXrOQItGTD3ppUriomcYYK/cJkg3rVRBp
pL3VlzXLXe4XATFfZUYeqOi1RzW8jW4ITQDGihFco53TZNb0FFKMahOyF/O/noVD
BBMdjbrlsR5XbsACoV8yucpOi50eY57rSdAV1PyL3tELJGyettLDhqc8X3I2paRB
WyNtSHu2J9koGbFH2gUjGb9tNMnih223gCvTV75MFGC6N3iHyQhsnV9TIRtcMLkK
Ud2BFIYh8pq5iV0gQSS8+VXDnKEL+Hhs5t3TnzSWeh3G4HvKplnR1Ejor7khMUVH
M+4G52M84Et48/N21qNcESiaG7m1YQTYcUildwdDyJhnWwPGPafpBoAQLv3D6yw9
ikGoKJSGb/f1QE2w0qdDNxcsHJ9UVgiAU/6YnRvIYuSvmj8h0uJ3V7wQprBUy1j6
2mf8Hn6YIEGaovPB67e23aXyVLoMoKtBPasjBk+zh1PdycdNZepgDFpvVHziEUcX
b9FaX7qJr2kCxfOyvGmRUxiHrYIQveRbGSAj7ZjnR837gLBy2rBKPfGVLM/wYeT1
dKA8jp+NNd7RYGOfZ0QpG+rs8kaZfu3JkJyDisFPRnVZUTdwzLHhpxywAjoJn92i
HTycZlxVDI0KOrSfte2ZR4ADOfx8o54+Cjg+kp1Ksyse72jxkGhJKK3XwLiLUKpD
WiUp9beG6DJ9PFVoNUgl5IqPUpGedC2U2OL5ThKSzOMvZWtEZ2yx1BrqD1mH7+iB
QPlfFR3FlDCgKbmzn8Zf6Plf8ykEAJT7xDk95ieIPFct0+4a86Sdj6FUDDrkSWh3
f43KXIVl/vN3M04el/Aw9qV4g9tEfW0kUqprjwOnlHBqVsfa7sVHiezRV1NwTs6p
aVc3KLhJCBbC+X0S4sZG5nTdq5cZnBdnhvwqlKjRCfyAli5UMREHimia1fFdn24M
QlgyxZkg3jYxPlEbP9fHHisHKmx0/RdWIFOfpQKwZcUeCeWoPJuy7GX6jkrUY2HM
Omuf1fqLSiN5qfTziv9jNWKy1+LL72JZRQsDdIS5GsE3IMcXx4AbwCPt5rgbGXXc
mz/YRnHcrPaTi221aVOJCxEzyUuYVFIc6iM6LZ6xMAQBd5po4bHC1nL5PQb2ueqy
C9vrnuOllRV9IMTw8xzvhrI9rDNBzbV95OpVY1IAWp7UmHmGsnH1Tcy/IfO7q4pu
Eh/9gCKV/cZFiqDiO8vMx8/h+UQIKo7JkaCnn1xDH6oWHrvnZ4SN9OLZmkmCc3f8
9BO3/RqvQwLcIWnISbxbqz1cmVRNw+uzeC7VNGZm4Lr5alOaJBONtZ3SYFHTFZh9
DTYjZQgRje+aupkiHHCf3A0M1lHxqgaj96aegQvRnrsqBt816WHFEowg03weOXdW
muuAaNj+dQylxz9Cpquussw5TNePCFZPWib380viyaUqGanHPJqFaHjVj2NT+HpU
gGMegEc9lsVzz6Br8R8m0QBgqfVhxhrvcgjzMUdOH8KAjhDjJdxXG86M2VNKNs6g
PXssa+wXr9qpOzEPaClzkaqOzsOpJHg9JaVUhIEHCx6FgYPt/1TaiOeA6I084kDP
emdOg0mre1QRf29wpoJvm2kaXlvZMQe4W6j74E3WHxKwtR6bnLlUCp2LGYefIFRc
7+vKnJkZQ6YyJ+ZDgYwlXDQYRd+waqejhRnR7zCg8R86mKGdkPRBwehrQVSZKEWV
D/p+d1y26udUGm+zgLcSY/ltd8axLoOh424uc/M1ZlqEJL9WTsDahUKmZMT9igWI
fqGJXqzwD2FpXq/CzZb7Q0oXUQMbSFX/qDzKM+QWanE5XVb7hgUxqtQ5NaEg3GPJ
4O44Afc9pq/rHha3FsNJvnE+LFcmtZZTJCg4Ds4N7MWFmMXWh58T9Z2+oZpKLCbg
DyfMpFxDcHiiexwNS6OGhc7gYgGB4uXQtYtjwXRjAjqyZJ5ytnPMh+H5Md+D/xKP
pDOfOGSrstrFHph/rzWmsTr0W+U9K4KVOCsyD/9jM3WF2hbWWtgR1zWYnqMIy423
AIH+uSvFnHJJZzFsW+zAE/SPYddNRJmQZMYfPiPlXogcunP7DBKHKsUMkWy4kp/4
q2WyfdY2VwOCmnL9xiWaL3dd50EGDtBG0OiOLMTjhGGCNmaxg5bpeclpm6snigRe
4v5zZrx+hLRABDGoi3xpDO0kq3L6ClxLbnJjFdy+/ve76U02RPzWDPd8Sroge3n8
5FwSKX/fg2xeDTpokwqhIoF+886YD4zLqC9zsTg8AQ1RQs1eaGybkYaQmzHRVQB8
iy0MTXe+nZ1r7wqA4cPP5yvH4FLvcxEFl8QIpZbRvqBfmyP4pQ+hwP0h6kpJNdM0
cpbhDkxKfzgF+uJkMLfwQSI9B/t58Tgdg1Ziz41CWvoXMUW+eR525QxUA/Sm7YTD
WiDUXHdkfIzoYlAmzPnEKNVVsC4sEqjkSkpy1Gp050uAtgz25Yr1+j6GB6A7+spA
t1+0IJ7sA4fBegBVhVo1xUhZZ4P6Id2P5lMNVGyNJu8+qVpmasPAXj6kbI7tSPG9
vTC9noAc9COioP0m7rBL4K7S3zYx1U/5NiYCAmETrUxakS26FkKUTgxOoguw7jCM
AUStt0IU7mXE91GxwfqI3hxM7z3lWwK49Zr1PyX+GF8C13iXEaGrEFCjRLRMnDRj
FVoahzeflmwdXX1vPPZYBSx3NvBkEGzaPDZCTnlEsLJ4YLaJYYChdzRAy1UYJeur
/rw7xiprsf+SLIVyKnlSitAQn/FstHz2CnfsoIFCMb3/f1eqBaKCISh3YBsBRZGD
nVs5rV68YW5Z5/NorOY/p6hSkUrXZIKd7Vu1DiRIBnmSkPNssXH0133xPKH6mgqf
81Q1Ne1J9OIu/o15ORg9vyEQcaJZiGeDUSqKh4exG8utlXSqIMcFztGR/25HzLfX
kvv7gOWXTmq1UAv8niWrTH5x9cni8dK/fkWH4EGRCLT0p50xlInFNO75Q1InFGEH
Yoe6cFodYB85SVGrazTai/WtG1dsAPgyhGfcI3ZJZQO/826ev5rTpKZXc3ouxlLB
FJWLwYi5f+7SzNaIPn0l+MZTDa30DKvzmBAAc1sz+lj16TAmoWp/WfgwaHmGrr+7
cCfWxBp5idPZB03Y82wHTkR+Mv1xkZHARfWG+yL/HGtkcptCR/FTgQnQjU+l+FBc
i9W4J2q/oOFik1BlY4F9g797u14gUlqkbHWDnGM1Yx+C5ZmayXLXJ1ryh2+seaL0
Q29m2VWGDbs/lW4R9aHLi4/tpMbdeHzmqoEqPgFm6CDecKONGkQ4eqeDyOOyYNuP
+MnEflWELadKJthNIAiiszIGk3RWmHRMlYaA1d8SSB2NfroUzjru6s6pKmH58hSr
y+VLj5ggzDh7NppXlzy7uSPsUt/MYoTKmq9USoxqPz/Htl1/ylEZZecuKLjcYk64
5aXFmh+H4jp5Xu7t1DmGR18I5fXLk3HDdpMctoZf5awfo8ASKCdSGcTMPBQVN4K7
1kmuvF1KRzXzJiORbPnfVNZ+Jc6n3HHYNUKAnxVWhZb0sYRjyp8c20XOBAJRG4Jq
hqsw/C2JZ8Sf6IXPv/aPHywOggrAW+HpXYHoFgGJ0y4O5b422nMfk+WXJjGII6Qs
aEZdDZWAzwAzHa0RlI8P7OfyQuJUIXEDXtZPOXpMDwWmuX5laJiTPYhob39Ym+Rd
0Ci8YJcRhtlsuqrRZd3P7qVm6jVuAhRkNcluZqBSzXiIReckR6HPQnhjhqs5Nzbx
xgcYo50DmZ7P4QADzfGK7H9zSQIr8/DNedWOzcJ1l58lLC0e9j20gvmYhepMZI4H
QT1ZT8B3TEA8G2KB1O6Be+sPc4okMWgQcuzC7bA+v6oHlaAhCMcxGTzGd9Exx7s+
PXTpiItzPk6i1hPwSvfrIA5QYwBFyhg9LaoGwraDHF5HIcVapJMqRO0WCX3wDzl1
6coE2oD/JX9CbBeakqUud2dKQu0n0/q8P23xNDSxP1md1Pe+oOBNbpAb89kFjy2p
rV/gYTb0o4hQ/jZ09IUK1YOvDgzUUaOoO4MQCyp23NzFYWNjpLBWLjW1LaaetDnw
5gF9cZHgZ/8jQoJ+RLSTtB7PQuEBq7E/U77Wwt/wP1yVEJgG2k6A3glkinBs+BLe
njSmGmfJ65fbpk+zDgU8SVWx/i4X1NAEILNL7Avwpt3UHGnyncC3pKiaKEwMBTGm
OlwKrWNFWpYo6bTNpa3ktvpAqLxGkbn/cUVsPRZhViYD1ruqu16iyZYF9urIcz7f
B/dYhxIbEt7F5pXZhrktEVd0+5jwmg670h0aCayb4MCSi0phTYVv61TBvZubcyZn
TfVEiJk8K1+Dvu/jgHYImR5vVzjzEqwO04p3bf4TEPPqPOx4db21gcGgABpEVVBq
82c7NCjE5M/D/D8/tGtDbAdCgYOB1gvkt6U61cwq1OrOZ2uQsTP2OVK5r+yiZHCy
x60RybZYJSP5RdhHr/FfEz1ldDTD4VSDLYlSz13mSmeyqpH3oysdTsuo6kPGZytP
1miJvDTH4IH3G5IkcTL46MKn79lNhTq/7fhVIC7zNkgRElpJE+ilHOU2suI7CDPt
4NUCbK5fYbH71SuPChkOe6oLT14fhdww5dfYLWR8bAgpQdbHN7mt8ZNUqv70DBxM
qqcXsnCwEiwceAlaR83CLw6AXhcJTSpw6TLBpA3nLAagBYgAb+7mrJW85CaHTkYC
/r5BGZERZ0jG6vprlzVcMMtl5s1L2KPxUqvPVJMWNAuM+sLnZ/XjupkgyJkbDDp5
yZpmUXhV3O6s9S3mBEScvudBK+0JQpc6xPX/uCGEJBeKZ/ooZXNBVnBjpc0ghhK+
1LZd9WkfXsmi5LxdsIMDC2Ozc0v/el+hGYe+lz3kdKLyviVGPEbOKOqT28NlgV8/
oeE0bdz/Ii+nDncMXPrHYeKC0u+fbYJTd07uhTJ8XKQF+jXuN74kuPJuB1gdyqcF
DN/G+9Iv4/rU03A3Cgwnniqddyb1CNiRszbNi2dq7/mNKtgl8BP4ToOSJWXM1Utl
eTdgnN5k74jff54fUh1EOSGzsdMIvlp+ZIdUug76xOnk64say7QPcnUzNpXbSPD1
3LFflYbWi1BcCM9VRXGzgiRL8Kv4prSlkOXm3gifjAnE6FYjTQNkKzeZOCB3sMML
FiKxx/OmqIGeMRB6o2Xg2KtQwVQGMZzENXnLJN7YtImSbmUpauXdhcpJ9n87cfNt
HIPmql3l2QhP6caDT1l9XJJuD5baWIBh6h67qEVske8qdcF5vDG8zYyjVaCiKi39
eVGZP0TToWGgsGjuDY35yvacWxJX4pFCsXGm5Sz/lEQedri9/lwn4mepBeH2Amf7
Ixnsr6l4HwbEK3bTzjEQBrjsSHSWe7Tm+iWdNFR7kkHdQNsnlKaODFYRkIlJADYm
8awZooog7XwVxA3m7ZN2ADR18KB+lmbj5uvEeqFgsNwtgPTQPNYjLuspDOIy52bd
uXpqkEZz1AakTgiugIn+jbiS8OktciqIrtp6k/S+igSZAxsq8omjHrdJc/ODtQ1a
btMFODHHzfsSqZ8zhrWmUovCkAfJoibt5y2rSkuC5sV9dM6OMls9UKiGqrWU2bgv
tqBvbgvg28JHP50NT0jHxWeIQzUdnxcp/25INd6wC4Xb3qkKlIrCIyrcyiKT1qaN
j1nQP0GGKpLzzH15kgu8NhCz2Wene4FuV8dYtFQ0zQ6spG2M5AjUmJiNd0uchO89
OoWI9ahVfkcxUCH3mgu2YLQQku06aIz820qsOsItvxPBA9ZmN6hlGnf7tOrazJL/
Ro2PzKMpkwbuyEu0w0i02/oOwuZgY5o5369IgZVL4z2bzP1yAIqFmkYEbABOXlTg
rqH5REl/m9sQhLu7k1a9SOXEgENgHCuYyoOpKO2cGD8duIyc9lXnrtxlQ/zFxojI
mAsJlpezmKHy4TDrjEY6cQygoffE6DS0T2Fox8Rmda09pEwzosgF/PROe6llXD9h
3p4Zrzv9JPHU58dKA5hxPVuFqV0FPu8sQ1SCZT+0VVWyLcwE2fWmZ6FXej/e4UG0
lgMCD95N/C525NcixopFo3vvyXAMuGo8DhNjWYcmXoIZsG9i/O4TgN/lJPgovhA6
0T2UIRSiIj/yVZKBbZF2HnuYhp2kwyrQNcsJl61DR4opix1pKj0q9e+ECQYlLkVD
P7GrzZBehqM/h+0wfmJO93/6d4DIMQDigMs4g5byNDcuZWRZZrqmHksEQvuVGWN+
RpbSJxTubz90lEDUkAGvEy4AioFFaxCk2BIBA3cTpbPjMGix2Dqx8lyVkkfoMxmt
qurNI79Mg26B6p5ug1HLob+JkkNSFrjFbzXAc7YRxmE+NJq+mJm6ab2Fl7gYbSKc
eogB7ybt5GNXT0r7FJGV04vtKuzi2fUAr73H8aibYPLXnKr6GkL66QzIMglcw4Ag
M8goRkQhlfMGVJ3IKJz/8znGJFPifUs8uw/TKOJFZ0VdydmG1zbvHErj2gmBShqI
dYNgL4NJvmDb+sMEV+Y5zv/4gNf2UaP+GKDACY6Du5q+8KOGP+7EdqgP/5FlG9oR
V/AMMi67NZnbcSVjkTe2fviAaxFbD/5kdJDDk3LHHaYUal4mZkZfgxKjZDnTdet5
nJX5uNrI3Ft2rjTUK04XTefsGUvCE2FI9Ur/hjVTHLR3LVt+SSS0pSWwXt2ZzP55
Zuc+RQPBuy9yPRSwsh6U3+9Aia9FRwCO/OKdcJBy3mwdjlfhXPHmgVo94UGUBwk8
gkLZi3/kRJ2aQxa7nafWdVLFAvMxZsvBFMP5lUe+7cxs7VAermQVnEGW8JvCRg61
QbL5Pws6wR8xmSjDRVNFCPdBX9OsMVkTm4r0xkNb8E7LDBBDUa7cTydnwCSqHSnJ
Jx4NVeurRUgXSzYfeXEXgR4L9KX1agVsWEwUUMaMNWoEbMNFFbAZWITrQou9+Opy
E1o9lDo7cCiekEo22Sqhbs45ZnzbtT7NYGQIx9Obx+jrg0wIIZNXkuoSbivxFPGW
HAaZyiihmP1cQLyTr88TEYE8Ki+5yHYeDev1um1y04gjkBd8dj8o+Li2q0zkgYQ9
2KMQTbRwacbLsdtrgFG+A4WuTmZHPmbCS+6neQ/Edv6Cn7ppMLwbbNFhrj/H3sSt
2SqvOmZjovgCRqNNZn/XH+G84zY9tvmzTP2sLMrJdDsiAJ1hdS8t6ki5anl+W7of
4sRPlKaVEgMc7x/l4xMBJoO7jcy/ktR6urXt50Eb8DIPVDE66y8j+Qtg19CL5HBd
GQkWl1z1VNFRn+7vx/9flpNloh3nJBZn/gGXJTKVosGY1979Hav6BLuOcgpHvJZq
tISSTmttfDs68UAwdrPh4y2LkmdJkD89aRUGOyQDCGssyNf3PaAtjbid85653dzv
QexhPeVs78rCm4GBxZOc0v0xScMLFpTspkGJe75HMABOOyMVzrs8Vnd46uwz2Tql
H9erzdwGwcv4XKLyCs7uarTEMVGFvReZM7isjrvU0rOmgUbw2RhEsoN+x/CkTco+
FtkA3A90JglRaRqONfkK6EWAfFQMRLMEPa6RVtOQgMpE8HGhaKDBDCJs67Qh7Yt1
TEWrZcnSIxXJCivkRfllvLUS6Bam8d+77Tz6tnVNKIT6wGmMcg1FTOvW5VRFkRUm
M+EvmYrqD4GCFm4O12v5eIniis3qzcffCLTvvDksTOzGJwfaiTukCGgSOqzLbzbD
8jBK7grklbzwfU8mati4rjVmBcsW4+3heOv6AfNxoeLyxhmPbDXvc2gJL1VZrFXB
i9+4WZyRG7Krnla4KvRk+0GvgGs8qpExndWIh2v57sXoSJuXB1Zg7epqxEEBRNKw
D8LqIBSxew6k2QVL4Oh4yJlTL8bbcNlbDb+WuK27dt/L8B91Ay809A+c+BUr4o5T
37qKaCJzl3bxUJBxdK14lR/DnhQa/8bVgRKEfe9qZAngRg+/IXd7tNVhYA7pPrL5
wYGanecsq5Ep9moXHr10L3wD4IlxUgNdo/pnr+sAJ2dPN7fjsB70sPIW4odBhrga
wI8oyWCR06k39oCW398Hi9p0LEbVmfXD/ZlTzcOHrt+5pqqssr/Z/8YJK3B0EOoW
cMTBdI9X3OVvEoMpAiaDDNB25cOYS01xp1qcwtfPttaF1cXgEQUfgebWY/fotz89
tBCbBCnlvcKFIf1d32BAsXGrxboDr6JcuIy4oe829aiat+YNTo6fgVdHjDnPgnuc
vU34rF7M0zbM2iVpuU+jt1d3pELPiwzx889aet7DE1uFpLG+ZRli1cMhhOTz2Hb9
TE2vK/XYB1h/y8EdDbUWru9xSybLVgv23MMUTB1l5LKZhC//E3/HhOZuz5ReurKy
vZCURGOsW0YsHZyWwCDu3zDJPa67yr7wrSguo9hAamNTjY7macXMIy4sXPdUfN3b
IZ0bFs+GhyJtbKz3C0uHQ3kB++Nr2pPW1TyOxabSXqPbicK6+abgJDb/lyU8p/+0
ENdJSstgW0JyWPVsiomk+KkV3ieivhnfxQvcWin6X70heOBdRxmNSvCsu0m9vgaS
ofs9LX2JYKBANjjq6a4N1EObjOhQP0Z9kwoy0KY4T0jsydHIIE4m43wy/oQcpqba
R0bWLRpmli64JsZENC60Z/+6XJnBNZ64XFG9j7o0APslaFwwjAubeSoYFyBAmIIY
t0/HFWa5fuc7enm+PNiCfABWLzDZtMhaZ2am+kWkGqhrpvRzkeemqGgr+6CdT2s1
S7u1Rk/6LkGm32PrQuJSMPLIPu3sbKwthXDOK5N6W/S8xPW2v/EGB/99gRHpVQlP
/2wgJtp+4K2/glxK/3uMGdGFDwWCj69Vnphz6I5Ktpfkx/SR2GvMov+LLS9iKi2v
2OFfNIl3aZ5GkwqFifY9D7sZtFGAfeWycRggw+CHJ1SX0DFoyARA9PfMXfLgE3oz
F1m1Zok0IYa261j9MeuD4uCuJjt1qO5ZlONnUrR4W2WAA7tcufnhqB0Ieex3A3hs
cA7OTYLF1QqJuXqDJQSXR53QKQu07ZXXcZx6wD5/2rDQzziOt8iagFAGkRwTef0z
Wco240udp5XE4zKaN3Sf5lYl5f1z+8+U9ybMqrkCQpGzvy9r0UkYS2kJEF+DsLh1
L4qC7Ppxw7XkJ3+uyIW8Hj/WmBXZkxAWvw8FAPf6fIWEicZd3JuC+GNMah+Vg4Ab
LtqBQ1LqetSxHw/t4oZIl7A4eCoWuAV7CsyGK0RzZiKHhnk83izb6jYCuk/Ri4mn
gjzTHXwovcyQfy1bgxdRo31C370Do8kV21Jh2X6BlBMZJhl66/c/jl8mSnWdkZao
h9DXAH5kTjzVtHh3jb7liAAEUK//ogHPPL5n3bWazA/PM1nAfT0NCh8nFij/MKhf
Ox2JnjzKZpgEwiXf4OQHjYERdPzqN6XGPo57a2KXc9ZVZyKagCJQUqictlxLRCjH
opjMAjIhJR2o74lx1ta9hcsgC/DGcjHCDSazHdgaxMkV5euGLycD5W07ieQuHfZ7
+lRqFdDuWj5I72epR5s1ys+uVo74H90SUCwPh2ZN5F7uC00ZSROhybvfZxweBKms
DNDV5o8vW0197OJMX9tX9Mq2cOsarlMYny7kWL0JM108Nw9XDOdbYKco1OJ8FXaN
R64Hh4hieBO50zrArcclCmSASydiReM8onrXZMr3Ew+WAjlYDfwKwO+Uu6SrqV3o
zV3hcUD1uoXLAsPCofg7Dq6h/xnwZI+zbSDeo66GSffpGBK5Be5apxfhGz2npK1A
4KhAw4IZjKmwKa7ndCbjYDrfzDUi1mFkfIfurGnQM8icOOkfoB3r4x6TshFQ4AnQ
9MTwoEAPhL29wUhEk03AiyKiWtO0gk3EQ74cNShJmUd8NY/tiIfU2uiB9aM/mytU
TGWSbkhOqgE2yZbqR+akqzCXSV5hc6p8IggVdIjbAsUNj49rX2ZAnXTg8KF7LG/U
xGQK9XE5TfBlPooo4UQ1kzBIqEVx+FaPXwOOVBbpwQEZLZdCmDQ+ifR1XuEbIWEu
nLT5f/32XMXufZyqjRPvIedtvr0hnPA8Tw7Ot4TdglFfM3cpvV3pSDb9AULZ27cz
WPXSOrrR+tJW+5uNVdhi0wWAhRLpTXriwt92nbdCFHrtmcuVqnIkXo8e+nuNV3zo
e4dGpOiYJZck3YDFv/d4E5LLp+m+9tVjfnpmx0u+YPIMOXs3eW49OYzx3ZWjJ+3T
VGnoaH8xmKT/nrBt/Q1Y4LdwP3zp/LyZKqvb5/rJvUQQNy0dDXfsu6ieKVFe/3J5
SD+pms3M1je+8x2DuQe+tx8j7hts3FvW6W/faeUedR+c3WBPObX1jX+8zNBPNV5w
zut/DrktGyhrPCFaAJ3lzK9MeyJFYwW6yenXqMj1Wyl2mecNmhYWw9lRF+FO/ZoB
cXvm+sBvJAF+9lnpT/6kf3lA2FEmue4jVxT8o9W8s3Dn8r6eNXLZawcMX3J2vt78
6aU2aGPS5IDu17UlZws2K+Hkg417uQ2yR1RiWQ5mu5D48VBfEitYRkbCiV9kh0+C
YVEomS5THItzPtgESl1miNJn6qglV+Fc7KrJ9b5OoVsGO6hBh/Rj7iGs6COYpgiQ
sI5K+kSHDpEczhq+Sd8zWk8eIwzTHMDhAvZe39zxCqFeqZAywz2dhp2iu70/6C5V
ByqaCiES6d2SLCmjE6iByKIRdY23HCu0mjJo/c4lCNlTdC7Js9UaYEdvq1w3zr9f
M378X8atfg4PlboQHvlFf2zN2S1M+dxauwBO/+2ogVMRyO20wryscM6+40kz/7Qn
iongj7IPSTQmS/J9JIhJBpJsfWPgBqSkaTeOQxYvk4OJ004SOMxxfWHleB+y3L59
jvkEY2iULbDkhS7uJaI2kD7NKlyCJw66DhBUsEW09xJ7oCW7sztHAYWb8VhRiygt
VlstXf3vx7TTQQnaQmXHyRw7aSf+JmkCeb7GcT44UQbxnfej/lb+tnMNQ4eLqSO3
qkrbp8zhsnNM85w3dYP6omPoR0wYeG5orkU85DJKNLi1hu5juVSn7xh+uU6D+AWR
EQuAjy8VEXcrzVuEtLIAM5qbFmBQnQhayzAvhGl9bQD9i6disKfreh4lKkHebxKI
+4sJyyRwDtLwpe3glg07qIkfRG9WwmC9edsFcz05oROrVmfF2/QZoJbtw0jawk3D
CK4RSHdrQhyDdI6vCyYeXy2g0GD5ibKKXK4V0eqZBvnZsWz62F2ksF1xeiGzlf/K
cFkVwq1azdeBTVMkim2K0l57aeL9tI7txXf/7+RvcK/0kEo7CTXyq/3mlUrVzV2f
mLD+P0XkTEJ32VMgEkMYZZkMau7vf4gU1wTCJ9N1+8RrmOY20lBUKjHI6iYqLFOF
VfcxybCDr1f2kyqe52rTPl/qc0v5sLlmODX48FgNmHieARHBRGJz6pxzgYgO1eip
DiDFzXS4cYT+5E0rcHcNYC979zZ89W7Lx5Rtw+tDF93BgMOywqt5YhW0K9kFA61v
BNG5DegVHuxUN8umGc2uytUjf3KL5g2qbtCuk4V3gIsP+xpV4xjdPqUI/+fat9x+
OvjH9KemwKj0+9fJ+WxEbsSGGKpAdgD9ka/Jh5pfL9znHalPriDnD2wFvWY2aqQJ
tWE8/5YiopnAg0qiSU13HIhjD79fAfRTNeAf1S9NtlTjfc2MA/Sm2GLMDEzkIzua
WqaRxZfeYq17VIZlNe9UV7jAW2U6yhjLvvLbeyyJ/IEKHJj0yDoP2O6SQKP5vsZp
TfpLdrI1vT9fli++56UjMsMr/EAjYzX7myJfeUviE0vVCXthpBGgsJQI4w6LRYcx
St5W9rpRN+QnPBkfTZZQhn0Wo6af4/sfOSF7wn963UYbq5vkI+HjPTuOJSxZw5hf
vIYM7mON7af/flL2Hp0B+XQepBUO19LRbYj/Ti6yaD7b16mp1YTTPshQ6rOL7WWH
sYA3KBUrLA6IYAk3B6InMkNRcdISNLMwrtC1ZZ380LgZ2RnxyDo8p5GCeqFCxJyh
IhNFMONLQLvDUqrAXdee6vh1mmL6HFgyDFv9HYiEfDAfqVa28i/OEyf+aVrsmlxg
iC/WR/VjUdqXIyZyK1xH3uzdqaFScBd0kNDxmtO03dBbSbV/XlSytUFLz7AeEcE3
QVb4ouZL0+8qZj+TZUQNy7b/HRVZTeWyxse2Jwpz82vFtvG6thhtNcTmOAOir6N8
/+gTDeTSRQszVFc38MvH1KVP1bsJ/qSfClb1d9swjgp+KhSBkZn1LS0OaJrmythV
hNXVoXny23lpzA43mCeQe0icAIIjtWldJ5AK14L/rzb+Z8iGsTZhUx/zlm4ZafqT
D7rNqE2oUQbwQnJZ4WzwBd0ysMkQ3wYZW8UXUxMcjx/9u0/Tz+3iv+iPMcIXuw6k
PK/tgbWjVXJRIhdbcCCPucUKOfvH8bo9yB913pkuvQb+9KtnJ5Dhaop3vMJIdVcw
GF1jjn7VeeubsK+rVdWb2zY7qdcmXTJkZ4waBusgHbmgkVCMe2Xh8GVwSSm1ex5W
zxT49sVF31kFxacGQ0CqMKzfog+ZYPx8USoTbNEStGMKBAsgfuryp+YlVmb9+DSa
NI4q4S4cPLsdJVuAvIfmPKC3JBj3ha0N+X9+dAXcLYUhxVTJCochxk5MotNesZGJ
rKQJDdI13sRWrwQzR9hyHbXH6Rsi1JMAnNxo4aZCLDJvXhlKf7hJCeyQZJNoe2hk
k6m5zbKmwVxalXAmW0gEUaqKIAHPsV3py08wtRHdJ1NwMrlVGInKkHzwnlFhEBI0
9hj/BdpYepVMAUQ29RCozCb7f+IozzovybGBznvqb9KMzU9tztTIpUgbYTmnUATX
nW9n2Ta1co3tEuOoe7pUPf0/JKzh66PDWqhd0ymBmy+XYG8QFmKp9/JIVEozzokq
05Wez/X2lEiYQxVhYqNo64rgg0gWKNIhQiE64FF6dZ4c4Gpk+XCYu8EDkK9ano1o
zuSACFC0sTbSe8yB364LEnxWil9oJRgCQ9MVK0boiX3im91tghNIrU24NeN00xTp
VZeb70a+OTAROKJwpobKgvwVOJNxD/4NSvIHXTIGXEFBbUadpO+ew3eJ3oydXFyl
MIttCj8AZFO6SQp64Y05OgMr13GoHY6rgLZgZt38HyJGqxjgMFs0iJOsII03raO3
HXlLZDzhYwoOrEgHfrbHQZyykvYJmLlHwR4D2sNLWfvY921J522/3D6NRizm7H7L
1yqHd9eLuJZBQer4rTNEtk6uUPlhSp5D/hvTfzI9pZYvhX4L4VrNJ0uOQceZl8Ct
xKud/ydmUGp8z+yqaj3TsHFGFQ21lO5JVpb8Plkykm6OeyPLLzNH1lj70ihCx5AM
OBdR+NLcCNftNY+GIAC+Yr1p4TA74S3oB+CiRd/lecvJpo3jeSqtga0K93cHTxif
wC6nGTLvL5w/UpiIaeuwMGE52/rItN3NRZ7KLEI+R3Le0xarCMabqigTUrK+VtLU
sCp4XX2+a6Sje9yTsyk8TEZuRUL2pKkj4+tGm9uvsEgUnt1MU/XEUkQi5E/wtk2C
qRWfwr5sPp5c0E0zPSrhss4y/BWsAG0Y7su6jy+PFVHUbcrJHP2EW8LlNbs8SLbd
vhzSZi+rgwW168Jo4ZAR+s+ilFd/N8p3BU+MRnve6/VdLVacOaXKGWezPdhAE/Oh
12LioEFhmTgFoIpMMivhRw7uLgS6TyoS+Uve1We9Ej6K0+twIPgtmWdmakjTgINu
cv5KrqxG1QfxfSI+IjxS9rx6mDL5jld8beso4mee5HuRtu+ZmF9ity/rqGmZG5ZO
fWcx21fhA3PACm1Yo6x7dq2PR5cIkHPJh2PLSosvdnpdBwfTdIj+W/eee07Ksv6S
6gTOuwe0df3wGKVR+w1lTsCdkOiii7Od5Y/cAOn+Uq4Z/woYER0NLtncXRdqpGj/
OjrWKG6hrSM1/gAZylLIMjAqZkGtyr7moWLHW5GBBFL2YURuqvPNLZ/17r/JJ+j0
VrRInzIgld9AX0ER+RYFp5Fp7Cvq2SEr37fenK/DN/Hoj1G8/UfaTdDPTpZDRdkP
jC9dI4JlG5EdsWv+J1RxpaHEoDfhu47NrJX3kjtdkLlsdcvFwQDIaB3EGSJ0PCvD
PzvS/U2bVd+SqU4XOfxg96ckG8CHB/yJWJAR5QfOEdH1prpfHv1BYsAvfJamgMiK
WSkyr+uS5+SLkgPq+0KB7tS5NsrszN5tbIe8LBU0YZ7ZJPKapjV5lEZIs4S9Bqo0
CPmKqDcY/9ab5+9qK8NKw0vBA5tTpEaudyhEQEZ//rHXTeCCZvBt9I1QOdxeO5gl
mJ9hFuqPF5jXxMlnx+chFWhwX8vny+WkpZiy3W/mH7GaOYLuH1y3ACZrMaFDt9D4
HLbMZOjwJo1w1xvzNMY2iICtYhwdTK6B5ev1/uiKcrKSMxtCHCepqoKXiXyJ9y3H
5r5WSKLKn3KDuDHV+pJw4gT5jwW8GEmUCtlyrFxA/TgZ0v+W4XYQ01HaXJgwifkL
NO1oyQUBD1YBOX9m9Nbe8wxP9vszXJsKUhESWRYh0+bw2T/2l1zXaqHQ8asZAva8
tmcj8ws5jDQXQMn/TYSHF6sbONE6lKyIUKLxNHHTTc/OXnUK4LN8kSh4DPqO2UjP
qYTmMJelUJ9NtidJha83gV+hKq4gM+FyntqSq9AQ7efZ9BVl/FUljyJ9872UUeIb
TiLRQNsU5spYlnMY61H1Y3qnlTPtJyhpZy0edms6gha3IrAbgOnJUtrevcpEZmlz
fePu/13lRhjIXK6ynlzhXt+KTxv8totJ1xh9izDmH58EUAfsHThzy5Pb1mbgzYku
RtUW67O2ShT8IWn9jBBMLp/kxrOgMb+WMloTkY6MmN6I6g22u+jnDihI5iJGGzx4
tSMqNvSGyKPf/N8hnsgPE6QAL4eU/j+xccCYkVyh8HNAX/3QU1Onc6JiYjSoR++x
stLbsYVgaGiyMBlg4leTm7M0sfTOeSi9QKrZBdmAed0nmidMkCAzLtVjrlmYggBV
EzyqXIGV0yn0MlULfjJQkXIQqNU2viqQTqzIKWyrCRuFZTuv9ljBoorwNRMJaTLg
gU2M1TtdaOwXF+4HJlbXK/B6uB3dBZmkMpmOZMEvoA+il2XAVBpKdE9EhzKvrHDe
GuDIGK/UNhHjZDkyP3TzEwrvetY/PSNTn7vIuWLrvxzklzUFx5QVjmyB22vUkeZb
CErAueCpzGVCkOZh6njs7b3SpMiUdNq2EZ4ne/EUD2Aa3/jVTG9sz/TFm5T3oYyK
BTEX0K/A5vwoK2I47MqKIPQu94p7HukENOV55k2PjrEFTN2MnBtIdYTD5FWLe7rK
F3DAHJnGvVYyXcOU8UiyroUm7tIhc+lqmtMtzFWUytMaeyNKuMdqiNwA03HN4M6h
EWscGY5Go4iNw/o8meWcqa2J/OLVCFrtEEKvRXfIIFLuE5MkvFR5k5qpQuRMDAbS
mem8+BjjgF67MzHeqLiDDHP/GTWHpAc0q67IybipXlKAbB+trKK+XuqDH0r4tbLj
VOGIxFN2BlgjH6h9EiM5KIUsYgCmzhjo/HA2thMwjSp3KsZSSP0Oz7TQCEUmQKcY
cgxywIi19fudDnct/bbRxNbZn3jWSfdOxr5SYdyM/ga/Zt0CvaG/qXuD6RVndPTE
nMH4IL3PQ7yxVH8VkaGCxKI3BFikXCEyzx5lXq+4OUGNkIXV7d1UZgEc+5l93WiK
s4pVJSlQQd+6J5wfjSYOsEUC1Xmi2bKZfwRz54YsyOsuScohJCdhQRmdfoQONA9P
Hm97AXIm1VqMGL1+PI+/a0RLlLZVKtfxI3UPKTM5MoqZS87hrnjqvi8I6wW7siaa
w06yTVcJ67sNwlNHt/huz+Wm1ipbGs1biBGSsCgAqwePv0di93Cdg2s6iBRVS0wb
4i+LBeBQsIF62yLpTEEuPypTQuI9Ve8Wx5K5J8bNbbYBCpaXqAviCZSMfcHjKL/l
m4zKRHFqm/2rD+dAoTV9YXhu+8CkntUKx/5LCBFXH9+AhqsE7lgpVwf6YPHpk+W+
FByDuQRjMQWge17BJRMzjxoy1pmZjISVbQymyqHoWk8xkUzAgdHDbck6w1BA+5jz
Oy2S6lyn635fkPaD4G0sI3+6UOyaH9Dl/K2V8mubZujY53G6ke8PDFPxazimQEZj
vvuht0jhoOhloMMtew4TJuK4bmAXxVoB3xUmbnVrnq1fDuIqdqAJ3XE7cja+f6xl
jBv+71iS5eqfJyQJeQbJ4QqDwv6satYQKhgvEVRAojzJEjrhrueNIogdf4n0CIgd
my5fSG9tipk0OZFzjluCOlJ4lY9iX9BEXgJ/0NsWgdq+yONZCl0drSDes03YheGz
wIwytl8kjVwAS7Pk0BsihraJmTkpVRCDC7e+bJI1MVMbUWYwO678VqW8TmoowyWX
Sj947duknvX41nORbci4SEqtmaHPCIHHZfYRcXnIi/6iMiYeQvtwbzpxWLq7tJjx
1mLTT/TBsHlLsCRzSP0MqVaUsyq7MSwKIXvPXy+xieyLGdYUNkN1X+AbOAV7ayCj
TVh917eOOfw6VpSW5+sgJbPp0G8Q3jhE/WkXZQdZbzWZDj+jGSqpExBKzA2iCmJX
sKj8Ld/6Yd0DX+cepaKSW2A1nMEy2zYKlWS0w3kXRXbxneitUuhHpd5UKurrOzS0
nn68rnPxfHUvgdRcxAhMxYRd0w8y0b4u3HeQtjNa6Qvyf4p+jGXEd+rSShHIsCM1
ivUedk409wjYn78UmjUuko2qpHI+RhLuDhc+EgE5yb9iijXpVAqrZKrPLqeonrCb
MIh7u0Q4k/96gTMwEvwFtelKVrmvFIhYCV6QT//A04xvb4JFp0wJ7Ypu1IL3dumW
+ToRz0HvpnQtwmySi85dxzQLf9HHxcBMnXWCd5WAwaqhhYn97UOVKPROzZ02Io02
usyN/cha+3psPR62p5uqF40bskHMeXt77khGmK93cdnQJq9t7VaeczNuHAM3/leq
ytivjd3YFRv8qNWPM2GNzwfqmGmFKy6ZI+sSQLW8XrjwG8VeHTq5r6pseWrOwOML
m87l5V5dXiHwkXMapHUJpa6UZX8HBOCFrhhWGK8asj2avwsYKcImjIxeLcUFEsHc
eApqqfeMRrua+LKICD6JFrVpmAP1WrygKIMTCusrKIXlic6mcTUKBvQQw/rCbkDa
jnKhUhihnSMCl9f609HMDg7Ps7P8zGmWeMuHDFjNevVak3EhYNM7LExIiFy4YG6T
6z3oE0fl0jNtpz0NYBUAwScPqJnzNbOXVW+dM4MoWeafHd9mFZxP8ylWQ+xZ+G3x
Uc2ccMv/8JjaJ7T2gu6O37XwTVn0EQm3ol+9xnPBxH7G80i5FiBqR7jKSZmib7bU
ioSxkFAwvIraQkqUGUumw55s74bXFZw0lbkckrrUMt4oogX1MWV+5MD6ftSsnyac
A5Rooi7FVJNGzyujCKKXV9ydlE1IN5JL/lY2934nmNlQo4+aZn9LBuATTYUzvzLP
9YOu+xvgB6AxqTGxAoUlp+bNpX8Yzq2wOuJ9Zmdp9hdyHPtQA2ITHAUlzXIOjbAM
mf3BmQarOlhB9BwUG8DNJNkS3YOPwIw1udjIQFQfvHfeCWVsZsHZyBaLH+BpR9Np
+lMb5GDzA++ADD5HMT8e6sy+uXw5rhaA1kGdLqTNJGgtyEd0BerC9QS0HoAxpfN4
oRMODxYBLM7eJ9+N6zRLR8vlxE/tAl2pEFoRZDShhclsEMZzQe+MLW4da8/OAFMK
udEQPBrSXJr7PGyjXbDAGJmr9+ltmVYcwoYGO5M3IvZRKdtpXTsk7xag1w3N3NjC
V3tq2H4IY1TOcbtiz2MW49mRsUhVYXuQkHbLW+BhQ1NOJh+wfkegtJ6z3j3ldJoH
Sco7jjZhXTB8qFuA8KErfNCuuXooXLqKPj/9EnH+hz0GyahHxZTHZ6G+pcJiYdbZ
5G++uArRyKkx2XyU63zj1EdZwlfmu/yvVrtJBjFb58ISagzcqRKbZW6x8jdmz78j
Zr04b1R0R1RKfCFlVj0RDpTB7CMsZfTLzRqhSg7lghwwcpAz9681QetWZWsIpcEe
w3l8Qvn7zzAG5M3V1MHBEgYsunzsVX8TSmFl44MJdgNWwYt12J+bTrSr/8I6Cpyo
fDCds54DbsMOYNkhLyBzgHPW14TpHRY1Hr1KZHWPwqRcrBC4Yg+AX09CqCYVNfgZ
ps045hS4q3pu2xhvo/eO5MphJqMjgAIJVPwzCigHYfXmf6mxZqt+9t7AvPNATclR
IgRSBU+HN45lih18j0jhXkcEh/lRiBSUWMKZ9m+4HGmFSs/Za0Mm/SHN6iNXnei8
cbV1Fk/woF5rSdK7395b1uWdIYccg0g6xTqLDhoRhJwsdDibRWU61ySVX2d04rtg
G849IjABSaAqDofE03IL8a3FnEIkdI+YEeOQgn2FHMQOB8foyrBjPSD1Eyc6dz+6
/RBznbwBWMZIz8rYx150KBXz5hXu3my0kjqwmONhhzQpb+2PItOyd6gByhOv4ul/
JQffW8z6cRQdUGjZ7y82SKtTodDvzmG6EqxouBVkntDlHtfWs8r0aI84m4ZvXW7k
qMUJOo0F9buWwqVMRaYP+POsoBLke9SsBRf/RomqcZJged7A2CNYT2hWaVdLK8C5
SsGFwQvvTuyuKetiLuJXODmgB4PRmEM0c8Pb5DajacadhUq3eMhxw/CkuPUg7WMJ
TvNXrvPLzTO3YESXir+4ax+rd8Mcn/3nYsZKUBVh0pQsgQRCBGvaF25lDDzu84ux
5iRf12toTWW2iAfNQYcthLmhG6e0UYWMGWrOQ+dhne6Uw5+Bn+4oLHwrKUeDq1PP
fz7lYX1cu27hsWCgg7hGbrdn4Q8wRsT3Kl5QTvo3c96BFC81fokghOj6dbPuv5w4
Ah7AujItpXZpPDerCTcg0ZVLVb6i5dTvu75LSDxqMAkFapC1gDmRUIpzOGgvunMd
Mv/Ys+ignJLfBu1WHjjzWO926XfyiXAf98sfhNEWDeZPmQFOmAqtGEt+w8cR7w94
4a1o4nTCjWI1vyE21bvw0ZdGtQQeaKKrGfAwGob1QIVHG4Z6ZMcxfRFNTNhpGNdH
yaGPBA6/pSpXP+j46oCDBihCDdSis3yRjwCOUV63mtomY3AmnxHGJ2ZKxV64sgN+
KUSPF7VoG7WtpUKLCTjiC/cUp5eewh7hVt+ZbQk90DTk3OOhXCYTEat8E7s0RCRP
7vdI7y3PAlozfLOry5YOJLjPLJ+J3t+j+Nlszk9k0HY/x6ncr6DyhZ/+kSgZOS6C
whGeGJL6U7+CjMMund7aMOBvt9o8df9q513R9/E2CGvA8BZMjr/sVBAArG/tMXDx
LnBG2a8NElPFSFcq0ZU24BSBNb7Dmyh1LVcVbeeJe34TEpGnACriw7SciS0ZKuHS
QsXh91uIMet9XqxDX9oHqL6+azRwjc49CT5rynmdzYIA3daAI2hIWGC2w+hP//oA
mHuwyr2EOVBRMAbfNnpyp1ou3rKRROqTgdESJ8UYp5N0fjNGTUuuJ+cm8OtrmREs
sn9sVfrljmyslUacQpH1BrRsZDgLwb2GAMJBawLlFOOBalxDeDlr6sLzCUGNYe4x
xcnpwWqe2GgYBd4IDI/tASnxF46Cw/SdkJbKdx2gImCFZ0aPenmgbHBeHXqTdDmR
BolPpTZFl3SxwSIxUm8UJTZ4xeHPuS9phGt/gcFH/pgAYohOwRRCLtA6hf1SiaLu
8LXFdXEsGY6Wn5VkbeMQZqjrM82Uy7aiJsFeTtsjLcfQT7LR4SlL5XXKByC4TUXL
Jp+vjDWuYZALDJoJnI+kTr+kM0MQG3n3AWqYY/uf60ysbPC+libVI6HDoz48Wiv4
4qPT2vrVk4KfqBcSZOcCZUkEOtOjWxx2YprRTkSo9oXW2WYP93HOdM2EI+J70sFi
BTPGLH7zqhDhTsPyup1ACh5nYk2HUi7zpW4kzKXoUzynHkTiF1V35lW06gRwxmy5
S3aHAYbZpV911UbJXudlk4hc+RvET6YnX9U9rpQJC4GUAfJEUqtE+SD2XZim5bq6
woGw5bxUT/8n9HcTe9qIJi46UElevijwx5ZXjEY8jz8hewQna70F5Ytf9nImHSd/
Ft+BxdrBJleA1b1nIa9jeRLR22znhUYnFgTdJbTHDfanwYnoRW6yJi1ml4TrI4tm
h4UcMyF7BCv8QY27JLbqItwUTaz4IXuBu+RQOGd/zKj4ZXUYZx6NctQf+XVGNDCZ
IUU6/ozXJ+/XBgLWcPQ9QzHrPjAlCx92/ZzHcEKguBMznXt0Nl8XlABYPH3cqCBy
VZMLdn2Jn3UVZ1fW5IUM7trkahfLTncuuNUs3fkEb8bGjoA3fMImF/LQiBnmcRDd
md9o7PxsajQrj4eZtZA+xC5A2l2BZ1B/G/AojpA6by4kkkyzmwn8vK5BiCxLzsit
Clfk5IG+jtTjryGPS3RBGAQyn6SeHN0+v2KsKmB9ypNgXXjGI+NXr79ZyAEKUuZ5
O8CryBOLSz6eu865/DUVjYV5Ekfah7NI2ouIMRvbAwlsMBlPTltpgFa3iibx5Vug
1uNL27QcnZmyWnYKMB+kJVrIiI6NoPiZKw5VB5BA/GTE/dzRrqfq4/flD7RshMHN
Y8RskCgTAY9nkFKRxxPghRRvXJm8pyZDVMJzC9mP0eEZeV3i/J+hSGFk3tOvomPw
gxHOKSlPJWA+1CCXHAZlA1mt0yTpSejFVranra9lyhN0JxnpMrm7FsOd/PndXZX7
lrxmsE3uUaNI7N58i5IiqmOkY1L9M6+LQdYuXEiHIcYnS6/BlEZjU2emTSAit2UC
8PM/wWPOYGOcsKnieYZfEn32H+pyMtZoDBNl4ATDahPdN1+uYKhRwMahqxqR2xhD
Yhdiz+W98D7l4DINBI++q+828jbrYbBye8O4Ws4kE9+eqK+qlc7GmcLmlDn4U3JX
yWMOTL/zvGjy3LrVQbxrh0PR5VwbF4sTmprlHknwM21Ef421Dl/OtDRoTCUJ/sOd
4BuZFGqSxuhMBUuWlBjhN8+mh8VCnMKacmdzHICYcDp1JEs+uL2aYsso3ZHVKcCQ
+NwLL0yqKb1TpMZWEsardmM0Zzxi7smLFxHWtAOK/0egdM5mCwpfweukRDeG0os8
Wc9D1lILTisZoxck6mNuNVY4R/j/7Gx42BhPtnN+85JoQVYexd+qEgcSzjTtHCV5
Q2Rmi1pGKXG2/0StEgj5mz0mwszFhmjCe78KsZr5lN6KWZ5heIoz6vbEqn2u3K07
rv56HhSA3XE1ypTi+x4kcaxq7M8jrw/G1MqBVTwmGN9RYuT4jOcP9PKKeQEEQxV8
jQiG8Lo5m4iHR83Nb5HRYoV4DmZYGq18YqgIavwXqSRcMsNKKJkjM1Rbg3Oe9KXQ
cMEGITCcnuQr+MMa4ZjFwxj6qwq7dz9QQI9jXQ6O4/kOLqwfjkw7Y8WKaCuT/CuV
/V0zjV3ojFUdMs3dIGGcXqB8QQUcMrdZICmOJNi+PdXg19iV+C9TaETqTR3ZDf44
UstbOo2yp7ek9G0I5iZz/arAkDayJMPbZ16CrRzFtvivKJpI5qB+w4qQdMvCCVFu
Av9OxRyYEkknG2AAScpOTh7kRURLINd+eAyb/fNh+xWsUpAEmx4XXZsln2Dok+uz
+BB2Bg1y7LVNEHrMXMewA5PUWnimENJiadTdb+MarloUbN6WRLeIsayMfR6ZTPr9
ULOksvac0ba+gFaIBLrikttIwBJag7vMvgUPoPEbNUYRBeX83PIgUOovJA0ySJdS
Zql06L8UTuKsNRHGH1NFO3W3NFfO/hiEnawkNuXfBmb/LYyYEHDMjYghKwpyS1o6
K4VJWnq1Q3Fs9f1LqGDwOm+WfmGmNCwtTUKMf2+9DfbPspUazrrHJMPfjTSa+UJr
gVqf/52W/eClefKibPYO70LNLCNVx3D1UKM+nJ/2Uk7cPeBzi05PSfuY8lmO3Lmd
IPX8f+zO73mJnSpYaoNBhKEeeI5E7t+oDsvldvYUzP48tKbwtHGZz0cvhrlWdOUz
lqwU9OBGF1SAhVAoDNTdtXVY6QYYm1IbNwVG2S+gaLOQvFp7F67r4nwyVlwulfEs
8gTuLMQOrMB/o8Iz2p4RL2c8J3sD6m4xEnlIm6Hf6ZpLoqrvQGiK8K+Q7uF01nQt
61+xihv/6kqXJeEwt85kIq/0sfDo+MwIsSZ4NFNAOhuC+5aoX2MaPbz9iO6EnrE4
gLnD1WORbsLiiHm9VNB6893ffMCv9e2nHswnORYY+/i30qkDymSiDGSDvEHYGQKM
Mv4mZ2yjKdq8eO3LPUs7T4hxtnYXRJrNlJAs4bC8/O2CQcvmACmOPUPE44h7/DjJ
hNQQ1oV3ka9fP+Id/c2EgYV5eozmeuxG/deIk3LNmj/LaHPKoO3MEtw5wk5tCBJI
14tgrdJi3enUZv2GgkEneo0t6SThEclMYfPyJJALyWoRdhuEbp6osFdDSKAe3USE
sz8piPnx91h9WZEp6lYoRTMEXj/tluaeKxt7N0ID4ZJLDbuzWw7y/sVc5s5Zjdnp
0JqrUU6qnDrqrS+MACsROt8Rpo1sy6UQnI4cyrYbczTro8L0/OYTsXKCWJ/jDQwl
jBHUPX3Qz5tMA8kR9qMocB38qukgj1gM8+pOAmLciBRkZ1Vuazh8vIS426ceFeoI
4BxMupYzVQo79WSTTiaIqVr/d3B2LqkbkCmiLbAjHfHVSWAEBNk6xaW1NoOMmFPN
izHcWtyFvENlmrF9mcboHJpv1tugqgGVCb85Zgb0fMXDUIV0/HE1TlOTC9fVjUCK
/nRvOnsDjH2eUx8wnd17vSsWJFE4z1MM3jYSjjVltSFuVotZ2rHU2FSYiI1wbr69
hXPfZvcHLaXrJVUqE7WAXhatjsRCV7oXJ0Vac0RQpg5tSGzvyJY3QXc08ac4bQhq
L1l3A9CaZr8t7IsvDw/vymEvA2hW28PfGx9zLdTq9MR2ql9NLVKxrS/U3PbAZmAV
6DY+Mm0EwYQJAaxfNZ+EYGeZI+q7bQPr8o5ec3sPzPTf69RkiwZrX0tpedKMQrrS
syBbTDunXLkyMsihj6LQesnBjA8m2OIfj6E5tSH8XDA3LuH8CCJQUlQREo43ykx7
x55o2wXD1wDHpNkDwnJTgad4qYKVaLrvs7EA0ASajgVTKa/4X1jKaRrVzqQTp29O
1xAcECyS4u3dY/RiHsHSmYGB1j6oadgGMIQv8zMqsmtLN5XfDTT0xPVpxXQMGp3I
Qvk+HfnHs5LJGpQKXmEEiENvXo7IDM4aSEc9rvAMblLoJVz+/UYGJUVDbHMZJVMI
Noumgoo1RAbJqasS9BTays6TkPMEYsNejKZSDjv7NxmMAe5BNMPcZPvA/18v9Zi3
4nnquWSzsLDSzE3HQxW6nZWb/FuSH931LZKPqDTC2JxSjGA4A0iidFkbuIG16g/5
UmtPqWWjBSBybJ4WhA8PiYhAi8UPvfroJfLBQHsuWZX8l3roI0D/s7abynASvoyD
0eEhyoEnJuQ7fVAQI2lVIRCqp5bN434KIRDrpuob6GZWTzSCMZSakkWZbRSM2wfD
gfCjKlA3D7J7NWj4wx0A8KzwSTF6oilO57D3h96QbQJCyw7uDi0mUVpgDA3r5+ca
03CS5nLlqUMk621RYf7c20nnwERiZb2uJF1IG/gIT44r68nkxgw3SAu5dwdnkkP+
QXWqchTzLQsdtYYfhku2X3TKl7Ig4p1U6wydmCCKd8vd2VkM4vKHz5RRVSuR6Llm
/tpVgBqXv1PFjqupur0J6+apwV+kGknCP5e83hzn0wGZcjkNIbBz8ReI6YFqHgcd
JVtZoTvpD+XwPgMGhAVBE6e7E2MfqKKHhIME0FL/qtSoyHfOjU9M98CklahRpHr1
rWLDbYkaWrRDXOhQpJUrz8Hy2eLWmO7zqAgyvulshvCviKzbsSTFBAi4G+dDcGMC
uvnjH+u1Nxw7JH6GZt9MzB0ivUvXMIo1+Uu+fnJnlKBBcNVTj1hbE8Wc1Nm8/YN6
rWCi1EurYfcqMkZLPCLxNjKIkZIwPbwww589RjHIaSvU8rZGWVEhUsULtEDRA2A/
9YFrkwAR08kQe5dWib78GfZfblEVT5Nmdun3zKxOtuphYcnQCG8p368ogQBwA+wl
01yRjdOPCWXGAHrYnSVzxboVFUOhbJEYrhcoup3ZBZwEpEt6gz8t9p/EXbG+KfFH
oFQYSnVs3L9/t7skY4hi4fY5tc8tQc0mzXt82+buj3gsp9WrM33kB+MQhhQ3jA9J
TIIB9qOUTVJsOmpiRiqeANS4HmOZq7j6Cz5Y4EesrxBkmJvv8FluMGOns+E+3N1W
3TmofThql3If9r2yzY2NMgotz7B/71ZQFVmDJIUoy+3NbJljnESCZKyaBJSF3p3d
AfGopYKP4WcbBYJOYvlWtcS9fLku424CmJ0BCRR7EIg9J3wxQlJ0GDbaxMYqK3R1
bwiw6sDt+elCfVOdP5kt/hIOVdQkD6fMU0OmiF8Ov1kT2wRqI/VuffXIsKqFFNqb
IfSboOJidTm40jZv5QkUPEkCbflVvPbK9eGdT4ehkfhL6xhyjMwY/JYP4faEWB8P
OShFrg4/V1wQLlxiAx+JCpoWksTTF3+6R/gTA9bfzic8Ra+QtfHS3ZeQ/vgjKkat
pyxo20aBcylj6TzQD1viRIWqReBusHDtIFRqSeCz5BDed03f2I9YhXTsLSkXs5D1
jOqYk1eOE7R0AG5nbM3Z8ueOwszsIzk+zjFCLU8ILjZa+XZtaTepEont1FLA/vx+
X8q/3LTNrGNO41ZteuY1WevjF90BAYfYfT/lz58MFnxUdDn/UpTOyOcC+yCDQN1h
fnygl9rRUoNLf15/lnjABq88gWcEf8Xe19uHiuOXW+8eW3N8Qiu92RmSVcQOfTFj
Agi4dd2BNVGb3E71SIzQvF3fymEcgJFZsPSE7WE8mU5l754//fTepx9jBGHVuxsi
K0arTrUA4zSJUSoHFmzfaqR5jSQ2o8Bg26mQYowfEZVdAYAVcHtJersG7GqmQF52
y2REntcDo9zIwjyd616kd/7qQB/yChs6UxuBJhSBkvq41TC44gtUjonUoLLkv0Yq
8iP7QYg1uVbtTZMqoD72BwF5Hy2VRyBRrNqy7ow/D3zTdsMdJ3Aedb5lDRb3d/3k
uaqXTBStrxDPzctpR3NeDhJfz1N4jGXg/VOYKYxvnjIB3gXS95JdEJjK2D4Rpzex
/o6iXEMvCntzYGJ3YVbAp9m2wgiq4TK6s9CY+1GVHCbAQ4a7TD/Z2hQIy5EZ4jh/
e79FT1ge5TEQQNwQsVLP5hL1pK7rLF4jFtJ0jNh29QMvMgUAgJ/XDL3uTBrHm80V
kRbOtxZmmD7t6xMBiUJi9igtAPC+meznFJsIkRxzxbpGamp9i17RV5NwCHI6EyQw
C1lonMfQbdJr0S7dNwtfu+C0vO1TmcyOwxD8xbC1nIfYM3EOAQ1a8Cf75jOpt/Gc
BtcqpGcj/SLAhnJyUfpSypK/CFdNJ+MZgolCuP2NahGO2nAbX/LRAEkQTO778lX7
ztY/YG7rORQbxrz0PIk9aiDhd5NsBOUhYx4BprOsoOonom406snOhVcqMLM+Lm7+
DPPulxAeP6xR3zoU9WT1gFTWuHBKTjMmOPKTLsq6CoDGRzvKX1luUMcby0lBXGob
fE1yErgrkfwdyI/zV6hlUBEfkJMR+RY75z6VCiGSjfmLIxPChfEIHbRTv3g31LKX
x7c8w1M6rMg9jWJPFqj6wkzq4l1+gYsfKqhePJCr7W5MvgqgJARDIvEWrsy54LYa
Y+etUtZ7tJo9WTggH2WF/5f2R2FyZWOW1dfGbJPMRKXY69m6bpby3qbTC7/ldD6A
+u/BsVLQf0taNazdQ3D+5uB3Pnx+8n1GQmCRwlIWmRErYU5nxCYmYZ0VQJctbM65
2kwUIsZsWWkqS7Is8l84NJwzNmoOYI628jQ/1b+UTsy+dCSZIEloACI6cRx87pfp
NcjLYkgyokpwqo/8XR/FhhYRX9/7aPpB0G/ZaBfy+/YOxvbqMXmE2k06v/C07Phc
qyT4PYIt9lw2tv6CaB+h/T5UN/JxAEMGVuPzV7fS839oVkuAlSRNAxwp4vQhmFJy
oojp5Ok2w5HISHIDSMDlJJWJ8hI/G1yiHLBbc2gtbdPO1nkme8KuUpSZ5CfEWi1+
3p9gtPBP1zk958ZUIJelt7kALBKyEz4qsWnrNtfl5BG7HBEJacfPZRDbkcIBUaTl
T0QdJ85OBxADaR55439sFDi81xWJWoJ1wczm/ExCoQ7CX7B5/rJm3faUDuX9C901
zvjVfE3hkCrVeznCIQPrB9bsiWP9453MBdydCORQIgsLwUt6SptHofC7l84CMIA4
qK203cO4zHvVAXCo0peZy57rGU6LEjgr9BagSxutb02VZSmrOLaL2cxItFDYVRcS
wxsE9udVDo1FVdGs7Gcbu1tDUPX7i2t99jtCss2ttqC4vyEq2+ZYHy12qFqi1NMN
XkmyxS35mMA1Me17Wo3kg1VhfZb/cI3iH6cN4K+VpTRxJjnr+tukkeriF6crGBkl
YaC1pFHRNBKRlzroHkk8J4zB4XiP5BfP4wJaxrbmMLCUvy/reHN1/BJO7jBrW3GL
8RVRgRhe9tQJCjvE9+FIE9yYn06Q3EWgab3IQSkoM9jFoIdVFiPmMRc/hj+4OF14
QktSliTkN54dCO7WQVpqAu3LW4cBmujWGLeS/54PCtSdNiL5yTkC0HO3hVceKm8r
JbOnYMxxf/HNgSqEZmlKHeIXC/eyM6VxrhLwKtwOZDji8035xhYEeaDWuCZ2E5ht
+VUkz1GNSxcK1SrvuUPZegTFnOmu5sAQbg6jSOMgMOJPLUgWZmldKsUfpaN1aAzC
F5wZMmoRrUnXF0btZR/AdrJIFbMQcGPwcAjJluJVdKGZz7z1ugCl9rWNbeyROXn0
HOoQsACMb2q9lCPTZMR+e6rbRXQyPwcan6qFxVXu0cqIKkHmoDF9qxIaPNta/+ld
7Ec+6oVwhd/Hih2MalOSUZK3LG9eKKSRUpjrWF0FZaNkcVNxphBACrA6hEu8/XKb
kcNoKISotUw9Gmr8+fORHq3A2mBKKfYgwOiCMWKAi/bMoGN6w3XsONiOk7MPnQWZ
MSTQcw2zpy7JbogLO6RTQQikCa1cFjTXDIWAm03lj0VTxpQBtnDBO3+WOSml/mG/
kD5Jr7s6OAa5wcmIjoSxL1JNPkgeSnzQ2u7c/5fRbwmgTJk62q+ZfDvkTKWsDGU1
iN51vTGMgwnZPCoeGqONxuR5ZhY2RN1yIdgEBkY65kCdxwj/mKUbaDHZrOHHBzFD
3zPYsKEqADtVCf52woCNChjNtbsp6gtCpg5U6Hy44Q9UsHQ0t/VN19Jz+e5GSh8R
aym6j9cBb5TMgWBXZyWVHqtqP+o4JcHlQEoJeTqNtN0fVi3sKm79980aO2c8a32n
ZkVy1pp4HlaDJzVAErjKkKnh1E/sNPinh5Md2n9eWVK7+cMpIdkFxr0YFjBgbxrz
h7wUM7hDGAjijx6txuxwM1Y5ySzb1Gk2gR6aZDJ5jC/lE91+Rp+8Pt31tWk8Ff2J
qBaoRS/n3uOIDmSszghxC3i5u0me6qyK9ZBvECvvnV3RJBwyVH7fwRbGMwi3y1IQ
xLDN//U+LnmSSbkRMLBWoJXEvYfP5B1EVcWZlhpzj/LBwv6NmdLHNLMw0DQ8i4k2
FRrp39sp6cnd/7jhPps34WEXnbIoTSJKx1qIh5RQnS1o8lKVtEAqWJvIfg95c1wr
cDlV8DxYHZZz/wqKep/pAN3LZcNk5OkZ10dbah8/x7hVaxfRca9lqyusnGzPMNgk
5EW61BA1KfQYF1C/k+/Uh6EZcatITUhNM2nUk8Lj+6GQ2L/A7TfQa8eldK5sFxJb
7xJxDji579J5uBw/sK5tYKMJgfj2H6sl1B73EepB8WOImuHOk0tWPsmxwkcKMluc
v0Q/Yw9KdqhaHi7U3UZUtX95OzjKEBojjf5eqs24G5Pl9MLSOgeN7WykWFuvR2D0
/Rib2TMFoqKC4Do4tapt09zIsNMWQ+52B7Bfp2QhLukq81LYuzwGSF98vCpVAuit
o/lIN+l89RDcFB4I0IgCak/K3+dHbHTrLWskx+9ZmYAEdS/lRc1HEeKYvCUnftth
lX3wI9y5uV52xe6m3kPx+OeYC4o9cxIzVkxbmQxwrykbvb24nKmPzJ7/1p0AShto
16rnH1fUedoKJ/2fL4UY2gYlbnJo4zH2aWa6XVyYlgipFatu/SgeZ+mcuSh5fmD1
RXCsYeTzUX3QAolraGzUrsds8mPwvdkNIXVokfO7w86tAn3dWl6Bh0ZM54kj8UNn
FpughSmsX1IAnoIqw5fRRy5fPsMIxwL2NGeZmOjc7JgZI82VAa6jZuytzWGiUoZe
iDvrfzhFLPIKPl5JffGvamrexbFfbhaOUdtG+TEpwBCrakcFWhW2kZQ5/cuOUBVH
D7euI2QoMjWgJ27Pdk9rnm6K4Tyhh/QY0AENWTm7aYoRu5xUV//IT2UkjSA/urs5
UM+k7aVIuM7tvoQr9GHyyNS9YZNaWd+Y6kRt152J+I6b0XNfm52YRWLyjzR6Iybl
D+wpnltlLn6WTUkK9GU+2x+5e3YS2ZYPCVlOIiIx3TsPXrikriKG+UzRCZM8+DuX
gJGnTbxsCDRn5s5+Kti3vOo2RoYkIOEfzhAWi3kNlQK7Qhj6fcY5AdPcS1F6qZit
q1qnubiQZiVy7Aj2i9C4lq4U/+U5ZWq4JIaLy3pXQrEwuv5S6s9SM82FPAU+7z7z
8QUy7eVqQWtm0qLLiP5MnNnuIs4IVw3z7SHrg5jSLvvAbECRnfFMeys1PQzw8aNH
Xlg9eEUGFO84BbBzg1/9q0ZfXAywxQS9xEmAnQwjGVf5cX2MEV+u3QkjpMaw3ShN
2JEJqQ1kn0XhhOduX7C2chjsbMA0GGJXZ2J9Q/tbc3aZTW2iwumZGfUq8cqidafj
+55SLoc+qsCiF2yN1HNi4uGMKK0dH5xRcGoaDpPVEISQmaAR6jBvao1pJuCzr3i4
DqHvn/D/Vl2oREbEQMAAUBSKOMOWf6HMO1UIvFIroQsX1UM6mJ2V38OEjPiA2TPW
3NjD1uBlYuOU9coXWdc/Tki9RnNdSPBGSGV35QBd4OAHloLis47kjrrcksXzCLld
pky7IBWcGQYtr+LNx+1UPexblRRwJe55tEjbRkOVeoZ/KQYE8iWx0BctLJ1lGtE0
SK7WAKcFYNw9A2avA+4OjrpCG//OFf3AYvfKpFGwYwhDyrfXm5YODCnjXEjX28mx
KIolz4MLjM2sozsT/2tcNQMwZemRsaMQpZQuTgN6jQ8rEiwl62tTf26jHNfTFLLR
ieizpvnGSaMsea/udEkpf0iBQJqJZF6XWRzC2xb/1l93c73aOGb28U89gi88D3mx
UT4odOW/avB+6aZUzWjZ4zeUueB+arbZpndVBwulIaIpYA6xu595s8iVahhmaWab
GJu1klNusyhhYC/94wy7roP8FhHV4vnZZE2+hJdCg1OZO9408m5EP8pySyq9aDxn
eNVE15DsG0ozKqAXIm7YYOtAE8YLaNwZk0E8p+ylDy9lyz+WH7A89KoLgQHx4w2h
tJmpo5WUKCXkGUmG6jY40O98FyzuCus6NnvobsOPbXmu/DpYOXLbuIakZHPrtGW9
alwg8zDrl4SYcKaC2SeoJDrzRf3smh225KOGRBDhDVB702P9y0s9o7dRn2mlZobW
yytkOAcqS1JLSbRjDJWSNOT8V3qPqFvBasIOsiz8T6txGPxafD6F0nGUPcqVMcei
p0xlos4FCEm8RkrE/cdMEXtutr7Gu/d0ykmyLDEZJPaQVfP0p5gFlltSRMdGoh4S
9RykHPANTDot94J1k4OpNDkFMmbAtUUKx2Jv0WMABCtPh7soznS4hc0oRN2AuaXr
27XiZgCoShivUjuUAK4c5UAMz5yFHxTOw6JPw/6onzKmUzobXXpHv8kJZdWg5RpW
E5HkS+WdKOUUb23jbkeZgkE3RvWqmdDByndLMxDv9pKtJm1L/rheu40brNLngF6Z
XEEKRWu1tp75S9Ao5WIwsmBzGRfnLBmw5DyI3mB4ZbUhT6T5Igdb+W7EkKe1LRQl
0a4IHmrI8eOYylwqSeOKtF9p66Hzdfq6Ryj3nxJeoPyw/Bwdt1o4kXC4R0HZbdTj
O5n5qhY2Ceka/VCOeY7CGJM0AL3ZXcthHDRix392QrCq0zxcbPHT3pfcNRcq+Nbk
kMcB4ftggoFN+84dd0AD2lhujrAqdfstn/CZ08eM9nkezsyJKNZc2kEQwLEASzPk
5aEEum6Gz5OcfIZbDypw51p4XPqK1HkqRitxEbsATgxE8iyBty15Fc0cJPKH74S3
iWT8KIzyffyH4BkihJ7RPS4esllSLOMv+MZHdoRbpiPS6Y2cgg+ONgmIw7z1VtuA
eCY9E56Z7RZnuK2webfux8efIthNeCGVITMykRv5t6n3ee83/pKk+f65Dng/lyuW
PVH0dStHp0588AQRhFdjxa+iQeJ5lfke9CH2OqVsanInw/HKNseAS1KhfuFGvFWc
ydmjsUXd4/t5pYcZhKuSamjvhONcAPyzq4eOEEajj/XOzVxmctNWcXFWXV+h9h2o
do1WY/n+K5o9Wd7y2W4qEvn9ptIvKlmHIgrNOW7bZqRCNk3zSSnYfcydmOt08ua6
Ep4ll8WxohYJ2BkORs8DWmMWeswsupr5YoiL+fl1M1uWhMJEJ9PbJt2HHfsBia0u
0uUBDBr81SESZteR+qIdDsjp0dGdb2ppuGQgTSLL1BbDQZIh0eUgh/9rHqqdH8Ev
pSlvdhqb6HWodfIuQJ0F/WoL7jBgd81JG5Kt0xukVF13SeWxvZbI6S0vG7/QRFNh
`pragma protect end_protected
