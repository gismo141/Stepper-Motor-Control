// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:51 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
tb6P1LrkwPaC6jzVr7hFL0OvcyqMerJl8D0EMtGN9qPxF/DeZLUAL/J/jaDF9ssC
6RHXVQ5iammjqjW28/pEGCu0NE4bYM8icC9Kobcf9iCyLK1BdNF5LUOEuxoCO7X0
u3hnfFMqRqsJG4Qec3NcBJMahZu8rvd+8Dm9Rf5j3h4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 58368)
RiLchdnhhXW+KDrfdCApNjAxm2Qz8L9GYyVDapy+z1SJhTzn7EZIamigw3SgNaIS
OuRQiOmLJaYwtHAXJlbaKiEFdmqo337Xhp7blG74lkw3DaeDD81SS2ixcDJGDkV+
IkQSz3E2hl1H+wm/LQbO1OeFlkPx3ko4mIbfsJ7NzfpiQ7HyC2moDP+AerfNPcOF
SOMQ3ryxFBU6a7Sp70gDmXlGexbwVGwJGVo1daiBI6NkNw7i14I40LWzMOFgEFZb
CzkW4znDCrHFZO2Y+0wiS3mHVUbsNfPgs7sE2lYiGFQeEibt5xkbZmhR51Bc+iNz
TzkU6xu02JixrNSxyYMEhMYQXoDQiLzVA7O2LLQW/9eA51OuxbNBvDATZ/cSKbtQ
rI3cRel+h0oW4nbQ355Rv2p+rWsKPZX0m/nSeo9XHfdEka914XG3ri9h3laaibCO
ZeqDvEiQ/xoQbz5HqEJaQAeskR78clXL6cHT6hpbU6b3O2nFl1wFcY+U1am3ypqI
sQ+4Rm/UvhRNYjXliyN4wc6c8X8Axq35YvvWfJpfpn6hTJ2NCNOlGbqZ7uRfjmCy
gysTQvXsO/q7XaO2AJsZV7OMKBcfJteH0vZY04PrP8aP6dp78LL+RapcPDe5fp/M
hN29cwk16BwZphBklrWunys8qEgVPYxAZdLKUYRH61kK2/QUIsCwLqjHFBe/Qp0i
V0+cgsH5jaId9CWS5bZ9niAMpNLPfVRi5zTsH9FsL62b5cHA3ffhO97uX3zPYvlf
VM2DbS+qQNd51bfTRU4t2ngsE5xdHhJ9tFuHjkw1KwTov1lkavBgT8xRziygJwo0
Z2GB3QKS9LvSQlfRKVZV47P8PCNlJ1DhybNo3eQD7M4s4838I8cRAC0RiZu7ebhD
9C7g/h8aC/ujfXGm1qbdNd/0NZLFieO3rElaC585ABAnTMz68mHQddKbodAesOz+
u/bmG6thSgFW0oY+jwT4RX7GE/Po92/6HyLxd6bVuMmNZIGX0L3keX/0JOrTJF0U
eLadwoHmiG7TP7PraGdIbWxMHJ3vZ8C5lyuz5JSKs0eVdnl/jMI2ewtR9ynvuSMo
FGQihrsrodC+oOqqtN6d7RXl3lzNP0Hc9xeLbzoTGbQRaONwBCXPJiabTeEpq7nQ
jol25Tvw5AZTgMTb/44nuIWJnwnX/Lpk4CcydLleEA2Fq5cGgrtF9ZjEM+XBdHD3
JwRLb+fw01pP01c0AWhlWG7akeBKJNL7vSapp90hmbh66uwP8ZyMQRQxNJl8dYxP
n2y4lfze+fNNL2cQ77GLF83Y6IdT4frJpw68W8cq0UNFbUEpFyGnFOHPkmlsDt0+
5VgijIVqzmiT5XFoKMEGSytq8BIorlSL1LFgg5eKWwuKg9Nft6q9gqholeVmBv/T
kLHOFFoFWZJRE2qP+Hixv6yM5NWBKVnykhMGJvF556Kf/0odQfzXBK/Qg48T3zk2
3kwNhClMtQuPPHFLfdQ6m++AE1RezeMSft4GZYPb4tPN3TBHRwLv8J/S/7XY8jGN
9X/7naUlFSBgIP8p7OMPtlE6htVZlsSZBP9LWyN0hvCjAAda3XSkiIjMXOBCIk9I
AuGtoCp8o0DZccatNc3HaP06CLMscCELcD9sUDBbyNf/E4mdybyZ7XUKDkyAkvkq
ZmjmYJakzSf8IltxYOxMDIfRQfWipdAmJkwLHTGhd0RFYlgeKT+6Tj4H28E8sD26
q/q+f1muJGgbaWUo9IhXQXy5VMV4R0ClR6kvzMa6wdVAnbaPG2dPkl3G0Or5KtVk
sxA4KClqNfTbuVnJt6jBtYVC2jS1kCmvS1qgbTJuCgzr32euyMOfAeXU8vphPbbu
I4pf2u/J/O56FXL6ztCoUb7NX9puJmltzkBlYIKkUTAfp1A3bYM60VZdYkdDEwDY
BYYYgfGRcfhoa9oCkdjPVM/IgXkNjFNJM0IQJHAc11sqdyQd4xG/9zq6ejSUHNr5
xkqdPjgtalSGct0YZSOyOgH3Ofnl6G0eJMwLWMn6NHmjUf3v2asfFj30P990iqFT
xkjrs/M64P/0jR7HnDG5AL2frJQDvEXTuy4oZPD18jdDVeJkonBO+Mexd/TI/1j/
DicenPylMUYf9Wxtx2DWCVE2Y2WmrzBxiDeGm8h2XVIj2kxCVsWXcqsFkeFhaPZz
ZF54++GbB6qJZ3V1qwcBr1tAacGxCNBfJdP3/ZMxqYnXhqYemCQ7JOQENkasdV+2
VmcUYC0Zp0NIlzH0SOjZDiG5IjbGyXMj26hkveAPuVKmNXBCY55bFaI5J/Wxna9N
NnBjVXdfl/ph6DdVHwEQCnUU/Or77O95q65lYj6zkKcHyt7/VUbjVQ7ys7/wCur0
sdsVl/hw517t9SV8LxTTtyCD/5XqB7ul2QskA/6nZ5uKBjV6keoZYZIfB8zUbHVm
yLV8361OMCzmsVG/+Mo/iHarDwy57Ij0l73Kyn8EnpfMdKIG+skekOBqo85r8Mel
H0kNEOL5MOjQSPTXyQDPV5CaUq2aT7nZNz6ErmKgOGGLHmikzLa2x7S/4jtpXqao
lrjeTTmbextNTZ4TISTo52tBXOwtBglVJXWPoDLjNJK7GRTgiHesU3RFqnFr9E5J
bgRzFarNMgxACXW8KwHIiOGs33lhRzIsBShJI6ND00ekGe9Pwi5c73iR820DfXLx
rWfV09Qjq7ch+spusEzIO5qpZsdBVh2va44BY7dbKzTsccUsLN3bBN8yPIav0xrl
gM8x6eg4Eraa6vFWJdiOH1kI6uEDhNNxeuht9RPVn4Eo+R0DyJ4l23FIPB/VSMRq
YLyRPm7cQWX0RMkQAjwHGRsN1cWJftKsCOc343Tdvd+rr0AylTuQIGkPtAQnbsMQ
4Seo3vORvMidb20a9Go1gZMSttIUINPfn+73z8pPW6Xtr31DNno2/uOTeRPMAv5z
EdXRpe0CKNK1J4me7eAM2u9vMEYYBgWI61Obcuj24eo2ZSCTTfSzd9G3ze0LLc8v
Ow21dPQezL992FuiY9D2LAO1gqZv8a+L23LmZi/WVG3CSfU2sxEHvokdc81zd9cW
0JIuK2GFzgWvxxAw3itR+LPdZlCPK/q91d8Sw9WbbOrNmJbHMmSNRg08y85PV7D2
GftlxktM9yc8Hy7OF7p7mr28KLjIYAe9a8/74aLLQbvx/a/CU/ekvr4uJUeWVuJ6
7AFEY1+H6CbZ7/qMEPAk1LwbaPPmQ8oXaW5koO8GBK71HzD8RglLw7+2U652U/gK
2TytKijJGxU/iBfbYjb8BXvYwHoS2oDfqX9Hofz2bV6057fQTOg7nxz+oPJenAok
82/nIvUVIBHuMvup7iOrlfqZ3QOjTGaLJElu25BlGb9jNn8PfhGdW7L4YsBDDG4K
Em+9MQSwSEZDUJXsyAVhKUSqfTvvBuZVP1FmJ8yuwQcA2aHzSC77lGh3I2im7Akd
mjjE+8cxVVOkx/SVT2Uh6KbeOwfLk/OTEqjtSsx3G3OvWzOnMPZkt+TifSxi5hNu
vdhVUrTjcaO4zYLENjIHtz9zcHjcr3EC6q9pPiWrjwRll+2p1OElWlzcwlAvRywc
mLQB/qallPU4fdCw9Ji0OzSQ8X7k9VWFpPkw5Yz1QJikiuEMomKOtn+M2t0ePFLr
WwOvZ7t6/ZG2YuHIGR03/0l3wKSaAsKJ5dyjjJDjN9MVCsbrjHbbwF9zW698soqO
1WKDztoN+UNr32PFoWO2K9Dma3ksLEnwDI6YzV7VNtAXt13hp3Po/XsTIjd2WaM4
MuBowKMK/rRdeJ5gyWRYdSePWRce7fZ5hYehsg3fYJcHGxUF/ym7lNcu7jp4993J
zQZ4AmmWBsFYoDWcRmohQOUQGiQbPtvSA9LFLrzugCMRrLG4sPmtT6uopkIbOtLl
lQUaF9bNA4nBOZYDPQMV8J4H/sBRpBcjRbaOX9ImmDD0nY/mJnU0+EJRtF0INWEF
Xk0huk8fcRRnbWW0Fgt1SD5yzsFqM7o/vQ9DQLI1iNpyREK93NdVXPccLUqUVNic
qGOgau/z/bILOQU6tbMeNksVAVugk6pSIh0sByVlZgRy2eV7oHqYPjliL0GMccFI
2PjYQ0KppT5Hb7B6DKHfYo6lZFFCUiAQ6mB1JzRJiqJotTos6NwKHOBHkPpyXXzE
vMO0/ZgPA23OXg35RiufqaTRXw6zPyCt87zytV6uWopFnfbwuk4y5AiKCRkLROYl
ZHhR8r8YzlhU8+SyiZZT7eloiUtbVdABX5VruxY+Xf462uQh1wWZYCsV6v8zu8//
XypWcfdeckMzT57HwOTbbbbEgikBDpG9qg98jfcnmuugvGuyFwO9dveSa3aqST/9
/YZGYlNtCTrGhSSTYf+AOKKAQn59QIgeldS0fOHFa5CfDnPIXowm7jmfRZdPwAAU
3zp8ra2QBoaeHdzwngxFG67CHzjODrchpoXgYYKM0LgnTA1scxRoOOUwk0oRR5Yz
pQMNZRd7nHu2DB2ypuJrwYZjJhr2cCGbeEgOXqEIWMRGbIxeUTeFmjJmHYbLXoMN
x4YZlh5LWjFc9tPbrdqcyfOV6jsSQrsLqC6xnZXfAXjhsTalmkWPB808ysFAMnxZ
WJFg260Mv21ZWfi67COf+5fqxwb/fRWz0zl92YV2hSzIkRPI0tSCOJtb6fzroVaQ
ezdQn9RXr7pJPcjOH8R4CSUOyOL43FUMWDOt1z43H5PhBlGW1CGUI+5OBJ8aGJK8
qinAhgY3m15f7aasT1a04vbOhM+drh/1+HqKvLUGPs6v+Dh1C/k/8Yw7ncfjrgpq
DW0lqv9yLh7+slYuS6b8BUUhwW22XABLRqPcH5o4x5PhHL8V5KaAxbA8p7LBdRvl
sRL8YbJyEjch6kt9baYLD+It+a/WFpP5/qLH2s6oPz5TewAN8NevVD/kqcnG9l7c
v+9xtgF+kXuzYkRtv9Hs4LSho7zVwg1YYA9Jr6PU9sY0okbUWoAgSQPk8UsAFpOp
+EBOvpB+eJRWOoftjLDUik7+2Ms7ztJwHDB7os28qyJOTrU93gIlTK04DLXHwrZk
P04wygjD3wgiJprU4fCINjwMqVLGrD76TkGAFtYxPUJvR8R6NTfsLqleAm6/ocJl
nq9mDbUZOTX8cCEvHX1BLS1Oz+AYq0+fyWD1uy2z0wXXNqTkF27UpdRi4t8KLBZL
gJ3By8Vy9brKXPYCH7p/bMZhMW7U4YosK+t+d1OPmIaQPGL7LgVYDscRQjbXLXUa
n7wIFRLzW9Ygj78XW/0IgFjTyN5UettCI9j3ezY05cdy+GrUwiy3Af74yVpcWrCQ
DTDhAqmk7F6Tqp/Qi09/4eih2wSgV1MPHJ9+gobTx6vxCgCvEnFWfEMgJSmZuff2
H9nesc6K1RL4/h+pVJdj4O3aznMDMHLD+TExUONAF9QXufKZpt0rTNRsn4KieYvd
hZWIOMSIcCl4BPk8rv1ruO+p/wNugvBVjkA1CzZV3m3+z0F3mMKMISCNhm3fUNkd
jRcRXIZ/OSGoYH95mmLS4VL07718QHYNYmjmZq3puSZAX6GK0Y8wrgWyrhtV2QpM
e36UIf8RVOYMUBjrjkj3DU0/tw0K3u1/dsJEPyD9Oo2ceUPVdEZm7d0nFlrfvsZC
FBnQpYkdsKk/bXuWydNn9JCOpC/vEs/drlvIMffRXCUg8UwFSAksDLPdnrYP11GY
ZlXKMVHkINbZYJYN+lHeaUHPo83VVpf8VQ2V77ODvMFr+HY7BNt4cmOJP2t97Es/
FRS/lVL+h8KNvBMFrSALEg0PCjQKYYCtvJELAO3mw0QzlD6s6ufZ1hykdRRAtnP4
wc07zwW2cnxyywxL3NcIA/JUBqzMPqmzo2jBJIUyB/Re7eCZXg1J5k0q2OU5Wa6n
ECh8nEaoU/feoklbeJRk9c3f/ARUmWep0jM1UjqWRkIT1u5+3Hinh9Q48oj/aMCy
apP3A5pIDsrBywnWlfokvx9qlLyhpHc6exFup7VAKJdJdmHSRS02C+u6dPlGkd5i
pCpp2T996iUmxh6dz335IciaoEOloVXUK5QWHS9E7r1A1YsiuHsyy7vr+5fYCOUw
Ldyp/VNzxLJkUi8PP2BDciNOQee0sZ3B3apcoVmV5JFZy6fGeq+p1Wn9AXr/yhYy
Yc4FnjQb2u1+AZuOb6BF7X/6xF+WkFE1LadM4sswcUMm/BRFaaJhaclrJN8Ig+/0
8JviImB05pO9C7N8LeCtnl9HR2JyJ/OOnxGayC+WxXIjFDvth933Ha3aN3Y9X534
hfJYSSTBIMXwFwD9CCUSfliDiEnORO4JI5dT5OGAdseuMYNJo0EJ6MitGLbSFJJB
UbgwXCSt1lHUsQmuO0EPwXD8fI5uDwOgKJ55tO6Es1GVQSvu2n2fnS4ItDDcDYm3
C2M36zInnyLfQ4Ec5xwwif42AzQ6O16GgFobb4ZFqbaEAFeuWeglYGC3BhTZ/cla
G71/qf8hHxXzb7QshKnReAJiwVwlTRu/gyRPCzs2ABYO86FOj+GNlq9oTbCMDH51
sI5eCjvvMLSEJp2s/pF5zh9Eyfqf8Jd+wTOUOs5M3aGdAWs/tGTEMz0GXEq3ic7B
JawieTZtWMLLjY4NBaIPtBQmM21BHtWxjZsKIenihe5GPPHSekh0bj6LfAYKh6iz
dzXw+EfRVl/b3roFy0msINbaqid0pXpg8c7nYzmLjhVL/ca6l1gFfxDQGITZjTQS
XAZo73AjPckD/MTUTDcJpJNTKV8Gbz1mbilXoblWisCbOxvoVqBfOP/xzpqPZwri
J6vxJkxHiB5QPbVqMaer8aVD1Gtr+aR2RwVUJHAeYZsz43gUxt2J7ozTb7jCIMDd
u80IecSwD/2mG3OXQTkLnqyhgVm26f93jR/x1Y1ggj8uedKSw3hhBuUX1UhZJ1ws
rsX5wDxVd7E9t09mP/sU619zj6p9OUIVmJxMuR6z8onJzU0gC7sggvvNcGpVvO5N
tIrTceMijXYQ4rLAdvN6uHVjt5PYt8KFvZWKPtcLENWOHRlIBjcMWfVA5z/XISj1
E1YNXoQ9e291E0rl2C9fr6h09ZwIP54wIcfGypRUBka8jb3U/EIm+P2m5dGRMYBF
FSV8WggLvWABBvjQ46nF9WCbJf+6dQTHlBlnLNPAqb6OtZvV/d9bKd6DP46umqIA
eDEfsPzmez1X96buOoMH3pKJqwOl9IJeUgHzRfywU1OKi3l0kV3E/nhtBQwEeVAK
GfHtV2CVXpVi6v37CzHyW6iyMA33MPeJ8Lwr8Waaij1uyRZgS5A6w5XwVg/31FIN
/yNkEjQjpiX8jSSo/Hyucm5iHGRetlrlUwrwBgQMJPPVkLazDkFhMe5YaXmhe5fP
xrILhsRXqeEIJGM/Jtmjpi36kuOcnToEvifcEtGdYx6gtxlvoVn+zuviQ2TXHXGQ
T7kSkLuvGKOTAniql/7yH0JjbZi76sJ2komK9IiD3enSZ+se+Ys44/UgarSgQz8D
Kce2x2PME4mskOKQh/sTYY54mrzGUCWfJzE8xTBptDVAgx/OYiD4nQdImvdynnWg
OaqArC9z7yNmq7XJ6YorNpkm47zROzAbV+MpAAbigCB7U6RoU4ASr4ZotEy9lhh8
jXBDjbp+d52FBNtiL6bcGaNaroZ0SMOiOLdOVeGM9/8w4/pFCvx8IqNgapW1x5cX
0GWUM9eiN8HdcfHMAWQXrQ1ZOXjJq0RUmq/5kLDHPiMozGhKkET9TJGlcIL2KmPY
+AGviGkqvfrBxIjzr0wB9VRKPdZl7OGEDu23WIrCY2pWY/8rYzXeZKGf7X3bO1S0
QXAVlGkfBy91qLs3DkMWk1ur97aRDZDy67NKtlUtK3tNUmmQQEsyAUfg0in98fR7
EKZ2tOy57pPnvr1NRnvAdUaLKnD7xPK7mzcl1h0Ho/ucAFwaRWrjuZEfjBtuw8xg
ERf28us0vM5uyPqe1v/fMjoDccLljCQe68CK2JhglN9n6nO7yUNVu1MZK1/h2Ze3
EOypfW+QsltSTnmG5z782uXZEwBuVDuH0QCmBdZZXNaqTp6PM8mwVsrTbNG+7MA0
n9IE53yliYFiiplo053+mXIl5m21ous6TrR//YYHwwZwcZhG+kjJ/V1/GUV6ivvb
K4dyXOMWgiyqJbwvMIuJcdDDDmG87DyXI2MLICmchyKhTcPjkpuEmWZKrzbUx61j
utFsxS0R8oRNqlYmdtAA1BJDILb+3qxTWw5RVioBhc6HICvYWRpkWtkkzXB9I7PQ
QKbz2ym0hgNBbumrER1z3OyCPkS6xwb6fLvNpTo8WDjH4VEbFNRRQA5o/NYUBNxg
wJ+zR/YboDxNLp4T46E4JgEWWYfN4dvTvZuGMgT/RGynkdr5TeEJGKzmMmrvsRVb
K+9EDGjLVNGdTvjEJV8CE0JTmzVAj/koO4y3ZgYstNwM9gwYZiJHDbkgS3jW/F3L
wB1UhI7zTtJXTNykfNqpJo5Q0Uk+m5rqQ6tK3tI9WqU9SbCC/kjZAWtFIPoBY946
51vtgSC4fkZZ8VlBjVhJcOBPptLttPKbMhbn6oXn2c2Qs57SOQDTMjYBh7eIYCV4
rEwiDMIs5zhRHJvDX+FNK2qsK6ZGxUJa3FTaqYavgPLoQKmxNd9ylRr/Sway1Ct3
NKAY08b5O0WVo8BAX3BaTPJlOv0gWep1U2z17cSJj1/s1rL7o7e3WYx6IIXDcGgR
LiXOzLu/W/kaP75zwRFCHE+G0Q+AegJikbvmbMo+s2/ZKtfB53gHXD/uzHa0l9xZ
nQ78JA8ig8f821sXf554beZxXwtYaGERzfJFp0W3S5ok48NRd5eWIntsNNPN3C3L
/WpGI8pm2jMRXJVEwPed50bpWiB0z3RF1hUrZs9CFFKVCcb+Uh/rnAVUYvxbzNj3
YFk74yISL9zIW1AwJmot41cIlOEi4bXzyzU1v008EwuDN9L7iGETofc+GGEIF65i
QScjq4MGUtuPavUQlKTS/u0iiYamC1KSbTg/i/UlAielKVOUkk7SBkmTw8DLcphL
XAJUFaFIxMMdpgWE+FC1XBj/JyJUIDsEck9AmthYA4/eUhzmIqqAgVnrzssgI78u
oQ0wFM+cCiafwwuJhbQRyBFvtV6da+ShL2KDeDG+cwyRfrjP7h5kX0K5U8EndeSu
WfGLejpETceyzrF5AkTwhhT4k193e4hwoIAGKlN5clZ92n5uzkwpk5OiBCLBpZuq
5pcm1j3oFrWXi5LqlBiy+FQ8E2rzdZoLI0samqPhMNC7DQNvMkMVhfKOdw7JkIKQ
NKdsWm/9M+OQCdeImVRZMpsmzJX4YLUuginEOJy9JGMIhh4dOk36AfVKS6uBzXkP
L+kL/Crmv45VbQSBdg4IyXqv/yfLa35X3TxP8GN/BdtnpTiBI9pvOCt3P/IR8akh
ssKlQWlG79eLDDLe1IKHlnXRHcUT2ZOHbnetCYSF/9jcyV68Trefq6mkBVA2LH75
LqmNKV054aovzkxGy07unBnvGBuhiYi47diJnx80xBkHXM35UNSXZGGhpwcDTZY4
fBZWn8X2OwdknwyFVqG44CkcOUzFa7FKi1jXGo23XQEGrVJX7wD3ZnfzEVi01bnD
Yjhn6WLPjwtcOuOk7tkgRnP3Dnw2hEiDJ3ZYZRaXXSIM82wB0BlZFWpL+6DhX9mt
VpbU0gAfzXtT95WsYscPqgSMgIJcwWOvvJWBrZ8Fgpu0vXwcovBEScflYc3wZVh/
ICcWbIdxurl4Q5QaAeklJYgZaLJUzdYkPD5oto4MF2DqzLxOLNWWeTmf3vne0zP2
ZXYNKxmLhWyNmr61xocpAkEiSxWpEg77OaokIw+QLCTxWLuJuDrJDP35J53RUpLv
Wocfb9HmLU7ehlt2i53Hoe3k6WP1BgUt2DR73B8Z5lHn5Oecr2kq1IDGzKD8lqgD
fihJc6zQcfZuctFseY2MBZkQ5bx82486/h3CLVNCY7AbHXHHGa7kNGGr5dNM9D00
kiM+1vRbGHbxzMShFejOcZFIulYNU1X9AjBAD//jia4KNVZbqhS1prsd4iJfEHCa
4L7tHPHX21DBIYl6DfFlURTrBEhnuhqLwjLx9i5wRUK6cOK0B/ef+z4rMfeqYScY
zs49tlL7NesOvA1GaPHQ6Nwga0RB8OF53Yk9VvXC8z1U8gvR4cVCONgBnvM9GoU2
QU1nLg0LMM9IMNlXAy1SCAazurAlLM1soEYdYz12qT8wL+HPnmBOowAx0T7KCaXq
PWgwWis9rtbC0NYG/1EVIHwHk4lh6n1ssC1AgPXUCCjD+B10+KemOzAlI8HoRoZP
4I+VzInrkAOrflK/hWE56Nv7Nvo887lmFUN4fisA1zDNBpUbRG/vkue8TjPyyiI+
JwT8qwyc9kYF4vML6rVxXa9cnYFE78zGkBXn2sUXnxqlVZpN+QWKTqPR2ENo23mm
OFoBtEeBH3AQJxw6OJSRzFlnUj1WojBjKXplcdy42Qzwqxm9eQcRDbgBm221dmiD
ZvgOGIlLR72/rryZgKeTznNceHzsNRF2bwQPSN9Rmi35vYJVYzlVymILZ3+8oFTF
7dSDViEgJVzRQRBWa4ZAMzDdxsbrdiK2IKXOOXuMV1y8EReqllqROrrCETAFW72U
6XWmpmrnsn9pBolSjO4EOiJ1HE0DsOyAUvbmgfl+32PmYwgERHigocfGNSKA+o9+
4EwgZmmH9e9R62wLWMunNUSkMWyiGBhuQiaPD5Kbuxf2Ky84Dedqj8QSjaTlsJb4
YVvmmXlX0UKphtVVH7bEH2mOo/H2aHaOeQnD2zvve1AmJ1Re/ydmeoKmSd0IOeUH
qfHGkzXJFu1jrRBqX4yyGxpTLXDD07wfHYFaww43aU9hV9AXUm2DBjeeT6a0Sx7l
pR3sGR/IAyEo122c5fr4p2Qqdjkhjp6q7uI+lx/l3gmL8TaNaOvmTzN9eF6ZahJS
RMSx1qJRuHD9W7gUu8VNruSKBYPqKDE6A0cvJzAMSB+UdGu7BrWaTdJtWyiJoQPO
wqC/S0Mw+lXiOF2PNktytzmCsRunTExDHUdRKGvA9+vvL6fDI3viuZIXjSD1ym+U
glC4CCtU5r6+MGMMAkATdy2t426UomNw5gQKJbQTlKCur4dINB04+m/U1gaNfbhL
LFX5EESHC8EE82fVPGnyiu8EjXwkw67T/yfwxV74OrCe4y4zKvoUeGemGeP3CIfl
GuML6ttvyYQMO3SUSNrdvrbFXd4eNO5/6WnTpDrX8Wq19tlw2qblK3Jx21nklCty
jbn/BHBNLBQ0Sy063UJlyY5S8nhg7/c59OB5GQFKdohf1GTwsDJ5nQGxf4biJgZG
iBhZvfwUDTn35m5Fkij8r3mCKF3Np1gpDOYR6ip2IfOXML2BVL0u0S75PezRyRww
xL4YEdJvWZQjXhZGF1sFzUSVmpumh+KNTz9YAfs2SE0ijgXQm9eljymCBJB+sgUV
7NpDGaibD9PDutrHCt/4sqTLar5yvCBa4DieK9dBQs84E7V1zwD+NzfjWfR9aLSF
TIFcLoqic9ZoMxBTkDlRhf2mCGRMwUWttnuMnjZcf/fDJi18NQzA7fGCYESUdl86
3aM6Xiv9hjB2G4LDxV6bOfu8XybXM46lSXE8XLf3OOh1YMYD+1AePilWFUCqMVYV
Bq+iNMGWu1kogJ/RLIHwgqdS9ehGLX8Kw+TN+xrNsxGzC+kkrdJDDOK1lYUgREnq
rt3+vrg6XzunZVpwm56kZMGPppf6pA1Xo5+jkF0VXnQ8K72zteZmhxdVwnpnyTLy
Y1dbKYucbabp1ybiSFuQvbDOqvkwNId/OBHoGT6N9wX17EwESIMBNORHEm2l82bW
CvYbK98lWuPe6j5lykaWSVkuMhUWxNuW34oY8bC2DJ1qkw0pbVlxM6WPBjkL7Le8
JwIWqaTMZIYHATgfiEmO88eYAVtG5Kqf3PscWd+evjIoWpawgSBf46Y+nuQkB9Yj
R7a64zTg32vy8jgdZSKwO+Ggvkt+SMdk4OK3KDkXCxFEwGUqGb5a+Fr3G9Dpd8MX
+FjsOz41fOGstYk7tEiu7BQSoHlcHmrD85OYgMnE4Ooz4dfNgBiZZhl4+nkPO5iW
FtSlvaydIUUDZNjodkJvguBTx/B5pwiwa7shKXhgf4QPQ7xbCSY2hY3MAKDUUyhh
ES+wtSimm5MSKkto19Xi8dZyw7ImTBzZDx5O5Uh48em5KXrZBW/Fi55WuNl+q45F
paFDR5ch5hM/N6QICFcTvhwkFY8fx/ZUScMWeYfBiqKxc1Ni51cJr4v3uNH0wErR
K7tbxH4UAHW89CH6APsC3IsgeG5PxphHT/iqcvuMLOmqtaf24xFPWuTLxUNaswQm
41JcOSQ16JriVx2w+r8EeeOTQEjUYDfW8SGoGJPyKgL26P4IhEYVKvyuVpFIrBJ2
2qOSJY/m4O/CbDiL/ykH2zBQ4aEi3xhL84ZygBfh8TdTirc6oakiYfJ6gsu3VDrq
EO0FggEOgSpECzbwGnkOybNNWZUtEEY5JhDKaLXHdE9Bg3mieb1BcA2gFc2sIZp7
I9POtf+CYvWN1Ovr8ODSFbvtOEcd7m81K/Jbynz61AX5U+nR5WYIJa6dy60WXnYH
c9LOY94+QVDd0F9q1gpyZvsD3Rjm1tdWmeKYuC2zzqgEx3qs/4xhiHkaMo9eu7vP
bNTkXSpKq6F90j333fd6T4YoTAtySAPQo4mepaFSfouy2xOzNIRz7iCK8OQdGbof
Hy3BexrE7UKBR5mMdBFgZn3scX9A71FWZkxwEur5XWpuz6KQyUtyaFvu0l5dzZu3
EAgHv4glgMS8A3KqY3ZQb3xHndNnN+ZDWY9CP10VeBZYmTmsHifp2UjOHhn8Qh85
ALOB2mv/CNNXbYeJf+NXDNiCsxnxp+DncFIx70zq+52ElRzfVC1WGggPI3Qs3B2Q
zpd8s7l9p5HBeC5OWs22SG8KFFT/QP4mAYwM1ST+UQeAJ33Iec9+k0B5gqzVvaYD
9Omy2iB+1gk74yK3CcT/5gbmKXmR9ykh4FgzmX3blGlCFjKqvVUWEDDTJCHWCEME
RuHUXwgZr/PfAvbgL8zo7rMvaTmixESDe/262l6RsB6ojK1rws+2W4XCA74zUcvo
OHxCqgxOijPA7S2aaUBzP5EV3CLzqFIAkkMOhy4NzlsaZDEZMlmURmwYafGxscHM
u8Q5jD68towVxWIuak4CS2sQGMYGRNKcDBfNVArV8Ss0GiE9ah7QPHAHOZGFk4JM
gh+hlDq+YZAjy04mgHxRWbB8ksTlm6U9TfCoApKuxmNqXhCgh1bFkKcrO6Mg8BDi
VXYuyK0me6TDp3wqqPVaBTQg/j6l9VmGpKENDO1/p1Bceapb4J55P/ePxCX2Uc2Z
fa2amN8MxFTRd2Dftvq3CA/LLdO47h4Hy9vJI0NNvbsTR/FYA78CpkgqmiQBw+1v
V5MHc0akFSVfPVtXN8vTnqJyTxLRJqdyq2hfLS0XMh4YV7LxhN8KtZtef0fYSKIK
+LfzTsAW+Y+/VDYatKCcb3Vf7wJSDWH0L/JjGuGDtWOySmaYEEPsttwrzKEFMxSp
PX9teQf2a8RGNkJrF5rhk1WA+Ckrf0ts8iXg+ezaEMc+NT7aSS9iXSTPJwGYh8en
DCpDR0Zia+p40C7/p/w/4io79cxEUxjy5Kbahyyrqg1sjq2P6ZT/pinAUUyPy1xq
6gJZE7kaRwrHMedFrscvrct7NDEFO/Mv6R5moU3vrMyv+0d0I2d8TGZJGAS5MdSs
Bb905/sMVv/2LSJORHdmHdqjNd3oETukQ4WnIdHoecJcVoNR8Y7+5Cq0WxJX2/sO
ZNtUk6Jyzul5YPD9PR8y/TCBBH74KCL/8AS2ityLfNPFAVzRT9cyxbSwZebtguyV
8OWdrqGcM2bhSNXoK+A1rBIo6T3uN0MpcZlHrpWCbdzaTUiKnipVJVoirBOg+j+w
LFy2400YzMJA507lTwA+SwCC9qu3NsvJfxuhYN/eXqkF4W/IWMuHor4X/EzkrYBL
1CQ3mFfR/Wj4e0B0w+cDQWnJxb9wXA0ViB6Q7wis42zT9n07ZCQasfecYKJ1cA6O
1aL26CP3KtFLCPMWOo9bASzBTtJeLTY0tlI0nPXNp93R8ONF8RZJQH66EgyODmaK
iXDG2olycfuXv4aLi2xb3v1dCgghvIMQxEeRgeMfVroiARg31yi8IwDz2Ef5x+wL
SoOOvT0myupEqzSeD94Fos4WiYZ1cw/n56DAEd2fINyAwk6BtCZfFPgSOysnP93H
Swd0RkW5+6ImFdoLurTEUTHrV9Bf29m+Gtmas4gcHS528Sk1U+SeVU0FtWYL6nka
DCO0mtPjGpOSpkxzLbxE9DFzk4RGblPPIo7Ib9ksA8N41K9fJqjVujA9cZs2zHO8
UaofJHVW39zKMJ46322uMDxkyWNtto2eDlYUkRK1Xuny6zlTRdwKEBDZ199mmLhj
ABcmPcbaKhTfkPpwjnCDIjcu+SJP5Iy0SRrOzFvN41gi7uN59mcMA8ycytN3URlm
FglX7Qq1ya7ziZCpR1BiPqXibnInxL1P0/U707M18uMTQiQ87eS29Lp96iKi43l6
zEJafJ5CaL6o8dMGmXMkm8KAyEdsY8mFU3XaI9v/8T0OAZxHCwGiU/wAXzuJpgM2
Qqsfg81V1azUOrjSbwpfaArSD7vU2HdNElwzU9jVgZarWmWJZEJ34quJh+0+Qs7p
LPPmI7CIg3XZmlXbxrmyVoeU53DWg0CZT8eIuNtfQ6lWvROYD/+yUAWDzpI0zoWB
UY6J/OHGhdlirgMHTajt65K+1cwMfTLghZgVBeNt4w0RlwIjNBOC2OjWFWJUc44s
tPFFziOe9XQjub+x/lanyZAF+phdG/k0RF9wH/p8HrAF6df+R7tTo1g3AOVTmILE
cFI9yyn7unWZikodNgSGQ01SAgwFKI61RARv06ANFGyRcLxGWJYTvoAQeznYenc3
KzTWq1JWMFh3llpMGYO1e7kuEB+2Hk9MuJbAWP+zk+VQeBrMej2EIbDEjNynhQiu
kan5IHS68o/vjsZT2qdlT5n3La5eOD33z8ZfEYklczvjaasHDQOB8R3FIYKa1bYx
ejnYvAuiZCCNhiipjz0W/h5FBzU8a6yrLW2a0nB0YE7L3mtFvCifPK6Pw/bX6iOy
yzbbLFHItVOznVL5X7N7nCZBQwg3vzI6sMq6LKZDhfrtOltjr5B91FghzFmxyya2
rAHPvW1P4YmuKdZuAzuKbAidYzDKMForvwK/tJhi1jXgZvReDA77Uhwqeyay31If
HoeGrNDwB7JVcmOKU/vseb/inDSvYbWwEyZQxxmmmxSpyRvyBrB8rBu7T4FN3mXK
x897nPCzEzgk6aPt53JxHB3roiYSOcnr+ytuwIWpUDW8hyhCqcfgae5wYekW8JxQ
NLCw3DJKu6j9IHnyUJfSwpQjLt7YfS+kqzisE68lA7vMbYjxMdaKNULEoR5LLt67
rmbODpbpFhrcaQb77pLq0Df9hR2OZEH/CN2tcDglXFFgD0fcZ73jVDhViRxN/k+y
lt417Q7Ql1jfLOq9Xo/6RgxRhclKhiedwgla6sgf9llE2zrNuW6+oO68357SWpt9
2x9gBsC141sXUK7rOgLbc2u2pR6w6z9CDTvZ50kEiMzTm1TQ8s3QZPSqVWcCitAY
HRs0yCB/grqnPlw86T09p7E5868o1SVUVE3mSvnlKXQpvpNdOHDag8KbcMnILgJ2
OUnIPB/UMDxVWdPiwZNX7MpG3wPmprsz5wg+bEj/vwtDCI0/hT/GAXpr+R0EpYx1
F66jPAJO0Hd+E0w1WT9SKROaOBjmMfjy+e/Zpc/HCFoJIgaVJz/VE/27KMoNcal2
Wtxyjjyz3yYqJQYZO7tmAhA+RzLOUAMtGfo1goFCONayGF2eY3BWWx/Ggx5xCBvz
2tSZ/QD/DlLg8A//BfXS7zDsf+anew+WMxKaXNPavPhAHzx+fJX7ODe7X4Jb0gjW
N9CJRPVldzhcMWqr3h3Iw/9mw1J27FMbKDfFP8tCmgLxTUD0BqhWvIvcrsiE2ztw
usFj+So8o5a3hYqcLVERevdSb4K95M08JuocETOQjUnE1cvpgQcq+N4WtUJlRrF3
PxkVgv0bb3yOy7pZjXm0soAZZWd+4jRonbUd3dxulj7b8RkDcjXGE9Rdn4SALxgt
kM4cMmMFFxNgwGB9tZo8HBpj+g7vPWQMnKC6ldrLcQQ7viPz5UMkWRskVHPzD8F3
7+EiuNJqm7ul2iS6goLK+aan5Mq3EluLm+2zz8VXKD0t5yaqsPV5/JMiDiVHOxu+
b14OP/c3eMq5xzEDo59e2J3jSmARYeVhL/eRo9mC/qk1tvQCwBX+FTGiX1cOlSma
D7lOVqw/ZnOWMIYKhwPh7g0F/vjpaRUCPFRnOzizY/f/Eu0dw+e1oSoQpbkEnLZj
MxQk0Oh2g8o8c1g1rjD7LvTvF1BcnnuQd2WNjHWi2419Cei6LDnX80lp/Riy8LCA
L2bHyip1uVMO9vJxbRU/+QNjgtoBVjYDyFCuOR3a7xpOl/gMQYPrwmdGtMDVLHf6
ffPo+xcFPxwM9Je+v56LE1IfNh+TaAmdgpZ0+BmGZnGu3+nRYEXQRjZ093vv0d1t
zZ2XysZ/a/tb2MRFWRoQR7A5aIPeIRicZdGCNnJkZRcbOeW5gQ2lDrRgwnbPqaAS
AJAp63Yj8xxNt+zwNhZcmhCdVp0HjxuI4bwPxE2jb45hyVO8NY+zgnnB/dwbqS5H
1MhzH5ex/QG+BUnO8Cajx8AlekU1y0Irt5uU7al4sWa+dZueDy+nV1vko7A2Gvi3
NPcbhuIekA2rkuFRM/xRb1a4duwFQYD+Ws2ytzUARPLEmVsphKkhg3Z2jVqjGgE0
43V0zLP7ZEVO2E9+3a4xndyWBJDy9kgSHdvgkZpVs0w6DDdeJgT5agZn+wOkPwOz
f9IA7zKWrrG5CLQkeSlH071Y/HY+XfvJQ9gj2tSgWIaR+bvgsrp0t9MQgm7lfQhZ
lVapg9YAGGh1TRCCExCsT5X2a/j5bgmKZ9Xsra2k/oF50U6+YfmmU1R4Y2RL/cxk
H3dYcU8+GqUMHPfgbP9NdI+o67oIHPAr1HogNkv7QzQ9PFk+h+1m9O0HVwN91q9F
/FSOs4gL+Mfzg7M6Yx6yyBq84+3GQZlei9pLlHN5MMZ4ohBkj6sbtiu4Rmw0dqRI
eGIvsOV1vDhaHsWQn7TfV7GS3CKw+vYO81TOW6Q3qI5M8OshCggGb++1Qg5TCWkJ
x9kYabVMSqs4mBsOAuTaNOfnEj5LJS+pA6rFzzcMUlAMuJMjnjGesII7FGmA2RgK
FZTYRP/7ozodPguEuQiPu7/G3B5d+9ANL8uJceatwt/gN+ExQ5IyJaWUY3wIaHzs
QB3CI+2L+mp6PLkU8eNnqd1jR8PZl0ge2E+eiV+SXbHBItzkO2FhE9HnZdg7QrFB
4fPV18/CMsn6P53mlXIauAb7vFmbPljQf5OV+23ayRgVtJYDY8gCq/4V5FpmFMrE
yy8L33KTPPMcQJHV7S0FD6hAlFalHoz88NsfwK4onltmsZy4Wt/O7otnDIYfStY6
n3gHBv6dpeE65o/VJoh+S1QfLi0viRUBrISIwjDG92x6YHfZ9qq2vPsMNNPkaPCm
Y0W3n6mRaIzxHizGHPXThhTJs2skQJXwYCsEdk6wPAPhwH234pn9ll3K0NeLaYC8
739bebFIhCi9uL5p8WMQeSaoUzP+lmEj2R737C3Blx232w5Gzx62M/whp1EYpnlN
+H+bAHoVwqOjia/7FKyjzz1DoZcOnhOaQr7O2tEnCuDuZJzsZcN9cRucpjCQHwIe
w0o7C/HYx/sxpSic21kuucyOKnaaXkfUqIB6QGMlvC9VI9U6CMk9UvnAZbKuhJIl
TAGPYcsemOp7rQbvop2EWu3kLmVu7pEwQTdpeWGpkDmg07unSiJjWokia/2fFI7X
u1vqAIvGzOhOgnjHl7jKMv6xp/yz0SZp1YJtRFNhFyEWPaU/tHttMhFKQfnrcG1x
tu8eY0OHnARjYzVzOOZnSR9mp7TJOEcOA9c5sn9vEUwvtecovErONd7o8TdSe5a/
i2BKbbA9puEScrhJPncL9AcEKthCavNCRJzZgYvcVyA/MTZ5FHeT+cdVR17vkcmJ
TdOZtklhXxezePTWut9s7eAk18fnHDO0TnBwZoNZ/gFyfrK1F5V7jLVpwjcXG0zG
lQ+6O79L7USphBvb2Hyc8J+F/mYT4cmmOXAraF2A7U6OVNxxhXnIUgQ9qyptc11A
VXlRFRiuFAg6lfbXVCzxIgbwLhnbYwX75H8GSEOkyTSxbHmaU3mMqUpvS1Pg9v6d
ru50Pb6WIHppzt1CqOZIwL0O0lmu43LKlsGKGDf35l+CH+4i3rVMfQ/N5Hl8+TRu
/Kq1vImnLR6o3IBiHHEWlJ+j1tcOe70C/LQgc126ElzHgsnlBiYQ7tuW4FF6BoUI
BFZ1yH0P1S6E7/xQNewazFlRP2HTCXeWf1nJJnzQ780f6fakEPeUtngp1Ag5KS3A
qAcZuhTWTICS6ipQIDS3Gf12RZVoqIfQK8Z6mj42nlt/t92gE+8f5Cmi/Hw5cpHU
DFh9xiP8ht44xHGcykUWzyHt69cFMIbAqzDMF8Az9ocKpynR70NXMA3ZBD2teXbp
0xdMoX2dfzQ5VbgnCs3HjfuiK0zqGPJzLIevp5Pd7wQzd4LDz5s7H8dnq9bHWKaw
2nwOubdwmdgu/YvBMOMbx1eTPGSMgN4h4VrRAIG+vllX15yRdvTVFKrfzdQbYY8R
RvbO7Ipfvj/0O/DzuizAU4eesM9F0ZhTVndNzbicNsrIuqnjGH/EwdwQPBcmV93r
8ws3UjwYdlbLJJHffGowVnjiVERhuCf+KczL+6R/ugf5h08qVYfW6M8+CUo+yWAs
bYm2lBNuRxIaRbpT+mFDDCLYbU+arXxuRXfRwrTJvx43N4TER9UF6XQdfNE4cxe9
4IZVTxsS9XNswLVcAoVnhPVvh8lAs483KVvnXjry1AWDeDPHY/ZGhAKec9aQzfSY
ow14qvMH0d1ZENtb04GD4xsDO8YxngpTC7uA7RSeemKYPo5HXLsa0B5pyJoh9YX5
5XXbUvFpBTWUDWMAIy2UCiVENOaOGj2RObsuR6NWWkNK1DmD6nTpaDFa6jeCmhy2
Xe/PQFkgev31nhLKT3OvrWc5LiPArNjNjhz8KiP68AG7pMsh+z0X4Xsoyf4pwa77
HrNnnyb2sQYbcCxfzdMZo9i9C0PZ//DviGIxa702EmJFx6KaB2gnvwonepLRi6tQ
Hi7aCcpsRvG/IFb76/MCCoCXxAVsO4mpEM7AF7uPQHxTSeyUYpLn5xv9Qh67peIP
jpM+qFirvs3WKwlDsmNb520ZI/AQ7xjJqN9IGaSt5pfLiZyqE8gg56b4r29rVkZ0
ngVQv0AXDx/jkJQSaQX5Op/RTiZJWjV92ww7b9eK6pc5mqN4m1gA213VMXA9G2iB
SbhHVScx6M0ZRD0CMpu7hba3RZ0gwzXH06Blll+6iDjpEkK7brEheptVvcUXkLrQ
cWhhhWJhTzLOSsowE5CuUB8o7B4eVLca21NolZEVQOiM7fNVONNja1RRtzAzgdbA
cRolZELvC1szV+s+Ps74PBQVoHP313JQ2giL3xxotwmhUYQRnHGBVy1PMfD77+4Z
sC9U547EPZq1EqoLv+H+7IXApvCZr3YHi9Su6XlyW8DvKr7UxHeCe8pUBeGkgDdL
o/rZUmQNM0UEcs7kBVph4tUJVTjmCKlAIaFFkSwL01Zpr7bZ8U0gctLrVR2tfZkR
LpZfBHlqJ8GZdp3bNFu6XwIbkss+AoRNfNYBzXqDBkSp6pcVQnC4s/9lcUdgWWWR
w6vdg4XIw8G663fuyuTxnC8IAj46G/PzhBXP9OSP436x0f5oP6WyqIV5D05aHy3R
BfFoFIz1y7w3HbBB+rac6IlMuvr8pfP3+zjqT1L+ocVKszYRrjDTIYG3aVjw+yty
WK4ABh2hs/yYxDBCwyeGmaWc48aSwYcH2ZgKb5eGX4JL1M1Y5xjwN2V9GPQWoEPr
jl4jflt5jDyxhmiOJLp0bTPgcclvRG8qavbMl5/mToBF5PyTCyBtU/af8EfBkmyj
HFqoy5+8CsutyL6r5Vpu05qo5GLL00uGsWXCEupe13vzC20oj5H8c84et6c27VCi
8A+TipzuuSik+vJePtwROprv3rRBObxORhoqHM7ystFFi5q4KvjEikQIQ+5EG4r6
qB95NeptgXr/NMq9v4bSnWSZAPe5jk7WcMi5LLi7zI+kuf5EXeOCAQ6ppQkj15rE
0AobdsCb4Rl+SNHk2z7FaNRf16rIT0GFXNtCyMx8dapPrB4ObriJBEtwEhlWEh62
dTi7ZcWbuR+4WmVjX1IEfs2PbX5dVXmQb4QqhFf3TY/9VYJ3rz509KrYqqEqT58a
yrxNst6qlChAdta6FFnxeSH+tttrDvYDd1+xjh33cIqZLDPFQGi47a4sWM6AYAFc
DwG6D+XWU+OtBwsWvWcjJ0+If+k/XkEu05lKsb4pRk7jFiAy2KLILgr/RiggzIDb
8G/r0Ex9AOCjATUSm8F8nShf+K1uQKwb2quGkml2s5oxtwgkoXiYx2tsRH2Rp+G2
vs9XldCN0H9xMGHrR1oYlfBJntE6bg7lxfSHwX7kSmSTl5h/cCrQXLWbi3OTRoAD
XpovVnb7Uk2mqX5Jhsx87Bol04ItKOpABWK8UWfI3eqmoKmiWFWKvCRicp0Md9k1
eAEomlOrlW+X91jkMp03QvlsQAWs9Ws1ozpOM8Hq+4DPWesKrnXZtFTatuUy/1Iu
Y1OWtXKE+EplSf9SvLGg6p/a6E3LgHSsMzCdPQmjJIFYDYm9pk67YxajLX0jQ/0C
vuyq8cDXXD+teG9VKzzT4vIrhmD7FtlD2MIzozn8ILGOVHh3kSLAwx+MsmRDA4OV
TnBiqApg72CigQ7SVuI1IwIn5BL5M6UmXw+pfkQtZX1nb1y7fCFGiz26NFZv1bpB
ic9+d3WtFGgmKl4z/7Dh84g/srY+MyGOmBXr/c47JK2oPXW5f11uVK+CJRI/BbYm
jGPZqgXFJ9OdX+cheB40PwbwcvT79s0vzEdDaQHp2QR4Z8IE2mEn40NUpSE0VBoB
41A07LQmv1dll59PcfDphfd7Cb0nyZ9f4GIX0ICoSGGQ7KKqw/kZufcy2lHCnLpp
3L+lietLMxAucwFg7TR9nasH4N6ffPM72AzS/aoVzTjABqd/jexJA1JlhJGgnpN0
xzhtUAPuyJLniy53uixkrnU6CpZvJMu0DyWp5xKIgWsDUEbApBiEfXXc+o+YI51f
yIDx8ohIOpumoRKECazCc5sskQvBxZSs/gx70smKRlxL3QyTitldeo4SJjJktgp7
XjZzdKfBD4OjQaMIsPfvaLDF4DVZEAKhl1YLJUyppmYjjvTX9GE6qUyTRQmydIo1
p+xkJnfbCV0fJe1Odr1f5OS6i71orqywNXzHtEZ4gvSBD5xsQmasOgMNG78CJvvG
qCC30XZItqNA+GoCBaiXfd5yiW2mUrt8n35isu3Y4pG/fJ2rq8fIrMGG7maVehAT
MDd8w4T6KnLJAA4jrPkqm5rWqAb2ZksWf/ke/zcP1b5F2MYj8XFkiwArLzFQLiq8
hojW9zJJlj3SdyYi3+41letfaVID55gRKGOUumcw2FiOn2gTGnv+vvFPCUCPMXnx
Ir4dvSWV6RS11TjFMOP7xKqi9K1nzRe09A+R8lSzDYRng32je04PNjuX0gYyFH3g
RJrvJ/Xp48fM+Fsjo48xiJ9ZmiwXu2VytereU5kaWZP5bua2Ytl+ftpvLhitwq3A
jX8/1fzCaDglK3L5k8jEOdgJIOAZ64/Xm4Tb5ewMtJyy64kISm5J/7bYHdUqCnga
9WxSZuzsvyOvwiEZrPsHLjsFFh9cnVTsMKQ6F8ZHgk9RPuCknQjghE6ck5/ac1X+
LT3yj/tC+TX87PTS8ni4F/67tt/Oi8q+6vNVApJ0337LFhTsOshmFN8omok4QejW
cFDJiuAwHghEqtn6eoaSrIQ/kHKV8++esmQ63XeltqiKsFdcQkYffIeihV9jdA6A
5qb1XCH8VPW8urbkU9BXrB9uc/e3lPV2XJEP77oRyyLEV7gqNC9mWV69V6XSU0d4
WW7Qh8w0uN14BZolaHH8/uciiaiQh/XcsizstDA/2D7nrhI3kesJ1LbJG81f/+uG
7Nys5wA9xaPLHJGx/sfWSK0Nn1v+lhi7kZ0HzlWpyUUFsypw48jjkZWesfmwRoz/
lV9its+Vm1qSbfuPGQ6B2sdErmhJ5JR9Z3Do9gZFh8b1v3uPQQmYeaPWqzRxFlVh
l3NRFbHrnHBmb1WwIjzbFB5m2OQ1v8A7iQj0I+XNXQdCuthDZQfXtD7U/l/xAwcW
29lGOFOKmTL6SuJHqm+XcH62n4yB65Kp09foNRPexv8pK3OHKK6Kc4mD+HPP4wKo
3Bb3wb51Gw3Kp7lgZJbCOQiwp4B9kmG5DlD65gd7uTIHok55ZcO20ozP1dJkSQPW
WAUdXjio5sZHEIFueL0xG9cGQe963hMqZeEB+4CkzkFZi/vVd06zTIi1hcmdboFO
VztIx2xuRUSUojfmjRcuvnKMoW5juEFX4VcT8jbTw6J/pS/+bdRycYBD3Su2Y3hD
pUCHbtor4b8C8de1Aw1rU1sWnld61i5dOYMdJp88ntm3pkwuyfIRfHzGU+eI6lwe
LFWtllnTh3TR6TLNoZ/CCfY2aCgabzeVjtyOxlN/TA8znGTLz4Dd+k0qNrSQLjVy
n0C1oy0OZMpq+pCTj/XpMQnqHoasZO76theRJtFaYfCWW141+UKfReeSRXix9l+N
Dkak7HKyd5FJuO58iX7ThFeHRdAC1Q0cXuVezbFEBlw8JvkaoF2TuB450QZFFmHv
6LyPamGqMBLnBLz9F7H/a5musIhmNM8TUYXv9s3MQ0SDO3p4p+l29UGj4TL7P/1F
ODS+rMDDgWxJUA/q8DpRGtWkq9T5B2qutI3uU0y1TypDemME9L3jlrjOrK3UgpJr
bSZG+8ZNEsDPRnOthNO0/BOgUidtkQSHS2vFFM9IX5/rCXObjQsAucgvwZbGV/2I
rcBxizhnZ0V+1O/q6NrkbjlqdNLPODDLL/tolkZgOWnoyN5mjmcla6/Hyd6LHk1F
exOi1H+0/RwNopDdlcPxUOvKJVbWxNRLqYauiCCbUQwH7bOzZRcXKY86wTorzSmO
PnX8iGcW+STLyEVW5nBECAL16irL1quO3mGIt9Pc5t6HeytXel3gFGjloEReewVd
yE5QafUtmFzYWKVl/Ck/N/hKyW5sYKdCzxXlrFv2Ze1w27RWn0emzi86rd7kx3ne
irBM5WLzavPsqyTnzcnvWPeRjaf5d4/VMrZZl8nrP6pEraNgJtTMWItlX8Kfp05+
31RbPcl5EHhlDz6eELSVW6BEmAjqV5kz/xhqe/7fTH5Dcw+xhc/G/pdyAY841nwY
BU+/OU9WWVB3HE040LFM/Sr76h+6ISNaQkekbyNqunn+qUHGS8vXqquekrrX7XOb
OmbotZSzecVWsFRkhgXZsXjJJ1Gx/3ii/UD/O2Ch7KR2QFophMAvZ3rbKU8YYpDs
okwzRalM+TLG3zDDjCdBPO6XSivbEgSUCDrCzzz5FzUCLPuxjSXJi79bBnwyMuLh
80ubbb7o/edUFWzwWnF4avog5Y0apmGfbmXOQ53VRh1k9Upzwqv1XyIny2LJeiqi
S25qCjAbjg0xTfUYrROcTFGXuijfd0xz/88bjE9cBxE9G5FfL+u+YXNBlsD0QJIS
+esrH15hdUIXi5pHPLxnBgDjNFnk44roWuVUlSqK9h1T2o24PQh1my940R+IVZQ+
Z+ZKT+CLyNlLIgJht8wqRSFCUBsraYzAjoZkcB51Z3WPU4bHaLyqiXpUhs5WRgUm
Z2yThLxKD63yR9jYko+bZx8yV8ckwhicF3pu2zC0/sBAKhjUham3h5+fVugGhnLP
8zQAcHqOHM5nMWVnofMJ6LEFB7+8PVjaz9hVkHPxdDw5fYp59feozDZ1vTJXG6um
tEthkbtKdbQfdmm2JKwEgGvk/DQh1pehdL23j13/vLj3LH0IPsgqtOTZW5MG4mV2
FyHKXARDbBeUaF5jqe0vEKZ3DoG1qN05S7W1lTzIBIhOLgY0uW4EsIDxcHgIqEYz
Y0zWEexsu/Vsm6Bxu5+8QNr9SvQwFgUWQ7cN+CrC9AEie+Nj5tD5k/3cAmR4nL6A
SM2RaOhY959aCx1VUda13wSTbPjMBC40em4Lpc+IpF/oG2S0GOuXmsGPIyIQUCWt
ZabvWgqA1dJFIne3lFmGHcpm17a9WJozAHSJCdwO6hiDJ48OkvgXLiY55UCFz/3T
m/qlGZTX7qwwz3HYMs6hah2w6Sp3vRqelediEp3xDC7Mf/ClP+SnoqJBS0X+WtUH
0R8qk8UGGAyPEAPHsx9qmwFOJDabi+c6uNXKJuKSPnGMGYhLdWk3AHDhNUmrpGh6
CtVxOARnTJyexA9DjL6Qp7XlmI2+yruXKsc/Ip46bGpeBqi540gNxK8musNVbAoG
TkptLwZUA6vGEtu9jXtetmhRCw9VDzfsEHtla8LnIX/CpaPe1uCoEdFS7yKzweoV
8lW3xT5u4Km9OQ0kKaNTvhavojapi832Sn1+3uqjnIma7JodDmr+2g2KUYoeQuym
abMvFRi6bYmt4Oxz4hMGq2ir7Ocn0WofMp6uh0ahjVA7GNDiYKUUiPsAiUY75bCn
I/1UgoPKM7xnQ2y6HJR6JVHmTjbQkAPWvqbEWRgZ4J/IorHCFvMUJoiBLT4t9S72
W/Oti71l43oY1vu0yPcCH5njXzxWpLCq7RuIj22SDk738Z1sr0aJcsuGP23hHdk0
FtewDieI3uSxDsEm84p5f3FMu6S2EfWXhSkp0bNrMksew2zDbP3SnBEe1f182xZy
OuPhRhbH3kJcwbmyyjQb/nH+pL90sofi4XcAP73oIqSG2WthdvhBa6oLWBV+aVsm
fW0uSnImewCtILU+6/0mTAnWXrotPzFlXjdZCINsnqfAYJXinghD8kxod4kEaQ37
VmIoV4DyrCiW4Ov/aoc2yz7sv+2C9MxThlntMPO2asoFK943RW+35kL188MU/3S7
R5DH88rhvo+dBsTjtnrU5Vt+KnzyFvugjDWD2aA+OjR4WAeuKLiBL4JrC3HHoeu4
ZmXfhd+mWAh4TvQHDRw/w7wzcndzeTLTPXcfsS2yNtlJodPy4SWwSIRnxboY+pGS
8vZs1YHRBk+XWOoH65Fau3qy7yKlctrWSRkSDue+see7ZK8UR1ouWumB3DuNC+nS
fxn5YpDJ9QDk37fM4sM/ZO8wE4dAYPJi88GtI9JGR7eetpjo/l2DEJxxUgRSNGZ3
iWkuaQlMqHIDh0iN4o9HE8Xs8coCAD6GCgy7KGffnUi6eELukrWLrPr2jRtsbk8v
Vu2HPDwMuDrhTJVRhYmmrXIY6/IkWJ9qs8T202yno/8O/ow9yGxn7nqdg69UXYY9
ED18HaTwJVwKrAhO4tH7x3OBMdczS4aCm3vLWG1Al78ya/UsPWEtSYs0lyvM+5Bi
IAxT6ITlFMqwRUyO5YYX4O9n0yW2Qye4Y9mvcFzYIdCYh1hqU339ZOXkAuExlz2C
la+SMjqZdwTu7gcUPSJq/kLJfHTDoWNRITrYftCDdqWz3xyrEjgzKqtrTkvn5Qgq
CgjSp1j1Xd7XYWFPGmRIu4SwmsEbh8uflSiMpSjbY0Z0+WsdA2t1I3KYbjKVlbt5
eAp9HS/vYl+weLOeVq5HwfBB4KLYETsm2i64TpI8y5M9zf9ALlPZKfIpZLP5T8QJ
xpdxjONb7p+6G2A3KZFO46v3LWHK1hqm/wsrkFqq/nSaGa7xQbufzIlqrFluwBpn
6wptOMsJ9FUBhaEZcpHBUUG3uEJmB2nbnD6c0lRX9QIYeigNTZGpeO3joFEV/ljK
vm8hBJPkyS9lPvlT5whaDAi/q62uddj277II9HIGpa7Okvj9uot4kDKMjNNdvHod
2D9b8qGab7F3AvMw5DUmXYC+RKCD2MIK2B+I5NtGC0OdpwmBkt0d8obkN0idO1LN
hT9snvDpAhsoqsSVF2qdASx7LwprH0Wu/ygLKQkmWk3NK9g4UXAcowNMgvn5Nbgd
tqGJ+zIMtmEOo83iaIwk8f72t0PE1LvzWn2W4rlnRFFNoSCcBgv2G/yXdoEhyc8M
EgDj+9A5QmFeccHhGJRA+2NuKdROwxAez7LHmT1NU+WjKFUUqnpvh9al708mjkJW
+dW2r1yWV1bHjPS3VaVgG+9lT3sftt2935pnt23hj2RV+zOb1ACcriwqM9XdsJ5r
LVrnnKOBheol5Gk/yTfoeTi8LIEnQ59xilvvYwt1jWspbP8BHn88Uyi9pWf5A2Xq
BsPr74GBBbJjScH0urZ9hQ/PolmhQ0ZAPeN797l4ktcmF1YhEZ+7uMXi+ESdUD2j
wYOVVBjMuD98S897BD4cDCj1q7jcVKQNZ/iMu/p3GqHdTLhD2FuDpYz4RxMLJFks
G1+lIRmPFVyYnWi9tS+USGTBHdyyrt2j+KPQDpJQZ+v213j1b4NmORPSKd9S6zXS
PpIIqO7hmZT8Nz33x1MGktnN//3fBy+TQXSgmm1cwHan7ogxb08bWi7VGH3Vy40s
Iq23RGXj7CVYYYLTkyeeD8BgXs6nm6KRhHQBh1t+BXbT8qCWxVff2FelRx0DT2zu
GFqQLUyv0E7ackeHJLwUW196CwC4PZgMpDr1UxQBbw4ovuFysjKLzvFu3XoEUm7h
duBYYSPpeAIRTt1pLQkjSC5LD7xYh7wLtq+3SItU5hYOIU4EkpdqZitaeDR+B/Ll
I6mWUPlJJYa3ojtUDm2BYSNdzhCXm0fpR1GTCI9vjsNSGDrWPYFD4K0R4C7nIsYA
spesNHtEIWzmo7LqcPB8YaphsJXg7rLymWRQwo4TtqwMdDpEaB179U4M3MGvifFu
1yA/bQM11jgGUWV8EZf8C0FTmCz24puOt0XbLCTBlbrByaf1CX+8IxnjPTI7RrTO
TTyvYk1LHsx+1vtRooffVWA9RTL9IiCxtF4jwxxAA1jvuApBRyjSjEbZu20OiXoz
EJTky8qnxOijBGLNX7P1fmKN9cWEWgmQpuKkOgf3PP/oEChEmjNvox54FrzKEzBS
k2w3nEHpj8lzPLet9TYJWxDhAVs4tyqIPWhHq8n245V5AMNgKzgpVKFz0tWp86CQ
PaByaDip2P9p4XaQnwPqG+hLJzFJIhXb0oPeTn7EG+r4bIsa108Dw4tCqzFpAOaO
Ccb5sgRj6ocaGzw/TBUMRhw4k5G4Gl4aAg3UR8CG4H/wxT/LIKB/fT64fesRcwVR
rLEaQ9me7LSsH9gmS79vFRo3DDEujPW5aS5VJ99mak+e3uH1SdnQjaTq1J+E1DiL
ZF8Y3TAxlWF8aUdJUZr51XHDmfEHRWEHnYFU2qYYlK36qyWepf/HgjWH8JQEWWxs
aTm/o9rgxSwqxlOA7qWEMuGJr8F413afr1+Jvr4R5lcFRV6u5nVzzPHqwz5uNh66
/pdO5rgX7tGmjLWQWGDOx8xDCsM+lbi92xdsGaFRapUr7KTfWcwN9emdrO14hJAB
dXl1+uteFFS4Xx24Deb9x8upAvca/et2n8yPsnkSGgEz/ZphUErxEi/AW21gwTm1
a/3UgJs108gh2RqHQvQw1Hi8u3AfPCMkx728g14hvwfHAfA4ywWogyl0P/W06idB
jyNwSdNPBlxERzacHVI3ANEJKCsx+yFVi9GzzG8jecGgIlXCUfrHgq3Hk+Pm9e7u
UKQbCyTX8a4rtYhc7eHxChS0eXPO3921nJ6moeOcV4z9qZusus9Imuzf7uJsnU0o
Dwwi/9thnd3F8Etw+tfskgwVR7l7UzDIBlX8vV0MD1ckaRH/T54AkgnxWkKiNPtp
uLymhp4h2LwjxX5iYphUOZBCMq0SdDfAPsYqPHq91yp6dBx23sVO/iMWXr4qjEww
ezjZsm6+rRU0CM51xn+BOb8405JigzJ4b5PWFY4JBbmZWXIgSIs7N41gyjXO+FPo
a9PzbuHg5e7j/3BiJ2WmDg6shqUYlbqRKEg1Lo8WBc2fQKszzP9kuUwkyOKR2rBe
HHf5D1FrZirfgVVe/HV7N3fp273BWsCL9zX59+wR/UBN9dFW8vQTHk/uTEesYFMt
FYh9KVRXcmOwpGmk1u4TP26qd0ActNCB0IM3PNH6+dHKUV8xPFGoGKFFZndYmsJl
O2vBmduqfHkbOncNRmk6k3v7kdKHX5DDoe5n4srHvnZtyLRGQyE6+c+xVSIKH01J
fKlT2JgazNFpOX6orXh48doak7AAaLEs/YsiqIPbavKsqzI66FfRyXgbiz/yUnLY
TII/66aElOjlQAmp9UYICERb1O2GUCqTiT2V+RgpPX3F4IMXL5VB8BJ/x5mPHYZ0
4eEKTBU8tA9C40jXYkCU56pCD2WS4EH4c3oP9TkBjvB3ChhvkcNz6zsOXgGtwO9s
bQMWUFGzRusFcT4dxRUn0fs6/5pUm++JwqAh0IFY8/8RnjPNG6UtB8fiSDCxFRld
Q7aQFz6XFYBDtQLRQ1ac1QevNKJVEDB2oxL1p6CE/Q87asGMln9ykHNTiI9NCL5R
WXtnlXOaW3l8/nhALOn/o9ozoP0POGj48jozP1PcWZ5/pwBi6IBxXjf9fm+55h8e
fYCacUPr0FcCtFZYuTb4ImC5AfA34zRe2+3REFuXxuS0uvm8IWODu1JN4Qq69Q/V
HPHr86sLb2XWsnT33682K7D0g66DHlrlbc28X9/Xr3eoMqgpec4ldWfBpi0ibKW0
MeHEQgtw+SlyLp6jTdX2arLzzNHKSeKOFEqLlt49P8Eqar1GEDmowmwJQ2k6bFLC
qk0wujpvOJcLLraoN9/jUNFr75re/EuCiIHT2Gt3ANJ4MdyrLSOTptxs2MU1a3z+
dXt5etR3Iu++E/CwmG+4n76G7xGBRYeWdsSQ7cEqnsRE8SLGWvnRnJ5a4EJ6o3PI
qJpX1IEl7Rz5OEkEJsIuyF5OJonCi6BTxsu7MZ4nBwh3b2v3EcL+hzKVbIT2nrFy
rAdYvKuEGlJX+KjuujHR/7CeMclDZgkiysjwlxlOdMUP2Yl3lzwqu5Lhd4ZvoGBK
E+2mvL1nJ1hknUZk1rh4CBHaxzl/C0W5tHD3B1MexKZa1J2RA1wEj4S2KnLxgl0E
ZoJkLE3U76dAo8ieyqdpJr1g7lEx4dcPGxnU1pk1E7eIYpvErChGkqS5ueIfo3RX
Zt/Qksr+SxcaIFxVuHtvQezSB11yL3diOICAMdfBIIJOhCMq0IlOPZ9aRVN3pz0S
Qx9xGPOwr2WJiS07WieMSEh9z/M/KsHY1/G7nrcpXWufAdCiljTZvJGfWCSFXVnR
wkzZVoCHuCtGRb5aIg7xCA4h4gFrm4oohehWUY82aF3PiU4fXvuiXiynoL8NacOC
NKEMAZiU+syPWzOWkGcsmpScBxYHUUZHvqvqls1yab6b0MVgjfWWd7EJXImD8D3l
wBbwHNCqSmTY/UGU1BZlIiqKZz7rYRjb20rOnqfMiS/H6tbxE5WcyWBpRgpe9WAX
GsjLwadc68ESDan1uGPdvmWwjofm09KlpaBVg40gC7oNBqVGhVnYCTv2ANKNoHfy
KZFb9aA/QUjzO3EsG2RoADNAWZkQYSlyHNOxrJYqHAApyjW3NQ0nddXi2URosoNA
QTwwdVI3x5FmlbRXFP8n/APwce1r7o9iDSBNscs3eYA0fzqHsvNfr0ZHR2r+W/6a
IqA6g4WCJ+BnhiECoWxh2y3xMIvW4m94ke/C0ZI+zm9LlX/yaZhhMCXXPmwT0Ohx
BHaZ2QUgVnD+kkKK8s9o1ScefokShL44d/3SsRHG5f6GSwDSXCXNtXZ6wq9aZIPU
B405ekULN2+6TNeCtw0MZOSQ/chRZoPBA8aj0Nil9lhH4YqGfGK3qmdBHkORU4u1
nbd6vWbaAhfZy0yLQHx3h1mhxjmAMDZKVPbVU+gVP/rxItJm3bAFBMqzZcy84Lgt
E3sXRZNcmv1xWfhu6G03EcxjaZzXRueBvK1HqSO7dbxHvUiDTIf/z67foAyI8sa7
1L70XSH4YCF2iAkqH4bqSUg1sHw3pYPB5wMahqUH1QfsOrrsH7YFQ8bvULhH3e0G
HEDlCf87OBUDpUFSIASOoBMi3cbp5Uvvb+Wca+MJyPeR81monJ2y/rvoMSEX7W+o
vllkhLs9YpvB5Eg9cLFd8jsQnnI1GA7EI/EVPQeoXpwEbirw40fcmfIsywLd3rnr
M/emQ+p7ruslWj/g4IBK0dZt1lV5f8CKDhIzsUCMK3lWUW7lDhHmEIt/Jc48suwB
b4psRHxdeViTItPa1w9NSRYwByw4Q+VeBnzGsWLWSYZUJ5C7ZETToZLwxdpR67YT
HcLfgkQg1MLiyY3KUT8x0WJ0FK9Cbq5Ubee6uScsQXrvvLjsfdZ+FYbW4+xX56Ma
OlkDbo3MolPW1XE/CwzNeJ7zyNCT7WgDX3CvdcMVNsYG//AyQenjTZcER9GF/Lut
IiDRGCxX7lg+10CI2QHnjOxrWYin3WnUNUqDPjZRgwcMtU9CrAgt6W+Wk2Qf6Mk0
/NcdzpcOcyBG+05espK1Gl9WTx2mkGb/i1D6oHtpJW+4iXHdl7ySHqZtVrBwb9tW
0z9B+9aq4o6orSdIkeIVIfjCmtMr0nOUlmK8CZYdNV/r/fhm5GZuNz70wkVn7b8z
AtAnoCxTpQn8t40VRm10+N58WSBttm+gxewlak5N1TzACwEJrdDg/oxV1NkXoJn+
U6Pp4jmw4Aqw15dhFPVt/gs2rPs9vKY/22/qmxIdb/ZLoOm/bbyQOOzmbpCRqfEf
UizKJp/kT66Ba+smnuQMemyjsouXmwz5dz5ZQfx7q4RtPm0KXQFhuHV90gRrbcrl
W7gqWYz7EaF2wPOc2gHCUEuTrbyn7jshWJCVS3VI8lmyCr7TDmXZMRpF5AAIiiHb
5jJ4xGHIQXEpwNAngNdSqETCRrg1P2afMqLS3aRI91taLtDBftVdxkAsuvHau6XL
0Uia3ZQEZrR7G/NDsL/JAhKNxQY4kPZWdyIKDisRGIG+HVTmPT6xFCG01lHMAifZ
7pmdAZC1nUXwUQgkYRHaZkQUTpunSudotWMJtXWoxUWTV55a6ZgNVAmHIeTErytm
uMI2sJXbtNxxoYleKVPJFvyYXxsDSA+6isGfNfDB+A4Y6L6d+jKgjRil/XZT2isu
rkuNppkqGB02Ib3pPerFca+7osd9yxORiDbtzq4jFApwXoGuu10mpQoB38jPKlXI
fTjfOiR9YnvFowkLFqoQY91S8h6l3MCHAufUy30j+wzvXEzbrAkFPr38XngwnE7/
x/5/dTmYS2WrFkBeJneriSnj1lf5q7A2RAyTQzp1Ar7bCpH5F/FN6aBccQyqNyVX
qtRCGBGD1c42kDEJfilA9fSdZnckW1rBrdWFlDJvS2b0GC4uE6gmI2gnf2u5gDRL
lqyUHW2cfeCAEqjvWzivda5SsEWq1qmlrbMcX2uAOvd2DZC9dvVFOKnX4Xc1Xlkq
+vU+07/Ot6mKl2pCRsfLlt783IJZYdwKrlf6CChTLY3U0ntfWKdBrsVe9qNxPeEm
aQvgbBCkEhFAvXK7AwidoDFoeAfxiuJq3wRla5zrfkd+8efwxAeA5rQfMqtTAdVm
oHIa0o5TQOQg8NxQilvmqWKyupmAH4qPifKcKJO2QRY1LHJ9vThtlyNiafKiBKAH
4FZbaQq2kHNqU0FBOD0937IPq0iXklTJVrjDnNqRCy6w9TjpGD92vBIpkebV2GNB
gJmLImoXMbd/pUQB6PAvZiV+DXj9QeicXoXo/Q6Nsuhfq6VPcq50m5nn/epE11CI
Xy/JfYbO0qUDZ7bj4UUV+xFMQY9PEKuiVylu/xGn004uSbPhxmLJeWxTS/Owx0/M
n3ivybnDEydW/YTid7ejIfcZNJ9DbEB0drR2LV87pCJ3i14dbS8mAfJDEnHKqDMi
30suGTCNt9t0N4ntWHrtqxS8agsk7IYSgzd8OugyNrRFkreIo4ZmM0B8uqqcyr31
PNGijcLZvJU0iUxN8QabuT193JyoePhtO+QIJ14HndoYpws0lccg9lja1jSi3fDd
/kY+U+CEyoH7wIFnenfO1Y7CK984jBD8ntDG4g19WpQIRqQ7l2Rpl4Z+k0VlCBeC
UgzrMoYT23V3i3aIhiot8Dvivg6c7TlTCixUoi9DMhm/T4YkvIdlylRAiMcslLsP
QmtINyseVHRfp9dYkgzIMWxhc4vSkHJAFQRvWNRpwBvxnkCBtu7cdAbsMj0GYMoS
B5Pwbra5d9uouVZSWvqCvrMldVXGIYOO1epeDbS0xRDva6lwkb1rB4ZCeNxLFdmC
kmz0s7BoHt2hvrcwO3Z+Y/PbPcEJlKlPlQX94b6G32S6QX9l1zbPM/6Ak6N+lpGn
+kOH/bsbNnGB46tE5v0t7d4TU1sItXWmTNU7OPtllqXvjOM+p4q9LHerOqE+gLvm
xq3gyQc0gv4mw1oCEyI027SglDrQtT3y9f4lEmWkzSBFmCfbEwD2X1dD8SuEFc0z
/i5+LzdvXV7gJOyMGo18ZBGRrmY86cay20tnlh/5fGxBUwsKPB4AHrmK1Ve6/HVF
XQyoTMgi7uuQh5S13234xwlQe8s/APfrA7VPiVZMKX0osYMlvwP83sfb45vGbUjU
Ntde4sJtBrUuANUpr5ntGqp2Zeguv+r781J102eHCTZwndfeMFWe9sbqn0oNME2z
SDFCXx88K5m19FuTMgPZODxyeKVGha+NPJJAgHiOAGX2+fo+na72765EPXRfY4aK
ikqTIL09+wDuBbRiZbYAcGY7vZXWaFJPmYz9/Amaf0CW8G29CrEsp1/e0fjWEXxx
6dj/NP/lhUxCPxMQyeoffJHAxXjTz4kMRZJaomMlrsTdIm5fc4hX/mwSvC0IpsdG
+LLoLdslwgsTU6rP+Bsf4wY50xtP68QTiUZc1ZC7CqaCkAHErh7dFiy5yrtIUiSq
XEaEiOqXj/AitpwLB5AXvjOsRzOiLVH6aRcikoDvokE87Mnz5XTkcugyqGc1AF7t
5LPxqTMCMONVqhD+xDo/Q1pZmBqlYLLDazWvJvNpkfcJZgpAWF4ml3kh+nmBMORg
Apeua+B8J6X6HU2Ul9zewQjSUxbb6ZM4LkoRpbsrJolljYaWIgOIqZg/TRYePLk6
HEcDnX8GLKkNrn3nlS4U9GQUAofWdGuUuLmBYf9pkEXVCgKydFQQhyB4FfPXfQ70
DVwFrD7l9PazoaPgLO7zRQQKcq7urXeDntWY8YL9o4kcKxZPJOtI5KjEm3RneUoB
GG5fdwobO5e6lN9wIUKxcZB7ANHFACP6vVD58WMO+EVokwHNUTknTljx21gU7Z1N
rFWooiSdBlt9fyoymt0WaEq6t8+yeGs5jHw+JxtGXH3U56gk+Ml23bTJwwd0iWdZ
mB6hhfvw5Iee/Uj34fSfelRWRqYzCb0YZLD8W7Ui8texV41e4RdDzVfwTMyFNzJU
gnjdpdEqy+C+WsMpuSHOiwnI1fKulnZhbDm8VvRjW5fhV3+3Zg2heTH6S2scwqCa
9MBRY8+q63XfC5PryFkTKKI76oGfd0M6IB/6ohcVSthO4upnHGVbj6Jca4EoFLL3
WLHmIi3//IvdD1xhNk3yoNOfRyc2IdDD9sfDQBoQSqj0hFPnCotpWmeuAwaH35Wn
xfBOaUzlXVqUFpcr0KKJkWtaVu0RnMzdU1LfknAFBMqmZhVWZCY3+ggi8/etGqCH
crfoh96humqe8nt1jHdmq9BY9cQkIz7Fz7XsBpt4i6zD+HgyjVSKROWB65kaiqgF
PaD15nkO/WYj+RaxrWibke9+fmhBouLPL0xtT7jNXmyfcAiaolrQghAznNv6W3LR
XD4E8/rkPn3nYBKSzARhuwxR0rK6XJSK7IBUKFswg5nln3xYSzCqJh+8pt84vK3y
avXU8diGshmO3Dpo02J0rMYGoL4gGaInbbntbdlKKJrZ3875JeMuPEfITkspl60I
lxDcJpeICSAtPlGDJET48aLGqfEEBCnxRTiJqqDRudFf14iURfEzYA+BTyzLfbaq
UtYbY6CykiggxbsNRpqcLQR8IlgbhXTpdyXYdb10hbDp3aRdVWdglRgNBJBgV9b5
JYqJYuPLUwLpTuim1WbvZD9+kbHd1rhMzh76DSlRbmuDN2pzj5xCljmBzuDz1WTN
5KDEiLXcaFeL42LXHajKDplYK0D7zjjakhRNdSkg96aoJZwnLkBdV0dYH2GKx21G
9OjloESACouThIT5DpIKxfmZODMwbgrXTjngfQDx719SYh+X0PGOBVinJ/BSGT2r
q29YwHAGcWrB0xHLyv/4325GNp/LQ3SGBhNXFwNC7MJSh5n6w4lJnGR6f/056PGj
Iv64rw/wOMBoGNeNsSn8gZkDu00TDazqnnSQeQJlgTtPKetbkHTRZaJybe+vOFsq
8gBzLlbiL5rPbTsqcvb4Qb6nUlvT+MzZvJK5Y+wb2gnFDFmQITJITFFzB5F9PvQE
jpN9U1UzoeJzHBqJSGuEmXwO9BO386vcQDRRH9jtpbouns8cCgtXhFxf+SqwlxoS
VOXvpWIDTXOouSpsPXsDVgfsF35mj//Ur+Kw+514hRMykrcKQ+apYr9CSKqZozm9
GJEene6xO2zOz9goCv3cJEBkmbuGNAC6tPL/qvpCblM8uSCnqwPdgG0cXD+/EgA1
w9npGSF49p5lb7wvAB8Z9KlYG6ZlgM9Cszb7ryrzFPcYdn8bSlgIiJRbwRoM2vWW
0g00hKg5B9xlTs7wjhB84bpU3QAw/p17cGIPP8WCKyxYx9c70tapXipyhECBd+/M
UCyDPMMKkYijD8t8yiA67s0eexT7kyWP5ua/hvCSeqQjihEJO9q6b2g70SPbfFvU
7inqxSfdD28e58Mdl2aZb9WzUYw9tuZ/p8Ezn34/MJ43A5Z3f2RSvABTWgzb3XFl
x41B6tWjMll+KsNCVeH3nQ1ctNmppsvRbv91mg5ck8p6YO+T8OPejFyk9CfqFYiO
ZKVsNOZCa1PElFufTucJTOTws8Yef6jo4N2nThfb/oXIuS2qxfht14l5Ca/tvr1N
mdwdhtQt4snoj8n2tybP+pvrIhoQ9GDhqNjaS71m6m0jPKjy6eJFJSAOOyJrciZ+
+wj/y1D3z+Q82XZ+jE7iYcKL/MIgGFzCxbIpce/Lf1JQ569Aka0GhWPEJYUHG18B
AWcBQCCtw25ObxBQOZAMTjSiVMwheqvatRPFWo1b/ipwIpRxv1pLckGPd0rhu6im
d++0r7/x1zXU6SYQAxXzbjycGVPe0Dk0KqDBduKpVFLPdm3UjXkfTZoZUWH/h9JB
bkeFs5VD9fxllIBXuZGZdHIhPLU1C+P0f6WLYFjKUB8oeEE5TYqNT+XP16F12L98
mauGHcsvivqRcdIKKnFiCEyxj8K69+Wo2ObT30VSDPucHg3jm1LyuT/5Om488XKf
YlH9gF8rwWLozL0KNoPfzuC6J2UoxWiqNkG7b3sNsHtrfjQLHOY+m6POqyqzdDvA
PXNYv+iFM5Rd72XPSITsZuKne7ikyndcqZd5tnR48Pby/QLnRgviDzAlk7yGrRhT
1/YMVbBs/p4wpRXAJTUThpY7ELY7gD8cV5R52qZJP6U+obU0HZxXEWiTGxtmpIr0
pSD8AYnmEHJJ31c9ZsoVGa3TElTWFC/6ZNG0LmN5w/l7XE8aJsYuVUEn729yGfB+
4IHbemNrqGhMuXs+yq65pmWWUhcLnta4tqky4a9NswvqQTJUrLOuYcz99l5OK4dK
r0XXPQtSDbiXPfJnmRAhUFb3n+4IYPFZDK/Sfsn94j3rcvUt7ghn/cEW7a6AuT6h
rofKq730wZjrFJZIneh19AKUiqVq+eYkSNwCsUjugc9mR+tldRqYKQy5Iog80dfs
I65ThyT0xDPPn0Gp9s6rcFl7eS4iHxgDfcuYeumipAjGbCLux5dg/ERTA9gdq58T
spQ5iuVO5PtSGOcKx2glqQZppTljP76MynLibEjrYcTrHo8VlqU5/TCsgZD5XmVp
76F9faQglC0vARhnW5DWSTcZoAOncFeJ0m5wLDd8UUah4UK0XsURy37yalMOnYWa
oIYHySx11b1MufiTNFMhcucnco35532XsFFCdjdLl61ZfRxApcnTg2rqacoxFhIB
1B6l/yo0jvtyLtH/MdFEIPVS7U1B2FJflyxzNA9xeTeIQxZ7Q7rwtNx7xr1QWDX+
iiHDVaxeMG8s28XsXDBNcJIz27MCIX6vx1r4KMrFH6vHbu9KhNHeXvQW1WRm7LCS
C4I7/juQo/QdpSq/5IJmGyfQd+2FxJvEIj7eEu8lR6UT7NR7TC9aI1oDb0frFBHF
RPbOmM1CYKb95QlNHZrJC2ovwTQeyh3LUqjzdOlgLXN5A3N5xU2fCxS2y2Ol4dze
I9D+93rwPpNKN4IkO+25YqdOo8ic3YB4gQEAYqowpyj28cETCydeL8hq3WPcoGNH
LALSsQB5OI+vRXy095XMf3xAkijhQeOvzhikkEtQCBMJbTa2XH4mppU12Wp3ySaO
IAuSFstxva29hweBMmbD0+0ov2n/EJgXT+gFOkJ0ws1cejCqQh6w0KK3g5kuvzbL
L/tlHs7tJJpHYqI0KUsbzzxGPGbq3u3EgzWej/jCbY8Ef9d5cUz/VIzGPIrYrKYK
CDXxhZnvuzLE0cNOj6//t1J2sxyYS6bcMHqtjGnR3QS2+TdXtJkrU4NVK2v8JC0w
N8vQ6M5aJzSrXpQxUgXOTbkzLbkt7nlhJsgvJUtInKXIMker4FzPQU51gRX+R5se
te/9yEDJZ0DIzdPU/twx1GzqCjYPKy0kNMdAUwrk32oLgK667vtzLt1TGB208I35
rLGm/bSV1yfgyK0SVsJcOqAMbgvUpjfgvtpXRMPPvAI12TAlEpdOFwz7lIPk4jju
gEvUAAT7doNbmBible5AEJ5guYkJx451oBn4m1IohnxcnTJKAyO9TExxOJVMAfUi
dGEIunjSvfh0lAW0tjh8opMsgDNBztMZc9V+oUIoVUnTaw0sbjFTwA1uJhQdzgSh
d+JS3jeFpGLLTt2EWvdn11lFTbOCm8noeg2qV659r8wojITnLIoNRMI3H76lSQUu
vjDbQXZz9Uy7tHZzCNmWePUItjNcJ05yt3fJ7MWc+4yaAk8VuCh+KLeHS04GsFEQ
wQ6qww2VvK2gvEjl8Zpzw9kYXM0vJs50B8KYP0vp8vHS/YOGdWvh73BIZ/F1OPZk
hNHqFVUl59zXvJNnVRg1v/+Sw47MwsLvbzjjLPbjqHOLaZgRQ9W7YbZgH+nAGL8u
oH9yDHNXTjzPNMhdqkYn6Gazb+/SahO2WgucV942f7TxS7FdOEgHyCugYpMTbEH6
VYEqF73B4CNvUuDuCYhiyiwM0rPGa7WsQILyEPSBPN/Dxja5g9kIcVTbNp9L3zGw
kH9K8Qp7MJ3KcPz5DDECKxUxiHopHvXkbI/QpYU6kQfC4zSJKCM6cwu4BA1woS/9
+g8ZTE7Qb8758QRNzpLfUtGVuZuyH+iGQthQX5y4PDyRQmx/zVX8MW1yJ7mTCXH3
WJ7e7+2GcNwwRPeqfz0/iTWIcNBmXzOiwUixMG7U8mt12DiUZy2TXwdiw5fZO2F0
VEZ7y8qHFkZ+2OlPLPwDVfePWSUUs93zx5uPCGZ4Pcvyb4BtQNl77md7/hGDxkP6
BezNJMJTJ7BrJZ+GExhiLJ1y0+zV5QXYp36UvoXyfJlFoQq7jl4CPgM83d+bEGFC
Z2rI7jQXZXw0reri0wkgSBNaxydST2g+P90YZQZX3bJUfPnivuEZfqp23yG1KY7P
JKiWt8Owyk1fi6EfLiUutHJjMmfc6oTiQFtFdYjoJkkZ6j7+dCXPiztolZ9agErj
asaOPPiDi6nQLB/+fgzkqzwe6wJAd+afiupkPq8gOo8T78O7co1jB0W3bkJyrg8Z
FUjEAdNQCIXuH1ItcBIIUK7jYx536/SpjW+I+kFtysHQZs2y7I+XqZ4IVwcfx4o0
j77pTecoKOymZtFSwAVfN+mtBIDfk+viwQXg2BWNKV8TtxlItmEO6KjIHXnL2J3i
vOH8pesPRD/HMkW0XfRwcVzOzZrzhoHNsA2bkZujCOc7UofnT3MkDmrLZnqJjFD5
a0ghPmqR4dvEOf2GbokYWpVWGV1dLgGGfc6RGMCtXSqb6iwWreBXsutL2qtmLkhU
V6pV7hrjSLJlGL82wYCnSYG2uJQj3gEGHoX7a2ftOeTLSKq8EBUfsRH0pIkr8IKT
Nlu+WWyNM0BtBZBCsCusPkXWlW6UP89j14ISwYWqztqk6PoERz80+JFUJH5eP74G
3ECyNvVo5lQVWOUB2PoeqHUNEi+suheCQVHOXSQcuR4e/KE7wvJeF3edRa6JOwjv
znzjmHOH1sXpIkDg6+iKouv82TOIgiQYzquE+RCXgfmECJcQ+LuB9hwQrMCTf2Ru
SiJSVvBMlyodo/peP6lw77C0mjutO7rIwpIkx+uEmlleniGGKpjPGS/Bs9W6k5TE
aKKQ7vhxjnR3rpJSvls9rMIkXxVO1C1D44VrR5+MwSNsGaPDQAk5o8ItXXOiEe8h
hseGchiwhvssmdJBcMYROlvIuFXiggPQ8S37EQBkSfCt5fWj3IkLXbPwpaoYy6HE
7cabpF+cgZf2ZaxoFmFGh/IYUMLXVZcjZqPEtZcSQ0z+JiyXXTfSn/NqkYj/BIu6
dup3leR1/TjLXZAOyZlBiXw9LS6VAVNZCxV5DjftBfqkzCSpOiVDOrDCk2iHg/BY
GdsHaXaDw37idIwqyCAsiB3lshIUEeinoziSyo0ipqL0yxrctVDY+hpbkzX5cAg+
Muk0F3eW43x1n2d7TzKDu2m3yJhrx1gwIT0EUQleJjr4E94iJHttBvFeXmI9Wg7t
iRvFlYlZ4+4fOz4U7KyhBvR0mLNsVK9KCWKFo9U7hXqiLIFRGUW4EREYXWzRWtj0
uDdx4x49U9ib6OL1mmxakdvHidi0vmk78aEtAxRYXNqIE3PQeAgg/Bnn3Hb/8z6o
0GYQQSNku6yOfSffCoA2vyPhz35UU1JKf+GrHlr+idKioPGk7jrInHkfLR2UWm7v
qhb5AmKca3f65H4mcHvtPtNIJnJbTo57vGVEviRjD1PANAONvUg6qErrDDFVinOV
URdgQ7R3lZYYwOSr3ki8uQOK+WxI5qKwRGYNixLF17Wyz2txT0SobjILPpaJDLka
fPEdlTpkVUM/bVpRJE8bblmglqH8NcX+S/E4oshqnBFoynLI7lU215i0jd/2C02y
Y+Q/oG9th2owFwQAt0TJFGuNUv1nnCoBErHO7pO8GdtjgS2ANLltKWfIs3BgnmxF
L5tqiUXOBNia+mha9qrWvTqqIJhsBf+GFrfw8nlDBC13UezEAWJaaCW6ZQvleiWB
NJ6Mqt/wMUd/qNRTrL/k+mMM4/Lj1yu1IiLH3O5TUMNwdqEK8o+OqSb66FPXXYZb
bfCzcUhRXRYHF4hXUOZRnI+q+xI9VJ/FCMY7dzEkYtNjokcJUzrMhiouwUnnWwQD
ReYXiVY0GnyPaPw7BYiaI5Zae7jEwtPho4vw+UFPtKc75vuElyVbtL67SwHFCVk6
72QLS3qEcMSjBYg8Qv4+o2BKTw7tLhFeVqLL3iYklonxD6Opcg6BSqoZX/39fStx
Gb45XRBi4jAu0BJekbrxfuuTBmajQqA6sURe9k5lmodgXrikDcRWWzoeJsskUxpw
/YCOvEvqfnX1zj3Mbx5Me47J2tAhv5B1JRlwwVh4C4lpuscjCu8EsorOlX02OwuH
+ykvy068TUaI0igVCGjxUxTykv+OmibPsPEpCCUrq2XUso8ZWW7USU4sjE2zY12Q
dGTcAEGZXMqbGd3ThahTtnfQDRJKjL4keMSqfBY/wqn8J5RSwTb+C2PFmKM7rfYY
01j/R8EtAbVFCxVKrHs2FQHRfNmsB1EFem4I4FQp4aCxpL+ystgk9/ll1/35wZnZ
iB+SUKJaghVYhXsKjtBRIl2r23W6ymVdJdRggjLSrzay/YuV3Wr8ePGBYSEPtzpU
pxOUcYIzPTpDa5mPebvlikAJ7cJ4HZbiFxyISLZvqWN/mEAkdOzQSpYnNhUwNlsJ
q9sUVL31C5pJje6QBO42uwmLKo3hrJzsA9eArzSn4HYME0bxo2bA9HogvHnNjHKB
EwMyyUvCz4FnygrW4sDENkWY/kxUU8H06Ib1t7L72znlTD/4aNAYugKGpA/bMFQe
S8iL3F1Kjq7Gs6/Jg/miPxD8Ez5aPFy5b/fovtnhffuZ8qbXamjTKALoUDtyqZbh
r+zkH9B/WXTumvAybXO8/z+Dt97HHcUDqwOHy1PgLpeWHJhA+KkMN5JQcya3bJzH
/wDzXyCGrVcfAz1FaDojHKWGLTPnEUJkxsKid0ILcHmyMCedWN5n6nkrPlHlxdsR
ZB88mrqo0VLCzI2edG8UeQ2zLGgW/bJm7TU1xgJ3yXZgt0CqYDXuhDSP0vb7tRZx
1tJf7gaQjz1ury+mrM7bSQCG90/m6MZGU3s1mXtew1LB7pjKtVPfDHqQZU58xHhq
925MITj0vbEZMCk4BBMJDOURk/Ra4vFHNfnLJWw6nH0IZFX4mIr791k8B4YdK3xg
KP/0bE1nitos8YAZc3m+QgSk6Bamkb8VXd+BdsIeL0FiBe4w2QbG0oIPWh9KCol0
jjbgK9mIdVo3r3gO4GC+9kQvxnfN/MWYRMDqJL//UgRS1fd08b2QH14qOI4jX54g
e2zVS+r5XnZrK0q0h9fUtqA9VMfZFxDmOoXCZJa6f+fVioC2FpFB/LJODZAYCifc
Gt7g0qIBvqqxyfH8TDancFAHCq0s9PAjkGb3mdBEIB3VVvcs7/mjBhIdYGjcKpot
hcEe1fqq2qyGm1uv786n35RQod5MnTXjjHo1FZJMWbxVIfQ+680L2LdNuxDj5P6s
uUhYGgicHKAuCaH6geH4U1rYZs0TbMsB76k4FKR3M/PRaS5ja9YEibX/10ziMUcy
xg6MCQCKRB2H5wxTv/1aKG+XPLju/dy7T184jje71O7fii0xAXvXf2gWj8+0j30v
1eLgvwUUyYmjRZDSpskDB3dJfHxq0kcU1SsVsXgQdo7ZbaMncOXG2mUdWWmrbdHh
S7jt40CHX4NQntKOl95WvwmMNYMcfQJJtU/5NPdEnx61Ao5gvOtdrDBEmCqQqlVU
PeM7pZb98o+0LWo4HkHit/Y1ksmJYsFk7jctmv/qOtInG1/25mRXS3Mdd6w886wW
hc8t3ZnyVeiHcV/cgNG4GwCcXG++ocPQkBi9v5EOuYK/AWdqj9TtPew2I7nPg+BN
s73j7965XHY+SftaJn99/8v26gSbEw1w8wTlwcIUqh1WbZU76eVuVzA0silivIEi
xJssczOsBsfs3scAHtPt4AFhDpxTzAmAhJRRDHCqTFRB6xWZ2iZmmiMEFAIyP5fM
jtptBdUq4aE+oLb4r/Oy6YM0Mrh2Kqn/IlgdC9h/FbwThoP/+2dezn1KjZdxf0PF
7fgP3s4ZtGUWRqgdMgWMiNlWjk0936261Mf1wAhf4732tZCc3GPdzHmqN/iBH6dF
p2LCoyQP+V7+rdTg5+EJ4MM4u7o5/FhAqnHQPu3SMcK9VVfwddzDAdMluJBbQ3u5
ryegyAS8AXw62+Cqi0IGMuMwdnLskHPTcAArttOUTwqBzTNGM1feCEj5BB8cWGL3
x7k4T9cwf0A/UBkLW5dZosno8wOChyykXGALJSeA+vGXmhTtOetYTu4zZe45Iey8
PHHlA0gdeoPwsGBPQWFCMiNMOFBIgi4JM4f3UwuidnxyLm3HOygOPRXisvrCkg9r
psvVW/CkbosZpTTmWy/eNGz40q+ygyVYzkzCh3k7SswJHEijYW55zzScA20YhKdK
SQwBF+kNUS8KCGHrBiWiygE5ZVnNClvatzKOrBlK1RgNlcLf/AcowHN7OXASO2vU
pEvQxSr8iqN5hatauwShOMOfSpLS3jor2fouPYVzkbvTfSHOyv/SMgDxgkexEV85
mPA4ucSDIkvmscljmmiih/7D5WKBDVwBvsB9LjsDvmO1ogZbr5YrqriQNiKBK+gH
M7m+KqMq6EhR/woROZ5cCKkObaglifiXR3aYb5N9M1MXVtec0WIVpgXXgyytJirh
H08gfGjuBo5Cyx9nr6P0dZg42BksEebApbraYNatoFW9DnEuO8HPx6X42eymMVDA
FlombbwHEwAwrfDl1PoGtkWeMPOTqWZWVwE+xZK9p3pp/472HggalxHUZTaVZI/Y
PXcsT0IDYyyXONQWku39MTxNDhrhbMNZzjC/defUOiYkkM9vThF5oAMqk/lyvBqz
FFOeAVEIQHTfFOZOY5jWmMSjhd1Z1VTk2Xt8xu/p9sb4Nxw9PCuBWfgGSpUVnTFe
EKrhq8T6k37YI75yP07j+eCW9QpuQM49S+jW6+SfJzYGlpxNFmp8DMmpHHrL4PkD
mye0AKV30ahSAsb2zbLaJot792gueOudZ7IWXzENFZ0vgLkxDztPRSQOVxrtRC+7
Vp5PeltpcfUJwRacIg9joXAP+b8seBKFxS/uoj4hgwFhhh+hucxYn6hAzKhQDvKW
wIer30Hw1hCenHSN+m7jdwnPSEse2Nmtu4J0qclFtnrrgzCQul9GMCebmKfudbR5
ry3iASBqqFQUY3KNnq1dWYvYQoSa8VfAK0V6lSBbo8OhgYh0uUSPNzyiORe1qvUY
iIKN5sVwKhvBz90RxnuR7/PTu1Z3vMwQl1/t6K31GQLfGzrq+4CUadEs+xJX+UJA
8GsSIlKSQM+0KSi6PCJQBkmtwJ6mKsnVP8hqGdAGoILNSzWpCG8yTMAa6ox1ueMX
bh3YU2SiAzzpzAHJq4wRw37ol5stSdyklPCctcml6IRNtlhQBbIYZGJD79VGRCoc
QUAsCZDa+1qr7Q5jUoSfOtwW89gHyQyWZb15bE5TE0SShi0xrJEJr0NGk2hXWZpA
qtjBJ/CKDnJ31vlCtcVGtMTg+YkYA3NnUgiXHbsI0moRU+YsqLOOoekFRTdxPRfb
h4qYfR1/TIMCP8qc3ImAu3xQDDHiZJTUBYePO0XXKCdUHhaHI4XEGAgW9cnf7I/O
KwA2ftibmopvDArplWfJouT1x7ZUviwscAVKMoWAmRFWvT8f+fBzjuHvHx+opOAF
8nXBXixmKfnqW6uABKkiLnKhk0NYh9jZGlTUXQumCNaCm8+ssFfMPScbuVxnq2on
pIWL/LkHIyc2GH8aShxTwo1RNtjhN6TyEXVP7vc7mgLvLRB4d+l//UOPXeHcb4PE
W4YfsKKCC7te1U88d0TMIW2Y6ovoUaaGEl6F8wIrsilvmKjRPvWBQO/Bo5I34jcY
IsuEOnWOHNg3BvzrwjRtCI8T52Szl3rniAniFd+XfGoXDRTyoyrfYrkLc2cU6min
Ao7onnoGZaFQq1DAjBUSsH8B8/9WpxnfXxLY8esNf1wQOXNnmzlmL8fUzblGhA/N
Zv2+gAc31Zv3XWKQ2/+IjU3IUF4htYwuI4GLwivE0zBox2scmUdbDWRN+FIOQAlE
V4YKpjTRwXDjW7k7V0BK5sdQ4iG8QBnHXwYVOtb3jItzUszQGA0ibEmZWTfwEO+Z
KpTn3CHUKmku4/wLwNZY7Bcrt6mWvKkO2K4JIjKRgpEpH2bkLgtcrgN+/aFrfYhp
95sLaArDdYypWQ0BNbBUUx6bIWfC0YaB4AXZ0SdJg5NLMwdncmYy0bYzLeOBrp9/
yCIFIUCvtwfynbKnmAnWpZkrhzjt8f36eWYn+K1IRlBTWqdlZ2hUaZsk/q4qzmYD
UggjmHzP8vus3tPbvAk+aoenj4O7bkOtq6h0GVWiJxWMm8UhAAzBi851U7B7DeEh
GSG7pEMePrdRZ5PjdSrL4u6rFkfQbxXRXvKY75i8vQVrqngNpcjjSvb/ZkwZzv3j
fte8VgDm05G8hhCQiVsCIyaSuITV2frqSZEZH9Ms3UJ4uxwbCYT18qu9MbkdlDZm
0qB8se8Vmy1P0bfGHEJeyPmho0s5j2Z1oSHmqXiWtcWE79N4qRRjqeoUy+mipWSH
evbD7i8MLDZ7xTUDjhFVVaWoj/PJqXi9InPA4gGvzFnF2Q4zD+RuOhocs3egLVje
ctxF7n9MGrjnrG9xiwiRq2UeJWHCDmF8HLruwNKeWfsVjSGfjfL4G3z3sdIFJg0Q
mIlsRoYU1kwmmyrXaea+cmV043UF92mD74yC0NiodDMqiD6Uu5sIAcdmuI/9L+nj
Q5jfzO4DPLWL5xrJtjsx9zYkZI2Te6SBtOtOwUkKd+fFTElfYBFaUqctGPvnDM2w
GAxTlr19Qq71Ub6uGz9Fjs6QtEqlHcm4UbKsCoN7H1lA6C9mQsniFm7K/Pg4PR6E
1YowJenhq8r4PJZQZ+9ZAUu36aNV/71LmLD4EYbSAzGRS/1UFqCy3wqmn2F7lbkY
r8krc7GoAzT3vdRPxXMWueRREmGksgz3Bp+eOXNMqr9G4Ta36y54bBSUxr1oOiAy
4dIP8+QHegWmesr6KvAKa8vHTEuoH8pXUmB65CvJxwfZeGM9WBdUNHtCrOx7X4Af
g6cBFH55H221wLyWOJVidYP2ubn7QMtB0nNANNvXSGxxUMvh0Mx/2n4dl24tMiMe
u5iPhdoOTuZNfjabARHj9Zz2RIp2F4HTyIL9In7mAUCrINCPqhdsb39en+/lSXtf
7ixAePlo8yweNFfRu2jMrnbx7oKPRqWv2Fb+g3t4GV00gDpsfkQUP45OySkNrXec
9CRjHnRbHxOlrbXd9QdNzZFE3ItTEuPTc1vdML37gzMVyQfZYjcrUPCKDIW2Aw2H
mg14HhGflvAg6UB3Xjf0F9iw2LyQLwq9H5OwLowOVIdPfm4cHXYvCTejYaL7mPmO
OO+iuzSavUJMIS87Q3cAM7Rl4dPAtyo7Tk2tUhcJpwixxDA5fIT6LbImsxk/Oc8w
nCSyH1byE7wMr8pXN1RNvCWuBAYMv+dQRR3XA3H11y7PgIFBeheFIILhiaE1vC55
DXG/z/7GDJH+n3bxD+I7M47MHO3dDNsjQ6qPa3k4SmndaX5TxC4euU8yVFQQYh43
pdVrW2sZAF5gWh8uRZKqHYSjAVdSamuXZAJIQVOmC9J9iCMAvmrk7N3AjBcU1/lP
YMJ01lYBmFFEFrutPnkjm4iV/Vefw46XBVsuL9Uh4s5cJDPM2zZxyAcQE9x6Ldqu
ERv7v/7wiBlXz3Coyyh7YM0SIXaz2Osb406HJEQK8nAnf9s6HFsmdOln6snFTNfF
tWhyQ4gZlLH0ai/JonuYfL+gEq65aFfB5IzKLzdS9eOpiynxI4X0cDHB9xln5Ofm
L7J7gJzNSaomLU8x+MoI1bS4WmtwiyXkPTEMGwJK178vhqDWHP1Um0KqQOGh0pN6
gsErb5icmsDRiiP1vzIUpsE1sbdhc71VkS3z4WppUS8oqcoSZewBcgvGgsSBCdxt
PilJLuac6/knTEs/o68DhlzlQDs6My1QGgVdmTEdMRTtAjp2Rxg9qy6lEyOraELW
m1OzBG8M17mBw3LlwXcRVKdHy4dMqCduqU4B6u46LFeQJJozxxdojZIEVFJV4izf
8Zp/CbsGoLQUOLbIVKWM5yuwo6vHwrXsrQOijvP3tVlD3//1qYZ3kPxI/pMHIufj
mkQlDgvMwp/ephKzlFcAb04LmXDnszNwlNXCi1fQrwCRIcCWZ9u6DRo9+/NqFZxl
fO0PoYZjrdtD9Fn6pAcjOzFhGX6SMGQ4OidxuBWTdHYewUevSWFI0C7txDxHeWnQ
x/6Kb1dqqQzm1m+E2/X/jW2iumV929T4Dh1YHWWF5IJbFltKHUs+oQtavqj5Xu0O
5fR0PEqDKHWuwopcNvbkEeiwXfbsJg/cU5MFmiy+VlT9BIOzZnzalYqzN4IWDLBh
y5xru9RURJ5bLAQAOLrPGudWFzcW1DucDbChi+jM6tByLJNgcwGID1SZ0SSbIwNz
CpAz6lHrSGmQo9JM6fF5LpwSx2G2Y1R1fFsthUC0cfQUsmWPCNN+7TKbghMPy1Hi
haMGf8pqTz8hUlsDDBToFGbyXudYW6rHdeV+hfm8x21o5xJQ6waFaKgVvhU3yYjg
XUKYmzDmpCJKa+PeaV/g2KzEf2ve0+AHiC1Ns9BjMOSrycyjvWHJVXocWZTznQOb
+N6OTzLKYcSH6K49QkW3mofOAB+U2W/p/FlUa9XeUILPsnuTcsT3xyfNZWKgPoOf
LqHJqM4N4md9AHedDLFKgWC2mZ79TRBbl4awGZti86cDtL2OZLteKqqnm6LgfCjf
kIhdb0oEj6JhLCmVX/2sYZus2g/DjvgyVYtz+LTSFqf3De1o19rL67EBlfR3xdat
JBD6dcpU1B6O2R++fmGxuggnSbEoyotP3WiUiZVUAHPMH9CcFlc5uHsaV+pnGUSh
A8IxcV6gQliN516wt23+FnA7eZw8lm28Triz5TEgQK9snUC4JpHW4mQoZoERdRrm
KcIr+ozKCJO8RWdQeo3XNMSWJ3BbvihMIadRt2x3ZK9yC17+mHo3+c5839tzcTch
deujW6pznsG0T/EgwRYuvE7hbE1jpgOOouvi6iRJKNofSWmBKcYb2ti1gLGh9F5G
aVYkBbqhQT9++fuwn+jE4yd2341zWKr72L2MyPyemNdj1nbMQe4FMJwohkmzbEor
axtdRXvj0hnyfbqKWq+vU//BVZqV7coVvdOjVtPsRXeiVGvjJip8OigKt5Ko0Kgy
rFveyxoiRGlcH12IdSFt/94UH4t150dRnzQu1GU0RKbfAdMAFiQDl/6G+pIPCORF
6YNKJeH874i/5Gx/I1D+puzoXYUNVPbtywitit3omGet/wm/BLbztL8qWrB2O5R5
U1x6YLq+qGrPN5Zo8UAspQKhn9cqIuxMa221X0RANtA11co5aglNLJ+u3qvKycxq
xg8G5fnnrAIZgZZ/39J4Y+o2D1NfjvIlwik3oSrUx/oA1Yk92laX/4yssdWPlz0b
aBis8dxThVpPe5uc1dd21xyJzh1awv3Hp3HpB80xbRxLHWTAAteXPQvVtCxqcKz9
Uk5bn3F/F+93g287S+0WtQ932fj9MeCIHyqVR4NOK73BiOs1M7EZKRMqEtUJGhRA
LbSXtJ0txGVza77rhHx8o+uEwZVCE80m0Kx65UxaB5RbIyO07Ixa88ndXK9asRL9
oGxT3C0DeGjYmCMnWchkB9Te/tNtqj5xHZRMy1jD5pUxY1LGmNAkr4e3ayr/VveI
oeLx5N/1x/WElTTI4M32xvMhwrn6VNuZ+gIgUNvYZl6Q12NmfE2xNC9VFJU0RtWi
RmWgH57PfjBnnl20Z5X8KU/RV8fJLyd0GcL0mpft09hQbKsprMcSHz2hIomFNrEp
dr7h3q1dO/O9/df0/ePBo6pvSztv4Z3ozLNllO45dUxzij7nG1ozXl/rar+CukIU
z8XtcILngteg6ul/+02Q68YXXAAF+bTMNg33YYe6MTEsH0k4UjbxD2pJ3jaib3zx
06jYnC6e5sMWZRTKZvou+qZ28zyMNxcy7e3mbx8hAiwCdcTd1C8TsVJNGAmneLU4
F3viU2trA6/3MErZ7wFGHzgFQAyib2Vfn10BQQkbCf7lRV+LvVmp/9qWvxHE+hQo
OX5goty7ol4i5VbEP13vII8dwpQDEs7/kV2Us1cyf03QujVt+6cKic2FXE3gq+B/
aHsFCz/CWr9an/YVyhAjjPD/3vdHi0kMFqjHwaKgU1Ws+r8VagBkE8wFhdoObXZ6
CvVgoOnyqMFjssD1qsqKUihLEM1SxjcbKk1v52RgAIpKwxCeej3ucliGPmrqAS/u
UggOUDx4IH1BV6k5PusxdSFKr2Mte9xHueSO1cBickflmMU3JhyLnFM1oEuPXyJY
npCilDqpgKM+Q28uLm4vWkEC84AiA0H3cHyy1UZS+4DU7VPBU2ye0/nm1pscw+wQ
3WnwfWAt7r6CBT8RKmCG1yKzJ3fwB45z+nUOXzupUfK7Hmq4NrSpaHjhRonA4ClP
hBesNQsrQbPswH+tg/5ba22j1ic8jIVllnP4+0mK/AUhD/HlgJor75ayJwDXqLMm
usV1DFaQpr2AEn82tdfybOruIYyMK9QnuAEkv+kih2V8tIaHDh5osiuJFWgng4PD
9ggxrj6Lf2CmSN/GPTuKQTvvgkXT+Bq2yIE5i805V/OEXgDQg4NCiFkX50+ytMay
4LU1k0DlW/YLKYW3vWKH5cJPBgxT1+sCgnIPed/TOW/CU6vbNTjvoh1j4ZXq868G
E9LNRxS3mHxegcFEnWv9n0nvsdLkhV/KHP6ZbXXoC/4VL3e/Q7xMQsAd6ZLfJ6x/
yhR/Lk9jA6KJ7XXuhgG7uXQO1xZJBgj58urxei1eq4h2ynC7KLW6EbkkuENMnCUz
eia7iBlcfCHoCoRyhCAbtIQmU1vOdTlN5an7WSlE8GbkmN1YAXfzjAr7Sy7KIraH
1YusRNQsNuYHU8k9l73cY0p8vjRYejGJIPCaGltUHdVh5DvmYv+AJy11lX+1QcQB
/vXxdVDdjtT5yPoJCMpjpjCkvs5IezthHk0pEW+KuEVyoEV1Gih6armawy0p8fXc
A7puYicFdpWtTlSoGBrUmZ7TAA/hykZTVSlSPcBhb3HUFIFtaQbr2frCt9tse5Yw
E22t3dHTehUmdc/HIZ6ebAlNCWgZXE+WwKcZgOj6Odra5Ioq0UfkkDWH8WRsXA6w
D+lT+kJHd3SKWiR1c+ld02iD3zyBzQXofgqU+iXuKrO8sBilcAkHOT6fqNUpZbKB
RVufpjceA8Wn+i1QFpgf0gVETvLylYLSZ2GBrMbLenVxJxUssXS5xxLeUdfV7T1l
m3PigjMnzrRpUDDqQ/nRp6uLjfWn1vZCpwgdtLrlkq/rt/zqE7LFq/j4ziJQREmu
9FiaiYBLZIjJsuv5VkANWYWTZDAKmptfhJ1pO/HDsGGZtY1YUHmYNOHQfOWBln7Z
6qZpGVdP0pahoU/J4Lwz+YmGWaprc89qqh0qO57hxz1WnVUgrzEZphB799qUaB0l
Ifu7Ko17tHXxcpZW7yyqcUzS8iRt0DGYqybCX5hYYOSJX24EFPRnPQQJ6EWfhU66
qTbxElK4WXj3IMri+iDWIRm9e5olfHFVz8iAcYKC+W+Y5sSBQFWU89D+3k084CIP
PpMaaWmSVe9tLK7cH3CDNW7ZJ2jR7NSebpIZe6+23tPZ4hKa+AsxfyprTnJw2Qc0
ChThTjuHmgDYyQctuy0EuChKrUShofaxgnc3+dC/UcY5yUcWnUm5sSBYMy28/pru
jOSu3lSxqT7cD3kBnd1iP9O7i6e2bcYGI45NiHi8+zh54N0mFYAXH54PzhOh8P3p
clVtOgLBbzR7ARDNJgAG4hawyIhi4dXSzo7Z9y0PA8Gb90iTEeLQsxcnS056mJ0A
iBLSk9ImI7ohf95ZQovyNXC3sytvzrhFqW82ClkMkTuawXJj4OA2Jv/3pTn7q5aB
akhGPNKzqeNFVGxAKl8nEkeHHm2XfahEmhpJJW2BELkzvV0sFH8tI6zslpPFMcsV
pD18BqnMd9xZIPDbjeYtknOxs/FQe0ySchHcHlrxIs2AM2O1rlM0WFsCCWVEfTLQ
lNvpXEX4wBiwhXcR+I1b1We0yfLlM9H3dSoN6aY7CltySKA9VzEQGVKaQVlQp0Th
qCbi4Kmf6+qxROTkrMEwTsyNr0DvR0u5Bf5nHkfNXIJ21H0xNvPjHuCnbII3pcXG
Jz80Z5x6w43qtove57P8DbuZ3OsIK6yZXVbvSPV6ze0j7J5QVlXFQSMLgmyRYM9F
4WB7fXnyDyWzGAAbnfQ9xQK9bpG6rH8nBA+vEpPqbYY+5Yiq3FYTshiM23LVwQnb
HchRCJxW/jiOnpMGcLWwCdrrbzK8us4vAw6QOvNLWtjcpgejfir6vCd9620gNYVW
BjQChCb5AucozRFcWwKpfODr5JY3yShEtm5Hg23G+FHDpNGYnLvrRlQK3+bIUcrL
fa9+Z0CFR7R6i5xbD+GXAgzsVveJBht+UBuh/+OP1Q1IYlGxJ+bFT83wQfI3zdsp
3yAysCuKZVRUFdTj+Y7z3D8PvST42JzWNWyCsF48QrTYeWlqJUUuNfSGvrAFQY7J
xKFYHre2nMN0dYbsZ+Lqf0avy7qTJYb5Cfl0gwpWJr0yY/W5X7I42oUN8pMoUXFH
OCD9VJd3s/vCO5BeyOfRU7TWsU8IbAfmxJCQSV2J3TC6dwdYbmO8HPKDgxlx7I7V
rOetgoCZFqY8ylDdXL7UuDwqGuTU+y5UILw7HK3zZiPgH7XxHyBfvS/IxDNswyDP
mcoUH0/+2Rp/H9BW+qOAsmCAYbKjxQ0WbqOjwKZ6lztkt1WM/2Cr1hj3ihlRRr+1
VePSr5cLjdHzSRbBgrJsNYQD1gVAsvL5PkIEZw5lm0uFgK1erqXMfgk31v1Ydm2U
JT2zaKK6345CTYzTb+4VTAZF6IPh3cVfkO9R3mC16V7+xPN7XHgg9zpVrtUWlKsU
k9qCBKPoD/heGQl2SDC0hF0tvmb92RBaLjO2oAzDk+HJDnVrLtZrxWVltNyUSEHM
oJjNzn6NxK+1r6Ft0yO0rvpMPJgoCMMRXl4mQ7ffKXYg0BysOyTnv7yfgO5+4Dh5
cwSof4HFXgYvpLkOTW9sCS4scvCCuZNuMUqY9qL7xYvPNazYTUTMnv1BoAeYDhjR
q6Y4WWLrY3yWMJHoH1VZiIZ+m93gqfW9IqfmBvXSd96yhq7VumkZEI5q8skA6mpy
8heGNTgwwNIMi0K+HJMy0gh1DVsAraT7W4y6OXQNRT1+6Qjknyy/kD5h3Q8T+21E
Zlq03c/3QUo7Fglr6lDvT+4yG6gHc+Ldn+3Zr1O5LEAQIPFp3z/ytY4z8CuWlgQk
xlJEuJ74vqfeJ5eEepiN1mGG0DYeBqRI+WzIb/aHZCibhftvwALnGFaTxmYbRzUZ
7tnoBiBzLn9yqj6ZnbwSzaPwBRURYIrJ3IUY8a6fMuXNTxGsK+nAVghbwV27Z3sK
oVmzO6z39rbwhs+b8304y7jAMlH9oFJYFT903ygueKsBap5J/dn8/FYOVsLJ4U4F
GKIJrVAfT/mqXiJtfOJL9DnOG7CmQWYAwbW/BtGAMnan56bT8u32D5GVG3/zdWtv
N33js67kXHtvjjtTbylH71ShSSGbjczDCrwrfojZ6Jf1ikqDNnyy7t+8B7wuPDCD
6JHRYn+lvM2tcdyOktlgveu+Fr7u68niUW+VZ7OF3FKkvbkZsZNZjRWyrihDsxmP
/8k/vNfT7/q9CIP/osqY56VtztHqsv1XA4S2eFBgOIDa4DylQw5PdxU3MDmBvCd6
4gZaiUHsyKH0rNXsXs+guORZj7Plw3A6Hhvlh9z9GXdIoqOqJ9UQY0F41ZCZS9MV
NmaFc6Jle2zuHm04NN+yePSWpsRuST/wDpXLCVqf6Eu7OAkgoYTQuN3Fp7X2CpoK
6C3zZNt8GkXwC58qHhAoSqUsPbcTOeD5P1KHsvdvRVdxXPmdYCqc+NQaZQ5bGTk1
2q2Io+EqCTAZUvXetBhHsLmBnSXE4m9K9/5HuFzTYE0oCeBymftFCzA7px125MA/
PYgZ2JsgArcVtdyTGZ1KkSc5wzrQQQNF89nq0iam207P8wEw8bhfXND84jUJrKsc
9iirHMachByriXpNIcldsqWCZu25EfwaO4EL1lmmDF1AsWo2+BzUoCaFjPRASkxC
sChCpKcBC0YFx6DjD8jfZCcpVLsGxNI8WzC8raN1SGZ1H3iKhTSz5NEhQEBWpkdj
gpBWF3yRt5DLn8KrsYk9KlfGvCBLnwenkMG1uots2jYBOd/WByDlLWZfP4T4j/64
t72L9wyS9TKjn6cXgkDGaUWM+LGjUWc3LBdKz3LGw11P3/TWwdYY31RmRjW7nXs0
/9a6+oD9vuDcWtBkIIzU8t1+JW+Psz0pQ9mSKq7Z0Ji/MvaIE9wmJ3g748RDCxT6
SIxNtW8L3HhqYz9GHqCcq4C8Ow1rurNURpACtarOT7cGUMbBywv4I2fZtp7OIrOG
jD1EloytQ3GZO1q2k/Ew+Ady056Srt1vYug+nRVZE1JJmrr81vSheUrf14Q/xED+
Z8IRJg95UuT8iakJBqtp/AfQ74xytCkmeWqBZb+N2Joz8BTDXecXvvRatSpqBy40
pPxLIQ9IGE1tFGuzyBpx7NjCRe0FlTm1kQbHq1VoONmymAx3UTYibcS4ciaPRBBl
CEM08YBkDS9booYZeGYDhghgDLt0dJuK8PIgxb88npz3sIwA5CXYYRInjF5L2s1q
USOxGupfvmyYcyEuQowRKjJfnIBF8Q586kVsVYNzqwWjFH1OTFTxhjOE7nOAbyTo
n+i2lYZzq2D///gCCfAMHFIybVMpr2wTcSHb2BOpihzT7LtlE2uH2/pmCiGWhjpZ
ljeAw0smbiSB5Y/kuRb0u/fcJAFo/AesmRpB8p2prWzriCi28Uj8lZqqIzpkBUbc
9/O87RWpa3bIACqdorjHkCjQI/X37QjBe7MDqpbPYjVqiqo/oZq5kAnGVUUStgTD
rJ66riIsqEOo8kkigT37byJeMoDfWxu4EJp4SM1+R09BpEDZsUgTUWafZQ8mATex
FR0SWChisCyIZNELjqtJYcg94th5pm51gNrxywGEz/IDy/zK4HXq0nrpbtO92KgQ
1j+WOYFD9rArN8QElKiX94AkKtnpG5LasMlyj8dW5sTo7NgYvNX8LeDQXIXkJBMv
loZf5pAI1gwJGsnSO7e6bDgemwqoKWE4kse9iP2UlACbk9ieUrBrNYsgVaBHv5cM
i1eMJ2SfK/mptecAdv+SF4R1LZDhi6SsZF9eCO9QUxtxtmigJ0M3JcDgFWKPfnkQ
P04LEwKPBynozrj0cqan14y9zqLWPPzrKOvz6JKiTIN2qZW3ogFvPar7u0iVhOgu
zIxRKXLfj9vv8idkU3JJKGcRCZPL/87eJqbE+fuuO35Y84Hz0FAazR9g08dPaOC0
8WWZtW0fLT8HOJ85RAgxfMJk9Tc9fGHoPO9/w52YI9zz/1H6kEEgrEm3/b3Jfo5d
eXlCSR+zyKcJibnffikbM3Qa1BNHk7phMK8kJCNF1shxa+h4LN0MMuXlkCbkIM0r
YrW26F6YZtGSR2ol6Bm5XZSq0P1hkf0Wt5lIZz0JYNk2p6QjHBfNGVBCxRCahbUY
rAxwR9y2T4EkCfbFZ/fM5S9Z5AvM+pjbOUdwegrrtEFyGs9uMlQbcb4NqH72pXwc
9+ivZD/5pX+hRNvZziwA2xvSutD9zIdt7/Ys9FlWlU2tbxrYl22w6Gpvfz2CY3vI
J2JeB0hpRLJ3jnrVtWvd7zXcDCCQ4oqApwVaTnIlVmP05RAiHiATyGVx5Kvu2X5n
ekok4r1FaSC1vLrwKcA0/LVUdgeEKa/4bPZj1jveLY7IUgFW4w2SjXFY4kfOJvoB
DkwtxawgstCaEYSKxvgOYWOV2jScmMdgiyC/USpDir+sf6w7Ej5Wj8ANH0sL/4eJ
/cg4/udDn4+LmSZgMIT83eCMTbbv7TxLcPw2zTO+ajsb4FKn0Ltul4TLiKTF+kbt
jKgmgiKpqe4l3pysJxFIgTrqnld5vZLgryAp7ZozqAGnsvCfcYcKDG4yPOVq2lxO
LxFMvmf3oMDuZSH7qGm9qQGMU8V2NCI3h9k5Vwjn22Y9VGIMpuHczcOMcPll0Y2f
X38ffsL50m5hwihWksO5HBXqk7uWqqrKXg0Fk59Hdz1CrKR3R7Pa9iqz21SQMACl
uvzUtCKSamdwMFGIFkda6caW93tO5P1X1kHQNvjoLmSPQ9Re0HRZcc2Kd0HRTWrm
3kHGSV8b/U0HCvYiUraZQrpEFpL45HgelLuukqGX3eQOR89G+WuRYeOS4yZl9tsd
Hw4MQFIPd/4ISwgimBg1+AhnIBuVQ5l7tUyFyUWIXcUpQ/KDP9PvxPNpDHhI3w53
9E6Xpjnx8pnKRP90JCT+TLkE+1y01PixepIZp98mTs4aXTY7iiCOljK1NRMtIHuG
ng4OcLYEqLqfYqEazmpCxg/4wyCLbVtF1ynq40T3sOgkeJTIGMzjJVtGxjOYnH9O
J4z10a/EIhEfPZp2c7NOim28CqgZKTqm2XnzY9rAhR3XAdpbL9diDqY1uCVQHUB8
bpV/ZQmi63JjYnhqe2L2Tvxyo3N5aMAiGm/TElpaVqhjKB6f2hzzpuISYb/tuVCM
K58My/Wk2ajsTnimca0GgzILwKEqZgn82xRHFnJa0CjrkDWx75FMFcVNclzPijnF
UHXRRkiLEJXVjxDbejcM+WO1l0zCNA1+51330t5uAm25gzDxSKZujdHx/Wm2l1xJ
PrItwJ63gVHeU29wAXxUAnaY3FZkNqpVFen6HRJ66I6W+0ucgGpvAqDd3JVIidot
ozb49J64oGEZnVIDXdLoIvQm8VMx/dxEQtDzFiPEsCvUKh1QZt/6b+ndXMoRdjMA
UlA65MX6SevTn9ede6QVRUR4Fq46t/kuksjS6GIj5n7ACWgeNRnUWg9mM+MsM+fc
QPIdVMzLpip5jY/e0Av9duvFSNBVfJFR3fi0Sakj1fEh6MXSSFIqAlZRFdg+jy7Q
KEoPz1AoxSWGEyNK3vxJEi2YJ1jTmix16KK/ZftMms5tz4ZVpG4kzckWw2hQLznv
1d3j8NjD71EWq60n6Vrfxo4R71xUG54n/6KEWDp4klLajvl73tQm19/2iQ58fq3H
i+khfhaCcUjUo9GLxO8DOZtUmMkrt7Vom+gwTC/e/BqbjTMPRfDqqLVqYBQ9rke1
1/zJ0zVJhR2pqv6Iir0zPOHqdNEiBFe9g6R36Xara07U13bFxS5wZkfbcRMaY8Pk
ByO1hGyrMS1zgM7ILBLZJI2HzxEwlJTvcROg0aSlgEhffqo+Ih7xw1YYMrR76TaD
D6B//GX08nKrzSdBjLv3kRD/C6zkaJdEmPSL/dofPc9eL1JZCihRmLiXTI8RX7UA
NEza4RzF+gTF+THOlObKtK0OBwd81Tc+DV0bXGJThzZS6z+8hSgu7L8ZydYn4WH3
7IG8O9esTzddHC7VJiBHqMr1N78PEKa5njlNj4CFOK/+lLhKoYdOcsx/NIoOwdAW
PPk/4i2L/J1GKueDX0qhBVr2nSNImCX3blzCmLGd9llnO8b+S2Vm5GeHo6vQe6jb
Ew80P/XJJuDk4XG7FUnwyqVeHEb56gP8P8PEQ4PFk3grcjNWM13uiz+MrgsNAA6y
r7Rqr2B8ZJj7bMgpi4EjdR3iyDoEPKX8FvVqzf4P4E7IpQxepEt6bBes0HQcgoEv
aaWAfHiSqgDlohzDrDVQHuLWui1ZablkOJ2SFPZvlYT5w3qwS3JL8kdWDEtj1EFI
n8/XYpjsq+xNZG4M7LifIEqsTCjdpk9Tvss3N6Dmh6m2WIAjhJgb74bM2gurTrOK
4og7kG+5AevpBrts70WoxqseZJW9rrRWdzdNv4g0uda4T+Aziqejr7r58u9FTh2v
93OLtGOUrj6oVBjWFtbqsIHpJG6Tbg5p/bYYV76P3GyVl1NqHsZmhTcYTLBK+QM8
rXr0elx69MwnI/roJWcpbYAqJuNuV9H99a5otUYLVYrC15AveG/6E8CNPlQvgHU0
azLUVC27WZTD2phsXs60UvhZJ4KfhoIuGIAcuWQL2whDerhnK/hIm7kP1Si3Exur
NW+LS4TamAtSePxs9n092bj9U9OHkopJgyw/IsgzKT7gn7QLolaP31ib6ZfHKTqG
xrCJzirJ4M6xOURGTVdZugq5xF8mgH+PBhg+PjpTVI+u+bh9XQLbGN92+Fts/8L6
sOdzoldmm2iRh70+teu9rFQACBAbB8m59R19vgP3+LCzE+0/oHRn518NjRn0dww0
hdWaAtoBWC3H+IWQKhSJCURJAc1wUPZ5HpxjstZNHi35blZTPb1V832FQdcP3saX
utCWe67WB8KILtZA6Y6c2obYRmM6zfJ36Lgx1Wcw2Zxsop4crdauRA+KmBfYTRma
sBljuDIMyAthhhZBBVh+7PhWzYEHKH36U2ZCHgD2/NgD+wafakbBrsSRQyOmZxFk
6s2yjeiT48Ad+WVtbRZiwaA1eAicWpSe3yvt7L/hFS/jI3TIarCZ7Ucsa61ct34z
7SmS344RnPVDZtonnuiaQjoqYjd9dvk4IOqSvFEJvDBRGaJgDNOLPl9FwbfRrWeL
F56Z+cL35Phh3APxQDQSf5Vj7MTtmysWWaaal80MfXSCZUSQQ1LuVFz84nCylvyd
y7291jgWYXDpd/nLYYGOiK4987wyH01gHCCir2CJTXBlElv1vN7RqPOR0x0+NKO1
Jd8ToRIJ/cdWcaVrO/TpzEEUvmaGOY8oZ3mpvMIdIYJI8TTzOfzI6/luFWJGTuDQ
DXRkI1MtOwQhK7aYpTIZI495nOPYTOS9dzkqQqfVJLdPaPALujQvztiM3CxIzbYJ
N+tKUGyM0U07t2EpF7qO7aPOTNxoZzwassZPa5aqY6K4bYnRf4E2HeTeCCZ2+G3Y
16UPBe6FwUyW2vgBfyn3cTCinRM70911KwjqnS7jZUj61ss9cDsvsUyQM6YFgPAq
h+fleaWAnaqtN/iH8wB+R4Xh7OiXsuI47UUvC8vxMUGEKMkqowhIvYcX7nswCuCo
Gb4Iz3MLxqw8dGKq0A53bF5M3CIkqnmges4Vu0Aj9WCF4mZmK8FI3sP5C20l9lXU
J2qiH06HJxwejZZFcvfoadORJ81c2m/ypEqYF+fhmk17t25Lb9mjYGcwDIZNXscM
6Kkdfv8b5P9oB1yIE7mXK/0OmnqW5flnLlsqIvx3uVtn1DLbYeI40walsEi/3y/i
d5tMzRN70bVejFMCRz718jmAPb1tvLv/MiPFs3D9zj4XyAgCI0AZ139UuRr0VruA
Br2Q2Ktf7n7QHt6uoPOZoozw9UYMWQOS5KuchgIDf28oRh26ab3+zhtqIk3Wr366
WmfWNfeR/TbVMgb5/ny+hTOitMudAxeYfOxwl4mX5XnTaftUj5WewTq+V6mKOEcj
OT2K8ifiB7OD9diriQpj04JjwN9l64m8MFPSVEFdVE4RF4+Y/VVP92p9h121kO9N
/arY/J8Xa3/e2uL6vBcRRgFUH6Cj18vQEos+2TgZ6YdFUQy3gllxR1/xZsO9Bc7k
B7POS28bJF7HxhlRhbVMlaBHm4WjF813xGfAPMUaxexiRqrS/1lXmReDt7t9wZvy
V0f/OvZzZQVdK6YEGK5ftpz1UKARabbs/QlrsLRpXAH4/r1G1DYbkWpS+W+uLUIC
5pcETFJJ7f9rvcFqZsS+Tgr6Hxj7eY0WE7I/J+nTfAgpzcTXImBRYdK3Jj0hnEQI
RzB6ZsLJh6XKfSvP8agNQwWh4zGG46yGVnY37QFtQ86vFJHhJFeCezYB7vbRyyHs
CB7Kb2rKHbHYx3OjXi0Hs8+laDspUYwhB31F0notr9P95dYzPU5E3vlPWoIbhVQ2
PhCbgZeQ+essNf+QqRlYwoVxSwt6jp6MCrHR9WWi6RrrZvBJikDUZ6kNbrtfH4hM
DbeVKj9rTsnN5CoFtkdRooOsqtZUf0y8TkrTzYziAl5wbocYKv+eTA9cjmrZ25Ty
m+zLkn87ozEmAncslTlwNpw3Rt84zxnDTyxy5k417W8fBuuzX3TS073wwSZ+yItY
0DiB3fJXHJvF3NONVZDS05ARRFvvTjWBNPRwx6Tgc1IQEUInRWwA+Yh9dWVjcQIY
/FtlsKt+PUkOP9JTkWeAIKUakI67T+VPERtfYaJNg97gGX8gzgjk6dLhi54HeZx2
x8+xRRtfN1jl6o9uMlyY5ija+iKrZ0xHzBN3FsRc+Qcp2Vv4DoCQDaVxjG52dpp4
LREHsc4qddSRu/1dWdowCIYbbpK1yrkKdH6a2u8Jy4pF6MntxoONVdRkWcBzkThg
95EESj8ggaiwNNhXbQW6Px/ijS5wpY1WhFabaVut8bjAU0T7xWIOSfKs2N/x6ty9
pTJY53azkyuU/rkPtI3e0Px+ZYcUyxHme3mPsw6JgqnRp4FtTqZ7BRqdN9KdxBGk
C6Qy1tqMr/p5KwKZ/vZFIPdTmcsIvAnd//tqGeHwymwJGmmqIWF4NGYWabVRFbqx
Gdcr8ti7OS/8c2fbOyaxTx/hpMBfT/h/qhfrJn1zU34lIpRDM1R4J8ekInFR/6cw
r/x3bVCmttP/ljPdpohMXitOXaIgBdStXsS7wmMvh25HHJopnaHNP2r+5wF9FBCz
hsy4ilFBEhcUbKdCQ3w2eLGWLCWoED4Psz3MVxU+/IV2U2aeflkTh4o9aI7QwIFu
HruOg7ba54x5ownWfW4gH0rRblHfzPlF6pm6oO3psvUyKeOcSpzftAaZa5cgTTzZ
z+kOSX5LCW6S+7z7fZYLtl+l261VndLLKnrvoE2f7FkZRSrp6gApokQWjsHz6L5d
tnqJ0Is6sP5GtgTHmhM3HppSUpfOrkvBben8/YD+yOCZK9Lo9Zl2wpklvMm0/D+S
QvtaAbRGzKPu2nsqLGkoH61D1CzjWRUC6m7FAuGhrV6Cl7RUS2uhMb2EbFac1Vzn
NVeeI8jRek6gw7hztEwwbd1IPZ+EwTkCPevTlfOn2uXp5uXIAPHGCA1yApv2yw4Y
NF22RKfZEqoxhGIcyg+BGJwaq/4MPuvFDqiUjeFXogRMxI/osAQ8Tf8BFiRR+aP+
IKo735f4kOaQAVMwZkjaBZbehO6sQeCr9FH/66kZLW/5tG6rJRkcoJ//tdzYM1HD
pYurHKsD1oaGhhEZeurf+5T5O6yf53wBKZqB7jc0/W5wMBo1CeWlXrkHsG8Zoakq
0iG9IrIHd4Ukq44sFuAvlMFk3VzpwWgnpxOM1OskGqMuEg9HEFMZ89R1jrr8yiEE
qMsjhoN5eVnRN0PJG01EMpVrreKute8/WM2080HoKCYXC9TmPS3r3dzMLkiNvAcv
ob7sXtk/4YYz10AFYF7AxZJQ2vx2AEL31AcfjhirKZ90eBllqzzUD+OMLYa05qSg
xkEdfr8M6TKkivCAPArPUe68UayHYZIKpUG6WGkbz23rz500FfXicvbAtOu3AtGd
OmXbm6B+xMPC5Yu0Zsj3OLP8kmGETZNvtysqsMmZgn1uZ9ZgYrKdOTyghllKTZcE
GMt4tYWuUMeC7BQNmTcO6NIdDBVRSdM4R1r4ndjVavZEKXR3itd7qz0aZI628l5R
Qowzs3VGnsDdIns0fFWoPjp2yDsdDK/CspY+BuY3Bcc4Wsl20/EGNyImHGSLs9hg
Q1uu25P2EjFsGzdishYnas9S+l4yMoREUcApC1zUp13wdbPEWSPWwTKr3CrYrjE7
jF2FmDAb06G+hp2pTvjikpAZB2WFuNSWXT4jEiWuUvBk4+9Qj0MhFezJvd68Rnkr
mNFOp2pJDA7fIvhsypwQWv+vi3A8lu+2QjtnKB9TXXE+Hi/uGIq1nfX66KSjhPW0
QmgE5xyLF0HZY/eCrGaRkE31bED1thQIlCEv+l+GPSJTgA3DAPs/o+6YEv9F+hou
VE9lrt6s/l8Osqhw0crloG6N1COLRSX3PxLDEeVXQtg8hDQDBCAC6OStV47cqfnc
O6nR8V0WBIEFWat/jhMXHrj2HiwN/VfFT6I9kXXjbfgxi4zX7mnKBnVHXJBoB7Yc
lhpyUd8FnEIcQDdEuQGEvDC1slxSf+QuBENQyxgVbuOzVZEQfSV65JYJtNQoKPsy
AqdkDKU/83ILMBk0m2JZZBjQAd1BzbctdccdEYmB7jzpyWV8C+FD82hVdXwsr260
EnBzDJEkXj6Irdx/v47XRodW8NcylDYqulb1NGumEclxk/fCs1b30LFgQgglKY8e
9Rqi/F218w31JV+DzZl25tItTKdP7afAr++yXwr+mv0cNFeRgx68gSmYGjpKZ30X
12waEoRveFktYnH+6jUq6rQtclgh9o00T7zfLCwXGXTA8/YjJBL1kqPs9zIXkPN6
+tqmuB2SqAo0U7fTxZ0S4yK9HHLn3xP6Y/a+pscCeX7ZsfLVU7mtdf5l4A4TlVZY
o5YNDwJwFM49pBst5Uwz/eDA3/caNOunwdSaCCiFh/fBZJG8afciBOib/owemn4G
DsXccRAXvOIhwmXtUc9kwnKefljowgDokAJ8XsL2kJ+xdFek6cm6KPAInOqayDt0
oHuYJNjrwvxX+EOWu45UZX3CQozfUgXlMsluoQBqmqYxPFNADottcMrHI5S7FArP
a/POcHAnFIwNF1/aXrkRs4gNnGk+t/YMEXPUu/TkThWDbXJttZOlhn/74OqwKZFd
2svJkBkELslViT48y2hiHDUn2cqM9+xWrDrVDTBYOBM/1/0vdCF3wfq5kdcagEyN
Wt8fz1KQnP1UERypyFmd3InVQHITY5CBuCrOVlnaqXUjoroFvryI7CzVEMZs3YfV
9I5QdaHu/O9R1olA9RWYCfpsTDNBjuBih8iSBceljWXL04V/2YYu3JuxmljDMnCf
/w7uqxHn1Y5UYz320WJwiJ2OUsa2Fj/ykPTLzXhtBwt1WsxoJ8Ixr+3Jtq5w7VTT
vWkKL1zKZwQccMeq04Og/HEFByV45KfD3uPpSgy2+k6BSbsQ0vmjOZptcMQcNf4H
0OFzonVbI0jHaGHnGIci49ckZHmVNiuvPuJuey7Q/2NG/pHKZEvlbUPNDXtF5ast
qeI/YGGRp1GtbhGnLWZVvhJYXtpKGgfFn2r6HgJRNkIx1RKQBU2MWQ4MnauzOFIe
PwBO9hTT8MydpROWYvGEQ4bqF0aOYEDDuOJbP1SARbXV1SN7R/ieERMhhZxGOT1t
DBAipLzXEs/reUuTc5bjcWLW/lalnCPzHgktwhRPSYjZDl7j/cDuMj01qkKgcYF/
aRWrYkksDS7OSIz5JZLSlwSzt74IlGLit5GUPEaAt0O2gKkvIWzTT2yVJl92vxPf
89wu/Ic5PiYKOmMII8Hs8r+F1TCmeNorFeJ6181i5uMnjjHayKbWntPpKSlAIaFc
dOaSzqSNu1yl2/aYGl4snmhDsSYcTgUPJaUpv8O4lYwrei2TB20yZBhUktnI8vX7
QsV1jDcmOCftTOS0adSqwOxYx2Nl39K1I/00QQGEFz3yQ8ju9eh3LnbSsh0iXz3P
P17QyglqiAX4WL4jvoWQyHrLhZ3gAPH8ZjcJ+PLb2N/Tul2Kg9vp1AhWyonxbjIH
6/g0tvMLDZQytGJcWIzud6QjUODI8bskG5PRWuPtCL7yQtnqcIgPSdD8pXK96pOM
9927ar44YRB2JZe66kZZjLHke4CBWhlELy3LHL0mINuC4zMPGjyzejIYAvx/eG66
USR0SrnNA+tKOpqALeFLtl20kGnYJjNWk/MxA2Se+YMqRK3WnAVvDVqW0jaxPple
peXDLR8mTAReMBWyD4poV0IgbQG3NV1nHftQXVqqease9J2baKeltRluRiIH4dcs
T1RbTMCjcihL7Va2X7p4QsllnUAb+7Cfj5slrCYcn0UwUZ9m42DYE4zdKzTj0LFL
9ax8OkM3dHe7AdN/IY9A7TZlkwYbtI/G5zAjOdEMGngN8ymqGb6J1t8hO5BGKpP1
2wQcMJxy04TpMxTpIKypyGRI2N5AQxu/UjRcg4koQJpjy2tb0BiWBTHgrc5/UT4Y
/tdMA1GSr+E03GMvTeyXDvWY3s4VtNf3NfuhLT3H4jc3BVSFZkfE2FYNqg1P1F28
ZTMhr9SLG/pNaVkF6fm14DmQpcm9FiacKo7In877ke0xSJN41sllrXM7W9t8B4VG
sfW+CZUgUdmwrlH3TOADCioDWlKPHG8wmaNxbR3K3aerWfclzn4naqUQezsgFc81
C6kOjgoIU4m1XFSlVtJCL+AUt4lqvswo5ywuftCHbYgWTCBX0w8EM98pfFpDrBMy
oNedOpx4XxJQchfaFrhMkqvkpE+i6bKyoF0nxS6WRNREWGGkLGB9uKgSEHR0LujN
t9z5aeiHYd1A7i6x53rl+RaHKiOcFTJGrc/rQCWngGA6CRhtVx8wTXF3rO66P8D8
RYcP9a4xHmKHYM1CWpQI4es3LANwfLEktlCgxuKDd8b2IcX26ExUqovqZgA99CkG
K92JWQm+FhqFR3ltNbmj5N/27SPXmWzKHMN5pfZBA9oyqn6fRP2hr1Z7qeoYXT/X
QxxyAmUTVGG0sKMIfRLJT7z8JVYLY3WQ4kv7BcWeoXXva68rcg7FnZORxQ4778Rp
1kz85XsFPKPoscPYw1hNKzIH2y82uzyg77mhM+oNOrsGr/9nrzSIegA6+LwC21ei
6Gan/SHqeUHwhIR8H09iOyn27CQkHOO1aoDNd5oSohVuI4pp7N3/8V0HZ/owle4Z
a74lpcSunQIDeV1ZG6UBR1rRZZ0+UNtnc0/Mi1h1EA4naWqtZ8k4i1eIT1kopkEt
IOQbnH/xxuWNwiZB89dyHB0KmWk8jRvMzZEwyXKAIE/6TcsziMJFnchf+lgyBZdo
ALPD+dfCHyoEL3+apIxbs+t2NoWIUFBrItuZD4Q6vDe1lWv8Z9Sa5e8sRzFOg1sc
HYeqGCmzSdLwu/mkL4H/MisVjx0YCCUK+BXzGI3MvkrclKJfUrEOm5pugJkjB5iy
TCnr2DFuTKBJqPSAQn7Wb8KavNN9gXjkCqzrrDu9qGSGNRFCS4QyTRsfzJjRMqjG
9tYxn0cm2lyQ8DGQdLG+dpx/8BrDHzTyCKRSxpGt9/HKScNi2i1vCmojAeC3l1d3
cXg6ao5zkhUM8shL0rYHFC8xv7lETBHYHRJuVsqs5C1lf5OMJES6QkupM398oz+i
clpwmOLa1xLRV4OmunpR87BbiM0uHN6u7BU7Ca4y9Cyv1DwSfPh/WQ3tXwqeodri
IRHWt7P0U3TeXjyaOiQLvTH5GpAl5vCdI8y/PJmxJ0PnDLjrg8VLDi6TA5jqaNo0
6ArR7gOkuou3PO0X92npL8gle/sSLrbtROsn9So4EaMYD5XjtIbNrucgarsHlGfv
aEmfjvGXVttHcYCYuApxFUXy6NrxcUMLySEqdqlj+19+SC3Bs1NqO2UyKq7zoWfL
CZwta/HnKrWRie5h+UemhePt0knVNCzQIbNcf5XhOxCVUkRMiIDTdErzeqFOESyh
FxM6csABxfEAk5uuPzBfic7NaxffeU0u0Ucs1UVyvhz4QGt2aXKhIxWy6Cluq++u
syu34Ru/CsFlcVJtPFvIcFDgXD9PzBzNLrB0nqnoAFBYYMgRtpNAK/cicfuZbRjz
FHYDBFLknHi8HmxOAFpiqg53Em32drqaCoY+X0ZD6ooauFSxkVP62BSexYxihczI
RnhQ7vlIuAXVGzTOBhcNI/1TwWL6SAdeh2vnE+E6mtpdg0I9My5cuuBUeavgCu4s
yYbR7ZAWiOUctW59v19ib/ScEpS91tjli4IWvu19rVQHziN5KkSfJmAGEvSdCU4R
1j9bij5NvrxGyDn0CUxVDhSSGKIQFLxNdIOdaSxkeQsrPRvK3xX3W4N9UAU+RXbC
Fyi+gtvWFbXYYFfyB2I+lLMHs9qnCiVIF5Zh0KoeirJVVNMR3sIKgVjqbwwPDPCs
ZtdCYCZSKAeZlT1zBfRI2XUuCbhBkaGFOna7HubNpDM6azMLuaV1C4k75CYiX/nP
9CT8vjcMyfpgl87pF4jy5ykBM43IAdah0aulEeyStXBleP+f/gMVZckQ27RoT1Or
VEszk86b1OuIWJYHEAihQ9fB00z7viK/EfC+LbjiSL0JYN+YGQEJHI1aza9rPG32
oqSmrtwo8s/tWelXljfgoObae9QO77qUqftpvoNcbuUzzNcSlBcuS+5cn3bapbDo
1YR9QUgLNGV0e9Nd67haHiiUNbHp4eIjCbzoYX+r8AbaKNvFD7E9Wnd9py6e74/I
f5bXdp3rGvI7zA5BVb1evl4cDCy9K/0cBLjyJDhgTZx0HESrNJD8KxWzQIIqOA/C
JStyXLkXpV4hkCOPLHF3WCzUWRLnxoxvioPAeS0GRnInzEv1ovkFUBkR6vWZviLY
LNuGN9QAlaeMjROBcPARO9zvaBwoWFtr8/XeXqLejEtmJpIwTX4HhQg7NteqehQ8
5JWJXpq/kCIbgkXOtLl8qjCc3ST+SJM3WxzbT4edRlR9hH4OdL8A0xjfaTtguoj0
+y4eudccNu/4RVkBm8xkCH9iS1ihbp1Yw58IMu0SIW6dDC8jzKk1SF95iJ4tleCp
q4PyiZGnO8liRtCFV6GTDYf4nlIlSkxb6I33bkocxIV4URLE8X1IH76VaGQy/+yE
9Ih75cXxkXEqplf5/KLGIpV4RccSSVavw6Gj8DticapJtjLBc/OnxXuYwN7Tl9/q
V+pykb03sVh9LPFEOz9VtBxWIgN+2A7Rglc83AkTvZmS/jZpzmgLKsdTcmKAsj16
qHsohNBE/tBLVXnvPGsvbReb3fG2pIiTIMThdcritc1hU5PAqUfcrKv1oLo6Ltgl
PTUZ+3XMQBWhGy8KG23Ztb2i87o3rV9ph5Ge7Z1FgN9jNw1gvMYls8+WuIDvJ6kV
GnkbypehsQbjJBiao/5oW/xpehLTCRDkMH/2Ph41LMdIO2uGkhQNXmZf+qoQX9/b
Jc0zw184rrfO5UJIoD4A5ZKUGFwWTGiwPX/XTW6txxVgYg35uBG97xXHAKA3C6XE
M2xG9DRLkHSX9SdZerpb5533fcxfKRbM0jg32aSZw3Y1gjZn0pFpRXAg0Dm5Yrsw
/uxkSbaD9Cr9CsaJQZ0ThXnqS5SClCbRr8FCcxaPCzYlT9Uh1TlLIHvG7CtXyQJc
vn2vBitFi7XOCYZSYKVyZUlt7H2RWB4xGWuZcBfrN3WYIiSpptByAv2fBXsJYkPd
vEk/MeBS9Csv/nI+myhFgulg9NY529yn4TRPDxfYtd05/G61OmXPYUr406iOmY5v
446pD0XtzjDucVGyurKkt42tPNA/bda8/Arrz5ZRy5rhNsj5Kvn8p625uGemioQF
MhdBjrcxhWyC9EH6iuGm6SDsYYVwf6HJfRuAyjqhDkVTHwOPEk4XTKUbSC4PqR/N
Ru6ov2j9hHcm1V/aU5G7ysnDInsT77lQv9gcYrZCF/zx1qFjVDO7jCHuKq7jgCoq
RDvjguw8Xxtc+3LHSjSrLR9BBPa+064tWotOT08kZAmkUO0E9hdSOaBka2oHQyFR
7w2sroMffWwXrvwJ+PaeiPJpMrUo6cFFF+siHHhdHPM/yvpVXY3oTL4Lsb+xs4Qx
GCiYTlHQ3hXBRiu/4Losjej8ZvjfDn5kGsv71Vh/wOQqQ+j17YeREHr6rSPu8sKc
c0MiJ3L88X4w5L9v2tCXTOeeAh0PuenB0QKE3tbTmr/99L66DHpIDhonAaAf8NLy
0idyGasJmHy2ZWCgooQDhI82ZMuV6SGHF0sxUAvMcUuARgFYTNbt/5wWd+tMbvaa
KDlKzWNFU0ZPvYPPv7cfUwQDS4+zjZ+9i4B6izAlZSCjSK/1I/F0Do7ykG7h8G9a
BZdj1bXqlP2PpQ70F6xw9c9frwiC9XgCt2cnu+NXksHpbB6gzW1CpwH+MrdXA2hP
zbR7vhdwMxxgbKLmHGRsb/fVEsAtYiRp72uvLH+lXr8V71k5lFX00R/dVJJM6y9U
aPOfzgKdStJAsxjNyzdV8R5Cykic8hWFcakK7vtTpxW66f45xkpH7PicJbYQnN8Y
/opZeKXQulfVJrtAtEcgL+h6WaNRjcjNr/xsfzs4ubJRHTFsbC3qtZKpMvyIFZl+
bO2/sJ4nOuHvAmeMPPY9havTbwH1FnU9mMI+kKEZFLHDN+TciyMeDs65z9Zo58Hm
nakwQ817ViN9JImRZv+FiF8NiXUhInmQ1hPY04pmkAkwcnIujmOX9csSGIuHrGMn
CdEt5UwA84UFu3J6PMQtsOa8E4lywS3TCHBQpSucfjCl6jXOudgiHWgSvISicIMR
Nd1VgFXg7LdJafhOCACnaaeIUmJwLvbUoSXmZx2KCsTjBmV8BblG64Se3JLb2RBJ
8Pto4Aoru+5TT93LuyfdT14bQ9Bg4rYuXX4QuG9Y41gVyObF09gw78frhNbp8uDn
hwc9s4SgRrfEUFyk3vS3/KWUYaj003pb2hSpupTOuqvfpQwlpnZ/CdIlB93D6Akw
q1NDWMUp00MUvkaRJMKQkoncq4pXjBaRn1INXSBk7hgk1xA15wl8GaHWGyEIuq8K
b7KZy5rA4cCJJOi9cXvEKOhHfh+1Mv/4lqQktb2OIwyRgimPuycRxnW/9xPmyJFt
ahjMkyr3JglCJaDy3B30bOaJahMDxaXJuGvXOMWP1t7jA5e1/ebacEJKNUx+s5pX
NfuVhtZZFPJa5Uw+PfIA3i+Gg1k8Gm6Fj+sKNm11K7gkgJ87G+YQ/ihGIumCIMZ+
bQxACHmRX3uU+Cu031eWc0o2AKdHwPAYUkfh02apWeu4QiS8L3liishCpcujV3iQ
T+ACgAYiYck2YTSlTwt0sCoTVJ1iohzKyI69b2e+myOD/XWHlESoPmAQqiNYBQpV
tqSDY6EwzoMA6MY/KmOzAotTOjfK6sFgDPbd+bE4NLTlM8unVXmuy/nf6uviDd8x
yzAZPGfzrURNEBuFKILzH9tf+O/VHO+baoPGAwKQIOnZtzWlO9Fdg4I4fAS8I6d7
5tjPtOUBrTaD6Bi9NyvCCENbIvuBwtxZV1zKaJ0nGdj6kTZzxc/Z+RjdaCmS6J9w
vamZQ51Gq0Y8aGQ9zNRaRFbsW3AzBOIMNgBWYAp5yb+CDJ9ShlG8AkA/vkMJcxXu
zSD9meLLg1LvrkGizQ+zf7zzIjdmjQl1Tnr42/q8IEFXelBpxkYMkbLbbV66vNH9
m5ZSvyt1qr2bBTFPUWvrU9QRfvsBZqZX27tdc3b00VnG6T2kls/b7m9ao7tGpnj8
0/L4rqlEBRr7IxM51eDeS+w2n+TocFH5u/wDu9wM/67CU/7YI5qgSchm+K71SXpj
WgUdOWXg7lljkQZweYkY9omQVZDjZIfd50W9zmPb3yYt2ASi6rJo1LRgepwNkl4a
SV2o65AisF+UCmAq3E4dnRrlMCw56k/y1ybpb20NEY0/7zFX7ATcYJMzVYMFecIY
egs3oVBX11DwD4Y/nKMjocIg4/Sm8cK2iLkPz8Kh2UsLPZUmupoqOMCNbzg21h8Z
TY/O6CmALU3K9zvAMhqyY2xhovoy0fFmX638unpmmh3Y1nDYNmfyrhka3Mw6zDSX
mQms9N2IGuIhZH70cenFPmwa4y2VzG57Ud0/q8zEajgjj24xedjQiPEt0DvXDwRt
fIWkhaIIJULtPsQi2BaBRruC49/jGriB0cIojTzlbrLK4SCPslNAxrqwjoFi6x4l
Wx8EgihGKZsc6dzg9pMDTilhHTb4tTOzqO/EVbPynNbt5EIemf4e368cOewa1y/Y
0qQZwtwZAWype9+/Vumy75DPr+vCs+Uz15cKv1X6pNkO+g/wnbTw84yuNFRYv/DG
RR10sBmMrBYXPvwjKA37D8g0vPX1pc9FjUygQyDNhBQXymgFmW1BSxJdou/qO3pZ
wbiP+5ElBe27YIdb3xG++cuQCoQnolYlzrweH8cG4gkcmLQmmovpRbemQR7dP0Mv
d4RceFgxv+UWifBimwNnYDb+E0/3mfaS+L/VmPwYQFhkV3ejSp1l73ZAQ38XUWvN
sHOoak7g4rg/RF+vx2rwtYxszCadeABO3V5qLsT5tcPEJnOxVToXhT5nH79jB+Yw
fTThpb6pzXqqzl1lg7+czlN35H1bGxBIbA6hcWPSW3pYER+6CDCtzs9uCFcLKlOC
ZOHoreSpwnPDdH7IofmNYqnwdNDuirUWDynrdkpfLuzrXJ7UifiQ3OZV0vB0zEd5
nLNuVDGBy6M+/4SoUoCiXzigwOqBG/klZLadmIjh1EFrZXB1aL0aXOfgxoXeg487
b5Br2u1acuGfq8d2GTq1JAnp0QNrCihuKVPk7Y1u3FjvUuWPLnjK3Z5x9zL4qGmy
dHa8MlGopcuU7nFtVsAuBVP91rBxVnRP7MOJmpavsuXBcbUbNS1SgVTJCGCpRj2S
CgX9SXNff+hDZ+3A07pJaxreLRrF/Oi1EPpxLzsuDZKg8LC3POHgMQxN+ytsBCyy
IF7ugDtQGfy0BKsvBz+PdjgOElS65c6/yZ04Mgc6keW9rGXB1ixgrRnsCOgvGb2L
mk3S+/bXj4iZcCEgrzc2b9VRGrAUBXJAO3ybVCKhQW37oN0X21PdKm/P5azObOok
rDwJ9/Gk3Z/EJWCJsi6BqWZX/BR3Ve7MRnMAGbJu6sSp3l5oL0n2gg6rGpCHizwo
Km8SB5GvsgQy8OfKBgsnTEIbqPiqKCTA5injkQR3JoAhsLzAHT8ZlwvyPOmtj42H
X3JGmzBlgmpA5bSH7mUqT2bWDrTHJcXiS4so35lMhFastV1EW3WmDHHICeIX5kkd
zl++UnZjmEpUqgaqxEcdzWCTkzgV3wnDsrAKci1Etw8ADJho7N0iqZwVeYkxsork
XMe2TVzkApvl0dbAM3otCRRJ4MILVZ6G+bV0nWKzsxk7MCpGgN2IKCLW7qs4ZGct
jH0bUTi9uLNQwELnjCIuLvmT7cP7M7q6eJhkCwd/6RPbRp6nS8+KJ0vYgb+XP7C6
puabQB+aECyk6YYwKjurARdPwryyUZEnNMK3TcpYY9ZgknhrEOtqZi6Mt4gZi042
Njn1Gqzd1Gj//00tZaFOA6HjsyWkMVL711hLec77IoHEBenhAbfSgBTew2Z76sNE
ieAS/17fbeSawDoNhfV3U7IChPfyS2MWm4iod4QyczTzy8d8FY4af0P66pzbUJGL
awTnpsDA59sZo2HgaLNMu4ynusj9x+4PQ5XDMUhW7ZMsWVF+UVG0oiq0Rpqyw1RL
QMWn4sh5BUARmRqJHUEekmuHs35p/3kBaUeeP7gpwD8uvyQK6d84TzQtOxZGHLx0
9A8nSRssr0GJhv69XoNKigO7mNffPCKm7HVqcbPfi6hTTeoU61VG/OTlzwKQBRZg
rmMIoRt4a3EbTS0ljPAyXrstE6lDNQPAhTX2iw2TiEpyJGUiSCYwI07gq49HL8n/
xznzrXK4sDHNM0zkjkO7/8y7fKd0xA++pvpp9FQaeB4EUhHngEPH36+OIF+FuHV5
pCLjGlgWi0+GPgal8r1/TpS4FVb/K3EPMq/54mG9SNKnrNWfGtEyCehw9/RHYlF5
V25hLq2uwjhyJlJ4U8ksrXIXd84PEwXaqcYIRXmk8tawAjMlU85uIc68prpqBCxQ
JPkm+zS2JE1pcj3IYeDASLXT8NfL50I1WuUml2pfw6v68daIvw1jGiFcmk4hBYY5
FMA5MFuR1xMh32i/JweTN2b4ZExpltasi6vCDGa8O+XVngLzmyUzVppS0BD65dUR
bYEkj8B/V7oYA6zfNARO6vxejDIMymrwxzJVk5iWJwrhhL0Z8UIJmN2EXdZQFEnJ
JykX69Vt6ZzsqHpKVagkLDRw/OLeCb+rGI0FrojHNBCqvFbnQuHCExDG3RBG3cNV
/1dzy1hVGYyMgfekUUQ16md1g0CRbQO4L7qfjNYTjFkNpEPyLIiijHMNntimG1MM
3X7HeiKoqS+OdL714RJHWr9f1wBiUbPMkIvCjh7GDUnY2eYuT5WWsvwNLIbTdaiT
h3g8nKZWoPu+ZiC2y2cuQDLk9qF6OkyjU6DscGkRmPflo8ZgQonpwyaNtPiNhYQj
s/lz7/k6M1oD/caayit9tC+Q+02DFLLC8haQY9Exjx3JhKiolS8g36iUJpfr7CSF
1Z9PYg+UcACGVId7m3oOZxsEW0mzrixp229Bcu1Sn2JImoXiCHE/NfGpJiBtiL4F
PDexPpXj+0RmBPhEKOZ3sGZGZMiKJ58iDV/ayVeX489lzDOOcvEHr3Cilh6hEH1p
jRJdbJLT3gAAUdnRI7g0BQZI3vS2J9YM55LDdLdBpg+BCjb0ufSt0pE0aWGQMriz
5WL107jLhNAzi1QP7MifSCn6LNOmthPWw6fYQ8M64Bz8WdmgIBCGKC/5yADHvYMo
DS/XWLiWLQcRUQYr3J/4StPRl/TeIigSZMBHHJ9b/UGTvX1X6F2wE1SSslUfs84t
vz7tUK2QzBA45f6t8KKeELt5XzbKXZdiV7/kNd4W8NdC+J5oVnDXAoaRcjOt+AXT
WQD5nUt01tI27jGBgxBHlph1yasFtep8YhO0jo8F34vadzC0Lyw8LBASCcskYzM1
/KFK88rPNv9QZa1UqY6SBhN3TbH/wzu3iFREnQspWOfhhoY8gLIowc3BnElOPWUk
FxYU6aMVbDxzrINF2xHczbdoipb8TYj9tCmCwpUDm2hDWApOoxkXAcfKjrq0ly3H
Yq/QPSFRQmqPPh4gTo6Ub6DMj7ROBUFpZeIwyaZU5eOMnalxmidSWLHSNjbDpkMt
WcjJCgCdqBLAmJ/PE89om+zryi6eNxAmIXAwc1W/Zt1rEpgBJvOr/+1omSXYIoTy
FJFGmPv7j1ePJnI3mq5OFkb4agwWy/RbqRXttTy9bnZ2oXzGsGeK2Mf00kJ9WHxv
JQbvuGAWYrgzX744F3aLc2WBvZnHJAQEqLn456TdWuWw/1cozCPks5xPh8LCKYyw
dLogJx/DujDPSesaTHxsm6KAE6/+z8gaY8p0xy7DtgnwsV/FaAfbA2NYN4x12dq3
HY+L8tSf1iaIHWMf0MUUWu6NJpF2ESLK02nqb9/4XYqgj2TAgRNbfEH7Vzvtj4MH
4WJF9JYIVJqWOYmKLh+PIskO7f1y7F+N4ps6f7BofM2jBPNXbWgmc3wO1krZLORx
AItPRFx9fmOPsmJch4uxqSIdOi5o8HD9QRTSmmyxWXnWAQXlJYL7xg/u9q9NyTgw
KennXNWazK4glnFG6sUoyIKbTk+xJVL3pE+Uy4u8NLw7aa+eHaHJDQsT2zoATem0
b/8iOASqzWDeu9sj8BoFI5TGYJy93OkNHJrZPzczetriCv0LhP/dJyVKc7DxYr8c
m1CRLz1NsEkj+db9/6XDwUePu0EERg9SZHXUsMGLr7eDbYP67k7AUKvvSJ/sZz3E
8y6EgOA1DKdXopRQ1JiWMJP3TkpqfnrCyCJ5Sgup+IAfdCj6vMFvjVRyNACK97AC
prV1tNoQx5RMVm6O5GIoDeosAAEOYv39ynHvSmZtAES5SRxyV37ZwGpvD9o51BqZ
5pGdhlcm9enDPYbhHgWDqHMRBBq7GlL5wm64ieV7orLzChoG3RkK8pajE3rYM6si
7KWOAxFesxocTT+R5nAZGFTsXqCPsdd1ZEutDxoXsdOiGxUJS+Ipa53GFSOAc19J
oOQvNjNblU9xzPjwuv3PcvJyBVRUOwOQ9Pv/6CF9jy/M71s68BUl6uKeEPjHMoXT
FcrDiFN1UWqDk+kivAVR+5BCOmmmtLyv2OWhv2VBxtwy5yDx9cwJe14S5z1Uvap2
p64nlr5nNKr0vJhloTR/y/4C5kDyZkCiJTLyvz17HHwwxxfPVTml2Ww62HHnPA6v
eQeiFTBXN2E6NbZyfxRiVYw4UUb8YICtyN9kzi20QiuuMVh9vn2qOaXuJnYNkeZB
IfqvEtEHs8xxrM3mzqEgjzTx6Ucrd4PhPbMpX5hA+dKYnnWpPgUgTF9Qg7MVW388
SSXzbzBkLVALbqJllByTIVhsUjT90m8EmoYESy36bmzEG6PcbjUHDB0Z/sKkbaNk
cbzZoA34XDAPXfIQ8yceLET4JNIrnT9vTvdumaXlNG/veN6R1afh14WgWFW04W6x
ko/CGUkLccfU40YULP1Mb3uKKaI0cU5G8DqmfqwOC8KrfVHz9rBdzupUpYSsVQpR
Fhmig81SLFjD/n88BiTkVP8+EVrqLWPYdH7aFHTBT8nF0VQ7DN38BA+VNxCoQzbY
zS2RRCzHflwYdQZriPnHPdRm4ZcAZgIbURryCbNIURmgajnWB1PmcKOdOxvR6cz0
D9QP68y9jdJd7bQ8f0PICj0Mte2+kx9N9GFHPOGNFnMHGkR1EBu8Ceba70yX2w+b
pma/8NvAFlP4fCmISinaEnn69MBdYr9Pcx9lSoipxZX+3LxLfNx6k9F/7dogjEJ3
EBWzdEq3+yj2RuasBtZvDfKizxtmE3tHJN/Uz+owA6uvie1s+t22zTiSd9arStpr
CSIZ0oGz1oVBqVUFBLAdrtwJWRl/zXnEon9bQ0r2LJ+0J+o2fA6cdg66YBw+r/NE
moUrB2K97hP8puDNpafo7iIqQMRtN2r71qDawX+HTNznsFsaUAxeVrjrwUFAuBZB
sQM+UVxSt302xZIPVjRi5Bqe6qVr7ZGvrgBpmsJS4ZssyxQC99KuhBMl9NMnPWcv
2P0ZWhdPcx33MfD8fK4sm8eGN9R8PsjIOlI6PrlJHpRRWQ+3vr7yMQNRE+lQEgiL
XX0WjJqeemNfCzD234jtOZxeiBOI4UiFY0md1P4mI0zzHDixolbbwdlLssgvjriV
YPVDq80gkZIvfjD8/6grrxwosUT9+AJcn96q2qf77yC5yjI8h3ZeJM2zXjyJvBxA
IGuaJZjXaY4TlcvlxkFJpzG0V7fWrpsINewN9zU8eRUp3z2yR6eG/z/leXo9D0fn
rGKnz1c7dmG+4jKBCeZACDFTqcqbRmSbDIoZOYqCpKV6eFE/65F+VlM9eNmAgBXY
apa7zodxz04c9ryBBfOctcYiYXOri4dI2POTsM3uesZa0JDyl4R+URATRoHmC/Eb
exCor8kLpOZkKgvfQZBpub91Q/WJwc8ml2dZjai15EHFMcn3xb4MuZ0F+uUi7w0I
94ixSKYPJiMg5vi8i1UM+J769zfbEenJU8us+SiQuGrQAt4wT1TOmnzcZ1WJSCkX
LTa4p4rK8VQguvAQL0sTFCBkuMTT/tqdjypfu9+ISqT461yzFLqxqt+RafNncrf7
YTxT6BmxbFFWN1kxf65vRsCzQs8G/X1wrnB4MfGmfHRHq26o8tV9X+WX09yFDhxc
hz7yBZU8TXWbF3r4ol0VxQ16LOp5ftkxlnn47ZfcoKyX7rj8wwiFawUyH5cw7SSw
l6JwooO10doMfD/Tp5Ur33XIqLv+mDnS6R7Wcs1sx4mUiUx73TqkzZxa/x7R8RBo
TTCriTWnv+XYBFqGOyhPFNVh5BsjpBjLtK2vHxa4jHYittICehbq9ulq6u9IyDXh
gExvcpVpDeOpqnmxSf4MSr725wXWGfYasgntakDHHDTXxrGePdJlaVOQIOotOpHA
9ZNu42FrqtjI1TlROgHWJsQbgqB5UpcKCKzFnKNl5itfzIHQ0fDODwgdPiCYkcTq
dcCLAAhpcje8mCFGHo3MVHedwtrfX/NaBO/UhZKvx1QPNyOrd0kGFTlMJeU8qnKZ
bY2Hy32esQVwmXIr9j3zi8zgEFGrdZ4L6oEBNloGeIkVakSuxlk+3mq1jBev7aE9
JygWUYWGKfDdKskmNssIDpfNTVdscygQTy2pshKqs6S5Xnb8rj4Tmy68VAROq/my
3g4QZkwPcTZ4dnDAb8AoZKpzgNI8QjwbEGjGUWCZGRJiYnyzQxP3l/m1TSe2bxqv
/0K7oYyserb79II+vQTEjwYKY766TV0U5pVYju17reUsOWiNM1SORpvf1wc2eBVG
zl+EwyIiYTxoxs6djttj7Pc6n+asWcwJrZ5KiGO7lbgpHwvAA/BpITrWnKGL48+N
hMKuM+0BR6KwV6C3JYMZQl+SQMbcFPnLY+TMXjYY9EijR5gM9kncem2eEtgT/Re6
uj+yTXXwLQpbi/veWs8KS59txrlFKRrADHA3jRA4rtJGFd08ViyDQzfpd1EhYGwg
nJQ4nYO8ZSnJkGAkO0W6eLhQkLyE1xwssLU4CMrUqYs99WSYiZEZtSrbvRDrPCDk
VEhGMUw6iqSz6zF+1fw6VnTx1hTIDQwNjNAkKdw7Y1de6U4UO0mMfmLKv+fYVtxj
wpHwmfbutZzJBk3gQluAetYMPH7cIrCJkbg15o8MB7a4x1H563ltr1ed/JaxtrQ7
Bk8SDMBN86h1RBvfmwAQhojRkD8jQRC5KtwgOWZAuL7rDcN+uq7jK74CHsxEprho
3k997WbvdVaTItMpgWvfbHQS7QIVe3Bs/Zxfxra/joG/FHV9IXjQbkBuRmBF0rIj
WSmqp0VhLU7T0l4nBWooTKWbCYDZRro090ZKAYu7XZ1Dv3HKV6e4/Qribbte5Qsa
eI5ab9hJBgjW24XN0eCMGu53xBnyiuTLmcxLrOsJE75Ikivqyb60jlzYtKkeJq+1
0SECr/TM33ENNJXMU1yeQFOsBjFZ0IvNWhg3+bkTE6QvRBSBfx42TDzOAoubKwxJ
T2bTd3nEGRjHsi/sx7NidyZui0IN4XTs5TqG1OJBFTulz39FGawv1Y0YZv3JoK2P
16BitwnID49NZfjFZxMaUa3NHiUsf8j5QUBwS4C5/RxO06jJk5KVcGBvh00uYyPH
dnDgBqsHyg1u8A4pqMZ+sytliy5yZOXpzaDI+9xeplu5DWkdzyna2L200WxgXuZs
PBkTspqDWG6LaJaW9nE6Q1XcyfowFXNAu+ccERArjaPmYXTN6xEEU/Iqs6dtqp1z
3GzktlqcBfNkA04adTYSQogyXClGZR7xv/J0Dam3kBhCMsKndkjZRuMoIw//1Vv9
Tw7qzlTwmR/llwkFfdlk7W7zfxV8g6onMXsB9qKmzoYyL0d+gmA3RWlMaanL9P1F
91zy5cVPKHgjM2hHgAcB8j/tM3Tpa38IkmRyNz6FqCY5EhjbEdVa+0cEi1ZRf4R8
p+jbIUcIvSotd8ydC99NTWpoFVNhNZeU/YMQt10D0mKZbAqQ8ScGUpdzDg1n2pCA
iz8KNfLmI1Mj6qJ9iWhtoSgEonUWiSoBiiDxU1r3U9aCrnV7pQDAQeGjqxIQ3NJg
jcW+C6UZSONULIOxJ+hSCs/A0OKe8ouX5FozT7B/fmvL6cMQERWO7krDnzCQFepj
Km2eqm0LdzVWFhURQwfwsMC84cUEqjkl24B1h4yDeerblz5GHp1u2gcGYjj1MJj2
a0voDJbnr1kaj3FEKVLTxfZx4G3Y8CEyewpJQpmkpCYn19j/GhOatkgg/IXaFKD2
/W4aebQOdK9mWVy7sc5yln9IlDLMuvK3ifXDNHhd4soB8QPPacBJiNdbyNj2MCWy
M7WMINqmWsXlaD9K6R5SWUY0oIWZ2w6zLIYS7TlO6OiUuLxvmclk08irw306h6of
bSFArcdI1mxxKhDGmN7yO4OCM49xDSz4TN0V4yhARzuTDbbgl+hUscC9LZYIMCAL
lvVNKu/uLmsEDmeB4MiM2dnGVGELpHh3gyzEBL0RBEETcdYw4UnGmgrhJYHLbssz
EkKxUM272oEJwsQ0tPT/J7eEzLTuKPaxin035LlMkG+Owpm9CreYvxgc6olRh84L
pbM1YFjuuhkWELHdNUER4OHLBHVF7HI1/UHiWrrqpXb7sevegzRe65NFI3D6SrJG
MhUG2xAh8+QwwZkEr+C6QGX45GnSmv7E+HFMBmeYqAM8TB5lvJWp6v04opKWwTa9
5wsh4fW7GGuM1AF76tHOhxyyWkUGaUP7UYTf4COonWNizZLMSizk0D0Dyr1ZSGSn
lp1q43zaWAJEnauKneQAS4qaL4sF5+dscailGgBAkzuj5BM8oAwUIpc6DrlE6jKh
3KoxVb9JflRjxnyaI65xradcqeCzks48DxufwScByXqF6todtMKQixSJmETF1n1+
KSgbDA+FB9a+cTfyvmHstupS79olg8uNaSLoByEt2qbF3OEVh6q1bdnLHfIYpSez
0SkmTK9o0okjUtv0lSSm+47O2fEettCT+gpRbScj3ttguOPvN4j3mW8riXVURgot
LZZGfzTsAfg/geime4uAE2RwSNwyKDeoQgGy0DmMP57PPCW0ebVG3cMRlFCeH2qn
oARMMVJf3FeVDXjXozoKJzIiFfVJdCDR4pHY85LA2VwXWo//6PSTXHsv4z61VQP2
bHYkrHOI3vi/s/gOKWceEf0+Aw62U2kK4rskW30UmA55ofHOXKuglXj0dMYIiXXR
D+gPru0Y4DMkspRRprIqNvmUuDwxqiiQX249dKmUQcyb6Yvo3fMoCvi2GUjUoKMv
6fbL8eyizwIqva4iuBGUBXmo83l8FCEOnBe9UksV6Qn4l5Tj18BK2nhxtL/T0PJH
HPdxpb3jZdHtw3hvvOEGZBUYC6MLWkfW+R1RJLIj69wg1fuwDb6kfGHJT1N71w0N
UyiqT6GKoxfUeJWJG0G9UPdKXe7qCGbM1k0sWmZ64jPpCSozOf7ZfG1BOnFblF8t
cinQmG5uUwwR6JHUjte21gjjirIaf+9s7IxDtrNbQwJsSf8VgPuPCCPAXAuMb4u/
wYCSOllFMAoZgVV+Lwo6v0PSlyVeK5nuL3KLI4juRAAQLggF+6Ko8L7VLTX9YTsW
7sM4hU7zgVV5RQ6uNngEp4DRKcXJPw4X/OVwBb9GlgHdu8ZCuPeazivByd0tNzgY
rcbDZoe1DwhrqbDeLx7mpSbZ23m4vt4zW1zprUS58mLF05Yb0M0k36j9SgsVecgF
4rI9c/+E7gHWIXvrw7T5qCg++jR2IuJEwkZUTHRwPpZsTok/aaniV595uuO1oYVu
6yvwQunTxg4HQDdHCQYy02N7lnsz4iJEKXN/+1aumVKwuf8kykwNCcwCgJ2sidYF
ZoZvH9I7RDUvPfFsMo5O5cMWMv7w6dpQBV0CnyL3HyZL4aa8PgxGf0H4l2h73djU
6Wq3vENfVXMfztaL93dWsgrOuGlwZ+dHGGMB84sT2W3XIPJA5NgW1Y6WaQ33h/3Q
j1Wd910ITbRM9BfOctpUv+vTyni7mWwc+hpy5oH5wqYBWjYmraatqws/hH15Gklh
EZiqgv+JvOizVasZC4q1u4MHZdtMqSzuMPIIzDk+J2rAojaHZyQiQeTmDt2Eu74+
EtKgLNVvIcR4eugKtQ+n6/jHSKfP0NVBgsOs8MOm4yZaKemw0XQ1xNIxGF8ePp8I
7DGGbjYGnc5s5qsqhpZvWepPYfPp0xqXNsAR4EmkrsxXMNTW6B0Xw8cwB/qPxwiU
OOsc77s66cP/y5+rgVEw+J+frtjGIw6QlP8KDEE4M4lMrWG5vQoWfAB0c94QaS9b
F91Ml4sGbqaE+scUxAxVwXghQro3pccdVrb3VQQek4VapTxfLCtCY6aEYq0xEH2d
pBgyX4WTZIeP/q1mFTJXs7iaWPN48xkdat+zuTtDN52hK3BszfaBDP9wTHjggVcS
CWxedECGB21yBZyo/ZRbDoDROt+tJFRWXazd35fmpo8RecqPf/WjcHg+qQVsMLvK
JT76h9AkCeh2EB8qJCh+PcVehgvZnXVGwJRHVH370Y7QKCCAL4FqKk2/x79o97kW
SBrw3xlqAHu6ynatDIVItENxlpfJ7CEogoUOYq6v3+9IDztwndWQCcJkqwnYHXLr
xwhW6idjAN52uf1vS2Vh0yhPedPAU9M/LLvbn2diwjDvq6gsmRIHCx41EFj/nYAB
c4HScyG+PryD1yVOn5JWb6OkZJSDtFAJtnbOowCR0MnFPfSZDebsoeFnN1XVv1XE
`pragma protect end_protected
