// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
s30rhY3cnsQw3ps9zPpb6CjY9OOfV5F0/6GfSpBZAYTO+VJLGBLG5TODdi/ERKC7jAF/2FMRyFF6
De/S+mr/3nhfvNWBvW5t94yUPHSy5fP0A63CU5WfU0EGSUjdyOl9augi3cdtTTgvEEO03F/QNuDr
pHityHQNJ//OHy3kCYfiAKEM0i+EwcLlnoYkTPSAnLG8+Tdpz14v8925ZnYQMcFrRWWWgk8hRBCj
CfK5cBEHivE5txr3jPg7Yj25J+NFaS1WxLohOuOs8yVfHhGOsSzWNqMAYNLEr0cuP/53gOwcQAB8
KMr+d4Hg4GhSr+bSCJsVUFz2Tz+e19YeWauJ6Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
mBXbYdPtvZTWFG27Rpt+xIxQjl/2jIkmLIpGIFvvqblBIAITJJJd+UirHOSMDxsdw4+jEAKLEW/k
WgPgVxPrRFFOXbT0+8CIXxCpMQ5I4Imhi71mRBI+uTEIBouYbuX0sARfcE+cTSxnIfEr8F1FSL3w
iVhw9LDzCzsv6I6X3pKhCCH86kBZgPBb6ENfGJXMz3sT+NZ8aYhZB3flXd03Q+z2GjnvBu8TUAoh
ZX1ukMqQ3WY/i/+N5WRbuSSlhDDXKTPOdzA2T6nyA27ZhZ1lGvOmyppoAUxpHUA38vtKhyE925bg
sR6FV98SSdarihnGPBH5yvST+I8DcXRDBfbOvZy+voM/9g0ROfARLNXC67OdQP7G/z28ff2t4kse
Y0csk+6WVrHxsVO+iiKya8AUtukpcQzO2xrc5HsDDPqg0cf3sUEVXHf0YZouhf5a057txlxTr2j4
Hx5dGnlUOb5aUL/RGFd2FyI9+QsG/FV6d8ddTMnhl+mVL2o3dh3eyMQOfLWxIqREMvfGH3qXjeCC
/Dj8KuMM6tRphNnynMVTvTxAX+5Cj+dkmVfCwv0B8woE2c+0XDt01PrQqJNYfOOyF1uo2Ok6Cw9U
v54jrWEo8qJg4uMVPayb5a9sjhbN23ZNEghJAuKPXEzLOXCKToc/2ibnD68KSAvv4aI/184HTLcv
8pfUYCQYg7Ad8Ru3JMzURnVV0vYP+utWiecnff5yCh6Ylv7GKZvTF/6ESb0vTF5rUGYKf4HDABGv
bqPhxmceZN2KXfjqJjg/Mlw9WmLdjvlJNgDpQcBwBI5MIohpRYZ9SLFgj9wYRHMhvs62XrcNjJMp
Av1azwWT32WFu4CsNxswCb+G4NNPzDSI6Nv8jNp3Xq/Pbl4FrLJmdF6WQTLvss9nuz/yzNsRQyNM
R04OrXLgfWt6MeKUINaynIZ3nC9YNzgbypfAwmC4xru9KdrzpDq7MqRtPDYPaqN1Jf+KdQ2pCEX8
yU5yDsx8fjlUZEZfFtPF4g8yA32WeiIsaJ0TYeDNtIx+z5oXskN3ETeWZlv8SSrahRF3QrC0AEI+
JloLwq48k/rGqgmt7At3DXRUQ1BmXe3neNHO4kASKL2/MVpscSdP2qe/a9Yu9gO3w2xGp98zer9V
OnzSkVsSLDTxQ4ai7eYO5W5Qp+ogtfXKSRbyRjE4m3GMRSb028lLom9XSS1SBCOiCTpAPU5TpH82
PEsWZCv4WE/rKCWbKjpS9vSmPIV1BxBr8fS1PzsmjDSvggoV5LnOuMI4sDfDEuT2oD14RsaWIMnX
DdwEJ+hjzhBHceRBV4AfI64LvScKgXSNGxOpJBy9Gis+BR0DyN/urqyCxQmNDkezJkq/6GTZnM2M
GHOen3uyAWI2fb/VqlwSh9N145Vw53Tv7YF/zd1blw51REczTvRqUOz0NkW1qD+tLlT1+cB67yFd
UxQWqALBoeG3X6uBmapR1pn6GCt1NA6vX0cVlZq+5E/ADMdq4qX0oBToEjbR7xJ1JZy7VCRhJYau
ARfuvX0XN4GPo2paDCDgAl6AlhVcEhz0dHWeZKf2InpCbgSqyHScY/9ynaJoIi01H3Dly+GI+Ekh
pEOa8TujwHLDre3Os1M5ZfI3xnOPhQ3mJA2ZmmjJMv6riWASFdXt5lhyI+16P65u2KM47G4s+oxe
W2HUTA9f9QI421n/n5QYQwi21lWQ20QPgIB/KfqgdGPJnFOYgNGt9o5C6dCN2IyQ5m4Oc6igYbIO
WsvW+zPGaeNRTpAC2j4dv/cdM8cnmXhF+B6THyDSERPWAsGVq20KMiFEI4vgJItuDJ0N+pTWfVdc
cySkwHeGW4G15n5loVx1Dlyc4omJDMC2ifTTQ6gFysVWInsgunYfzczbdZ85Naw+Sdk1rLUEcNtW
dz7x7jH46eDc3VyIGk29fjr3zWGVzKNznz2t3YBFlRfygJRhlNXJ5Z/UK+kAZ7+oYfrdLXsaJDPd
KcyGWzbl0OHRjiUUHute+DvYGfXvjq0noCXr7u/J3Pu7TawBmTxmKFvbX/HpZ5uQbu7RI+UlXP4a
slGWxPOzuXNK/eFEhkbVfn/L4NM35qUpFjVejMgCRU3wj9BYgYSpmuF57OmlDYzQgVBEHaaSsOfi
uA+Maaotxfg2BvpvPSXtkikWjofauHiKxf3gRzTTBCMtn7dOm0v6ILg48T2T1hhzZ/Did2UKmTYu
wbE4I3hd1evsTQJLH3NSJ8gj4jNya+xsBtXnzmtrFi+K5Qhig70adyUpqeNwh4sBog4bcklQl0uF
PQEAlyzkWxpIialoZ/z2UTHldOwvxmj50d4vWzjEZ8YeC6iyLKDkdxDrjDZiDTa4fP8bYQSdhDCm
Ut0MTXXm16pvYILLTI0DuwtFuxjKb/d1wRzrjnV3Gc7XuufB3p8BbMeHcIyf5FSuw5bIn/HU7XxS
L2Es0+3ALaeUEDcHPOyCxgHqJxqMzpyo1lL1Mytd/x8JvRUb/5kUX45MRyUl37Io8X3Sa5l5FqoZ
0JFRQN3tnkxKlIU1cCiAXZvWHT3TdAsMhYezyMTxt41bLvYuVlJhlLHzzBjm6PtuAabHVTlGnx/H
2JNKKV8Py+1thK1QT5Z8j3bTG5netEgWWMkvbiXOEZ2w4Ep3K0lzVxkFjrkIszBMQw3k6sReHGb6
0NgudQKOH89H47mmSmYUXJ/SXpK2TW1EgOY0uTsTmn8K54jY7+eYLcgUfV3DoI5RsDIgnU0pEicj
XHhGmxnA8ok7RydSRww68zI+FhqvktJGENP85BgZvy4i3Qt3VBcxKExRlRTQoodws5BnFiZzAzLo
WBgyRu1bA4uvrCBAdPhPRVzHSXHWTrUFm2zVK0mMm/dBTdXq3bUjXHdaIzSJJYGHnGMeGHAXTpQT
28V36Zl9NOfMABvnR2tbiu4R3lkIMm+6S/0+ScKTp9bleH3xAItg/Hxhfv02xdJOizXACkb1BYK/
EaYyTUuDJIEs24eYg26gRHP/z64Y92CMYoWEUPdF6cAR4JjrAtY/jvYckkeFaBf1zXZ7MeDWgJS3
Kw+RoZhK/h3B0647AjBI9DUfTuunAsu5eDhUiluamuaYwQHHj8uMJ7xoyVrD4Fmncxm+gctYvpVn
1/FENbRpRJ00p4PjpOMU4DGvIUjj7TyFD6KVq9P3AazuJkimjl7PTe6lkA01wYjcESlkwDfdxqqM
xlbb7OptH58RkumIUnVCF68g0mQhsDecfZRf2DWR1qceVdFeZiPsO7x7OgGVokudxCwBBrG5fO2N
KJzXbbg0Xq/p8L9OP8V8wLG8RYXvFwcBJw4b5UOR6eVEyv/2N3sjdZJcpBkAw2j3xuIf92uFtaUM
eJ1Wny+Qk7x3DzKO3KMySJKtqmhaUGo0FXtZTTVJpDbmF6iESF3Wu1tMgIyVSGqytubY6d2NNjUH
PP9sNQTSFORlf+idKbor9sMAw1ORt8OrfBv/mlLbQ2TPma4SOViqmATNkencfWOq25m7CkW3wWct
yGB/h/LykfD6kBLCfHlWQ1+aYGfCEPmpwWS1caBMAjgBOhYvjHOiAwiMjP1NCi3YLL6gp8Iv7Nkh
Sl8WUUNensgbE3kSXcHGwYajx76g0oWO6us2oC6p3VWO8twUHvR6gY4izdTa0XtXs9GslB19Ry0Z
Z6UT/r5jdy3vXVfLJ9RK/WdJpw1ifUFMHJwdy9D25HNMSxGsiHKpa9Y01xMwTQBu89RGPwqrRuJV
SK5YQByF9aIJIE7ArrINCb6KKVCzrblQv/On8yJAaH0v14dMC4jW1l3xMuwqTMfHa0HllrXfc96Q
48Rjx6GYs+2O+kwkyx2Y1Py5+uN1/7DG9zUx2HvcN/0EQJ/e+kOJRDf5wqVgRoTb3DBlMWA+1g95
335bRb86o2kecfpprIspMSS3ZfRPXfUDmD88pIyUhlihe/luOrghLCDqh3iVlcK+hovCN3XFmBwg
nOfj3yohE2/j0IRUB3fyH6HiM0nCfqKG9eYpXTdxFT5hzT9mMmDrsdKKKtVg7uNR3bNDq6ykEZWg
37cFSv4Q4NjFr0lwI1iJnGOH4fwOkI0l9xjbAseO9bkyJOoj3V5y936IYrue9SF5DkL6Sz7t+MUt
WXQlXNKmT7CxcOZbEagEGAj2GOFaSaiSIJBDYHikO24xhFcZE8yutSMTgOdF9oE9S9hh+41B0IpC
WpDBX/FFB8d/CqAeF+p0DfXfKAKaVe34mOrSXCxpc5nGUyIpfAxn8osYtn7PdnZeZp/lS13otEG1
dFd6s1CvZ6xTkSmP4/mj7jkWqjW9ZeFHQrb3qSjowk9tscXQtUyNwIPB2tvrvmcKAztB0RqaQ7rz
wssTbi5o5x1L1Zg/lCUWGulOb36t/gZqCMKvF/yO3o4i54mWIrcunYhWsP8za/8Ya3FMwTtRlEF/
e82plijI8F9bIkma6OmAWgC9swlqinHj1bpbMRNqitcj9mn7FvsK9prb1+6Bm1twKFGnA4lAzy11
Qb0BzvYztpovV+nC5q6o6p/DNxfn4Y/G5b/wRWhv47liKI0ow+N1JvCIzzsXz/+nOlWakRZhrKMM
WPqZp80yDShl0cSX+8s8g+aGdjk5I3/5wUosjUBDS0Xta/2ndHEwUw6w+sn7ruwPYf6W4A9uVGmf
r4fu9qjYdwm/Y2gG5feycQlOnPPZbUoHdphzcCWM1Y0UVQVakX9R9QR1zJ/lL3122JEqbBqH2LCJ
aIJ0UNuVjOVj+AI/GzHblzoYmxqUQt5UjmRM/a7F06fr6nR9sZJNf8SSn8LII9AW9CRLZWRoEPPr
Duov0dqbmJgQ8FDoXQyW18Cm7NTu4OhVcM7CY2deruxwMitJ/IN40bLE67goLPXWwxohrvqIZ1gE
OVCIchGeBag+Fz1h69LkFBkZgA3Yoe8MYtoJQHnAznp2LEab3aWzzWgF7kAj0+zkOdjl9yYlCqMB
ku2mwG58nOs2wcsBnL6+MrRIWXw04SNUD5RQnVTJqT9FQaEnf44vCqtNs58ff7oephtGGyAUcy/Z
Psr4TjV+Tu+C+++d14HEagI8wcKwoO2spYDpNpWvyQAcd1uNYDPylQTcdPGq1YZUo+orbuHKPkuZ
Vh+TsrEsfqmc+82UUYbsaMbMNoT3BTWAG9lb+r9fmgDGm5LiwyWTxmKzHwBHHZKhUJfOOVkVmph1
hrPm3cCBEv/rxLu/a/Nzf6u7ifGvsNgYAsi+6kKd/BavKFjK1NE2Np3y+FBtImIUMPZoEKY35YHz
rysPFwTu0DtYxnHUj7jZVOlaGiOY9u+RnUrZK+3fsxzypuBovh9xvlOW+lO6JkLRqBQGFmQKdby+
tuWlbNyti3sw5PXT7nXzIMsNuVdYS+qNGB4ZaWb+hgw6rPCx+wn4JA5dASKgFTVcBJSQV2679BF/
XZ26qci+wYZwlgjAsGcPF1vPijVGr9hvDvTyyYXLzF4utgzUHVt86Kzbgf3ZnpuYZuLsEEIjdpwt
TWc3AMo4HCnTXOkANyYMsiwNrKrlznvOwdOmQPfljAkgJwuf8viikBmuVM4xdet3VyvGRwSgYYL/
/DjmCNcTAHo/t8PV96IvE/K5FQaR81rV+ie0nDC90ItqQ1ewTCiJea8h2ihWYO3TaQFKNeWarH/e
zY4ihPbVWV5Npi0cqK516uAiX8dxygvS9QSse9QsOzFa+as+bM7PF7phO2UObQKkpVdSGsILFVqk
tLYONrDZrc3ICehcu9PfyE4MQI6M0SBxjCZ12wqgTrXJqDn3JonuAPgy8QxUR6KhWXgdQ5VDGsCg
z1+at7KxFFhhtsh6nyFdPISDhBJrXfcUPJsNuvR0jskypMD/jrX4LMYKX9rkwFfEUly61meOnwSH
eh97biwV1AlGOF2xyvGBUkCb35sACK8Z9VfUpVyTCg7PJfTCowzoDdTPa9Y9NsIWPl9W1fF/aImF
IK/7V7HCYtjtmBLY3E3Nf00kqjuv9NPj+h2HIlcObR7sboqzL/5VealY0aCJAhP9McQhEgJY0HOx
jrVy8ggkjJXo1N6dUv/ZTde78eTl/CilJ/NmHXUb+aJFIGADu8wW0ieYwKxBWKCR3inuql4auVAb
vwk29YUjZMKOGQIfObkGUdIuS3adpnciStwlI7P6Rgq64S7da+YIgQdWgVBMWpAiBXOAeb0/waJi
ui9NIqemDF/4KybY0Bxe6pNvXlwH4QFdpjbibHTRoB5Joh+UuWynUQXNmJ9KXXcAX1va9YKZkbfT
5bwolU12lOLQBK2LZ9rLV9NTKv2lcLLiXXE4epShshwwd1wnZkGNLbLaxBf++p4HKBPoMyZignbg
FpVSDNyEdjyXH7zFQ9huFcEvDdZm6kKS4Wz0mn8cg1m/zakjuB4cZcHnvB58wXRem4SvZa9mX4+g
aiI0+Is2Qr8nqblUQHmYtCnI7+qon3to7ePg+PnAWX+hmg3UhrH0FvOcHe3MtCmjxLx1r/9+BejV
cngAAtnxQLA2t6AhaAKprATvYvMzspsRtbc0Z8eoxDrCR55Pd38qvBFwPykafXKzaSY383dyDmwF
IbtHB7mu3nabtByj8i5fApf+58/sNK48wdoW5KVmrNcSmsqhMy+2AZeLauunE00V42vtQOrmTjNS
Fdl1EF5JZ7Hl/k+4P/XRAVHJRDPmIddCmvR4IqbAE0gSELZn3uk9Q5dd0H3x5i7zO4q5NtROTmbB
bQUnOmju/BwkiXtf/ZJ+WobR9zwl1AvcFjETBAUw+YAxIXE0kqmzTag82nuutDTDztBPVCLrCiNa
JvvJld89mgDHt/65umFf3vkjwCdFAb+p9azOUIFzwi5xOAsrrpQiLvv1wmaH/k+wJrMTzpdydNxV
L+nRD9fUnO3Eu2isKj/COTa4BVRaGR+DNktP2KM7SzBIoz0+SfzROlMYlz1SiFZ9KNwJSc2NQI+X
+2FbNWK+GSdHvxptfFTJAbC+aTWKI7UA035VbsQTscuyrRQhksouJGoVHpxMLdzamARZGQawrygt
enjNSqLZ/oSnFO5WNXXi47KgCskafA5QdK8Q/5kbegRg1vUvFUHjaEi2qUuMcSssjfXuLrTsVJJm
+HwRPS/RhNUDslg8khC5p9JOAZ1pj0nX3i/JQhzUYADovpY//p55tnP1eqbCBvI6HzF29DWxub5+
qo8atKarFwKyKV6+RDAojLWPkyP6ELt6ewC1MMAbYkdOk23tBD9hqW4Ey5GcGkzMRIp43Inf9+Me
VZR3j+HfqZ94zn39Wc30u1nCoovIKEYD4AaskgTVwqKh3MU7hSC4p8S4tBgodHJJx6EvVQpnpcGQ
ORyg+Zyq2gq9XXeQ80a2718Kq/ImBkGAXC754zQHiKFekb0SIj+Dp39IYLm5FHKL3xZgnubUWMxd
Pbf5CWa3U3nfQiNNXkl4jBYvElrcRPG5oxW/Dmq/0GYD8a9cUoHa2TV5XA3alV3w54UYb026jl2s
CqX65hzBQarFmIyITvIQKAPOyP/4j/wPk2FS3rt9NlcrQAsRQ5kxcId2pH+51PQaTJAsa8qbtebd
wxrKk7Ansq3kA9s3VNB+SJ6fkEXbFNFc1BZ/aGmCy8VZiE8adSYkT8B1LvdsG3Jg3lhHi3zfB078
J6s22Tr1U+W9FYirvHXsYgY8K/ypY3hihG5Iw22Oj3UpsNRtINy8lG3Dyf6mmKzHmF1pjxnBuApo
rcYWD/eO7moqQw4rYE8sfRRys4ckJpi+mP2sPWbPX0ONd1FwEiWTIg3Tl0RCR5YQgQQaNhiFtIaz
IzoyKq3RrDVzwFwAMMmWp6SamslvVBAshQqx3vfvAJRN8PDQMlb35MLQfl41aGyyjJrH6T6xy4WQ
8zPEVLzNfDAEDEaVJ9rnW5uffoH2rDab5BgKw8w1U5n1LP0BV9PXAnRkjETnZt54TX7Xd9F53og3
xRcXHSCgISqN2L7BwtsrLVCDy4iXtebMOfKrVWsVfE2qqsyM8X507ZPY/xZLqy7ntyY3LI1MbAue
PzZDVeQKANQPGMKBCPhtB8ULLHrYjkVWGZ9TuN6bhgs+Zh2icnB6qAxyHXow2ZhdTB6ll0421sbY
hJjusaD+jZMWO1s/qGFZxrm47rAQL3zN0087qBILKYwYSLoxiqPC3zJ9RHCKaMTfS7Qvk5eo/oYU
rMSLEx8Bv6+BWPew6cADZoOZk+Si0s7xUPxQ+si1jXZ2FTq0cBWCWBOoZSLt/xORMBFyjHBw2QtO
yizT+1hBBZLtSaxEHpwdfRL9T9/DWEsxsE9sj5lSmTFQJq7vciqhZUjH842ScsgJ9DcniqxRSIKk
HzZJTZAJJ0eBZU262fDYJaGOtofUgGOniuvmxkKBZd2t5XbXLJxsm1IvsWI7q8LecIiPXVl3EQxq
0AUdFaGbm7unbjcqchV89VwGX0PXYwb0WAjrjlnOa5QmGOMYHU+4ie1fisJcAV+F3U44gOoiN0e+
m30Q4ZMbf+36aUuWEdmYH6GQpKwDQlovpDan7k6sIwOj1wVYty5BvkzQmcAXatVV7oDIb37cIyZv
pwZKe6hwt0IjFCVmSf9MaIOhOFu2MWQsA3kTlCyaIKpch6Ww0Y+v1LYu1LKAPaXnpPpdig6e39pu
Zzan5f1ZwsB5VOIe6y+3O6s2CxLjm7wAFh4E3kYlK/xZ62R1xJQyiDyrX9DlJcxnNPytfjv1HSUC
3HtHB2oMg98Khrzl1+SSgsVNRPSiQPpWuNpZuBwbzEwRFZLo3TYvTBoQKXPyyH9Edj3SdJ2HgQsz
ZfrDD1/0kBP/C+Nthso3XRJJsBLeIMW0DjJWDeqthj86Zsib2JtGbQHUo3oOrqzfLSlsvbHETdn8
MkVJaukMnlVT2YQybteKvcP0BOvfFcZtzmtxJgCL/lmYPEOC+zQ9w2TXX89/GN7iRpe9Evq13bI4
C3bbRFIqcM8TCJj1sjIFP38NbOryAKkgZ5pLbRIGBb+A9I2iN3fbUVlMJlJ9fe2swsSsJf8/IcFb
cEk5pZrTEtl7ILcy0cVQHqDiwE/GO6yV63VbqvMTtBGCjYE97q5p8tJL5ig3r6s4LC6h6Rn00mcK
HlqMHM4uXYpMykPe636QlGCPUaXWxTJwtaeYGWJEjfT2d1bP0jj8pU/3UccpV2881I9ohp6Mup9Y
+206qH3oEcUB1GRtPuQMqXba69rJIkRoieygM102NI+BiH58aza3WUiAlfe+y6qib2/byM+oCkeO
LMRGrYDMlZjEn8n1+LePngqaq9OrktD7MlUY1PnMwlktsyQ6qsAIIKS2GS+8anV4vgScnsSjQS2t
DHkopO2i6XXSkHxBUMsGxvqy1ILMnDn+kRTgbBXPlrceeSGUhgFLKpDSzhyC91Fevi0xBmY9orAc
hbDMRcFU2Toa/Ttv2+W3BgQGrsUBL0+eXTM8ZcrLdMntgvwn6rmVtMfJ0P8bPQkQzCD/wQUmGyYi
IWeB1aEb9mktZJyRB6ttmyYSLucMB8zyWX/k0R400mh51hom/+8YnTU8lbB3L3JYMuSvrQIYiz4j
EGQExyJQpbM6+7sLG3Dk/iflEvdYCX/AxZzL/2YlLB6AQXDhFfv8JxBhyr7NvM8lEKEHHYF+z7Wj
uYPRfB17UiOkGhynW+oiHpKftUvJZcri0/uD4omIoMfkcDgVRrypc7MQSb/ph9OxoljZ+gBjNZ5q
3/dVAbmG5XOpSD2FCTX0b/9LMoGHHvBIXjRw6C8Ho8UZ3aUWDt/FvTG24nQb+2mgfYjFUDEGjaqo
znvk9cw0E8Tch+ovwfaRt0ve2byW9y3t1vGdpM1cCzb7ggH8YqBEBaVa1Ck3sfyKX7CCQMIMrGdz
KscykS3UM+/3OS+CA/I/v3BVZOb/G+BbRqnYNB1w6mmXZS4n8c9BUca9d4LWgBPoCyPDn4Vi10MK
C6YeHS9uMYxNuaqLYTOxhP2FsPJsPYpe4CBREIaJru4jr9fEQFfa/wvLREWPZIbXJFUHm8YBz0Ak
QflmlRCxStbt1kgaKX1W85wc36j21AYB2tDoR/YhedDdNJFJ+QHtkRk4KzlWzp1QoQRDqxpoEsbK
KxTe8dgxZNJsvc4CZDO40OoLgmgU9dFyccvI4u4sQKcwZ2f3rhQkbtl5841lzMsTHgAFipbXXQy/
4R36oNS0nd3J2UCOgWhKaZxq+Yu9BMac3ySyGOrFKqKVQb7fosK+DCzbnNTmwuWknfxqmAU/+R9+
zNi0S0tQAAEl62JfkuXRCawVnejND6WlFLSAuu3AD4AfXJemQzC65rwv1PkYM5PQWEuQvIaEQs3E
evovVb0R5i7QleZrW0UUHLyQEaXfgCSvBvndK9UdzqJjVdD5YI/sNWmEdmO8N+InEhoS3pg6AQTu
4d7OqJxTrp2v3vBO9kNvFHjiEzJ+Qa6EBX+AZUidYU/SQZCi0a8DFxZQF3e5qV5dReiSsLoZw0D1
fEiMykVpPnEyX/V2Pv3oEg5QV1pdAQgb6zxZWyfjklw+H05rezUBDWvIMWPfC2u/4hnLOFn0bjFw
pc0po4g4uXP+2AYLeWvhGuckLKiInnbMBFfyXHB3mqCecXWIwUdkY1FCO2b7jV5IeWCFknabWnfi
YFXkCi0adosP2qJxiBjIJQ89rr4bxXtXIsp27yfMBtvNiFz+RBFEtmnpExZqZaZnR5wMW/1tB84S
gF8WWLnk5HeQfAtMRAZWcR2F2cDTi5eG4LXt1ZNfTUq91ctHDNj554Di+Ff6ztpPC1JEvYY//u5L
9BsMF3jQefMxhRMxdMBzFqKtfCv0d4aeqih4ImxIlfsn+oOTjvIdRt8h9jnJdtTaMg0jMdf63rb+
emM8iGpOLfieWH7RB3w9DWP022O070S50dRvjpGmjeM4SLJ41RAFHp9T1qjGyei4yR9Kvx/8jUeR
WyIzJ51YLZS379N8uy+J3RZ7nRwVNVPMPUS6hK0273gH3yuYjLExM/vuKzIS+jtvu8g+DyKeUtlz
R/lfyjxsVLGqkjkidvKg3ByiFY1XA5nisEWNqpETMOLp/qQJgpy/Z4Mg0YhR2EVI9KuntqZuPDhH
YYq+PXOVojlOqZFYrg2Ph5+JMi1/5XNuSfd75E+/I0I5rGjf4X1F8HLOwV/ye5Niwzpkv41S0JZT
+epWn4atyXpcIPi476E/9OqtXn3YJKCELRVuPWSAwnpFvSZTgYaAiK97J+AGJe3yZkkfusGR850U
q7793rGyT+dCgr7+99P8lJ8AAU+wKw8Lxsy0SXw51j8AjQ9k02nwQIxK9eB5DeyYjkIWHEsnR5k5
rY74mtc/PUmsuNBEjZTOV1IAEfVveULjUcWJpEGmwl/k6kW2chcWdoVhuvx85pxoR0oiqYsc9evS
YTIT716o7o2wgOMMUpwnIdYy0l8BFoiGQF1nv1Sw2QGT95C2xom4wGickib7T6hX+EvXi56xWbG8
SOuZzt3U4zOTzI69EEIRlG4Rv/re/e+8L2n8tp+g1+ffDJjSHl7KaIJlP3fKiolmX0fetjXaGYvg
S1xIhZYT78Vho5Iv+ewbrFv2xKnsZnNxokQn0+7Dv4FhAHpRBkn+aytOQ0BbV3S9bfCQFNQy/WHO
3kM637WvMqPe9szzO4jCY5oR4Nw41VfwA67JZ0JWDvM79PebpY5tRAtfqwm7SWvDYqrYaX7vqFqz
0/tBo9aMGyfyNj83YHUqZMrHsElz5vobf2G5/ziJGg/rf5evx8Cjo8YfLMOMEK2rvMXQyan5MDiA
ZZEu1eiiPt5kbKg6QsjymDrtGYFxIPaWxhn9BffpBq6JSgVdV2I1ln5mTVCuhuU2KENjn+jChiIW
k3XM3LSzIaXtkUaR4zEltRoSsr/+PshQcT6XGWdmq5q2sqaFD6SK8eQgnMA559jaILYHNKKbM4k8
qyfQQA8F5hEg5/RBZKh2Iv9ncRIwoCbSRVoCebZmV2jdGCmSNZ0pNVcZeZ7FcqeaeL1vLHRrph9e
y2hQhaaplJns0enT+U+49nkZQtuUhU0SdNejUpSnX0RsaTO8/MEEvXleldhimVN//RfBAudV8tnH
LyRf5Yw5v6aQ/MiS9//R/EeupcouPm2wdkRTEFa+snGbueeObWq/kf+leFsBA61DFLSUAcEgStio
jTMMvb7RSifettnk07wFnRSm3Dwp5Heb8CbzVXMWXszDPXQ3BnpRP5zjW/kp5qQYJQJzv3nL0FL2
d8idtJrjgzDEkbTL+PDTMvXCnueo6fvaCmvzcT8b5TRVTEF7DaMvdkEvL2aJ38xm2jjrizlA/zAK
BpLT9hBVv855CP0Dmf0n23+DGWCdvfbVfqfosBem+54vPYT42FU8PBUPHunIahK/s3JfrwZrb7oW
2bkwlMqtqNFfageSVl+gfoQu1+KVinFyIKIFrYFDKeXkhquwphAypyxe5SrN7aF75wTVv2Pn+ly9
aAfUwud8XpI4X0sI840asuxI5sl/GjgaSI6g6JO+VN62REHmPjY6A3WlKx/sjgnTcKzFC95MkvqW
uQ8qyaNY7IxTXYibe1+Oj8Y2vAxqAe2ZZfkyoS55uN+bZgMlzY8RhSYCtNLRbLnTzRLAoVF4obuy
ExytjQsBGVlLdHxEQ0gdVHosKk3IsRmG9Xi4QQjeCA9LObFQAVb7vuhqHE+W+sR4Br07KMv7Zf9x
SIQmN5S41aysSKtCWU9QdAbAWcpzYstu0gn23uUKlrQvmj0t20aIeT8av+dXomxVaP6ow8B8DCxl
7Gv+RafuhpA9cboXq84j/CP/EKC94wZi+2O2qCE2EPZb4AQBlt/pKjvrbLcraiD8mzzXQGbig8t3
70gmwEmqetWO5GcMjW3D4MWz9JTMQL12ETpWDu0W6UeklbUfiGw8jEKLuECguvmX2+ez5qPm2St7
IqUjjgyw+b77D5UOePBWa1tjyvdr+jS1Y1Qfm2S2gvoedwHrDyb6/wejWbCC76az8ph9oxEt8Yv6
Mu/pznJ63xW3eTsAQMLd3SQbq9RYEj/Lb9ssmD9ybdZq2kEeTa8k1URHdfFEFKa6tzQyAcWnu3Ph
y3CgqKQ8NpUqNZYxwEKmZD+cM4T82bBJIHoBLIJUT4v/fZ+fkdcuXPNmXIGdBptOEJIITCDgI2Ax
iK+MR5Ka/MPSkWZIaVwEyu/6UnEhy/pSTd+JAoaWrXHkgiBfoJxplSesHlju3eTa548EFEVnbGTN
s8FM5pyBvqDbz3f5jhrHjmZBKHdSQZMbbXfaLq8/gb4qc6uQcmDQmwHeY+IbOhkzVfXRzB+pz2wE
lOy89QFXjMJMzsowLGZ1zUK1PSMQ2Ksx+nqRSmukbEqoXEwVQ3VrR+ZMwKlpHGD0x7UQeq+xWOTY
vaoAUtyPTkpSSpssxUJWPP6ll/Uo2l06hV2hGDQqeUodm+5BrMM6CGoDCKonYK+w7mFPy4ZelXl/
XOyxI+B1xg0dVPBK896pODqqqVCiB8CSKf0mw3S756Bj6XDOdwIdSVoa1H11iRrwAD35So/nxW+R
z9RIY1j3I9YtEIQpPKU998deJ2ugAc9UT2kAIKoMWCivkiRChxSi7X51HQ5YSJo38TS3V+XnG4TN
FdLbTVRGjV59z3klQNoU8rHrvB6CgQ9yeJN5M+ppE8VeJCr4Cp3Ml3S7B1JXhXMT7QWnRvS5IhDF
P8lKpD8rBhwAoj0PqY3DQ+sCtPyoLacfC4mZz6o/fEmtK0xpTtyLdjp67ITWdTBDjjgsxDXJX8nh
CimK5tzJv7L4HSohRAxA3eTm+u8okK54QrUUhd7Bqwty/W8Au3jrhv9mmln98jZFT2zkYFfz/B34
tzF6hZWR+uJVoo2GbUZKjANF2YQKHuPzG460fLF+ZGEHBMJUNpvXg8+VXIj/fcWQewURCFFEDd+R
4BhxGkUeEyvSuAkBNYsRZ1LX2R9gzyDz49rVCcftLXPDJrL7vREE9ALNDLoaE8GeguIcJG8em+YB
5c065sR9zQSuZQucnOuzQmv5Be8Pbkf7ZSV8yUEU1NsNo2dXN3eue/Q1khu0EcOIGLb2W0U/RIbv
ii7UKtVGpcLJXPXKBfShGz4dzmoSf8NEoEk1ag8cFfjjev23R3kZzbD8+yC0g0ZrlWQkoaBriJ15
n/z17huKpgvJezKnMVZtOPM1wuK4LbU/MfZzyC11Znzpwc5cUgpu3cNc4fjBjrERfnFU29Vq3xTF
fqzG92ZtXDreKSMnJ5S3Rwjsb8MK9EGI5KQU644/R3S05fBBMtGn+UvThto5jOeL0QgPPR7mKOzv
ETaERg3FRK63fgSbIanhFooPO0QvviWv5RrCyo+EDUJdMmwZqer7BSSjRtAo6HQx1Oat9ZfT8KZt
k7GARdL24GGPTRhNzg0JsHBYfkA4RkhODW/HkfhhRxt+ZdY0tnvUAzlN6kHYbZiRed3qeDNa+mk9
UpF2gXr+LyJhs9oeJ4+MstdyrT6UuT8xtamR2I0hOhXTDh+aSh8oLUVKjdZsqzBTA9c0LvSeYqRk
qwSToOCmTxTU6/eYjWUcploMd+VcTHsjC14ETgxmqFDVGf/7mF2bwSNIICq273VskOdd8LJK4yXE
P9uzm/0pvOk5OvuN5aK5yYeu9uDnsckm7aQOzHP6EbfJdnc6quckGHIzJGf20FVNR29d594dW0Yb
qXEMAtuDxVoP7D8FkzbUJT+SBv7/bnwpfDng3BtK/z5JQFyLSvgtFl8U0Kk3uN6jSIftsrrBJNvr
wI15d5MLdj9gJYHDtmAFLZiAacakAxMykiKQm8iyJvrzW5uBq+Px7D7CemZrHfbrn2giafaqc4dE
cAHd7HODcit+w9VspjNCCRkTOYuK0zKy5sbqCT8eS0zqtk7X6P04cvmFcLxkYqBMALKGBCbqopmY
yMbUaOgJuWnxW8hyJoTnlx5zt1JHKSPdixYHVkxyyi8wH1z5D3Bw7sK7inOb8J+3ydCIzIHvsegt
1yJ06DtnBD4sYj+VcBN+CcjpFzo1wvVTecxjhDgVS38KnCItXdIFNmu+9nZ7g8pZGdCi4Lx+wtcL
hjCSwmEniSJVhzPZSicJKcnhOPycsD5Msf8Vz3mEDX4E4K+zfkqCdc2Nbxib+0QHFy0r3VObl2zZ
TBFCSCojc7heDzxoIiLpCR0K7oagCozOlHs0iq0ttcrKqeCuSrPAfCZ6ksS2MB8xN9XfQAjQin2e
pJdRfByjOrag6bTYuTukXsDdw0sf3/wEILxkaBi1NYMEQ2S5H0zmauYXMavEJp5Q1iz492cjL51b
e3SaoGDUFf3yAFe4hEdXSXTxFrI6iV1ZUDuYTUWlGeX+7zj6suCEmdXiZjqG/QDARTlwSLZ+trVz
viAYu6aGiyJyLYj3rNx1C74p6pYV686+cP6lO2bd/cOa0bOrvHdOXkC5Sb1Wo19hY7Q3sHC7SGOJ
GFDQtyZzEUJTEQoibjhVWhzqhEJZmn2v4vqJK8J5vmGJSDEFEwduCT7dz5jcSZwjSQ/fesnqGGII
WnRvbMv4NKe3kOsYqy9MSbL9Bb1/9e4eVGMqQSce58T7Qi1CQVHUXLxHD+YyBUm2DZ7d1mGKch1J
KfycHA==
`pragma protect end_protected
