// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
dYtFMKmXJu1DdmkCQPog54cIbV+whiHMpZHkfF7l5AUe2tgpt3ok6shm65ZEQxyodHCo6FSy+ERt
Nv7ityb2Tz7rtLtx/HMUnSe39qJutvEUjKr3HlhqHKZwA0vzcCOVeEAuQ4LDsk3u5c8L9NU50Ar4
jrnjm+o+j+ZiQDN1oypjz4/tIa7T0ykynHRuU7jEa/psu4sG6OrtBY0Wluh8H0DjU2GQb/EBEkl8
p32l0Y/fJ+YsimF9C4aHMTWKQ6j0f4rXZrUCwuEmHYYvApC3O1fe7NlrK42dX2t+FEQm/b06aILX
I2RDPzhzR9hQV8vFz5vOuPjm9HzBbnTVsYMBcw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hHh9q9x2pFWgLe0XLKV6AviUeLZJqARX+XiBiL5qFN4e3BhL4w6GMr+rDtDfdGMdxJr1hdzfm3pr
1dYAnupiT0qS2OHYcr1X6tImEK1LY2pOvxaNK51ZWwqzLQbWqVs2sISeHHtxt6bhtvIfvqqZLL3Z
pndfmhFWpVRb6wOTFvYsR0ihNMtlC2TU4P7fUDN6SmK145j3tjL4yV02LR3mtgTIDbnVkrsCZJdq
/t7Z9T1UE5r9z7JhnRU0Sb6JugoC3hG79ziuDCNVyUhNZ1/D5hp5r7hUw9lKnQbCvWycQJrcfNOO
2VzF0WC2yo2s1aUJmMyVU0CoxwKPGnDY6qodvrl/IxRAAb9YqysNXwA21o5wHuM9M0cvSqX4QNKh
J27I1tltn7K0EVcq0sMxeCmcE2d+56LM3fwlD/+Tc5WR1W7jpbQ+8BsUrj4r8zy8M9vQl117Nr11
btOWek25EMT7LtlfR7k2grvIpJuaa/3A+g8g2Ccs417wN4SkT7pzd6JN0AuvD9wkTGGbqJb6/17b
i2GVmwnSoggV+dt/PsjSJBwcafzie2haY5Q45obqvKvk9swyfMlQxvfHKiDg8E8A6FmEGAA7y7gs
4/sMlMS2bh5uLsnoRB5kdORKUtGVZAq2NV0K8dRAvAy44WgmCvVPJ+YE5cK9Kfuv5E0BBcAOW5/R
NxRxf6DBdoT9b55WFww9O3wQ9nY3p4Ed0y0rkUx7Or6smQZ5WPAE72ekVjWL7GHP08D+EzAlLezh
pfWoQpOFeyessr7TmCwJEse4hplm7rJSRYY/TFlpC+X+NKqN54FyECkRKMjYQ0RxfVyQbCv08BAT
ouu3mo+TBSQcSXEKZbMRAFW4M9r/JZW2Z+AU+2z81lkhZz0XuzadXjmNAIPOYZYeulr9UZy4dgrR
A7fy8KBjF/5cCVc/KCDdvd90EbbYvWd3pkPBkUpQhANnM71w/Odu17ZmjUpkHOadRqZxgntQde1i
8AJ80SnYGXTLQB5ckkl3BCfJnSPoJwi5uo5ICRvsNpgUlK2QMGD5lL6PJpe9ajPoPnXBAmRsuqQe
16eTA7SuImFV+gxSoO9hakWu4maGpdq1BLh260g8lWNt0aAwHaF3rCUUAC+Paq6xhvsN2/V+Tpoz
Bbh139lp62H4A13+gMK2B2of+GLoO/0SvhS4E+084nW1LABZqPK2GGq0mB0SoNQo1AvPrByaZNUS
jZxpx9tDJwCdQVEMmxLnpuIHYw6FTD6BkIOhzz6MYnNc7u7aQgHALXdB598A8V5AiY8W5ImdhInO
ABbPYEcMOs4NhKqtW/4Wf90JmWzW6aOnf8cAKxxzLFJkZZvkgS2V4Crqrosnbk0lxH5uFydoWSf7
+gbAI3w6uej4SuxEedl8cvCf/swnXqYGgWRGr6MfdGnlOGWKz2D37IoJo95FjOcq4/uREwEMM16k
cc4DHx5wA5m0OuisubBKZm+6H9RdV6KEYSVWWl3s2eNLUvjEzpkbUGVu4hDB+IrQLRu25TLSjRMJ
9Y8iIxLeV+st3D3Za77fd1SwF9sA/j10bKyv2GneLjE+ZqU2q7YyVike7I/KuhMI/gqdW3uZnW1M
UEOdmkWh3s71p3lYd9A3vXhT2cwqF3meS7yQ6Nq3YVYeaQBOve4jwuD97ZP/XXAJuqM4d6EgDLPn
O9YJtFef9axvwiSTzgDIHpzXA28R4y97CYJDFmm+pLIUegs6tFOQuSxu9uYBRPA/dzUliZUDyKSE
R3YL3H/aggh7ie+wIAInSr4gRqZ/K8grd2zl3H5Up9hQS1ZnIbncgBRop7q5dAq26VuwGVwfJUnN
Gt91p9dpTlV0/DzCfa84/h90+2Ua8MpH2Of9lg3qBw5RnR7a1urhIbM28KFyw5xRpWjweLZpfPuq
HjgGxAHk7FSr7uh+XhCxva8/wuotLWBZcnMuyUWoMp01sHY1MOwtd743zgsJ1OhJPdEfQwrqz/8X
RHuxa92XBozzjAjW3n4DkOI2i7X7Cyc3wN80FsHY6kvq/ykoHchHufKWqDvf9XCvlSxAeuRs7dft
YsCeL3vZ8q8UPOUE9CunNBkpZKEpYuPkqr4eIXUIZC6iW/Bn6EWGVhcpgFT3aQlXwrKAaOP8o1o9
2tSQCwBzYAuMwhLOhr2GDuOGMlysYUtk6Ug9yTHyZDkGuVqDgGLnh+E0ivUHMOclJp1Xhz/GQQIw
L3e/+r5aCkugUCRVolrCYEMGAgJsPSe7uZ4R5XQtJWTvc4niof3C8KCLDwash0x0GovDdcgjCyEV
06Aq3Pir8mD73sgUe225ToO9/SNSkz56QxvzRxVgwjTF1vH317H9ZxE+qNz8rZhDPjWG8NKtqTXm
hH9ulVKH5Q7EWWjJOcjZ0Tz47y7bM60PiaZfstCzlr3m8b53b/RV+Wp7I46uII/ZqlPOrhgVhxd2
kJgEThHSqyLp3P9Bun9NUquRSJ2ND2Tg0QGvrdcOCNfXJ8k0X024UyX++cqTd30mG3OXE2yg0r74
vwLc0SVuZdqq+ZS1OKVCUsWeLD3CzZzwtQO6HU5fn1hvrWCEnWbpsI651XnAeIIWzeapDS7oaxJ3
JxEYeGUh+uh0p5WdNbugyLXaZTuziNUc/TvomMcoUnHYfexoW5eJ22xBgENJP0DcJVsVrKPDslWw
8WQEjDWusmfVky9QIsOgGT6+IJshXCl0a8XvMx2wflQ7/0hpel4cokOF+hKNh+lV25f6iPWWX2Xz
4uMlAHOrassfZFd8Y0C5B5N2+422WZC7jhOpkP0aBbEXwBQc4LVGBwasm3rI8L869pCNLkVReIa9
c0rYQ9hvX4u8SkwqNRYEN3rP51fpBSzKEobawGijfNaqthygDp8/EsQpzIuU9fkpOxAlvTO3PYxM
KicPobyKc2i9CH7txUWQzRBF5NU3EUD6PgsIxyzk6xONx8exZN7nwt9EyrVva5phVZp81XX/PTki
J94pnlzhZ27gE041osZUGe5TaGLBUAZS6s38sqJNw5S+skcIKcj3SXm4wRQhFjLubb9B5jq93K52
qAYj+5/8azcf7Q9wyj7JuPBmBaZH0qHE3sBHbzQym3QAGgXFF7PtmHebj7FqEtACbFSYRrXSFJzu
+SSHCo5hhSKFiM0Q9K7bTXDUTMd9/LkHOHAHaa+OprtdSSCpVlzWTaAtUhhl6EYseeDSoygPtqMo
ktLzn4eOhh1X9hTl+uaRTGa+0dJ0oNZ0UI5aRSmaA9Jzth1ZYQFDw8ZKjGF55TL++BDZBtcrLu7+
djMEhmazeJNGO0LSYu1dGIKPtsAURTkQ5WlrMJb6W+0349t4k3n+EwIfjoWHsTNZ51lCnJ6WG7Ax
9S4YtrQm+dlx/QtnC4WoFjpOCDWm+N4XMS6x8TkmLnej4Jwx/DD6A4n7a+zqiz+m7QcrBtOf902w
rNptGfodC35KE0tkSVDX6dk8pK6chULjw4KAl0qGjas3VBOkPTZplpzyLn+Zt74GLWZPbYEkRZOj
05dHM2bb9bPKTLmDyzWOBEFzqqfjgpI4g8DNWwNco89bcBsJFqpb/zZNgBJ1TsXqIV4/PJUfOivl
EdGsUiO+Ajl7/8wag2qZMsXSiQYJU4oecvdaUD0+xelR7y6sgW7kJNEQr8VtOtCE8OI7vxUMzMNL
90Ho/PZlqrgguCRlXihfH1KRRHpF+vCGKb/TonOOje3TlOiWQmTDMq2Ij7HVQGnhKVxH350M8fKt
88e1eFpYY3tBDkEOBVwohBPGccs7QlVkB7p9T11nMQmeLVztac7z5QzJa7N58HkzncJLKFlSwDvK
CsqkJ7usMiTJZV0cASzsyUiHsd/FmlqQF49niBDW7m4SNo1LZm5HIlWdO0lHblC4oSz1KrVZPd9j
L0eflMs28crdEgEPpvc0LwwPVdiD+JU/df13pVeRjhdZmghk14a6CPmUmesLOoPdSF2nTd205pci
a708RUyqlFkL1PP5KGFiYLSV0woNlshBxsuvDwzprfBYZUyf7CtBEkd9eX8RIJwwlgnrinr7D4Fx
GaPOHkXUT2+AipQHrpBfBtj8PVsnC5iFlrACv6eCXv08Ss32dM21i9SQIR9TPFvWHCzuBe++WIT4
E6uoa8pBlA4eXNvJEAFkeV4i8ZzmeFy5bXZEz3KIMdfFldmG4QBqOStzmJlrlqsxz22rQRyrTmsV
rgm7vMF8zxABhDQubDHd8piFQB4EIZL3RHCfLnuPuKGXPiG+Fn7quQWsBXAzedEeaHZ7IEPSedZY
ABj0tivNVm5pjWS7mwkB5WNaRDXhFcTKBZS3S9kFVS/bTSnCFclxEHtkCIGCDDrAYKVn9Ql59Ei9
o5MBpVafpZV8IBIFp/U4Z3Us+nJWm4vwjvv9GiSewiqiIuPYj3ltcwIah6lCFg6Kp+YEvhOHuLr8
TFVwxBvUnrLwGQr3oHHPd8kWmJSKMvGftsBUZOVy91ehC1azZ09W0rjHjESJ2e7N0wayJCFZwVue
lKJQsHY4YrojBhnIfCHeqrU7bzLaL8UEB3J0n0c4zezRX+wtAIzHlPJTKBrYb5RSSQmkOdcvQOEz
9Aq551I3eqzqPyaJXqBq8WhrEzn5Ce21Q/dUfERQwk25t+QZLw7M3L9cFLqUNZ22IBzjW+vkXJms
Iin3K5mIdM2PQv829sSaxnNeBNPVq3Q8ojvUzIJt72eua7TIGER8yZUe5kIYbkg+yG6Xk5KbaZZ/
0VAQMLTJuLaxSTdrOqxB690B+oa7d/zFUiStOP41i/WtM1E5MkXDClW4XY+aNhQ0pbFqmm3mVy3T
siUC6UqgyiudOgBN1gL09TlRBh9E8PE1DdlEh41xfEZhOgifB3lFUL6QLhfPwpafs4NU9qR4D64o
G462cEuPqJ4UhlFkQEQ6kLbX7UKrFlGstuIWvlKRj1X5tHsh62Ma/trRxddHFZAxcNYHX5iC2ksy
/5/tptQ+0HQv0OgAwN3Qs5u5o+gdhjoeP71DapIoAjonPCYoM+BLI0sT3NvrNyQPPcmJC8QVLhvk
kFG5wVVmyK2E8IjmKgC7QNTxMUP9xbi8C4ArF/SnngXhwQWBwwMgcvbmVUAxV+FguV8BHspKOCRo
1hQXAQSy1Td33FCPVRnJ3rrd750ssxnPnw6egRR+Bzn46CEpJ2xlWADz2CQntSo/8/F+KdycOzti
XOaR8dQ4RKBJgOTt/Ahmsp4tS6kt7Wb9qE3EdOWkYskg766zDaP6fr88yUe/sRSw6ZRM3STFCfxV
cYJMXSe+ebDK+CiW0ovUmM+W4T3bOu9M5EZrpC0GiGTSRHAOzLODc0/dsqRcRWTJAF1zwYz1ncst
W+sS7AwJMCGp76v8+kWQKAIoePfhJn5n/JGVVkMZCQOfbp7fyK0Gw+c0839AGp9/ebKCdwqGKcz0
l6+KcAucSs2aceLTiX+62nn7GQlz0pclk1ixwrCU2FuKaoxPxrCEVwQ4G+AAu0Wu6MhALuUb3w/V
apUz1g1DdwcIifkcjU7D5mOUJZdlElCuW8At1usrtdKmCufybIT2UD3spzqYAqv9CSWvUJLWKb6a
sOnXAUGsj2qWC1BDW/9bpF7yEe1lzzjl6ZtD0DnMK0LkdtOJEEJ9XC0QADlcA2u1VIvtpnkcOMX3
gY4+lcVVqbYM5T8E8byYO4SQmUDL8WrUPlxiT/qHC/6sORiwCtTNLu32TRDSLKku9soQuYZr/E3E
VRsrKEMQeQjL+nrSoYsUzmoRB7PeG5aThh2DVwxwQteaPhUYow28DXPbDDJDsfyiY8fJgj/IplPT
uDbfCJlZPpCU1cXyorIiYz6wOLe95XnFRWI93TDTMHHIamuthhi8Li9jyM587oDhsFnRop24LTzb
qCjb9UP5C2Megd5OzzFvY78+UxfNy0FX+PdO+Ex1sXrSVskLjmoZELt7KFS+JRSEH/KdlPxf6eMD
Ecl214xotcu3YrF9/XNdWL3k6molgFQguBnigB9+lkGN6m07fw6mgFnEH1J5bzynjQC0ayHc53Cf
o5vdPyH7AO4kTc2HvqPdwcrJtqh/XHMWadBWdvURUBF+9BOS76kRqn4y1SuEBDRTG0CdKThieCiK
FbIyHlMFAajZsM3mlm60OjoAindSOaH87bX4JHU147vhpDWDxmbCn2L0L7oDzjIN6NxBELIy7qpN
QkdE4aCco54/RYemnV9e/b6Y7boW+h5TOiEo5naxzKVZkAqL5ad3zfXHuv227utRpcA045ji0KHV
irXFqgJzLBIUDE2552fpa8UqFYAVGmZ18YiriRO9/glbRk++69sDIdbBBxOP0dxV15Mw7BcgefLG
ibaZ0+v70VSmI7ElqM7ElYCqcHWuDAScadPF66/vvYgzQkH5AlAtyFCRnQCaPeqlGks4IEhjyKl2
P0tj9vbnhwr150s2Xrz7TW9WKRMkr0+dHVyg3XivBkOVpjeMb+77tCtOUq2Lsi5hZyN4CRbmhxx9
a1lOUD4bSMitTLEUpUR1XOkqROTrIhL9ldqV5pjYsyfLqzXlijrPfRfmQVGjBKL8c8zf+/PKXrIE
N+xh21eXQmW43CMc+QVgrwUCvA5Oabtl3YUXkujNYDxkmxyJnwqCEr9pTXgf7Wjxj7eCY6u4PZ+N
ZOtHHBTtFHYi7jjIX5TIPd2mXX0XkjTYxRd3HlrCN1hhjhKZvzWWEm4M2ZJsmtDE7/TGPcRUZU2E
WKN5NdS0zHHjfgHYXKRAsL8sHOF4MbVnS/C1Ssi0lqX5vLYxMLJc9Sdp8/4/Rx2nOFznqoYdR28+
vf8uOYhch+LC5p6eUhRkvIbJKwzE1YjN+L8IIKWjyWE/tn3qK4s64s69tQ0Ytduss3a2xj+lTyAb
LKtl7Yzbz/BZs4EisAsJIa8q2lGchf6RCZxQ6RxWGS1w4a4LyIyt/nEAvTIg96pZ6+SbhtgMClbT
PxzoHPvoe6Ti/3zX1GGhnMgfaYWMlk/JE1sSL6r5na6u5fDt98CuvtR2s8M6qS1i/kiKOr/BxtAO
trkEhiJnoXbwMT+dYDH7xJ7+OPzZBnHw88A5X2uCgDX7CdbOjE/MO3DvjphbUZ2tsAvBYCzd8eo1
roPyy7OR3ZtfEycbDoFwo3uIOix+C52pA2uN6j8vzFi2DwUTnJcGkz2Nh4LVmvtPCabhQ02cEKbm
jhDycG87rZIvV1gwmo2YHoLhlGTSsv9BUlKtip7aJR+OVyeDKUrMAXEFZZS5w3Rt7QmveHsAPKT2
50BZlJwZC12cx6PDlqtaKRr9/i14+1oCgPxipIAj1XmcovZ/FYCo140RU/ix2p3ju+IHU39tvnP/
wmh6ztGIWL3+hcbTgMRxanWRkhqVw/ZH1VDzOYK5ZnVrclsptsIz3zHxqbp4DY8SSE3Ei7S/ko2y
6+QDnw2990KEACp/EpeXOaEtUg6Kz2Lqh4hJOXPGm2/zUyxYDnO9ZwhymUUUHQoOrxUWfM+Q2mhD
91m6d7nCypiQQ+mD4E64vjfGMmB0aMoWOCCAJ1dWgzNLlDcrxyjt+RcYzQhKaq2q0IommO6Q/Lff
bqgyUWEVONphVZTkkz9nlHEdYDQdzHG6eVNrGaiyWU3/DQ0AgRcx3SszVa3+1BngZbbZemEoaXtM
Eo+zQtSZu00S8BgIB0nSenTptC+93U3LO7GIXJF4Vv+6BfrUke7vuIwO5pDdfGnu1WLpTPokEreW
DKZDVAap/AUzSPE0KtvjTo5QbgyTh6oIuClP2pZgsvvGgk6MEEe3S9pgh/NuHyS7KuNojOm0crvh
xj2Ls5eQSTJX7cZ5dviKkJxHHzLXnJ3uY74mMco+QIg+O63RkZPxoFbMZBtne+/0SEgv5YMfN/SF
KBMGo3v5MfuUJHckG2oywwOXaZJMnG7BkDN5cIcRf8c0tEGvbaTej7RL7VLQxmt3ScWtUvNSJVme
5IPSfDBMsECuWln+HAEatgBTAE6FSkDUGclSIoA2Nx9g02jWontSL6S+JiBAASB3R/AqMxzPsU+I
b7ZRBY2TI1EwmCma+GefohnpY/GRU7kZkwdCnC2/lpdEDBN4EzWGl6VT2nFVYeQMemVJsJBPiLnP
Tr5bPPlYtHQO71tWVmkNVaog5SRwVmiHOE+bZ7TIsf45UuQGzLrQOL17OYm6BjaL7Bwka9EE9DN8
CAA+vqp2yp6Zf9kYiaaPIljQhHir3pQJMRLK9hO7wRX/AncOKfJ5YOjZfN78FXMkSl1GKg8mV34I
TwvbdIiylhcHI/DM08BpYaIOmXAYiiA5ZdRaP4bNtm4f5r3Aijt+ufcjRVXzovc+otsDSQSLfvWu
TuSxlbi8jPke/7pXxX6rvWIHFkgZtJUghv0NQEAikFiS+94kxTlfBn4zSRurHK7kpSx5UEYhjYiQ
Jl5tXPTpAp8y4/hROwdUckcTLZJulcq7FU3obHmXpMfreY80X9DgUENAEea36dHVbzQ2YnTR0OZT
/7BXXnw/TJrPr5i1XmwPk5hCoSZ6QJeT3JIGVVv8QHT7bltYt2a5cOw/in7m8m24dTgiLHsjSglP
hDfaH+wzhuW/EqPQbYNoRKfkdTp9AmQYvYFPoNAb3/tE52LR0HEnl57FWvDL208TIsF+O4yVhXvc
VqghhVwquVGTxEteScEQ483Nq3URko0q9vKuUeWJA3bMMNT4PXljFhwv59M4cjG7bm2MgHcifREs
p6XCaRCKiHbLhpBE9EKKYc+bx7O1NGWOguaA91nmB04Gjc3ZZYt3bsysnBO/rxi7TtX4dqUb7C+Z
GiUzBsI3nlv8h+7t/dLa4Pm/Pt/UvRtjfKK4j9Izo3tyKWM2ao9zO09sIyh5B9Bi24VNzzwHAUNm
XRoO+RTvcDGInZ2BJW+TvnYx/PSq/T/mHPJGnsPQhyU3gH/oiwVWKLI7C971rswE1M43LSGfHRkF
hiIN5cvPWD1c/7MIDeWfUogSXFxXw2Ft79HfJeAd4HEGKAra+Gh27eG9kaVcWXEBYMziTRM2x9MA
9DpqSZFwUtuuZzj/CbKwVbiNlaHwLaEfPOvF3CK+wQigRIol1rLbTM6eoM+J74oOzaXxPwfufC81
z89YAQRS7whSqy+z0wjO8EdNZkp84NpWO1CfsTpVdSiHdWJCMiHlja6Dgl4cC2C9eEB9RYYIA48u
Zv9vGiJF07YF8UY+qE3kzaY+NW4ObXa5sllh/8j2EpnwG8OJN76DoCSRgYDaD3Yjd3x79BiWno+G
HjH0cnwzArez/4ev4NckjEauEzS56yuIQDMrmwlnrgf5IqjHOxl6ibsr3LKKGwJ45meHGN5LEm3q
SoKp6kmwHOdlOIgtZWsL2MdevxwDHgnfBrCqKqKfu7E2SFQKDm+BhwLJGtSK1bnIAo6cfjRL1etg
gxDTZKfBfTJ8QkoC5NGD7sReUhvRB1f9ZM59EH/J6AJjPv5JNpRj8AUjumWGbOuzeZjcSUgaik/b
gf+XivDGmFrsWvSorOYuX3ykB3Jb572hSz0wt9gjTzBRUhPnTwxqBm2malIXvy/1MiRfff3EkyMa
8bB2sMj0nhNC1uphoMJCbeEWu4L3yOHKsRgzUB58bpRVCVCF11ZqZnrhSXR7LMXg9T+rpnTvlTl6
5dZ+pFp04UZbL7H52V8ee+NXtEeXsWH/WIasLmYaJ9vHhXfQRBeFrHFfGi4za8jYbUArgJU7vo5W
tLKgRIbZfF4q7164RrViRXu7lvHXFk5czPudgpz3TODObZMGFstjOxcLq8Ik3QrGzrIcctBBfSv6
uV91hPY8HJ17iXLHHvvN4iDrTytY6S7aQu+U/kFiBh6APbmTg70Byhd4qo8OQY+iuVT4MzE95m9N
9AT0dc3SrWHskGDt3W+JjDNXCuiuWmkJlZjMzj4J49Oc7ORXtcSIRb3kChfXehTXEDx8iDQ9kpDp
CGzbzzGTAvLOTU1LdJOLa0pJB+dmlpkV3IqBiuNAJNSs60pZn58YCHRRLITlAw68hM3HgDyU8SZp
OKjPL582CguqKyxjWdv+iiYyyJk4RPty2KwQKQcxajxRsVmZduR0rC21JlkorF1lcizuUWByXhAC
fkubHrhkJQzch/FrH2xqDHqY4gFzJAWeU31/dFCQfsc/tyEmW/whT8R3RZugM+OL5HVa4sqqpsb6
Lmta4/id5ll6/DaAHj0+tnesLj2krnUapKLaXbH/vHUus2tNsUlQpegNhtOfS6CIsBh1Fd4JPy/N
w0GepUAkdayd2ZPcHMqwXnWN88TCLT3J7IX2pw5nyp6SwVjZeTkidZRUoubZnj2/xFS3wvFJQN7K
sdR8P2nRJDpWh6S/uTuxWN7oDR1I6kThejhRJaJcRbZYQgRzuiHeW1Q2EXygquAySHLSk2iLWODS
QaI+NLniy+71gQutsxtPFnhhMIhZHY8k5Uh5HE9t1W/Qdtb2jDmg5iWNVDHL0Ftx2o8qC5HoL8Mx
R2jhhZfI0CwqZX/6YT2I4sKzmbckp2DW4LLMZPtD+N59r/z6ic0fovy4XiXcX2dVIPBeV9TLaSSH
n8CYtgs1CvW7a2R9VzTDChhX8hNedDhnXHHlkzPPoaG8rc+ewP8fQCWVQLpry52XAQRFSSGJwiAx
l2Yc3z7jjCI0LzjuTAF/urug5PsyiMEZxDY0DQOZpKZndbMjAQuVxypYP9myjAhw+GPd6s3Qb/i7
gL4/d+uOryDN0zuie/6HMuWpBu2k8BanNCJSyxZF6oRQXK+4xizDTn+vi8gBC413vRkeyG6Tf2B7
Yl1yeWIRM8BWkHeX/iSaA/Xyhwszq3pvvJ0nkAf++w6lFjD3BYXi6eY/2Dv6g1Kow9xZDXVJoOH6
3ev0McxsiNYTSK3dECXKXKkGxL7NTlR+yza++iAWec/EyKYs4BO19Xtyk57+r7ac7/x4fGrobHla
x4uulXGTkrv3qflgA6L706r+8Cm4ZMpoGCwEabqiwwSAMoTlTZ/aAJZ+6zleGAMnY4uBxu3vz6W8
O+QkmboUK4oDlUnqIUUaZO5YoR0QG3s+8QgrYnSmz623KnJnhm/LkNnh4Uh8x4XpFlKIKjU/JNLU
Yr9cBRndAtAM7pcc87XFsJFkHBYkZminUqKwM+3aLYY0q+LDeUTsFjxwBtNMWJi9o7W6T0c7ZLQp
D62Bm3ZB1/n1++rQ08zIa2K4SMOBn0m2p/rYBVOJzASW9HY6XvUuHRwgEeK91yZG05BkdbeyYnFU
YUHI4dQoj3O1HOc0OROJ4b45+gUnTjL5s5iQcKGN8zTwkWOGELEcD+c7/sdRCtBHRAF9ZF0XTwei
+d+56xJmXZJScUjInGUi68pBgnvA83qCYrueA5m/wVwGCleIShQ3GypWJ+kbpi18hrvWGmtTGlSd
vMmx/F6686ekFreFLxOSx45/gm16orEg4xUKHFBNOjZYTv15pLT/qNvlrXYSHObAsj358kcbGG2+
3tbhdeS0mNqKZscQ1VgizXrpayGFvjkPXdyuPN0cbdYrNaeeSE3Sg5PFb84nvruNZ4PfauA8u8yg
x2YMpBuPZXD9Dza4t1nxse8MB7i1/CgR8QYtkCJnz6pG/mJOQ+/+lEvTfR+ysjWdVHKvYtnPuzrm
bDcQGjctvGCHCV9EYl93k8QHvvdU65cqi29UXL/nOClg5ZP566/NEgux/x1NNwvK9chVpfv2PfOC
8dGqIldIB8+/wGMRkDoNfIyg5/Ve6Z26paSWmYKmwMFR4iqI71OHlZ4WGf9KmQhXs7YTiZfXfVvw
u2lXDf1qdylC6Ya2rvWIkrdXb2BQRhWLq9dc2RIPbQzRq3MAavtTYqDrybBXosDBdPWGN0rTkiVT
DFeCxhgRm0tYJioAnDz3yOj1TuXnzdE0X7JgloTvO0GNkKMSyQ7G0X5GpaMEdN4Jt+kixReXuM16
U/XeqNxHF9qjQohh87r7NIdHVNu+zI8dF9UuWIO+1CcNAuWDUJaB9SYr/nvpxEnMwM9kgjtPZ8q+
/+VEX8GTBMCI5YtzcwcZ1xK6WzQZHCQIgSsXlRX3C5FKzQ4PNqBN9TtB47h7fmvS0aIuav5e2bTF
Mbum3QHWekS9V4F3ER+Nu0I4IwFwRrFngC4M9ri9NQKXtfGsTp2B6oXLqFz5iQgZs3m93ljEq0T5
WgmxOdYDO93wswfBD7V7rMXsjCmx1BBcSplFpqZme6EwqYgXFlpAO++sxumssqRXzyZ7wD0pQ+mv
pn2JpGsb92xLt1NOChdg7IVf5Z72OOnzMfr3JGrcVVB6LuaQUhe7Xlx3bc10+KHg+WpqzXnNIjwR
o0r+UsitG01/w4Z0F54PyP3ABuepWdgw5E3zouwPqdeCqv9BX8cJYs8ORoq9jVAoJuvh2VlHwjn0
v/FMfg06AlHMXhgJj9nNECP8na8SGv5H1TQJfDRSqZ7PuiYPLwjd7KelQhPy66UFfC+fji89IEVx
aMfq/8tjgl2pNospxMY49+rDQLtEbldwoZCzCp8X+Cs48Uo0GKJcUKaz4voIWSA1GQvMzehqxeQt
Kx0GB0qkKKQrLZ0FOo/wGTeU3LmbCckPD88jPlKhetmlYx+jNZWwgz6JRJSQdbTIWXLWbNiNUCQb
Z3fNwRFoP0FsUVOsKOj6hk7YM4tGIZcBAkoHiCII6JQMwc4St88tmtkuCDjApiA1AzrMLNpiHZ51
c0/5Jv3ynWTKlYm7YMFm1Mx04BZFqxdoU9j0xrZc49lrFraA4jOjZlOoIDRZn/wpCU4rOINKaimf
1H2PHXzYa8OWE4q5j/aAp0zQssblkjiFtq8MnJzWKo8B++CFNLo1EMHHGJyRStjOqBIZLFNzfDe6
sJArTNnTGi+XPApaWo/lxXGpFAQBxIkVzeIqNk2TyF8W9LtbQkeg6y5PCD5T8TkQ30Zh/3bwIVXT
nORCIDBtyPlrflMWcC+8SxoQ79xIc2xmuOV5HeKPTVfOI1NnMCjrPYNi7+2Opmeg49gw55yYOXZd
x0tUSBpaHf0uXgadJlfm3kZ8uAG+uL1yv/mi5YsnLCG9fNRjLo+bbtnIbtoTX37ujVaR9XCTO7/3
Zzax8QEXR3FsllIQ5ONjkxEh/xnYuJaRY6c/mVDiqZqB5SKKCvqUcIp8+DOEht3zVLJfxusZGJTI
vZdAQLFoIEQXbDdKSexjGA6TnJal6wjdqQ6VygrHKOOQtBk5toPSb1w/wpCiNXj4YKBYrmz7fxfk
7acNaixz5nV8A3P4rh0YuuuW/r6nmu0i9fLJZ2oP7Qn3nZCuhB9cmlGJtMfrIS4HAFgPKrdmeyLU
u/wqHLSTiniGOEKW0Ufbnmzfoi1z7Cl5sV9NuCeGZdtCA/UrJqHJTOZvzZHs/+81Bb7w65uxcZlM
G+ii6F02YfHIO0QAmdreeAh1ENICsTSrunY9r5HVWLzwqzBd+0AnIn3dN8JITNnK/L8T50VACw0O
53R2/n2QAOXWnIqbo2wnPMHN5GFgbhVQsv8PCYsAc+2qamtAqfmCXNJUNrXooMdKVdnsa9iMbx4c
zGzoc9K952yaq4KTJ2Kx0Qgb0X5qV7PCvyYE7AdSujMe0kOQlT516VohdnQH0ZOx/SrPZt1c8PoF
ejQxkWBqEdxsg+4KHQZE8gzSQgwTfdsYrTkdOwZBR9NVONX6D4sObmizL+CHZIIS6dAaTMWmXu9N
jm/9o/1ksPO1qzj3VyFQY69kebgheuxNraFdRfEvS6g9IsT91Zv7eAdybbQaG12qWM8KxO5rS1lS
00IlVsRxAaArYO9LERIQTsTe8igHZN5mMlzkMAqSzBPHiLFOtgsQopv5kwtKanRblel+11w9PdfX
vlcJsTxNYV9yJJ96sY0aJ/EYLnCfz2OgejdbM+5y7a2pW4uMNYOvolcd0CNBxXvBkf+Tdw4AM6jF
/bY6a4i4SCFWWOUTsVZckGlPDMhvcSpFCtt5mOilpEzMGobAJQkENl5em5ZDBxYGwU0yyR7knMT3
H652Rm5JnOAH13QciW7wes0h5q67csldw4Ifu6SpsrpSBjb8DEEp2IW3HGc24s5F410y4Gvcb3RI
d3Czm5uZTMwcsBEvZ4YUnk0LNG0/KrFjZMK+Kj2B1c0lcYYQtlsEIlyog92OK8v6pu1Uw5WEUTIx
pkHv1Iwgt3UjIG2/p/mCbrEW+mKUEe5ax1zsYsJorjYovtaoH7L68d3hxd57WNdLGgoyL1l8Np3c
MvKtEELXB9L0ddRJoAS65tg91viFlpe0vMBH8T8LHA1YI3ZJA7eA7diy8d43r6QSAxm/+k4fHKEo
p4RbZODJchhQH7p3R5aMAigbQDBMjC4knExSsgXrm9x/vRDFy9aayvxLD+761Hu/VvngaiL+OaZE
qV1SnmJzUzrgE9intkJFrR/R+KopdFDrQBrOnMXSc3KdBd6OpEJyenxYqB8eRFGobC45EW7h+w6I
9HiQgLGT1LxIq5kWc6IUgpelqxWVW3VPCiQeoNFQdJkRcCZ+zTO1EZXwxvOT1hcDJ3sezq/hLhQ0
ru91mKlt8yAcojRNMXgsgNAgEmM3/lMhUEQqZaeQKCVeWeu2hhJRVs0rUzVfpH7vsWeHxDguppDC
3dUfY6CDqlMVy/nI1F+i8hwuHm6LWdukei+TMPukV9TMkNcjOz+2NdNoHe3TxLCxyDaCXCd0E+gA
piURPpFjbdFoU05rEIoLYA==
`pragma protect end_protected
