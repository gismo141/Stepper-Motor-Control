// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
DGm9ALnw+3OP9WDCYkKDLXI0lEVAewMPuFGcO5pVaH2+0vkmabYFMzFaFE1Xfwub
wrMUtmnHQrI5DThC7rWyB/j7vU64nFjWcS5M4O2nVET5cXaC1NfwsvTArR6To6Hs
UTJdJoKsZRIALgNISi18P7BaXYKLX54gaZm74P8+3JU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 21552)
98+juKswMVdvXbcvRHL+4etmigk3G+BVoDAeDFeNqOqvXQQdMznG0i6DOg4CaF5O
KCx0sSIqE12RL7PeV428QrmlzpUj2L92Si4yXtBR7duNTINkgy+mrNJRxXoKiqVx
0FBJ0WHxf7NaKUGVZPkPjgcI92FnjJJWkGtrABVVCFNOfZbIwQGkP7U90Od5HOK0
VRpiaJKrBu6hZhzyf5Ux8yhD3CjcACmlzMpzyzebd3uy8txrPcGjWmNMkDUV6fsr
TCQ7s4PK561PJYnJ9tLQ7PTO+77GIfaIhf1IQKv7L0N/Slz6M6i9WCztwnLAatG9
OhO7wxfpQbcokExsqbS2pdBAeAFn9SxbZQWLI0TE97G/SDa10dXato+zHVk9sReF
gF4BL9g/tKOyblrAyWD2Vho9G7uc9RXeNvgT4+7tz90fPcGkknpwbgFCTBNT7up+
1Kh1LN5h7vocw3BG1jUXZrcr3D7vSPgQ8RPMzTXoKTcUYdb3hDJbgdzuA5A6XZ08
fr/xva8Cl/xi9hinoUXGQkmjJitksx6HYUoEXuzJVNxU8eDwvGLSwfjmulv0K/iO
Gu9uMpsUU1d3YhguZDJr2fs1Ml0qCPNE8qLnhJycHzBYSIgu5SyoIsoqmHUWh2Ca
/j+2qNimiz4oiSZgmN/q52dVrnUkZCcJZybYzQjMe8jHDrBHccaOZyc0GSTrd1Ns
VBdEECNSPP0Jc4pd40eBeMtRS7a5zcpZxkXVv4WAerSsHcFbqrkkZ8t17/66dxZg
An+HrPBi1/QWjvVix8HS0duVcJAkil36EmO5jQ5FfuUIkHIPbVA/fLKNyuUcvoD7
uuPB0BVf2qUkeWf+C7ru544j3kvzJ52PkS9HZZhvRa7itCJe6WVyoQFuFyynDVKY
MSLi2PQRvFpq8G4OfdZSXqD2phryyE/Rs3lHR2mRySyZTX/4mTK0mHi1oE06NSYx
3JBzQESTzkwzdqMq2Q42X2sPJgy/6LU+XXEo5OC8rjsfXdhbrXMlDjCVvJKrikPb
A9KzTf8oDVlw6IWTm5o+R+uNRH8xWUzqg0/16LTHH/yakeDZvqPdqyYlV0kvCgbb
Ggtme6SYLCIO4lc7UNSrpuekdpynhCeISFctt6cEv3uOKi5dTClFLtdoJqMPzJyL
1O1OPhDp21jP9/c2LaGxlwZzSQqy+pvtXDyASg23E9PxaqbxPNy7CJMgQt9xZqBg
I4owal9Su5+ricBq2xj26MyXF9UurRCYSfvQrdCWSuSRrTX9a80BkBSNOHdoelVN
TzR7WUy4xE34yvEZwmmZwkXEgsI+6prtqwedH96GP/8I/ZgU2+tpwjVmhOp3r9Sm
8Sv2X/+B1a7CS1C+Tj28Z8/Zu3hWnlSe4diTTGVNuj048GiqMIrshlrwC9cjXmv1
hMgkGOisvwTREfsRWIjVbmZIAe/vWImmdn/grqpldeFoIsAKrzYAkT71Zbt3VW+m
WlQHq0WddJWFvSNgySKpMo44p0vKQyQtV1S8cMMmcwcv7xpkIkmOuAOOIvpB6bw7
Qxu3orAP1zRJ6zW8/1nuPcw/Qlw9kGYa4w/+moq8nDhITI6DpZJAzU/TDHmDI7dt
hiwBD5a6ZhSy9dnlv68GZbPWCyOVfXsbe8tXNWmvAdI2lyPxZR++lSyV7KZAdkCs
GdmGJifDuiYVIaNw5ceWuCMqJWEAVguMAGwh6un5IFPazbU8b7/mGAZ6/+TSRmwa
sp6oBf8RvhKIgrX7UDSUIN9d9y1fek6juXCBnRw5Ns0lkb8u71HDvCU98HXaaLwI
/13Xz5UVh3pm+xD8zHdkSez9UlK1YzmCSl1WJDhaOjusDE2rrWB6O2BS8RGYGAz5
QQrPhEKcqkIlubo/kFn7/djbl393+Bpt7bB8G7q/WbcB2bDAXFZyfnYni+vpFxm6
hQMbzF/EfRQlAf5qVKTwYCrUHemBS+PIcDudF+DueJjgWWapSXZ6EO89iYArf8vj
N1lut7V/r2Lz27Owhngr0dlkakxh3k1DkfERdTvQC87fsRm+dEKzSUiHM3S19+9y
GcbNvHK713MpR1i64AOUJETlDtZL3LcnIbbqxf279hY1hiPb4maA7wp8Nicoy/8+
grY6EvaucVYBoFyEt8mLzuk1BCpChKZFj4en5xooWtFP9CiKaESlTLAvfe/qzph0
CVrZbGlGMDZvZ3seXGnUmcpRTIz6ksFLkazUs0iPHqyQJ5iWefOR3thsljdzifQd
Ugq20M+A/wGcLBFHmMxN/XULvigx6EmUJl1m0FX0uJuEE0JV/6H7cnuF2iNAmq58
sNsZn1Yo/j2f01IF3cSPoWoSakG9QLSd6eXTPUPI5uL6RgOJhmH89w8TFy6W5Gdo
qx4U18BoRXICbrcMhkkjYon4v7ydoxcAByLRFtfDj55ADxcJ2xfrG17qrRDpFrDw
ioyB+Vl9VuE9vZ25ig1Hxd3+IhISYJXX8B7lCExuNLKxot9EAgDra5/oknM8502J
1SJF7U0meeJPFT1vgncTkMO1iW1Xo+jJYhBP85ez/uAH4N6d+3/6KasSpqN0w2Ix
QUigspGFXgrgqE0KHQCIafrc84gyj34grPwxAG3hvJQ9MsspLTgJ5onv8TewWyqX
dsOLk+l+MUMYlW+rkDh36vTp4SE5ZfFTqkmj4eIFjhoqMAzsbLGgmiihg901aOO9
X3agSwLJmJ42xaIj2yA2UCJfQKlc2HW30WrP2i/XeqaPZf3objxLEbz9zU3tSuDL
nV5hAPW3FxuSbMQNzxjRz0WdVd6wjgb6lDHl6BkcCkcslub3+lSl9Os3EbxS9pRV
RbdV98tsbSXWxUUNIOQRWWMuZtFQKcaR2BjaxEth388ixYGz/UBdeNd9k8zd0Pps
1i2+v4OWf8L2ZEqeI4IyzJksqDyQ0l9gQCL7+bu2LfBXPLNFQu09rNkiYg2ZBelC
OXlmgPfCActBTKNfmMnU/ixeBr0vgZpl0X8E1Vbe03eXAzHXh7CNJvWHUA8ts+/F
UqFK4jdJkNh8kv7lBBBkaVIQBnXvfrwAtrFbD03+8V5Gt3UsMQmlpvERIijsiL9y
+YvCes/2IOwMIIP74PH7tkDgymm9N4B1sCT/Wb8OpGzx28ra5jjSCXCGNyU4orZw
ZfIRTHjmu9ALX4qSp4ZW1ScbMWlSZgMyg91tdSnAd1A4BPkn6cFlDT+Lob+YEt9/
vVOZJr2A+FEk9dsqoK2gKbrOCISBtbB8Kpi6Sivtd/Uj+NTlIfiIe3HZQGNDdGsZ
L7v/T8DH2Bs2OZY9HqKDtvmxV+kSqQAOyRGMN7x5aKq3ncmjOQeMjpKgdr35nAKm
VRKv7TbElWu/5C6ZB1M8uRDc5FHPebhUiqRiA+7BL694Ycy+LIksCqCv3QhTFabi
WG67ujqzsgKKZt8U7x9t6pL9LIHn8ZK3TOPCFMdUoiHvg4Jt9EmyfrMEYXCAyIBu
+j/37TN7kZZ3cjLA/U96fGXRzVtldoxRi4LcqpiUTkbk6ed1Rh21DmN+bpsgvama
NSb4vqlwefMCOEEdCZOUVGh2i/AF71lfywxPvyee8z75RJsGt2FglXu4jhaJjx7l
rIIBgsVIonUNOVKPb85eOmKD/1qCTs6L3/QXItKYyq5+0PfYq/dLbKoBJ9Kc1nUI
2NckMNJEBFIMSVwCJtlL9b+L1BuCX4mZAO49PcPoPzziG2UkUQ/3Cjh5HIoCCkGZ
669OMpYDRpe8DSR2TRvby382pSC5USTro9FM0YvGSICmNiaGt8ZVaXA6nKrNMgLE
rkiiVHU03Zyp6HQqEL4XzmdZcGxe9oJEEngDOwdyFjQmIGDyIFPDArxuz0g/X1Ad
cJREeg4T0eI/EywSUFgGMW1VM6wIklJcf9VjyJBzvkKzWbjTIajZHATHs+uu+1Nq
m+LUeEQZT3H0LKsXN60Ut4Hggd2IaFw+zoRvd3zDp7/G16LSuOAiapaY/VvDbugZ
B5y2NBCmP1ZLcaJYW5TcGiCSsTj+4nNKbpxn7kDj01fuBfISSMO0TbSvBFl3bH+Y
8s/4wDWzJ+aSC7IEC4ubWTh9IqORTICqBvzU7/B1GH10GoUvCnBxqT1emxdA21Eb
4bgHhiegYUa+VDOl7DJUXbB6iZZRXCmiZJkoydAimEPYyFQJWSQrSIiyicoxoNCN
rNKPx3GqJ/hASnMQsECOIr4hUs4Hkysw//4eJFdV71AnH9xalGKIzL+khsvYYZaO
w2X0ysR+Q/M6Z4BeyouF/mBPzSw9smsQFO77MVsWy3NSjwsa2l5McPsku1Ajfc6a
rvwMj7x8lfeVBafcHl7C1Bgeg0VK+EuyESvuKdETn6lintvmeEtIyUWSvZ91+oTh
cGFBtwBLwma3pYR9+DNH9oQaZJcMXvW48MnAg3j8Agi2xI73nYevYDeifUUOLgEn
0WJebxSmZsZBDUoAk7gieHpah6dASTRIaxL0zKd5CZlLPDeO8XvOrnRppU5fJeOi
DSaueb1S3XUlQ5phLPrtD9F2VQ8UNeYg225rmkag9l7rEWnHW34tUzsn8+53ov+7
DKGdB799xFGR3pbhMk65TuHKBoRHXOvT/SaluXlSbWivch89nRa10CiPK6W1lmFD
5SzUHMhyeoFCQGtm3zljI+IdXko7gpd4yTaZte0q18eOCb3tJrBHFjmIp0mFpjXE
WXVs6Y+y9lmrzI5HX3Xj6nonPsS5J4z4VRfAGLmA8la8PdhSk8klN78hayNpzJsd
uYC+mGjEKw0K8JCjxSPwZGR7FbI9roKe7s+hfgpMS42uSF6DsMzP7z/xYOUIN4DX
Vyhh35KPvxe0kqM3w5ms3YZ7NwgvKPi3tbeoTXSyRv+GHdwe0/NuA22qQHgcLOCV
xEljuxa/YI1rQ+1UUB2tv4Ngc1Cko0A3ZvM5B1GNd/FDszzNaG8DlZPTsllv2w9P
Fm4iTLgJNTsN5GHXMbaG6jXkZPtEL37sjlwuLyePT3zuuCu/zRZSCqFSW4nobjR+
fNPLglzoRgoRFXzV8UB2EDiR97yWXFgZsWqAf+PpgesfdAu90LyeKo2c1jOnT7SG
f38RKoTvx1NKhcDYEm8SzLC2G0WwEQ/pCyQJY9VYJ9BHkzj70poxpl08Cqwr0T79
7z+f8iKuWIBmR2JweNzpqAbjh3cJE2xgFr4sK2ARcYMWGK5Q4Dgm6LvKCREOExyd
XGtXG156K6hPdWVESd6SkYKf7XnlYHSVFpudPvyEaL++1RELiKKQNIfKxVgKkmDP
/Ak/ZZCR7t+1ew0DLr7mCjDhf/vikwR5BlST/a006Wqyd4UjmyJgu979P/XSh/rm
+5KnA7grggxB9+bnekpW8Nmuya/S3tLwKaKQ9GH+dG6hcSS2QJY0sinxrQErtHGr
Hso68WZ8y3febjVrrGuVvpcLsBY9q+2nJV0eDcqWhokxeMDfadrJmbveRAQclty/
feudeB/Zx/18O0j/+DptyLRdwb5XnU6H1jn7lYePh85p7K5z+gBiAviXbM9M+M6y
tpwYFcRzRnKOlzk30ij+7vi6DtmV9H43pQF/d5PP76WXkKFr84XqTnIgnGjG/rhf
HiK7zYru/2LHa3SwmMi6Kw1fgAnkbI0+YBd7DcaeE7K1rpCNWnJUZ8tBr1BF1ACi
XVmmDHL9m3GwS6Pxzkb+MBTSwZtQddCZi91HFIYmN5RdQ/dBRGNZQiTbbX1doG2/
UcybqsLhcWiDaJrxhAmkhT9BtnqG3w8mhKSeXmbZp3RETxQquk9KKER/xiFZ5Kwr
zEVVnbhAeMy2rztQCki/GRNcpsnf1bJWjxV1nkXkVQaHUf8UYRgyqEoIOFr3wh35
IChdcdeocoaSgfhS4QjhL1uRk7QsKPz+c70yzblgSHTGzG4XfJ2bRkaEqRW7ukgv
YzIXCl/4jWbQY4hQaPSnlEXRsDF1QzqGdpwhzh//9ENQVBPGF+IqUszURl3OBEbX
4/7oJkbVnyD04Z9d8kO6ldaBl9HJy20SVbVy5lL809sYZRWkzXHbpKw2PRc1cxUY
imzs7KmMYB5wru3V02/vVLBuWXJ99fYcemf76ZsMnKmpDl9+5WdrJ/avmLdA/cVH
mwz3gBDJ6XXmJRoNRvQeUrvfThMasJ3ZFFUi6iydt31G1DVjiGXNi3hZjOHDVVQE
8LUjoC4/mgXYiIt1J/NlC3f/jQRPdzQK1Pt+/5vKyFHwNDRi7FWFHf54mfRcm/1s
+9RuzGEwnVtiENB0HzRcjgZmINLFNBOAgBcf+Ht4jRdzzHCgM0TasqZvpM6d8QQo
Z5A35RN6N9611tXQP6E/PNShkDvcsMl8lCk2m4K6GuZlNvnaOuuysYLWqCYFgfns
O0j4pT2oi1+tyCA0VUs+e8VXlxE3pAU3G8eOGSvoNscrIZlCXqswwzuGG+zU5fTP
KfkzdMzW2/oblOcMIeUSZ4207iT5H1TnvBpbhvnVjVuwc312yqSAkNufsf389kp2
brFOaZKpFa+tiliozFb0xzOblD6ltQO1kqmnqIn5li8NYGXkZp+TWN1iKLVJVs6t
yA70LN7eAD6vcvyxjF0GYyopVhVcDIG1oAIpJhGxp/Zcbf51i75aQ4TLieYiq9CS
BgBJFvTWSpk+wv06kng8Ia4osuTvNqvVcDy/gqG1KO4G0XxkW4J2zxigkfeRxx06
n0wqiiIqzw6GkWAlHD9OFV/mXwr94Z3eBKkpdxfR4UDOyoEpxkU4CdwM5gpBXEWF
ZiFDzFLUK9Ws3Sq5AsDRJjpmdZK7eKNWHNa8H6rXql3ZgWJqB0T4vuwepmPLyhnT
ITZn8wVP6hBq7Bmtc9eUEh4rlt0s8iniZZ90tNIMzSPrEDshnZfE/unneYGWvpre
i+//RVeigehObiHNUZg4dvobWc0IKIqDzg2wKAM/qAArofNe1mT2KNXLJ02LqUhb
3YN2diyjJXe8Ga0gEAMCvdO06zxPNmjGN72IHtqnhB/RsDTBkltlkP/MiHEQDsMi
p0Z+HHxe7NMPoDJyKrILrElfloUQ660k/jojSOf5v7ApiLAX0SeBxKcOB9DrIsBN
IqJQfgNlXlwk3S90EFPoUaMXzxKnh+CHbqiIs/edoz4Q3GyW3PS2Zvh6/FD613XP
VV1ugouwxw3HzoSfzlzNduGn/mIZvp4t7sZJ0ga1FB6oCXhtGR896hrvquG+L2nn
ZDIJk1aXzvl5HRbVdMEPCQAOKnZd65HVBDjHbJ4onNeHBgFeF1dxOTOj9NXCnlea
262kd0hFjX15Gg5gbXF8vGK5m4pG6AsSBOSKzPziyq2fmimFYyqtQCbzw0H5yj8y
5G8IW26n9TIusANq8IeYyqDDGD3HbC6kuQFYjAFJim4NxFa24NLgXtkfRDgBJP/5
18B+sMDHuPUdaGZElJZjak3eWWnnMRtryq0vUepYdrpf4kZoqcCEdBRggtNXssaV
OjOmPvzKIbqGa2qLsq25fa14i542/HWDG4dxoJebrsBn9U3kth5+jrf5f2vHmLvK
EHFjxAYsTDBgVAmc4hj1YWKj5//WYEHTNt2Cg6HALV14mRPseUqH5IGehHooQMVr
j0kvzKlCa9JhHAlnkjaoJF4Nd1xDeDBhEy+lJfYVjSMC+Nh/154YgkZs7BkfamVc
AlfY57bLU0gap+YFNU9aV4P5VmYTZY/bSiCEWciKgCLCgj2diKv9hTw5ekQaHiqG
JrQ8PcjzKj7BXZ3rGqL5ZdKYkyqqQrNILfBe6UyVFLJlATbUEjCvhR6SL8wMfBBG
V/5JaRByeXKij5Wue2YIWQ9IuWdrls8IBPeJinbwNcX+/QmGGRi3PYmOlJ9py9IK
ZbWnkvvZDmq9oIGfOlPPpfOVUb6FMxiyswYgWr09Z4yz4OF6UqQLxmEylqb/tHWf
hHGZX4astQ6F/4jPko2UnhWbmJgAjQfZ0nha4nSJOTfAmZhw8maWhhuxy3MvKP9u
d4Nh8AcHKdyS3je1vR4BzNS9sFcXM2mXgaWR7eWvzd+iaCfd9FkE6wbTUqSF8OVR
Z2SB/r9dC+KEiJYOjokSPXOX5BsldobhBIpYe4QMmxUeCltCggB/Rtiy5XI4eKDb
Z9WZ9H2MSRHLVl0TYdhKwRizKOH2qzLVZ8lCruGRImlrJAsSWeu23CU3KwdG4voH
pHrM/OytDUrWg7s2RMNhLEdCzxF2Jf9BdTZgCn/uV5q2NzX/433t4Z2ge8R6Ap2j
cQIPWQHG0T8CDRj1nfsbglKieSRmqu024uct5vxwkxk7SXFlXszXylGdd7MQXOmj
JXdc0KQ5N1IihFy/CfNzhuWVeJIyCLQgsVoEqb375Wg4DBvZdYyUOTZYgIMBNErA
eUg0ZcoBJk1xt90G4a3Xht6S0guaaDa3Nu+JnyMMy+IltvG4UcqKbH6oywZsMpRE
xbU1e6G0AT2jCcqZAn4z+eZNrtavyPyXsap4UfMlN/r/KMxeQ1XjSOLZQxZtJ0Fj
xT7G0Y+LWHK4EZtmAO7ZQHcfvbGHvHexffaxEvRzvshDj3ZCKCp172EL4XIqheTB
p7KoRJetHbAc5uIQ4owi9S1YQyLAlrjWcgS95UlFhHVqPhtVK6sgwIOpWKyfajUU
niZlPeEqRAERqsIVK9qfHGBleBRlht5ApbTv6dOzpvcXPXwf3rZriOOryTeHVIjQ
wGrBq+DnRXgAMrKi5m69XSJtQG7ltiQ1EzTCxsIwVWsuzDERanI5LRzYPg5IjI1c
voJuZywbMIafve97e6Lldd0KObB7QGYHtic+i0Oo7BeuE/pMdGCh99MsTWWkVm7q
0pTrdinaTT/hGFwfq1ceNCcK6oGYl16dnQd4uVKpqY0Avrfmxp2URMLkrNlrPnIs
dX4In0/sBqR5r5uVd9J3KwwQOYz+ocz+bZ3JPJ9/CRdektQAFJZ6u3ZkjuDSo29D
RoJ6xCQvAFF4zf0weAhCXts3KI8G8gv9vaJfONobwqFsCvzyLCoJKGQNMIqPsUxo
Ti6DeuAVYCFW0uJOHzHw26652YfofG3NxT6RQMC7vSnMHLKJmg+C73r1LcmCt73o
fQ/cIbzSzHb3oIl96ko5qC0d2lh3LWsXiDNQ1vyxYb3RQZnlRnzJIeNv5QlQu/Rm
lRAFY4Rr77jpddh97yNTOfOBBIYkFA3h2nk+f/V2m2SM0wl8PaUzT9ndi+D1Rg/X
W+jgGM90jvwtN/dF86IVrQrop99CfP4w4DYNyIAZWNRxVLErL0i0jWWqzbxg0wUw
x08oh6oTbTlKCWA7s6LLJXNgs6rY5zhXfYWMSTN9UMpKN2byuG4KiGq8HdGgVyMC
F0yYnl9ldkm5tnTgfdB40uWZ3BaDk5aVqzbJUGbDKTx5lNaJ+AsGhTgRsgI3Hbw1
vQRquo2R76zALLebQ2TPqCAALHeHemd/TufmvRpTRbJxRHo2f4Cs3FmggdDOTzPL
jFfI4XDK85Fqpw3dZ7+s7iAX44crbqJxpaHHeFxdtF721M6kI/97j6ljzE+bnGhy
EPsAYN/ZYr/j5hE4G4p4CFkeVq40eSNVJ/p4gBVMjp8SYYB6ktXvTh9nDKEfqg1p
7nISdbtscBDNSdpOtKfeiQP2EqZjjH2gQaiLUwcAq2V43uGkHAlx8KPr/MEh5nMs
RFRDK91RwSsu/Xbe7HwURBAhmTFAOaZO26j7+63JCj8oWJN3AGgMcWFus00XyTrN
jYU9LyCLfpbbWrKe7UqLDGbhDx38SpF2oiecBLgSvpB6X1WFHXlqwdv1Q093v9/N
OezMy6xTbq3tJrg2bCfuzM+WNXE66jW2GI6lBRpMa2TcCpmUmHFCt7MZNPPEoOjt
KIQ67/FQgtBTZvwLQ/QxTh3Q3EQnYksSyMcDLdzO91BuscmwvdOJN/r3cNAKVzBV
N6T628he+IqLayMBV1HLs6h6bh9Tjf6Xozt2hkEFqZZgyXUQg5+V8pNeq+IlFc9N
wsZDOlO2FxoybqG4IhBOCWV9OkbGTbFH4PbjdQjesKXFuErOyBoGW+kvmYknf6kT
L3l9uWIF2opOhmhMKSAkgoL/gI0U3HrrBwTfjEuJAZvQDrfgclB6CVWzsYBFXXFo
/BSHYESKe/9XaIO3d98qsp1ShomwsRxDxPkyh12b3hZ0aBrIvfGvioGdKy02+FVT
cFEhfU3jNsOgzeJrykaIOJDxGbV9Q5JK0OP2v2qwKt+zHYMIZxgA1mNXVoOMB/H7
3R6vS2UvOgo2moHOnf+zBAxngSfrAdS7wrtk4ZVd9uoIw817TWtwGm1ROAA4Esh0
6LjIFJQ9Fcxf3p9aTqskBtKc0BwNWgPoj/Vo4BeU+MrO8dYFikW9CcoahPSsEaoS
ZPTSBnySW5CaZRR1dW26kJe6CmEvu2yj7/qxxiavOppbWXCCH9Z1wJw4mDPXTCCp
kIJgBYa/JhchIfSkYc+AK57iLaSqRWvt3UT7Ld6NAFXr+xeugcrc+3FQ5nfb6QNo
5TKv0RnpB6JhsuWwddihqJpmdN9NSAIDGnnALTc/wEtIyPX64Aor9Rso4r03MwTi
HZTqTXzZHg6njFXHSZa3K9/IE8aUMwWnsEPardBT2YIGTBFQSQa7cXS0Pcfg3KsB
MjffWM9lhbHxhL/Ih+bE+QeFp8Z1fcMRFh+7/wbnbCrAWLaK0Wm8k1qA/tOYH1I6
NxjxQXA86utviUx/goPuHzCNDWVhZXeKi64qm3fVCRqKLxoyaQ6sraIqY+yDLVQ7
zcmU1rVTb8t3gLMxe0sD9Eouw3U3vIhRA3BKXok23JxpTYbyVHoGFr+AZ5p0nUab
h258WhNu9EF8wCji8fIm3OfT6ARZhTf4PGHiZ3l18Xuybiad4kvPJcYirrg0La8d
b/FziaFKWD4Y5VvPkDVrhWzqMa8Yq1L+7HV0nymKQRnGmIUwtmmGm7SXpkDsZKb1
+07Sf1IzY9BfoCALfU7VpXReBGnbZ9+EWs0HaUv+4YUNmSNm+xDCS4xDUqsfC6aq
uE0Iebgb77yrIqC8yhIxy3yPUGnEkecOLn/4GLmfL9LLuDEWcAZXgWcYOYVfGtfg
kjMqW65QL7QgpGvlWIbKkxIsyNBoh/x2KAmtsII55yF4BnAdQHy3ySJgqTn803xp
ecTWe4v1hl4+EIPvZRmihyELv0QenY1Hjl+JkCXCr3uTaAPFS7I21mVMTQbk80kO
e6VIyu3on6UXOleEZ3WVdDikPpDZi/PFYdLGp5O/7Q9kFUBJa/u5R0FXI0BP9XyR
DWm/Hl1/MiZ/Y9FDo6jvX8pdKq781kRC6SecLsljoPNfGwW+7/+YuArQKodpNVOG
1cWaBeNXCD6DBwo9lZmX1WvYTRDcp0hBnw9qz8Oeo7GRMFQN3q2z5OGhz3FFbbZe
jxfkDAfeuSNtNos62EcgfLc/ZqPUYtzY2RC57nM/Pe+dKgciVu1bvZzSIbNy+sWe
BeeRiVQ54fxbRueJXBk6VJ83Bol9UB7RgwG8VaRzQ292WulM2Mj/0Gm8Y/8sLkaY
quFptnWqAkBNiYnb4b9BmUNBN9Cv4efDljYOqXTE2lOgma/a2kZw3mYRDcXpH7ll
0X839vZCsKs2JBg7IFgWWg2YgbA/cQWiyD925YgsCCgwzU1GAWl5U8hSMPRxE4g8
Bwy6yNdJPl3DNiQJBKbS4fuLAA4yBOKhkmAmA1WTQ7Yfd4exVHHO3QgPU91vAc3j
R0UWcm4agfu+rMq2fy/BcjgCkG50+92veDqAStfDNy4MoIfLsZjDmYHc0cU/mQiC
Q2hsjgdt1OjVcQVYH5ffmnEMXbxafjUWnI2q3/1Z73e63yXxYDFOEwgHwhNWkKii
mc4Q5evGUpt5frhRTdxDUqP6rUNallfkJGmKxTsX+Pie5UdJ4V5s+Mg5DY4W+QD2
iMzHsnJ1y8pp0XvF34PmXOnV9RwZNUwk48da7SVMXC7ooe5SMIdE/6GnQ4spbbMD
q1v6vAxGUnwDiEbAYTFr44IgQTvg6v2nI2LrJs0dtWgb+l+jp89BhVPDoxQh9q0d
4Ydwm0CvotMkCRLXeXBQLZOhQMO/iT3nI6vNk1NBhVqW4LQWhhMD0hYGsXF+LCc2
IHB7pAe/k2ZRXxihuPm5kCYwQrBeEkqIxq6rM0DZMfMovREwhdfUBiFUo8BANEYJ
UlZpLXIS1qTnwmcU3Br3DLoP+HTn+kIg5Z7VFrW9ZnTZJk1/D5P3bpxB9ouTXi6R
LUdb2OIhGGlH9WyGjRJNwUr+sLkMG417XoRrWJKIv8Jev5U1n4H/3r0ln6fx95cA
gXl8BMlJbjUvtrlMqth+MfvZ4ItVEeWNnyN3VtJ07fW8wiHJvugdzWg8d7TimJmb
2Hi8sp4XXavycI5Zw5XQre4B7zxqY0nvI10Ux7kwZjj830t550cAxdWdGXlY6TvO
+ACbdV4dyu9dCa+1V2D7KLAWlp7Rma13rq1ZhQzXHSYliUWgd+iikTzczGP5LmNI
V0lG5D+P4c7j1Jp4cg+rcwJOzLymv85BNvdV7a/2jnqmdAIemFd3ZaJ0m3uTgtz1
VR4FlKTQU7czPqmd0TGDppH+tBBpYhMUt00Ad+fNI3nx8VGn/IoKy1x/ed1H0YSJ
hi/HpcVlVJEKVGMvGh1DMBMAH8SRa9yoa3nOI31XwihHGTH0jYv02NOlqClNOth0
vlk0Hqd/rOLcLODIx7W5mprIRjRFc0oGWzvbCugxBWU0CR1ByM1/BfU5gQPBpbbs
Sb4AYsuDzvqYy6dOMH3JkjKRGR2FKbntSGihFncvU9aAqOpTbogZVhjqgjUrTtxi
5RY8Cr+wtQlJz9cSpOYmEQ4LbM3hDrSG48z+0jquVHRS9s8Nk+JHdeC6CostWx2h
cBEDYL50Zhx6/C6iR57zqDS8mTEBBp4YakBCopKOjLRZ7BxtPByLHx3yCnq/0LU5
waCRsABVolHGDPZzEHD6dJLjpxoruxp0ORTxTYYyVPnd8H00azjZYlDn1om7r40V
CL0+SmvlgALLcrkR3c2NJqYcjYy4llRTvRESgB0Ukx1XxQ+GlQd2B7S2FoRWfm1n
jGu7s02n+p3Fps0VuULFBgd50TX2y7mMc8iE86DPTHi7Q+2oaBsxcPChQzbTnn2N
mMKehKxopXCIZQcd3yKwXILL0qj6XaCoG6T7UYtrHbN67Kw1VUtB99pTzCuY9Kk2
BtLZGgDBgN41GooS8CRk5viMRC0KEQaI025kXFwDT4udmg/NqLUynAzIq0SdE46/
XsuZV+j7BF39KsyPkcK+XhXKND4an6/9jnPtzv5n77eUckcZ2YIEo6I8n4p3zDRb
dMFP5jWSOqRCUJvfEDRZgi1w6JxSgWKZgFk0q95H3/HR7+GpsahFLYVGb9xzcfCz
RMdCVmovsiN7XhHrfQJdmFqbR8MKDPrdIvNw+m5jMh/KNwzI+KrUQIkUpzBi3r21
2JP1Oozucx0Nlo9OE2E9wWHx1sGywVCZfEBIPGXvlwK5T/HYweB1u4hQ2NLIt4Th
H7gnhjVVxyhOI5JDpPXYx6ubSiCeiWJKigNORDRS2jvjxt7X0NcUN+AuWHkl28vn
R/sl7hyf5DXFQPsHc/PQWo7mPd6pPkiwnbRaiG3UT3Ga9LuQE1Etkpxc8FNuXqlF
da/6z1ZvXJK4jNb/LPr8wxDH8+7iyXasOE8pevX/7s8N3mVvEIU9PG4kPeAhdEIO
QDotaKJJV3T9aChT147zpOLa1DaSqT2t9i2OAf9O3sPpvI20LsWgpv+1YYCEUh7A
KdmRvYTjzbIz4ZxJwKF5ZFaHl5Sa6Fz/7RSzJXQs7gTMalEJuKAhrKKjDAS/MAsj
PWLedEucKRkYG9QvBc64WpolSGNQLCH+QBU0+RZQGrj722Xx6TNe2Uc0apj1NNkY
W88SDFGyPYOuRMQuMtydAdhjyZsB8gVa0TfB8kbsdsDX+U03eyjpoMdAp6YdJ6pS
u849+BlNJqs6Xv/PSJffwEUobFTyEqLJfQ067GvLVeGCr+QtoZ/bha/rNJRzwner
nLY6nGWBp6yMdVVSz+9wiFOBNYPqhlpGG/N737ucdlliEaSqhIi6r3nzSnQVaTF8
46nfyzS/7ISWsZy+RCmeocezptDfBJN+2jec4tZ4uqajN7srdUMHHC9fJ5aSSEyZ
FEA6+pRdLvVE25SDrOAQiJ6KFrcWQ2fMf4p4hhIzoXwRb6dbLiRj6pnTVUeSen7u
RbRWl+VhJTlMaCq8H1fWkMwbv2dfVtL84YrbHga6RAh0B2zSglz5SYiJSD8nijTH
+9lQn7S3GTfmTL/uFKRFR7j7ncM6CJSJ0VXoad3AwMfFY7UmWswxD2iJVi21FtAt
LgZgZ/ujDNC2OIQF6sH3DUYBqg+Aj6nYxXqVPMOQXAH2bLgTOSUbPm8noNjJR5Ku
IhTV4vltPwMDt5zkr3OroFkVMW3SmSS/jR+1dAqPvHbzhDOej1m4xtbPW2h2LgYb
TuP8+8n4g5V9kITHP9fIWCu3gGeSQJaROXVj2qD3Dg/g8a4U2Ysrl4j9pv64CZFR
rbycvOQTEdCymmq/E1az5vtX7tLItVeauv1w3mig7qecDdkF/m0h1HKn7ZFWGb0M
ccAoLp6YAS9tkjHSCVHoUe/3NqPD8C0Q6rHIy0I9bT4fBLXrvPCTXPr6Ac/tjAOV
9H3I4WGNxe+Dt9kQQ1ZhNocmbuhWG7yyPEiJSBTQ9zdIC17LF1nqOoiQNCLKjxEK
aXohI58qCpN1sner8tWaRBSo8+7qk48znQhkx7jpC60jZNwuxngxU0oBTW85589o
7oV7ZIhzwHN7FEVnb6tDciiipsPyZIrUt2UO5GuKMLvSnKwuMrH2DjPyuT4npseD
Zgd23ZroMjv2Oudeir6WZCPzys1rV9w+QhsDtxo05MtBb9XbaHYU7EZw0VhUNpev
H92OVkVTLZDZJfk474K7BERGAuoQBRxXxzTPkMw7lTltg6htJt57doDz25ILqkQy
obhgAOd183GxX0zvs7hmsi4sAg67tcILsQzlX6wiZ6VQQ6jGaP88AqeKYYFzKhdc
C14NRGzf455PUm7HHS9jT2txtYYbljKXia/feLcRtvzQPOY51Ehzb9QKkpMijXdw
9mxjQfYCBbpAviC9Ze81fiHfzq1Q2MaswXhC/P4lZ02RSjbCBTXeUnYr/LrUiYyR
E8UQZse9bfi/6FFjtRfvy9Fpo6wQlBpmCWLXXxhEnRGsBN6wrO7LeeV1AaHgcfH7
ufvHlK8/yDqpmGo1UMVYyR76fmejtcbtH9Tyjc72e2Kg3FFZepkWTcGH4Bct3okI
YbmehdpGtCsFMLi/hjY5ErmmDkXhxv6zcq0i4IhaSAke4BuhnAIYrQOhU7i4Z5yw
JOmj1Psf7JO9UJ1y/vOmMx7tE/9VDJpuNKSt98Bz13q6bNFK79DRFWJzIkymXFKG
3Z4GDEsKHfV6zd1RRZSSFv865/V6czAxNqpUkZ+4+6XfT5V2o7ExIOzwir5/SsXQ
LxHpqJe6F6L9Eu1Lm9yIPyifRHur5HPKLBaxVHygU5Yu7BS1QGDriVlnugBTecS6
w1uDwS/0kYEctZtdYkX/PeX9kEZNd5MhcynyNqY/NKfjqd8HLChSUkuF7H6VJCqR
pEtHqrDUwivcpahPC6JyebDALDODjYQahlF5o9Cuvajcs95mQwD31WzmtquhRSja
XXL4GBAO5SlxdY2iPaS4MQZhrv1+64hfRHBqNi9VUgXXB52ss65RtBxaPPFQs9GU
seU7R4E2i32vYK2SD+GYZP1L5kOIv6P/lpjAyPynRsUaQcuEivplusE6vcRkZAwN
S0bM1rk+fXe67l1H1FoOkOiqLzoy0bQvdv/03dGzHcw8yYHoDrxy0Ej7x+cAE6Sz
05m2lk4UBalb0ES23F7/8TkGoYzW1cVxYUBiNp0p4dwXwLlLRk510usHNacWTn8q
ZPb58Cr5MaMzcoMCteR8WrY7/GTDcl+kwkmxcPVkA3wYYgRY9S+Dtw+jH2O2gY84
+vT8Whj2icZYb13tShPwiWGO0Pbz3ZQQ2KpZzE0gHA7wOJ1NiA8hRT0wdAZHbpIF
x1OXlFUotZzMQ+QZLb216+0T195RtLVoLhes0HSsBRp6U334Fvtkprz/IUkNirzW
kvBnQdS7OctIcfITBVp06LFyPk/DSoNYjdDkBeikfXxtJs/vqDdwIJCFFAunlGnA
ZAq5SWG2gSQvhDnICDTCOFp3vt/uxZzLYSY/6bFg3MDELqQNGT4uSNYiz/ppC+tL
B38/tTJWAXM8SA/GDGL0jg3AloDocOKiCk0r10CDwI0Ho/6BZfKKx3NK61p84eSV
Z/wjG+0+uGLxMg0ePI/0Rf7NI8FljfJFQMP7VxM30KMZlqu46BE9G9mNV5a4PmkU
bb1hpWEQvi+xPNOXQtv5uJroRuNS5xVWO6J0wz7AeYGBHQ+s8XgHnuXedrMsP3cl
KeO+0CkjR+oAFxKdkXbDPVBdkjoGBaF+gNPnH9HnD5A02YTOmc73j+x2dAxsMMcM
sgCs5wEC2PxeWtdx/8hzeZN0o7uIap3RjmqUdGvo3ps71BjYO8a1/l9B2CZYusKs
sgSIDse4lr/Ybx3Kcb6r/9dppt9VFIurcv7yS4VPEqq9CAaNEU+tsdRunTlWQzt8
jvPXxqK+DPjcslu3H+Gk/FzbY9GZEq0otTWFc7y8qlQbYoY0X4SjWpPNQlbCUmbV
oSR43idwYCJn6OLVNq+YetoPojRmMCb1exbH260+XeR423wSo/c4eWBmxIo7q0Qf
9U6bqAJbVgKmk3OxDFBUhjFW9jFqVy3ch+9xEvKfHid3KMvKFFo0lgPSpm2pyByV
73ubRjUWgKnrXeiseKaBwRssryzHlcrda2za+ObsyUXI7wiVyJ97WOEYMQ4nysor
L81DLnUm9bISvbpttKlhCbkEhptDRp2PLnpG8KlzPTnv0cyoT+lF/q0LA2ZxjM03
PzZNP+ax+98KwBGSVU6LKCG45gXQ7+oZ5geZxG5IKrSWqqTYGj99s6UItUXxxlRO
IUgHtx3WqKkYj2l/HrnAUOnlHz5yYhK/zOegsE759JG6DUtrb8eHcakfH6biOZi9
buj0yeoHl2vdHK7ir3lcIjzk76VI0tJ0hIqmL0eXBwQEfXaHfAPqEBuwDYZx6+HP
Xser6l3Qp3nHCsM8fJ7k4/vHnZH/rhi+qvvCQ6vlQfMUhiqMtiLgTjCNxEXnTGlP
JQaZvvBmTn0wSb9yKjvhGxeKhSiAR5oEzvEerDfF6CqvykF7AQ1KQCvkBzNuQWM4
v3pJiWNx+Uwy0U3yUBIBgIaBclX/PniTvh3SDFiBnyt3QPTnRGW6fWuaZ8xX2OEW
9Ir4PAkK0onhsOQNFSh96/KGT3Jtx9NxDf2AltWvO7/8MFIrvBft0S7A0w0VSgmR
na0eZgUXGvuCtqH55f85WMQHgx2ZjLBwWuMYFct19ELl0RNtqDn1sUgah6uXCNuL
NgBk1S4IC+1NFdnSFVOHoEoJQW1kKYcLRSxOLQZqZisdwVsNl4flFcsLeCfgcIl3
vejiMxVSSCq7qj7TG1eq84/jOcdrcw5h75/C8WKyyYW6Rq2Bp8KjDWS0YxYuJcYB
oOw0jpLP3pYnKsjQ5etPjy90VDfxr2KRWOniXF5sbLkf7eZ96wNK+o52lYA6spZx
evFABrrDRHmhOvDGcwxXVIntdSf04NnQhKvH0rp1rJI+DQnX7h/uR4WKqCs7EsW/
hGLTnYh5dBjEaRHjtJ4zuOdFXbHDuVNqVkPmSAZIhmoMEX88BOQnvesFwEXie+jj
d3WmBpckE2N7lwRheklt7PU0gpMblrktckzLEMtoLHFS7rIvmCbS3S+pGToNtDzz
g46DdN+u2aAaovxVNTIZZ9LURm779VpC29tPznDYJY5PrS/cteoaz0DYVypIfPB/
h8M/bwGqXL6BwFkSAsXFf1htSRAtUw+gmeUyu4LRZm1/8srl3HSZe1OfapLQfowL
Tkvkm6L10IbykaBS3d/iHQ8uPCjmjQc1U2L9FDk/fRTK4ZS/aXPheP5ztUTI6jcG
5K354qx+ARnDEm0y8rEF91J8X2eIiDLgFBGULhqiGdQ8Y1KgSp/5SIqwLUfkePKI
+rJjXpUVOEkXZ4JWJfvpFIUb7zbYH/RB6jgV7P8D38gSH9rS9Wn6V/Bnt8d2VGGT
tutFFiRT4079I/MAltr4zwIGinhUeGDPLpp53wTi6JYqOGLnpInW4R5F2UxPUsQ0
yaj7CEAhofZVE61zb1aEO9QRlff+K+9C8mkULj3uh2sD+U3/PlhqSZaFtmRB3B4C
S3kFK4Pt1efyXj+SLqkiP9yN8LEkoWii/PL8hxhseoxEEKTAhCc0TZz5ZgIStYLR
LOBO+9wLCO6kHKzoFAhe0ST5v1xmHDNRxPqhhSH0PA9f8XJM7YPEriLzmLt8nLgO
wOybmYL5EL1tiOaAoFgGeDhhyW6upVmXNaE0+35SosTK/iYmycNqfLldOFyS9Mbh
LqA+xl2IU7CVa6bqwJ/MeHN4kO0oUx9xEGHK3CeEHJNQ/Grn1vmbbrHrHi8c/uQq
/zUH0ffpisaxsHMFVsxns2uQXzc3RfmsIxUl7OKT+hi8PyKMicHkRRHifVkNNlW1
yqaZeH2QhKuefVg4E57BAHd+DU86mgM3HnMnW6gDmuzJuiOB6sWzG4Qmm4ksqJBV
BEmgrELS6nWEkIR2hydAlLBD6hAWikCfzhgSVUM0zRvx4PhnKeD9mhk740slwR/u
bAPbk1Skw218I/D461zhNO8A2/kq+ruIx7oniuYEE+Ygt9SbX52ecSbfaysi2NcD
RdAKbLG7iTEGPFtnH7M6KihHsJxGvigO/zJnr7nPIVNhZRIMzVAUhU9vbvejeGHE
U6BMX2Uv3HjUByOCB6jm/XgWbrYTCUysa6oNg8gldkK7qpeeUocoSvkQTk2RFIBW
+NZHuOK0UVMWprQAZXjjNuKjN0o8P01rDjGUjwhPJZBPddkzJStxOSkISYAgY7xS
I2t55c67aic6dab2OVFn81V0dvmksyO92cA9xVs/ZjB+z2FXWjmiU9iPh1xNiRSv
vjHVvPLAIMQ9AgQBtK+nGsc3Dj9r2utVsmmpsR1oioKeWcr1A93+J54fZSRFfzLr
GgDMQtP3hnzLlJOfx0AzaB2YEiKPuSawcknzp39HpB7tpMPqM6C1Mw+wVLc238Pa
q4xbb/rsQNRQodKJWi4SxwmYGZ6gJJ4TPpRXZjVcP2unxRn+Pj4qH7SenN/72lxA
Xs69W94oMNcJbQToCuAns/dGnJTGl9h9zIZ7CJknTSQH22j946XtZEqIsLDS3ca6
UUDoGV1s7K6eU90iCbGWHc5BhxlxhVr1XbW6P4e5hllZ2gEw8tlI+KrNR1by7mjP
IN7mitlXgviLd+AJAAPOaLDMdEiEUro+ThPORE6QRsKqSXICHlMJ6b4xcod+rBa+
ZfNP7lzyvj5+uYPIR7ucpip+glNE2HFbwNDDUi6ktCljuZwdQZ3DYqXwGOJoYt9K
SAhsQ2cG4CCSEuvzurELq+mLeWtYkV9C+k0fePQQ/Nva6lggjpi0A/emQPtzH3/v
sJpYyxWzB7To+JVS+Z8alaH3D9B9tvMBDGUF8aqsrfWu9wD0Vt920YZJUsTUp2UC
hhU1nz3U+GIDQE8bgT+E8isXyVnFdhBakdNydfb+xXt2FLEROVxo1fY4Phz+YPVN
3j1zkjiJEZPn+MaqjzKRjVkDO9Bzmv+jpL+B5SrzUSrq1qkexugD65Q/L0J6A1Z3
YaJrWL8bsFQkRLsp+hSbKovdU828V6hoAfpAhxw5J60srDiOCADXb3ZCmKy3liVN
lVIWnGPT63V3yB7z1FphgYtRNz71bBNq+5fWB7sRzTQr2fAqQsCqYAbN766XJn3t
x4e2DDST8iiYnLX91c8hXXAwUXS3kh72eJRTtT0D/v999thtZvGuu4Oyxt3n+hvw
AWQjPqMINqhZiHzRZteDJvnkD3sBJexbGkEBkmvzI+G0cFHbe5SiPrXVJDidxzy2
I94lW/O9uhzSQocrZyeYYtg7/V3Qst5C5V2hIt2hPDG/72hsDhP7zQZF5AZPQrG8
dgRAHueF+GB1T2ZGO8V7vw6Rl2rh5XW5cRg/U+Wrgh0RuMwghRPB0qNIj11ZD68K
TBuDG/s0ZU/wWetHFYchf5s8R3Bge/Kg/gqaP4dnfqO2vJyWhD7NxJt/mmtRKfZV
TbWofrY4nbUoRF08srTMT4RPmbAeNEDxq2qcAUDcRdHEpuT+q0WN98VK2b8Dgjir
cu0pureCG6JTpd/G0qqv6/02dT78R9pbM9EV+ih4iM+5yDNv4lKsNPcjEFn6mxbF
9dvQJFMeyt61bitfJP1pzGSpnpQflk5QM10nR29c/COyv0LFf9E0gFEyJ5LrlcyQ
MPkAppjDbYm/x7zaGkn2/hzofiLjHp8vNz0PyqrQE46eX/muymZEbO2MpVnHEM9y
fBvE2nFj5LMSEeq0qoR+L7UfKe2JMyVriJcA67D1CLTFwJTSV+N+TvW26nUrDuWx
v7/QEU5kHIEzV0tBjkN9ivz6s/3T+aPKQdp17tJmFgi+NnEmXNCfiNengeR4+vH0
NwCCi0YnoFQy02HA3SFP+gMtqv6RjOrGJx7SYoPXx9g3QTlVKv/wWO+0HeQO2o9h
EOa+/dzB2wQmkbwwX2Bt2w59OHLY5HRTEKDr2tP+kxT97cE6ivwAogFaFHDEm0IK
Eu5cGqVrS6jJyvSar9rBcp8pMEJ7nt8CuuKVUslAmyk9t5o3sRokfFxh0iKGoE/0
JSUF+u5BH/Jf7Ub2ekwuKf7mW1HXBop6KDn2hKL8AGEcjbZ7Tc8WLMVeArWUm/E6
DzrLX2pCgrU2TN/tDhUb6XSpkn48LkleCBOn70qj+qxnQf2AGfusuqa41qX1MHIp
sA2x/z4ebwCgejkTH6MzJ63xrBP/0XwqIXfwmp8r6ZaKryiKjB3NAxptxBV05CFU
+smyo6jR6GP5tgqQPA0PU+/yTcnnlscEDG7nYC2z09xx6sY4UfvDhjWsKCUDVUvB
ovj+DA8UMt6GnT0EVuzmGt80E5rFGp9+bdSziisjfwRsUzYnWbfLGk9DcB9sxHA3
KSEqEtPZZZ3Sr6F57yeadmBzOor4WWf0xgUllWdAh1rn12yQ8g05dALWPlTz2wjL
c/nIXufE4i9qOe0s2BNaLG82s2X9igoCoplqd0m9U+sZtxPI1oTYTN6llxsjFky6
olxcAgydBKLEVKk4SVZvwGLjte/f3XHB6MH85IpWd60At06r6+RLrJFItZ7soLTl
jayU4Q0iZXla0iri9OckAN3wwwVXmOqEKbPKJ0eaMc5+4pKcrzZEnCQCX6uiixhF
nCswaPHzIicWEp2oqch3kCEOfFNXIvIs+3ew/e1f6d5bWqw80tE77scp8BzdsIj6
9prEaKGJc8wuf4ZN/95dzYel3wtwSTAeRX6plintPf0myyE93WwaFE1VglEb4xQ/
Bb3drCCEd2Rk+eH03WW9rguTf/kgvvDhWZCo+do90uDiPRDS3diUwtayDMhdT869
ibL+vc7sy25opUfnFnnqKybEBCY6nKGGSnU0TNszlNqztF6zLDKa4r9rhGdVWMyr
HTTnMEvyTiAsQelkxjOSJ7nUNXRb8W9UEBhjM2xwF/VxPPyJ1y5q/fwJX2UUF4a6
4xtS3s1MUMpsl3NoDKa8I7Gu/5e5fO/gGta517vtWza/pSx7gVuz30U4mpStjEGt
ddmS69V3/JNsUARnPxZhGoRzfHPo2l7sJghk85URrPOzHer28K3S0aoIaxC99FJa
n4VgtQxTynyH8BOaRrLr4VCfMVzeNa3tvs7yUp8l3BJnTLNsJ6zMGPNzJ7OlMzSw
AmGl8rWqVfDCngfqKfvByvMos18MqK4CsRXsoyQfuVAKJCd8thFAUgZnWAFq4o2z
7UbwsZGSjH31HM+Ujzqcn9u6/hkGGRx/DxhhO5zvB1kO2oaC1CYEF8xrGjj3crnG
5j6j8MGOHuaD2Dum+n7kkhyXcBErDopTI17HNCuKrxZo0zq/SdSi0QfydCSc4Jth
w5lbSefYXFAJpON4M1hNnG0JBrNLWSTs655I8+dR9i1sjfeWlBzMxkwdkPDHGMAc
MIXs8TpfiQnRiX1ibzcFSQhZljHaGJYqP5AHbomxUaubq/r+v6oQ9l1RC7xOAMWo
7WnbuZnk8SMRdE4nTNtsXN92fe49taMl+4a2ttfQ5FPAeg4eb65fKWGCQzfjuXHM
VF2sT/4FrER3chtSlWazF0cPQ+aeDfJWN+A5FzXYyz8/5jFtzgnuL14lg7Q5BAGX
heiJxhjfnkvcJmVADZYLlDv8jWqpvMfYnrewYzOgKMqvmcdz2L/y7OcnW/SWKBYt
idL7UfsNwfOdbGANVlKUNtw8Y7zudXI5bMYt2pSNCDlGTfL+ngt7KJ6kRCD5qI2n
ShxgoVAlt2RmEfrelndGMVy8qrlxHW5if7osaLLzpKRwuTWPDTO74TD/RMaa/JP6
GWE5h8XjDkffwUNfgkmCsYtXJAAw9jlo2reSH7yimGq+kkx8RY96yekVxuFthIL8
9ev1od4rIGyZDTiJAPWej+nF1f5a2hs6mfhRzD4GvlutkeHAfWmvkUYmRq0AVU9u
t+BPbBxHWg60ovXU7VtElWH7h3GqCtzs03lEcu8n3XhZIRUZU3bSnGaSGAsA4Voo
YVaIyprrd7W7er6MEc6vyxar1ySNPbawUf6y90arWrb4+JP7k5aXfcuz5wMei2/+
BZnVOPTY9ESD+3Bg8JzUoa7k4Kxfy4GER0lVPl7XRLcs9RDsugcNuwhtWSST/JLx
xy4AL5KRZldfenFKwlTKGC3whf1Dx4Ni8UVuEHF8PM6xLP/rXLhpb7laU4DKcmpP
u3SouGZqUhFKJR/R/lEncMijnMJRGHpzNN58eetpJSToSnBZ1gUTCnmmrz94w+7D
m1Iaw8v3TuMHvPvVwAg451pIbgGr9sHO9bJrd4OCl5vCeYwmhhkxYBKubWTGFh8n
3TCJwhVrf0CvM5SN1g0izDDhUwlOHNFmRFmEIfWZ13JQeJJpmU3JBjHTCT1a1aw8
Fp9AuUrvWgT4V0f7O1kWdZIIa7zAIi7Tp5ZlbOesKhoX8+aETV3cPIbY8Ll5hLJF
iNHePCf3GZiYVT8dinwDirOPTj7qnyd7h3eh9qBpTAFCfO7DsDSj64OnGgyv5Ao4
beKYfiY2F4Ct8U4Am2VkFTTU/sJxL7LsTfV0r7xiFs3rdAtk0Di+R/H57yVVebhS
mxaU74BWxlUchSdORWR3Cjel9lUI0resHauK1/tDLY0TkbGd2n0qmUGEkgSWnHE4
qJGHHoh3EdSj3VmvT9B5A9NPp2xby0b1AKtQDVqenFQUR+bLfeVCDaqgUOcIOu9b
NfqZyQevFB5BrV0yqrfkzjKeflu/lfwlPkv+fzEImI9qkpAEsPvatlrLt+RXRu0o
6qbO5bDq61EwXJu+5rhmZI6jtt7vVorZ6nT8c86FNiHVi13l7bjfFuol4XUiucat
F3K9rOkE7OBIasVrc7W8USP4dPn4kjCfttyYWARtPE2dxToiwo914lk/Wha9Zhiy
kz/ZQHFNSCFUUZ1ySrvHZafgQMP+jYqWhE5mnkPcxnMuhpfFrqHnUNDlzZMXVsrD
9a/rWY8+qSaN64ks1mnDLOOC2pJUzLw06frGJlekJ0LNWsenRYJtiLyC80CFlwZO
R19IDecKNyTmajw7dRK7G0wDDt2yPCz4X84H79HZknJ6EZYpfV/g9677iv55JcwL
GMcUULN3ptzzFE406c9qs8rsGLA78gTKk/x5yu1KrvZ3314ZL7umgRML3QlJvGAW
tFyxAThiF9UyDZ4nh52xVqsY2WewNPAOYQGjUlZ+0XHkt/kHnedJ8QpphYQ9WIe0
KgXSmpsZ3emglKUBnSUWnZzenLNENfMd7kYU+fpf8RKyBXBCyx2tLlEYtpCSdquq
UzUFJxvP5md+/DCLBbWWVI9ythX/xeWLwxamb5UPr7MEh/4cN9MiNU2tevy3Z4eA
zeZXd1TLqcTYx+SfhcoUha7J9ebu14jNQE3g6oJC0vDDVMRiY9YPKJCsKDw5PkaA
kkLasD6zVzY5rFVdWBQuF8SdtG0bHkNdzcS3Mp/d2PqcPvd59ja7qAnef1Yoc+8C
kV4EHKsyq0rd+C0olTvmQJV6UP5D7cSYKwM0b79ZhuoxjZruGflacp1Ybj3HDrGD
N0tw/SzY6MlKmwCi/F4yxEyJwVJO+a19ZZpXskVI9Pd47jJL79lb2TW+qk6zONYa
T1mvXCxZA1uLNQ/2dPf4/MtLQuD+tFT0YqHlVbgWKcUPWSZfHVfd9dbyBoWjWD/a
AKDBDkNcM5IcPExisCOjsklsmOT9hQ96vjoWxwpb6oTMHJTPIin7drzps43f05sp
6e3FLL5HY8SjWbBsS+8EOvbWWqwuBv7rsRJaqjk7jM6qb/EpREtUBRAQBlRG4aEu
ER4Wa7D/bMM//FpNeqIO17UsRXCbohrEe4S/JGUZlwX/15/ztzYbspIUa5oxby8v
/lkioUH98hFYv3GaTR0OUWm8SWhQTcV7te8qcNU/OZqtZdRYckrU4hfTExu7aFZX
PFB8Y/jfKHcXhChyZHFXtjbkDEefRbQrX082ul9QW/xSqOC/zT0rRZzlo7rDNE4y
oTPA1kf0piZHCNkdJMKeWVs5djM90H4lIq0EYwZDKXVJ2Ye3AqvdgJmjjtnKMjc/
CmO33CaE4RVPJBYrIEaOAWsemjZbhJH6zrCoYhOuATAa+9ZKi7zGObHHnQRlWg39
6uHFXDWkcJqwUcwGPReKXoSexcEb5zPePDzSBRZIYlGK1IE7fBGwzf6CndnLU6h9
e5M2zpLz/q6k9SuveOpOFxi5BICAM5gB0VNGJ5TDx2KE8Q3nPXS8jUzvi9ZC3z8M
33i/VKqlYQw+3jkS3mdKBGdkiXVoowg3i+6bayZU8sr0R34f9TLZyXc/mjh5lrCV
/toxMD+Mo9+gyzkjcPeHs29bEnMK6bqNTth6rKNpeR2/pTbAR6hffawYc9vSeE3c
BueYJVi88ZxIUVcHx0MiKkJB2B04yxTHst+Ij7BLlfxkOVnvIrJx5ok5RhBrpvG2
6GlkJleErk/Zmy35EdqZnFTxawM7+otbXM1qhkI3z7F/pqKgbJEvURGPX/GaxvIp
qvHRdxZd6Hi3jaiu5eGrypqJshf1KNRP6eh9oE0C+qdnCuh2WDyOYPVO1xlgpBkz
YehzfMIugvhT4Ol8uLF9u5mIx8g+KZklHaCtrH6CtScJacj+/7SxI+bSy3K+oo9O
1JiEsbsrjHETv4NK3iyCmCiO4577IshLP6oHc3URtX5gNWbNnBvur+Y9e3w4Hp8G
2jW1hhjD9KULc468VcV09Fdl33umfH9K2I4+9GSyW5wsNlOAF8JI2weZE8iklRpG
jSmd9A8pwR6QcATdZ3SLaCNx2kxJzTRduZQwWoj1YZtjFpDipTUVgVBs6hRTtmdn
aICUMNQHwA9SpXfQOpobCjIM3n1XoW0pwvQH/rnKMFcfqy6Ihqd0LMdsdYYi2Hvc
2iUL4UyzaCExkC8Z3zsXE80P66mnyHaWVgh2sDLd7UDxLF2t7hVNaqKrJY1XVqgb
haCkMi1sNnYALjwN+Yoi1Zc3dmllK2RBPGlHWJHxU8NqsgzDf6gadvfucgjTHHBp
L9uI0x47DOS68J+M26wPR8OhQKkXPOhcC//wO2ZWJqYm6TGEG9nKN5wuzO2ThrBU
vPP9uUe37XYUhiFX5OTb5IHnVmo2XmqB/zUkanCBNP/T562F4TVg26he4S8cbNL5
oRN4A0QX4CJh3UWvyXhyqj643u0ERBIl7QJGYCYAYy6yRd/ZaZ6Yoo8m2RZZUX1I
OQX6YUVqFAZVVewhizBLBLYICs/TMlknHLTQYSm7So9XB1cHK0HfYkts4PmpV/tg
r4mEsyxaq+SLiAvEEjjaKboQpVBr3DXOvBOFfxR86RVkj+FuIdiGhBDVebvI6Qn2
N/ruo/zTuxFzhdInlgls0OhFrPIr0XNnEeUm4gd5VTTuhyhLNvL8og6Z5vuTUyS2
9C9rvEdLemi4H1Pkpwzga1W6m7kmBk08UW4HcIoogjV/uBfGeZaHcRunPCbSUnpC
T0XdLeqJzNo/DF2aEg2zQcSyNjTMgzqhZ9cDGYxxrUm3T6pVEwMuc7SYS1SiyAri
AeL1H0imLVo1KmW2gnjqfFhy9LbQtZZU0USCWBwRfDKIntsyIFt49v87sxi2rfop
qC2O/a1elHEQBis29cd/AwZkLkr6/wyL3snX+8zw8UYDl8OQcGXbWFLCzxq2J5fu
/oJahXyhsgTlQKpue2+uTpOhjJp9O1UkCcvCJNVj8P4W1PMrA/U2rv9EoZ8BpRJf
2k79eJZEdqBxblqJ79J7hlnwAdFvaW3ejUmTU5xLI1Jc37bhn39qkt0ecgR+EKbW
4T2yItbAa5E1KPCM0OWCsl71JCaShqLq6mI1afLwntjwnEMSW1lXctBsJza5lDOW
tDiwG+EeQB5yyY2VCThWIGa153k6P6Q/5/ZPg7XR1Fe8WShRF6RfO19IVFobmHpP
7B4Ux7zxr1uJu/A4BBBv1lsbzV4sutPRjgHndM6aqu0zWYaEnzc9QPm/aeS0m0bx
PD/B+sqCSr3c96WXn21QsRAakYN1ftV2itIbfIshiPXwE3HEtD3g08k835sU2nK7
oV6IyKsVebgt9BzLOcNFvQRU2j86qSp2ioO4g9J6O1R0TdNvCBCmI+hCSYgtIRSb
2nliTK7hjc8gTqxPd0zW6l0Vm31juLBXKRynvi2LeswG0ANYnVflhBqBYIlr7D/8
nuIT/5U1zAyGcvU1+/xO6AoMAmvfnijXLe/DJaUngAbcIW3xymU2Poe0fgbHGVoa
BYMgYrlc5wo+zBeRHjfVvI48Jc5DPymcn7xIutgUGncq5iaaD+zNXDI544lDsUyd
akFCtACRSJ+lTQ7H+6CHmPWwXyLYzoJhTVEupjCmkjBBWS744ZcfULWRpRYUM45h
KOque99Hcem74W77XwG1ebBmxkI4a50vQ4nvKoMQliSYmJ98mozRerXQ1fLYvZAH
ARWC3V2DEXxyO7zO1lg+NjLfaZ4pQfacQQGbMKSLNBtHID0bbKKa7/BLINGJsn77
HRiUcQADDIBdj7QTLKDqJKa58GeQC2WQ43C/+izogNhylXEHQ20Mdg2SB6O25Se/
bQZb1fWWYrAVVKJN5HU6tIWuEgbOrt66dAUlVzdtIrmXIjDuY66OFTB7dIDX1+33
Twd8HJZ1hovaDf/gtkTSamDAKMdI3o/ZjDKnSxRb3x9Lv2DBUSI27AhIh0S4wyy3
BRKvhvtkmabogdTn0g7KFuX38ptb+zNQxSnYBLSM2FWHfiEStPnLGYLZGYVyHkiM
LO+z2u6pn7relmdtxBDlWeOMkJK7/a84JZO7jpc3T6xTppE8XM4iqsy0OmZfCZCu
hyI7NBYmhCHWrZEYumdwvqPGWwMeLOOMOuOyZyhTD6+vRUd8qY28nrexYJ/Y9Og4
bqsJ/sfZqfPtwZtfo80BADxzbLyjRqGWPAMD8+bBOH8Xckv1A1l2GFmvSSfrzdA9
g6sI6uKMRCo1H7JZiHlrP+OJ2GRTFCrkL9DJb6Pok0XDOM5p6pHLyLFUhAaqzG6Y
qUeIFY2J59Yofoyi8VAfNmiqxhTZ7yZq7NaYl8IqKZGlPANgt5IsLweM0r8+zDH0
cwpY7z6vdFOLX7vfyOjSqBdjAaKxWMk7K+hbBlN47m5MAfXjAEjIrZ0eh6d34fjd
Bm9hbKN+4Tsbzdf8G3R66oYn33m/Myfb3sTaiTXrewgoGORBbfHi1dW+zvva0iG6
uLwkG3RKtkT0KZRG7faa6Yg+uOcps3sbRZZevgqT5pr3kxtEND0BFQJTSpYBc43M
nJX/3BiqrDDe9ItAGk6mJ8eLgW2EtS131ZjHFaszc2IKBdoROhCU0EmH6zyX26yl
RNSA6QZcz2eylkL48mt4Ypot5O/LxzU6N6qCK7muU74wEemAt4yaHYNdzDbSgFhY
qFg56RFLUnN3iLOZ3XypjMZf7C77HPDXknG7vlzIptauuwRvHHdjyhljNXWfFJPf
SkBjYX1UKHA1YDw5ALnCVddtuLSY9qPKkai1CqecSEElI+5raqbhrIKZr4qbSfA+
TDubZEYUB/YLK7OhJxVLtmvtGFIcRI84ScwuhzwDBThj9a1xFFp6/XZgqemuhyl+
wmFfzo8zlvKIIIV9JJyxZhzKFGgco3kbeeEojTk7fn4PmKKcMvwzymK59NiezWcm
OrPVyVsgltX1vqfMi+lNFK2mQkdSTp900aucx8hWj9w+OYDAu3KSgTC9J07aYTpm
gXADvNyOoj13uV4RRLFPoqjK9vudvfCPg6Ly5V73wXnE+bFlDod07n08GsC4XO7f
gdvYGA5mRUXBh+fc9GQ5lB0BwL+o/PsZtaTvS4uOaC3L27tnT7KbMxGws0B4daDB
r/Z3Fn6MUpX6D3iWQYn99RJ2ATTNbIG8HT5YtflaTqDUm9+WcOu0N4nYS5Vt0XTy
19HdrvVpJ6y+80f4kzt4tiPR6JTa+9KlcTn5tFkg0GkzRHEn3ama8D1Xvus8o15Y
IGSRnTaT9mQFrreOgWvwRBLWrDZMKwi58wHjVflsMIOiKPcXB353aYWks70lfcnr
conNtJKs8wmoIfmh2LXMmPqOWEQj5kSu90bMjofyTW+fwRLmEwgOUuBg0uQQhRSW
`pragma protect end_protected
