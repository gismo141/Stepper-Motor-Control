// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:48 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
P+HCoogF5e6nh4QbcuDuds1ojPta2SxCrGy1h0OvGvZipkGBE6elhnAGTmS8ndqX
+w4BlkgBGw9mpv7h3A7JC1UWddjmAi3iU+xDsQ+y6drctk3FrEr1XnIzLBp5T1yQ
Xo4r2BGFdwa/n3Aqo7qzVT+ZGlqgPmviQNWHWOb835M=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11168)
hX9TTcKlPKEINYRX9+TBj/7bMoiUNA3g/zjL9L3GQ2ueUt8Lg7Q6pzVTo0kO8qDX
Yj6+TfmLz/h/K4R4FgC43d94MPSr7fKp9gzvcbh9wg2FS0IJlfItlQi/x2GrRl5g
oFetnpje8JWdmrULoWJMDFXN4NTcoxhqMHYQjSBkgm+6nk3F6TK9ZVCMQTTMMkbN
f2Zc0vdWIJD/EBt9iOZ77QNib20qeMSR579JIS7lZb8U9m82vgfUNMBzswlxQS1t
hzvJWWYk1xxeb9DDylVxtBlacyIddvsqSn1388wxqJgS4dir3kyzIII+HvTxNclo
dgB9DVJx3nV3XMpvNVWvw7ePqINkz3KASuwyY74xugZcXXLnHVF+zxVzBUx/fUIa
OcJtSfGv6pZaVv8iFN8oPOug6sKlXy+DpV8J1Xp3006sJFGZhcotxN/xRL5XHaxV
dw+QHi6ld/gi+6d/lyIABq+mXHzRhztY/6SP5DogyWZcOh8NzEJZbC62/TuxLIZV
IgqM3Hr9IYjda+/K/ys3MK+vX8bMH6EsvwxbR6e+c9nRuC4i1tktifHUMrbeNt2a
w0lNSmKi0545E81S6ZSr8fRYhRKITuvAh4HlhVoiRm4pNxhmogdmKaCxixTQ4dyS
99xoI48+vbiz/Gs0X8/mHEzJKLD1hqSxl97Po104B0kKzR64Trj/Qm8hofZYaQP5
FR//tbFBp3be2m4kXi5j68yeTfTunkq/IrKHQlTMAMarksINMXDgv62M0YSX1Dnv
GXBCg9uY5yQM7qjzDoa1vxXJbuZOIqYa9tgo0kV0Tpn5HlguEi38oy6vil8Uj2pi
Fktwj0jBuzLQB4TEZ3Jn0iWyN40gZ0R6WmDt+S8sjmfoNZHF7j881T3STfR1c4nV
htjYh8GdN6p1ON+f5LG43cZ6eFLv/I1xTQgI28+HUrakQDObfZMRsPrq0PfuPQ9O
CiULOrjS7DA3Nz/Jnv7KIuw7GqJJwVkriIi5XUWrDVmxLdOX7qltVEaA+YcgnFax
e3Wbbv0tEoUeSQMoFEkISGm1lEgcivyghGQ51CnjdhQcL/pZN3U5cOVzxP9UGbuk
fBwkgL4sXYM4edXE+N7NzeKKaOcQQFAnTT+V103tXkAut9g/WJrUp+cqKigzKxKc
nhAdzTxGmlQHKyqcCqSC1wqB1KtPekyYU5sDD6oxwRMc9JdXcVtKIrYfALeQcrQw
Nr1WuO4m/6XITmJ1L2PeuTrfH52J7MEGJm7vND4Eu2TdpAusgQKoi2rkYoTjh2hC
iWT4+xC95NgjMmTC++mrSQJ43PreGP/UFFlKFSVK8+oCpe+TaTGvn8iLQv3OdnSe
pwNJnyFhymqssYmd+49eMsGkAhC8xRdCXJ9MlUhZ5liC2hqbVCdgkCsxMuBNfTZK
FtnqoYiaAET26QBNhaNr9lLDk4VcACt2SQp+/m4x5QbZN3L06a/o4PVkD9igAO65
yFLz0cSZNxTTPirlZnw5b9pNzB2ADCabcPMQeJ6lceSyHBZcOFv5tAGtSdplVgVH
JZBgHqp8M5UgZHxiGSEnTQObDh80imdKaU2ZzUyQ0IDWDPxFxZxzazhgfd37xEpt
4IXHfp09ZO+u5Cl053P3fz2+TagG0W6TH3upNwZkWQRCw8X1M5uN/rJfS1ZC9//R
hhuw+1cR+6uisj/jnDuha7EU7bte5gQS0VzENtYhgM5BFaEYdvq16EGkM2CDdG4o
gV8qos7cS01ppxKdn3CclkPjpNTHO8n9dSTmoHqwGtdR5cQfRkusWyEiPLS4+OcT
Ia6rWRaOfVsoNTBFEkqT6UveZLe9CgskbeIcOAhBBSluKwhObBeq6V5l3QMBaUGy
GJTjBzflvXwK3gkxRlLqUSx/nG3fEO+vay5xtLzbyxFXshMZwGuGsbJPbv7fTgBR
33v+4WX9PuefelA2FBnsq2RcPt7yM9Bpt/GLyFwi9Wz8NKBA03V7yCpopSRWK71I
EPd+uPfLQH9WLlNnRYvYxFj8WH9QM7VrS/qUxuOxwuLBQcbgxVi3TGemykJj8vAj
fOWF+Kx/jwktI5ueX3w3lShtCDXAUu+AosZkXlvaK20S6Go5LP22U9umsp8oTSZr
qrF7eAxUjuB84UDrJNTIdr7fs6b8QwPENQkjEAhS+slH8uq/EVD5icclBJoilkhH
qlP39t0GJbV8D5IBFnjo6AT1GuFxVemqt7Zst4XeAZpYofpeQsyybUbkUXTahOpw
9XajhmKZBmNvV719spLi4CgHxxjHVk+FLFFSSuks+S360kGsUMzfqydayn9clm2G
3vVKoaQEhdWbH6t8PiGeFEUY5prLSq8UNq+PNh+e49/pfvZQ7pyiOU1tLruBXrSk
8+/fdknz5misrcQLI7aiLIADpTAOn45CoWskw/uPQyRyPWRxpUglvOOvZnX0sT0G
KA9IMKouwllh8FPn8JnCDRDl11ca+HFF1rJO6qNiLpEaA8WESVwOuQJlMEZwjoP5
JMox91apBJm5AfYjS5N8s58CCGOLzJQH0d/EvfAr7w92ZBekAtGwZi2H3DrFhK+a
QYt4fAiV53CafJ6JL4nGUrNd4h0KhHcM+Xru5gq+h7o1LYMEfVHMOeWT9u0me/KP
2AUn/L4oDk1nseoSAeK08dXrcn3GYCwWPE5SJPnR8B25jekEI7tZlNXfKoKyF2B0
G2RAb47TAcKzifIxwXHTVpmQzU/zfGA4LsVN3sD4TF6YO4OXNs3POYNmEAVujiVf
551OI3uF5fM0HvSiQ7x9hx6I4dvO5rOy59rspewtPvZhBhF5DbpuBSIuBjixZJnL
44E2SiJp2Rdu/ZvneHWF7d33EVLT/nyjcqx2bIbrRk2zG4mc0T/bLEeQRh7uncfd
O6MW0m2AwkB0/1wNsw9kKzDm6p99xqxpScXZvzM5Twz5x3EpD+GlLBVE+AZBnkl5
Nyb2eB6D951aUQvkckUUzqdGH4e+lRQ2vTfHw0GsxUzIXYM3jD5Nwj3XhHVFbnhh
ZDJffTCeATtYEDWuQtGzz2hByYluHKQkNNErcC/gs504fxS/b0Ese58xvGWRoDiJ
vFgeIJABnjq67FYwAIvZ+MT9PMi+183rSZVlKZVcroup4mSVQ5C29/s8zZYqsHRO
KBi5u+XzK59DppAjiAmkPo2INpcB+wpAwyag8LyFqRzxJD0rlAjVdoqBIH39l0Jm
TjxizYFnyyQzUwlccNn9CGLayUirFm0swlBTik9rTm1z7lNxR9bpnXTwHHbAklZ1
ETex6Mvim7H0zBtfW/DtI+5yK+Yqx+4eR7c+NYJ0j7q/xcY768KIUR0dAvpAlGl1
4baxeXnXdVzb8TLJPs71i6RBTfqBS130r1vYzA2EpoJeMdE8lyjMFk2uZimNKb7i
syc2Kc5wjXEpqh6VqQVRjKtW5eA3pCChCIKjYVtwBcClBoXTEBfV+jVQEoAexvwi
2IrQ4ZrY4mTVgSOTXw0rfxtaBTmND6/fjSF/GYQWAozKQwwDDbyTSC1mVxQz9Cxi
PMyPaQaFxLEa09lhsWGN8MeQaoYghLoeFzZcI9RK3W6k9pg0CnEsqh0529ib2+bq
WwA1QJrruuVXCbMbO8LrxtjclG/p7MUEQBgjHhkKU65uea6FhHUSi0sH3qsUz21L
w1QGr39+pIVLXJkim//sv1zKmsjzrQUm6vyCfxkY4QN3NSx5VC2bkJaIoqDoy9pj
mHeZvwkeGfhzRLOWmHycIpOWEDYCOKk8bMv0jk9xdP65EHDxMgsBjmaX8peA1uvT
QDHd8W3tpf1clDKahJ7NiSWPM8S9YzCcrtd1xlE53TzNhcWf/IxPKg0SRlNBRj5A
K0SXuJ3s4NcU18nRYXn1Fp4Y9B6hVzp0iKXKfYa5I3jGJL70I+qqzS7arJ51Kzq/
F0CssAfSHA6NUGF58J6hndO+/ehaFZeunZyHdkB7wYGFA1WGmi9SoVo5n/H8sZf/
JFb0FXgKr7ZaVo9ecobPgKHBpK+Gl3XMVIkcQd+Off32/F2vjWwvUvj3l12Od0zv
Tw0D6OlCtXBQG52Mt+N6kWTHPNU2ip41iLb1j6MymeZv/JgaQK1gPMIimnmMQIBA
QRChEMUL8ouHhIbLz4i52vIq2e90vNZ23xq6rHxS7sMaqkgkDu2+/GyuiL1AtZPP
ewsL0vW05oiZ7yXvugBVrAICWXDug1goG3VKpWL/RJYLPEaRj2EucBQwTBs7ZNOY
fi00fLb2Aw29tZAl/VujeYlAuiTMfqD0hM1HA4nNmcFRk6xfjDMaINF51QUiJC34
RY0BMdOUTsq0lTZaasbDcZuDUW4cYknQl+u1IAjCDu6cPO2HfJfT5nR85ABmgm7u
44s/4krJfo19A5wyKLN/YRU5dLqlwo7LhReab7Q3cRizdQGkOQ7yaOdCIHe6eJ52
uVEyc/aLtTpTOoNCzyD1dUTlR5nQsLbkmPYHeQ+kqi8xUxEdx6CmI9S+SZ2IcEWF
96ey2gg6vrWJu7BMSp8Ks5CTXhcWIQW2kAW7K7Jw3rl9RpQ//zBtT5Z64QXQUQ7i
cp3MP1amv+lEdgmeqFs4ksH6+loS5N76/d4B9t8bqFH0w3lcvrjLL9ZUmQc5oYdU
ta75UnZLjPOxoAVblZsaDjOCIaNu9TiiHFdmdFZ/ddBwlgbBiJ51yAuE4ayq/VTE
iUOPz8nPZAc7pGWKMAIalWhyB45as5DgM5W+8gt3dRTrhd1hVyBStKSjMG43OLez
YBfZl3o0nLfpWEEQmD87Fj9my0u4AUEP1KOFB1f/kDXeo2Wns74xKnU5TK9h2ELn
F2XOeiKoR+6naDX8DD19aj2AK1emvqMAwAC3N8zqpZ/WSszMpGwmafTxGIp/nQ6n
fd6qfnDy4sOFsGkKys54AHgTzxb9q5D8cGTKC12iTOEq/WwQjtadxgHTKZgCa3QA
u7NUoNsv1ixsdh3UMefuUMZM3cEySyhAVTSjqXgNmQkBBXo8EWkV2q4yGddM/U/P
BCOy3A05OlUb2G7n5Js4bd+64LdvvSUBFIYGKgWajAEbQocX5RULr+0aRW4hKEtx
6svJbJH2JUYzrziKTI8XSeafP/BGxSJRyPWwnA2ijFR6N6Zr15GNeuZHABym0BqO
H1wl/9XHDvVMuDfKUUoRl7FQ1PvT540e/+sS695sX7uT4U2kq7v/3bzFCHPAwAU8
4AMaytq6C1TG3CIWEc699ii0AE7qW1Uno2zI8n607hYpjhWh2i49KP/jhYJTcve9
8PU5Gs5lcqrIWEzLLs8L7CAraxIhvyGGt34G3OUL4O6hAdozaRxLCb/gxsjsUmhg
/pSv3+EzGm0ggw52yvg84i+qfvCk0sNCV3bJ/nLEq72muEa3i5leqSLV2iRJSkHz
MX1gZAf7k3mdERNVZqoesYvvZydDuWVS6PQxFJdHMoxY+0uHXEt/MpPbFKrLJZi1
lB5ZzSaq5s2EqvYNsf93nLqqaEISFliWiiBcFZEThQFH63WYDgnvM0D1tYtem9Pw
a3j3Tsf9x7zfk2NfvPVTzNT83fL1dgqZyRxyDZxS4p8ICYqo1cfFxhVnlN3Aok7c
Br5YVNMyPEShgyeqIYa1P6DMuzWqBrdgZqmGJHVuQ4DO61FPzAhl9bhb+LP1zbVG
Zy8UK3t4wcvoDx0B98JVgTJeKYfKyLNAe+V9ALK/vjB9PHcNqQYUg9wvogKT98lj
9kBO9BZYkxX4pY4gJAa18FJ+DZ55eu0M3+qBvyf1KDIh2YWtWDaPxVEeS8rbpDeR
NYs1BuPgOtFmK4mYN6oSLd0Uz9x5bKg76OpQ2y4zUAzVyasseX711JJWkbe825LA
QaipflWEazr5NTspN5AeZ+XfrlyANgX28WT01s4RrWEeK4Gkc0RxXCMO2KirdjdA
i1gYlLQ+TB6csXpzsq0AxkyyFRubSGSY5ixbyOxm3tB3XdzbQXV1vllo9dYEIKZP
tp2AF8xAsiSR5Imm9fcZ0YY0cS5DR/+ZnM2IC1fA2lX3hg9vBzakPrGPkAsBpEd2
zEhJukLknAPzmawPsG0RADhf8dwnkUZvEkigLN8cZxcfAhHITnmT1UNFeNaW7yva
SqZ/u+xnpCfv2vXky+54Gk0f95m5aTcIgmcDy/u/JszWv0J9+x9AXgvsZG5IthMO
Umj3CyiX4CZ8ttJTt89MLXziePCXgcr49QkWo+7kTEilSRniu3SQfVw3hAGMXKPz
prPdjdUSTQfB0egMbQpGFAgfE4wY9L/x50IdicHD8WF6hY36zDHIpzwAvE7iLpdq
t2ct1Ufb8FZ1fvzUixY79HVhHYYv6yoNlpJ2jU314iAXYzBjXgD+RGUi3VPvXPbo
yqDem6v9W0mV3vCnT2hnUbhBnhVtCRWqMWKuS7pIMaWKGhyScOHguC+rv14ho5sj
BLOFg7WFc1G2qT62mLudkFkEItf6Bq0QfeYkTsZCcUpPEZnEON3YdqP9ZalQLQtc
hyZ1yOkHxF71vRt/AOOu+Or5wA2fbL5Mh6SlSj9H32N7vEzXfws50KOCASk0+TUB
0o5ZgqIoSNqEe/3f4Xq2rJ1RzMdpZTZED6a1wIQs/hyQn8k6MKZ3GNKKVwcUNWim
d8EDOdpc+o0OCSWS4DsBi1R1VZphkaThx8gQ7jB5q5OhFKriE3znwGE1rngVzJKZ
4uVxSSo2XyB3AofPWqLEf/rd5ECXlPQMzgFHuyoaGkphP4eNYHWAgdP8j+1DDEjw
qDUZW2cLAxXPwQDSIqgp3D8Ut3vk3KSLeQBrtHIFZ0QteH/hDGGz2THdim0443nc
aDRvbadnsK7q4ElH7vuxdaPA02dIvr4SzI2s9nY6WClj0pmHFWybgTxMqbMCIPnM
PiWWgZ0x+FE5ihvCxi3SFQ3RqZRm+F1qcfGORMXKZ8In1ji3UowRcJ7CHwKEC4VS
btiTmj+XCqzxTC/Cnldvv5OuFibUv/mh4t4BCfXUfcXeb4smLRo8X7OrSj7PhmcT
F9I/d20IMHX2z1kvvDRNCoyVx+RCCWk4/uXHhs8akt3sOfpcVUEUN/rmZkNcAWWr
dZg91gnl4JEo3mmMrkkDowSI9SvGJRgzprrmMIt6l57mRCIZ+tSgKI/3crs3O+yx
WZYHow9+U4PyBJ9DVYCATKLDSaeqDwZouCeBDflWVDvMYRMLlDg4fgXmwzQj4tWe
DHkdhC3QD47bCIF+b1z4fUqDuW+nD3imHJlPh87gZLWYs93tS6YOIulJp5Tea3/Q
AbokHotj7ogq9wJqNJHzyu/MeQo5kKUseE+sCrJdwAts4sxsfdSNKpO5pKBqKDVK
BeuadM5xB+KcnL5ntcVIAYHJUMjNa4oyNqRGdvPXOcaaZ77q3dhpaqf+9+I36g7S
/pPaNDKlg4ryyHsA1liT1L59r0Coaj/RTgmBlxBB2Q51OliRo6XEu+lsonFfA1SC
Ap/29kOwl/qfq8MckOhZG0wLr8ibZtEDSCoDcwHhBPQBroelrlp7PR6zlk4vK0El
0W3jGAzYRsduipn+pAbXjw/m0qiOAFqZuXDQmo0BwTthEAZ7W0JgqWhBD7j4PPOO
LGDv21elV6xvu84Oa3Lsj+ShkBrW5bJdMDYRk5ro5OBQtWiWdyPQOcPnm5Rlg+xP
2D8rznNQIyjGpOoC8vsCEqmepInrZ6jkkHz7exXQCv5+8oIdh+gAyx8hSBxeyTqo
0zfTUPO8creEtjjtixRLx54Wg0ZwUWxzCicAQzEkcAPXA+Sbv3+tChNb6mxGNbdA
8FY/eeQYTB4SRQI9LpmCYwpSWwAzACpkDPnc7LdCkSLpYHreuS0DMlfYBI/yZS+N
Lj28EkiJy/X9xRm0AgiAcNCBnMTdqWQcdtRVj/y7p0p/iJH6gzlBo3/4xEbO/leD
tRVHYBw8dgvUHdz3/8TUtwnyA7BJvORpT/mr0LJS/O8+fbtzAZsMA2bGwM/zrJV1
OtE/9S7DAJKO1wAMo/SFls/dmokBAj67HM1P9TFSl8JAIuMtvsAog5iPTcjefP1u
UnBks64hONIMcX4kOSeDFydT5pELQSc1eiHotlh5CZ+thkdrmtI87JILWFvm41/C
Wl2h6yunsKghksHIAyxp3u5w6lklZk7AIlHBWd1GhXEgsHxUrudIu2l1Bi3kIZsR
KtByoM5uPBmUvAfqB4dEPNuVSmGkm6Rf0/Tt8jNkTZl9p/qWscHCiJtRsWIGyJSV
HTWncED5b2XGppNwmd4bPVab3In4abatIdEY41X7oQG6KFJGcAWnMRFrIqpUCWsZ
DFYqh3uRXMaJAjrHoXiVRwFqR1MYTD4RTWZcB1K0LAGOK77/P9Jj78CAP0rIfl8W
i8w+uXLm/CnmZGFWhTq8otf2E5s57TcOLsJngXZk5V8PwymsqSn99WM8vJWHto5Y
Ux9Yde8fLx3pFpwAgoyqfPzsk6cXfqJDzlyeBmg+Om4rcclhKBAFvZWbVfy4FLc7
PzqFCXSfdqtLk9qhYt+p9XCzEJ3mbHn+8vo31/3cGAPpwrGnwf3NK6UXcOX/85XY
Sf3If4RzYytDeeDcgJGDZe8h+uoQhLEf2fdndKaxfZxyGoWik+NUbVyTRVvmD+DZ
NoZ6mtLiYGLx7YdzMxnsroOb+a/pkMujunhdd9k781JJbKG7xt4+lxAYZYTOPNB7
o4AJY4CSS6XFsEgOJFHfogvMqQjlIKonBflW63xU0N8nJc5YQ+7M3603eECQuhVN
6/LZJUXKulagcEEvZRKjUTtbcuUwB8SS3wvCljvPHlOS/hWGaHkwEW/5/+yywYAN
7e3HMCA4SQ5pi+UNg6yy0yIBE/5XZR0/vh37pBmKa0QmOeJ+fI5jVWcVQVLh2Zod
jQVUisfZuDzBu/l+43SFMlWgeBy8qK0d4XKTJLC7aLUn9jPOk7QIK7JNmo1sxqtM
MhDeGWwlQvxZ7XBjBXLvcYkZ3tv3jOLLzgGE+izGaZpdKBpKmyV3BLv8wvYIw82l
haih/GyGnzsvbtimJ5nIw7pi8n048kUwScvSQhBqTJNi8sNDyyeJUfjoym4Xt7Lr
qKry+S0RH2CBMNrUYqMXwNSiTnrQRwSuFXrNVz14trX+wYKnIUqT/u5H/zR7I6NS
viZ2zOAN6iGb3WEPykxBOgC3JGOSG3Cl7nZZ8PO+USmNzyeIDePoWfpKyFoUgZ26
ENP9/ocsbGfP88gHSosSJjbGlGHIn2RHrxdk7TAn4Y9Sds6b45bolng3Bo16OPFV
YARMmjYhQF9J7lCTbHcm+Yd1NR3vG0i0npEGjTbMmn46rd4EwsyONOC5YgT4KJIT
xvie4RA2xGLBzP4mp7JQeDoxfjsTVNo0tthlQONeHzAk+8LRUEQiJQUWdQKFOuAM
Vt/yl9J69VcNJnYkWcY3WR3moQFAkf0qjeLCWGt+9qxwBZOqGOk+oZ+fkd0RoLlD
sB1t0OXEuXoMLdI1ck5fOGeCcWjIsILC0Fc6QO3iCmAlQF0sk1m02yhcsimvk4c7
eAAd7Z6JY41slD28FbbR0dzilaTqbahbU4y6OA+ErKtfFtYsncqrK5n9gt7dzSCf
WJ9MDx/N5snnCEnDiT7D/o36L9gbOXor+rX/6eg2epB9yoQ3eXWE8LCe/5uwxpiD
RUbtXwNe2qbY+1to5CKv2DUMfcPlaFTjI9iiz7Ah5yV+LySApUcBKb/xMIA4Ie0c
a/IpcE+7r1WnU/52RpARL3I0MMPEgU8V3u6qkKG3325F74BGlEkVj2loZljFnmPf
mc03SpOlJxWtwy0lkW6qwmqULbR6t3TuyOKc9WgLwqf3Nx273NldGKWe7MOLweUq
GWbq7LngEwXSY8+BjXF7FU6vulaGomGGDuKqBxZ1eRTiT3uH8tLcUmw38N57RHE3
kHsYsF163aTvtmzOVFUOim8AQ5eYQV6+qah9r5PARRgATVKER7MsJJKSchfEEt8S
WpAn/IBDZ74kbY4yxyn4UI3mbrN1kR+i588dLnWSfn7asHEg+EIfc7LUSflVdG/J
Bcxyx6vrbBH8QvjQ2KutQeuxXWgOjDq35MMA2XGGQ4Uvd+jJCYmrorSbwJnVwZv3
dKnrEDYr4mQuqphz352RG7lLGb95LhgtUHLJTLZLNhWJrUi9zR5gYOLKOPlZ70+9
ntaw/0ZSxgwIcYyYfG5b5ImJA0w5mlZN5tW2kxneSyJARkUwSh4ug7YCdjNIqebj
ffYOaLWkNnyNQosgc0GsixC96r639KjMsCLTjYbqbkL2D4tyPZoZEUUiNf08trr0
+uXj18KFiSweCSEKRr9O0SGP6SkICJb++OMH1yn0IwVrWRssRAWZcAqvOfhxlEZO
BqrUOT6r/klbDhUvPuhRVfT2yZTfdTuQvwtd/fLe+eDNhD6Eb3NbnxQfYAKU9ulJ
SXVSiMOoITmRoH7tVD0aLNgzntqvJSBU7d9xIlavclbK+thIeGSLzCW/sU0ml/Bc
nrvTVeUTlArJDDocN50EFqiokF9mKcJ84ZHuxsz9V+ec1Z02hFnTFna3OWhhVvc3
Tf34//MAuuOWxvA2jvvNTUS9uSMTxA9JTLYVIfug8P7Tqx+ohqGUJL6a7nFg6JKo
9gbRR9SjVJ/CxurCg8FHuLMCeeMn3jPcZTivx6s9P5L6h5WP0sTXx+1BQMWgMW5t
la4AF8NTc5V2hV+aCDUoZwnerLKFKWQrEQs8bbO6xON7zSTWl/fl9qKL16ph5p1S
WJ4pz++fioiqc8/qoNshdXCRu6WW8SkhJ1AWXvsUrvPtyBVuQJ+3HrDLk4wdknxl
Q8HIhbUwSDr6NksYNun6ETUg29MtMYn2GtREnNqnRDOafwflTZaPIG3jRvzZJHK2
F9YtXNXzVAMurbNLXGuT3XEAvV8JgIMw2LvUbQdmzBzr30ZVRNNOMHtLT8tSW0G4
m/TYGlRWamsb0ST9B4oFk6LkNk36qkDBHp68kzuGWje1Q8QVVQ9mW0QdkBULye2Z
ZTe0Ekz0i5kOOHct1ugsaBuiE5YghFvIS91aulnqINWP+OJOvf6/C+DM3552qp2N
aHypSEKDsFRiEYHyUHBnL7LA+hVuboT2ALcJmyDyWkP234KkjBVVpZ8xUAfL3Fyd
9i8jtNYc8kUSvk2k+t8p+SYQB1vxIZ2TyxbTIV2EydH/Ap8wfF+pQd+r5Z4ysPn3
nyAGjBubd9Okqlo5+x/1ZhfPxAfJNpuJkqm1ouCRMzqezKQakTTqJKnuC/ojueUb
gtaoqYGlC3yr1C9d9GwDEN+GO6b0SBwKGox84ZAZ6xa8R81bguYDtPduyeOdbbvb
ps88CGEkPOINggCYMoqiBPzdjRKUn2nOPWFlUjrIbl3wj9nP5n6DSo3E8riiTG43
z4vhuFHl4ttOS5HDg4kwlnSN7NS/NWkACbn01+RM10g/f6NLizqM7O/kp2aMOPsp
sXcs51+vFmUWDcXlDNIqPD6e93yUIhlTgfkhTTGDNV5H5EDoQ9uVnJcKtfSyZZ5V
CRMhBaZaa4EnzGRcL9hlkc59QT0HEXRFt/jw4ctl9QSDKgzH0IzcM5GxXgWlb9Ao
OoooRx39x0Dz2gLMak2++uSfaRr2Whutco9qeOo1ypV/4+EANv6DZVagu0Y7kaCv
Pq0QU9AzZzU8L0qM9bXs5zfkLiEpQ4DlbD40V0JX+p9Vs5jIIWm+E10XqdW3QY/0
poW9cMKJD7A9xYrcx+/F58zIC0B2ULFUyTPXWv1gIhtWA/aVJaOpThGRIUkywM7R
UTiXELdoCDx0farZwWLh7lwnbmOIIwekeSbpLTKcvAv9guMBIde1ISfUfyX0q9SJ
AeoyPOGdCnaAOFi7cLDEoJr6tje9XI3LImW6FMzfzThfDJigjQ6u+LeYCIi/tMtb
zQSszJSuR2PQWaoExivlwx5OUb3DNbiurUdP6iWkHHLq8pQnU3c8BgeAa9jd4tVG
vmGkOcqRLyYtLOwgEXi5koTxeud+y68qSAdDPg+3gMJlQbgu2y/t23GZnZgmZtRN
rG/VTXbBo/kTMRNI4BRxGzMgaFyBM5/+rqni5Chj/DOFjdBpIH/dqogf5C0fmjU8
9WNtm3/X1Pj3R2yh3zuOiXSmJxyKKIgu4/4LUs62z+cgXVysBapvuCcXjnvsn9rp
NejNBujqGhId58GxlNJuTbzphDVKIhmfFH/YqrEwJaYIc/+eD4K4pe0BycJ3YVF+
4eoyvmZykxMYwIespcFH0pZOkynFKeuNXdJS4PLAyYWSmyUIUcGnkTJCYpdKo3Ao
wuXdERXp5V0UC1bRYdEOIN/D7ax28txlPOXIB8dalXKXY1kVt9aguiumQ9rzM3Kq
xVFQrrfjkskHjXBo+oohMdCGBzGZvtYeJJ9RTFPNgF+ZSqzGBFuZnGDFJVdQLVK1
rV/3sfnb5vKEcWfOVAy/YLpg/uK82c2SmTEIPXVufpBTzjt7NwCE8am5TyRS6fmk
m1NHHDjh/tblb6AJDBY+rQdnqmhG4vPgRZkA11w/Xm0wtL64itWVhq03FfLKhR2C
rd6O4O3/uDlDPuucSAbu08NhDtMLeGiEZrQVLxfqQavZsbwG1Je8iWLeKoLfBOPy
qCnA3tAD7y8hM6VHV8b6mo51nbQm/L4fdOkJj+j0mlPiiZwWr+Ni8Xomuhk7uLO+
rdWJ948/O9MD4InFYbwJ8v9VlXUR6mtYcX8ZuxA1AyA8EKLgDt0Rer07PS//H1MZ
TaIc6mCISj7lsiT4E+GqnsuHugIhIvRTTyW1tPcc4v+NkCFo3r7DhmSeHJ2cTuIV
J2eX9F6hqHWzsBP25o/zqAqHc6q9dyn8p2SKF+X9uXo15uk8LUuIJ3EZ0v8a4CFp
PMo181aEIFNAWm6SX42r+OC5tm4w1iagW4NXoMtBT5JWjtABTxdy648QYea6p2xx
zWNVDD03zB3XL+R1goKrSic5RdGJ/AVdXjl8EB3n2y1a04P8kybh00UXgOtfmphV
vOK95en61XFFw1oyAsoITK6rKQCsOaOgYHHJGwGLn/O5NNothuwQzBXOaTh/MjxJ
VO/XrklCwFErE4fItpLewFURgzYzlhCsZclBSCJi8s1Y5Co+DpCe9G7Msj5Mnas9
n4ruYifbBSaWKiKNREF+W+x6xEjVkhxwtmNkO/05oFsprqJHy+QczjwPjK55axuS
bPGhiFB2pVZvD1vHsk/KXSPjX1ekri24rA7hKr4HTG1qoCauEZWAXTJya2Vq9MXG
m0CTgukvoicMhNzObnXiw1icgxditlCw2kQ6W7xvwboz2uB8pBcMnahycEl9aYvQ
9Biqpx3Qms4sNnfsHEhxiFid8CfcwrpLib2WO+H4i6oAqoUAlSB+3m+Cryx5BPNU
NUvD+mfMv7yieGBOS1/ldUuakiF8t6pTe0qcntnMN464GOT5ZsfWL9AMj4ycKGo2
shj+qM8xhWR6/76qySdyzPEwYH7JpSjKpL+oiuh+5NKR53QewSNWOJsHcBgjieb4
2d5yPV6lNkj/c9ntW0iA4Gp0gxP7GquMqbDzyX2M/U/8e0Ipu17XLMxwjIl+wNXi
CdbyBfbwhilY2IqfDW4qd6xXszBTGPPGEIPFNEPSWFt53hateBmNjT5Uq7JeJd1X
Eo+bOpN9GnwQEyiMZynj/sKZ51i3sHyLlHM1ACUEehZiXx2ymRgdNlOS6ILhDUzM
bovA9kI/nv9kpHWi3ytze3l9DDFZJZApE93BreMPoPFbX/+DjMXCwKb74zcxHhf6
UkIwmihYT6cMfAW+iPtrrpWqOnZj84AR2PNYgBnPuhSaea+PnOH4FIUIFCYKyIZA
cxowgmYvHG3jScbBfyxXrQj9iHb5CrwU5fpEzk0GbHUIgbgCWf12+alxa3ikkdi5
LubqqtA1LJmjWqH33hW7J7YgrJcuz2sCgQjjRZY2EVyd21hHPsOvl68CZ1xiexEF
ZuUD7mE6Bu2sonaCZroSk52ol5xou5j717Cc15AxoIWtnDaOOGByPmMiMujbWlCH
wcF8Aeo+G/CPx7KsSwNEgJzXV0XSGrxeL4iucjv0RW4+EVAkPZVO/qEtfMu/LCWE
bJILODbohI3iC5t1LOMd0dRgd6Xxd4cF3WpcsgvwEMmPCUdyENLpzp2hZDUIrQGo
AHNyv7tACQJdBEDjlNzw6isCrog6w35Y/Ulxqy/XDzA8eflV+fZLYB624Pla494F
fbMUPsk1A09gZgIgwtpMcoLhPYxv+8RN9J3wMlMLsIX92B47IVECU6Xn75qR3aGD
cW/O2f5kRNKry09Whgwdk2buHXg5oFgaROPp8lKnSoJFs5DFA4qYEBKRxYAcnFE8
eI69OXCax6r+rH1aHeHefYtKODVaKXhFtX0MxAvli1t7lYFBn0o/+ZXfD5HrcShP
0zyqpRQYwxsHjIESV0FzNWCvlB4Y/b64f2rbZP8x2txzHNX2yF6zTFxdQuX6E4Om
xBRJq6kyyaadloRZJmfAtlhVWz4rvBIW3lKJK4IZ948qATcHICZ7c6ErrLjeHzNH
/e1h+zIG12GrDaPxcwXIaDfT1hoypScm/tVtzgevawyLM1IaGMRBajuQwQCmJelV
7xLcHUXJoRLDdkW3u1qJtFfCM8AKr+A2qlVlIX3B3S7BRLUFrk/Gdo6TZNWtBJgU
37SrIjKBJVMfKfu1kmHi3oCMInF6/gCyOyI3v7VF2A6HJBpK3zSwmIE7ZVjqPhdp
SSTMGWrj+CVw2y1+f1QGaO+3CZRadpPm2CVCTU0cgrIHC9yoxfbVYdxMZ5czmP+u
8tYn0lXNbdQZgpXrGWSYA4VNyh11OFnYGYajf9LweL16VB5HzGR+dPPaLk7U4xQf
c47YH27+Kh1fX7ZA78ZEtHUplerZg+Kxa/ZO+XGmVsxl/LTjbvjkgDWStVsF+KPo
zkRzBUVDzv4faDWEL7rTUdeDO1m1IYGMq2bEtVUN2uQ=
`pragma protect end_protected
