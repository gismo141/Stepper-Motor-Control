// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
V552xbWNcOFnEDww/NOUHLBpInV0926PBcBFfT2wA7SsmJDt6G5FsJXBkNWybDoQqIc2z0nO1PyE
7ZzDWKcnCbrAT1pmd90dZat1knLOz+g1VMfFgW6kGX5XADckeu5XkzeX1eDPe/2QYB03gGp0/FVo
4D2vNmr5vGIp8jkwJ3MquYIU130Bxo9G3xbjfUz49oI4zFtZV8Rloda3YKl+4iVf4NPoZCXvqMQY
Fx8jC2n4YXmInZ/W5x0JFUM17VD5x1C4ibQ9yghbYm+9fpBo8kgY1nIzY+iaF8fbO25kgNn5nzvo
a6s73VC+Cvzl5dSvq0xdINBOuHxGHVNWP04GYg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
hf+TlQloxQm1ZoHwJeouIvSS9dJqzq4mzSiht5v8EFzBSe/Lp/6o3N8cPz4fm9iem2JEKEQ2DJwc
BPhbFX1T3GPyuXirVqTBWbapSuDj9U1ubaDXyfjiG9YDNsoXP/9jzdAwuryLFVkaZ3kvYU296ZeE
QHFs8BHvwhnTvS7r4hDI/bPR0pCm5FbcGlNPKl7S/m7qZkY2t3YXoEXgrPYb63bY7dz4/plIRM/i
xkq/UigO27i1lJsMK1x4WJWaWdFlSG/RgIYJYeEIiYU8ZkL2O8JjWQWNju9zS+TccDbqz8mWlHav
o9fkPuhp+xGT3tAoHGCzb/ZZJot7FTT+VwjtUGtADw9aBRi+Y7Bb2tgf0a6/FmIKKXTWytLiOak6
QfyHZmL50tFneHZMSGQzempQZIWHUVLrXp2WiQ11UHUI0ApVT5Tgi73GYDmsCP6lndN+Xfu8gBg2
7P/tCSCebvnud5aHh4ZCNC12GOJg3sjEPepyjrR/6pByHMnuNFsihl3AKf6yCEWdbyG50jjpyWZl
R/4keCLo5qL1VsZqTMhmPn2U4HIEG+4A3b4BWB/yOFyndT+9X9uIdWC6yWKX+yB3Og8IBbYmnFGt
X2Sf7t26ZGslGq77zaQq2uyHUoYKsDtrtGyzN9YUWPWtqSFWyzrf2jNInOR/s+bIdwHJGaBceP7U
I6iwmTBxyOz9ZGzk6y4rSENxZZ7CkoX8h3+h7Y9Kmv/0KzHgjZ5ZTMVAe8ntMjsa+41QnXy6SKqQ
Bgrf8Gczfp0RaVKM+Z4/PQ2+IonacGxDXSyfJ2GGmwL+9yyn7vMBsC1Zgq2HH8lobUGYxXSk2Uby
0xYm6q7rZFIPCx0Wi5j9hpnHYrt3Hs/9a5h5/UT3dcTYRk7k9pcB0bVWEVh5mGZTe3M7AmTXpSL9
/3u+Y8ka04WKcy8/DBOuLiXG96JZELZ16RWolkDPxZXTLmw8dWQMsTlBwxyBv/QTmf8YgfsLCggg
/j2wpMTmshWZU9RlQmyLfYuRA4ra8RZ9w8CsMpqodzXK6g2B9e+QgmiTG+o8H7ZQKZK+e3VqZMjA
5HwRtovowL3sfK+b//VOrl4p0SXgV588sLV7WFJXJBYCkz5JWF+6oNtlBnz9b8m9HJMf2g0xCbLz
S7c4kKYKlrlzempXGVU9OxPEpUXXqLTjHoJtq18H0TqqrOz51FE78Ap1iTZbWmS33+O3cAw6luTZ
OS37RSpYwRuX48HWmcvHvlpmG5xcXi1Xo2UsfmAOA9vn4T/+QHOgZIngRe6VOWTtsoh2d/AJPeJb
8Af4Yda++1LvF+CqX6lQIscvsF3J7UmZutcNFO+0LX7rogqyNMRD0z8km721rG4Z+jT5XrM0MU6s
+tL13O1VHLWow/n0h4w35LrkQjuJU+UEctqRmDaePJk2uOjAxAawVd1sYto7NOB05jlAdT0JeMq9
kcLzWO7lYye61TfxZ4IU3jZHJSgq0DUkAsS2CjAB/578Pmve3ht3BwBAZWhAngbBWS4eVfMtuvUA
BtnXanhN0mBguNTAUw6HhUa4g+bBYzlJfCFJNd7XUllQH+PgaU8m7a+Oz2lidKS1WZtpkGP+nc4g
jHnPh8wO6kmmKfGFE/LQqK4EGAeW/F/Q6g9bReIldgjDfBYvsVa/bO+TFQOgm4/wfjJ30ymr+cfQ
DLPQ7PPUiLgYjXiIMy1rvPsueXs4cDsG7R+hLn7vBm8rTAUyWAXa5BXGdRd5SOQEiCwebTFLk9h+
JkYD1bMsdqk1T+3jFeXzBnv0TzClGYaaQvd1x5z4UE6/avc+gzPzPsY4uSUTHG0QtdWhVuyFsHZ8
cy5ctantSy3+wT7FBBB/FJIlQnUQHGueqfBUBbDW5DzUqj4FRbolOtuySmnDPIQJExG82lBSJ6qb
jyqzYIJuG3ueBlnwPXPtcl5VmBc5KTjURsvlMIqmzNM+xlBANmAAOcrHqUkkeN3kSz0IVqTFG83k
bIs2/Y9M8EWy+HsVH6IQu3kyMP7AKsnsvh7ieIH2rsnWn5Aib33uYxSjKm2N26IhhOuQVqsCmIX+
yYjQfm7uq2IGXFeduT+McPPEne+JjP1El/TQq6IQhGWTc8Tt1+aJ/VNO+iv3A48cAZtoQhmrR/lm
OLa4baRriZfooYbnRSpVyK83s6dABJNF3KdUEHP7/W+qNOfJ7C7J68IVEFmj2BoeaDhkHDfzngL5
5F0gQ0mkrJBNKv8OWKG02sLUZEan/MaBpN7hy6dlusG5oMaDUu3lR7S23OZSh4bfI8JUxtiaAQrL
YwUQ6zlTXV68rKu84NCrr2DC9DNoSnnn720rzKiPdEWwAewta8SdwtIO9peOniM5V2X8c0bo+5eV
FiqxuCtlt+xzIntCvVdJc0dJsudYnktj3IKC7JyNdPrz7Z/xQJfQeiZ1Jg8e9wCMSZ+hNoI7aWiw
zC1795dlS1KzC2SOGu3qMlaAl3v4XF7SBKuitW3GLiFO6bE2wqBOuahHFr5dK1VpsdpGytSn6eiq
AdYWQ07cvqrJ09YEiyENN455aqyJPwfawujbOIypzu86yV+YyFanMv/A3A2q9VyLR1RbFP6P+ru6
9v5xQxpq9GFU3rZ8t6AThIZrTawGhnnJEFRRYLok1sW1R+Bc/qwgpxrOMLy1IuJJoVisjBNLPca7
PpFuxk2jO54VzePLQnnuTIAHUhZKBBOHW8S+H7HJa3CP5XDE2a3DLcVGOVIo4Ok4PKZ5xpj23Zo7
1CX/WErXcDglL1+VP+WjfDADLBIGFT5fIQ9rkXK/rGzWGBWxJnBeNjkqMDqMJT+6hHJbX3bFnXQG
T8RO1RHgkUOS16xlNoAaDONeRM0ZWIhnPx99qx1VX+cP4bKf7xavjKeUbd2Hnl61KzsOdR/aSeg1
ZeASoqXXPFJLCqbrdV+xmUazwyIUoRxp64CgsPpu2KSsN+Y1R5U2arq9CHjo6Ey0ThlzH99ZgBUR
90Pa58l0PAxdCByCc/i1fVb2bu54lk9buwqT3YDeSIQDirfmyNstaI2xZpAXG+x9fxWZI65nixsj
5nqY3oRnoDzY1aHZDX/E/fAhvw8kLq5abG06+MJ4Ryep9AObWY8Cyv/uRLhI8pSrAX+BmZ4aFGVH
V1kClB2J5ZoZBiPhbW1UuRBNu3YeGo8EGIXiiG6Q/s98bgcP5L0FUJZ9rhEECIbHdegRnGf5VnFq
lEYsKbfgp4Nbwvi4ZR/STb9lL27gOxFzfQsflsE6jrVazIKbcJ284vM+fQHEJT5JBLGJi4yVWPkT
6KzzWEUc73uStvQ3DI0LJjnaW/Sx3taPlktg7t66uROZrZKhi1ZWIHr9keoDmZMo4G27Pq1d3KOV
avB0o5CBrpP0kGTM0HOfITOFo1M7FJtkl+bolU1xe4tocf35FyQT/CUUaLmLptgRbUKo7Ax71kNx
KD6j23Knt7Gn8aoqkE2EeDA3vFWzRDms9/Q21Ly5zIkdj29y47O/1H7BjlN/rzVTZAcahsDVBd8B
cmvxV54YyB8pLx07hxChI5F+9jnkwlWIOnTSud7sBjISjvgdhkC3j39rSKjEO5mNH/djNlSFpVSn
xYIkEY/6D/XmrvjXxC4nUed1d8dMQODNm6fH4bgxkKP8e5oT2ZAWnix13yiz6llpwaR/uQ4cIY1+
lLeMqsURwnMhb+nJ72f1yzS+Pwojo7/0UpqMMCgDwclZnO/FAW5aGCq4a/xCzi7Vad4/fEC3tL56
TbWV0x3eTEdVtbepCxPz9gtGxi0RxXX64e9i0csNqE8ZpxYzkrUrCcrL/KtrjCwu9RPYZN6aMaqp
2B3BzK6K69GKkRXdHvBsYayzgQ23QQTaiVGzWkRCbBusQVsyi4Z33KmE1QRBgUV/epDvnHpFq+8S
SDxdm3ErnE6N/x23jHjrwaQBqorEgclO2OPMauaIfL7VUmBdNyPLIvtdDrbCnw1RhHERwd5S1SWL
kcTtdsKxPSYiih18CczLmg79rtqWHH4ZWHfIrMT8rw7jwQU8xu2Cc7SxHBjL22uEy1Q2n1FCx50X
Syx/A15gbldN/NjFx91nevc9mW96j1+Z0FASiAb5KbBIivq38BmEI9MeKALz4t6pejJ8lsOtXAIU
PQV5QcLb7aqMPev8evFKxcMeZsDW2q++hecuF9o+nJfcQ3v88ibFD1IQ867HWgDNTNE0csBsoNk0
0d4FB3/zeeji536TNjKU1NvFoCoSUlFuND//ddn50asFc9qTdta6i0oHiIGQ5knnSjStnAHVx2Hz
ZRVVxx2+y24rbMW6/4U+/++yKC6uVeo6Tr6qURg9AghOWeC33CZurkkCNG7te6rADeGKYF5RkeKS
pzORX3uStuZ0/OpP/SU7BzQSSoq6z1akg6DvHSt0NzNiIdT3RuoV6rjZIWZtxyORCwb8ZWmovHRE
Qu2ZUiaiCUuK77xmrMU+A2ShW5b6IA0wUpe5LyJ2yhhBGzL31MYobVPclHGmC6MYqB3QrXGn02g7
AH73u7WDRkp1/noK7DZihxamrvB3ahL9/OMijFIGuCULYFjT4LteSN2rYEAFvxTMwY012h5xTg8P
Mr1pRR+XDna7rhMc3mpmY2y2zrIq+kSbiOIudzblFQQ+9HP4+E31erS+76f4cpuoj6stZRBqtuCl
PR/2xYvSJ+sqZOA13IdEmY58pWBID53vblpqDtHt3+9CgMUBU/BZCDB21P1VfsdTVboenZjnZGqu
hNapN5Y+G8KD2SXVqujiWejpqs6ZUesHiALK0iBBBxyekb4D0B00C/R1HLbEB53JkC26sbCTPgii
dJMIOpsEKZ8UFO3gYf+rxIXXwG27qKE3wEIAvvOztzyeYZ/uChiRdiRwSI2dsgyVlMDjdXm7riP7
7BYfaCufe94bmPj7ZKmZ7r+1qoYQuonPfPCxtFVbzKFBL6G3Hxhf+cVGQ211OVJ12P8B/rADtZQP
0aag+F3hPsbHw2R0E5d4/w/CzxMvk32aef5+dr7Fg6RL5GdXMDzRuTP7u2RqiaKvCLyBg892jJfZ
v+sEwhA4vs9t+X5ZvEsq0jlKiuUnQzclqJDVDRJP/q+Q9gCPJw/tr74SBPGr2KuCqjzVJr7c5YXa
R5CwT0KJWKzR09iUEdGBQU0WsdvGqe6JdHZk5NF18OCdWbyV9DGqvwx6VLgfS9c0MN1jxeIbn2Kb
O3N3vA31GLrBspnp/z/VHNF0Ytl/FOmm5KT7Xv9TM2RZod6QWlyPDD1z5BKvqKO+azfo1olsQFA/
T3ByE+PX9mGPakPObr65XyygjQtXYv4IlBk+TjU6FQ6rEFHltwgGhtd6rjUa3dVktxL4KBEhkAlz
UoUacfxAD14TzW93oDxb75jKfkUH189FbY+WQrhLND+Xz6bc4S5NF7FH4woHuBSNxrVg2s772XVp
ZjBhZ+mrsGsj94xIyeubpIAXbmsmZVpKsGRTEH61HeqHctwhPS6JtkDEAO5hHlrBKvRATjD1LPVa
iFTj8DF30tpngls5FabC4ORKYLsQ0P7grv1anwW0nYudkCZk3gpEgjpfnTrTtZBgd9LMR+bpxj+I
EaYtf0fc/c6orlETHlzznR8aSc1Q3Z9voM9E+pp7rz2zvG5EAwZK4cVgrH8wmK43oXulBz++OxqP
kgKwuLAL9onfDz3Cju1LrqSRAAm/o+1EsEPGxeXUX4hDPtTs0Y500lg9zBYEaO/0oeXl1Xo5Gl0k
VdiidCxpl/rPDl7lB/UxE4Sf+AwYEGi1Q8/dFTDF/8/y56Eynz0hdvqr4mq9PyJmsP2I080Lsar+
RRfJAgclTmuPsO6OWBEqrF57z5SeyUhjhvCkmGv/CmnqvkpfBAtOca1jBJr/zCnFbdx2mvqVPY6J
fcKMtF/2/K0kJwi8bgyXH+92xHww3LCp6z5Nc3Y/8RRBjIlyBezo/oycTg3SJg5CAFmQ8Hwj3uWG
4TuP5okxBbHP9RzUBegXwz9Oy1V5ZiiMrSr080k0y/IYsj6UgJvuJGHwWpxfjISaTGCr1Ie3W8bk
XNvYhUU91Rt8/l9uS1YFd3rafaoeNPhonZFEnfIMnb7kkCcL0oVDwIe7xXKTamcfDzKZKscLqjFp
w+xHnp+XgCnCrnDsgrfIE30DJnMmCwC/e9JGXjyZmTTVin5ojbQHYqGz7s1/3VNxxuEwqGYSicSV
4yrQ8EpA/t2xAwk384rZRnb7bt3gwgKJWDAgbHh8bc/DaspClbCJseu3PqyjREQ0gZGPdhDX/RLO
24hvSnnXFl0VcNPOOX1v8H/YiBuy4mQMts8TNqw/0jRnsJrFPqIphxel8XGF3RDNlYSACbghC4mH
TNBiICcHI/Dsebj5BUHfibzmMDWBPS29K4wo0ArW7hD1OPZiX2CoztitupBMMQ2jFHU9MWhVCmb7
uWrmKYEIzjPnP42w18EGtjXbWYEnYPXSzVCT+qZln6H8v+Igou9oCuwzQd6MkrTMlp7U7bDog8ff
WAWUpe2jsB1uWXO7bj4QZmFdg98mWHPNhDDNsVtlF35I/dX6m6iL4KX+H8cIsQjGqzFqHC/y0cyX
9Q+gADr77y+DCR9nljfSsuTTTeOQfew309Ls4Z601ZCV8bJh5vKPZBLyw6nT53+KfFRupOw72VLs
KWgKYMB3al2PUNKgAtZHmxFkdycbeR1ZdfS2Re+XieSVTL+pd09UcJyBQBs3xaJD6tpAEpXvANaM
GppZs9qFENSZmv//boFuAZJPqGSwrDyes6aXJgU4YwJgYpMUNvZ8BAPL+Ai1BxjumGuEKs7hNrYs
BPfnd19zFFYBVrCL7fs4T5JirIi6LOzibWzf33rI4Fv+m+LMOK8HsFSIjtI4WepjWG7CoVi8Zzvm
o4F7td4WkHv5UjesSL+0N2li+Pdswq5Iw1ovxwYi/d3/MixQ0nVH5umMYS77lOCzQgMjCmZOMFom
pdN7i4eNCG6nMtmOVlKOHpLlajfvf1avtbWS8MtQufB0/F0P05UxJtPSWl4AQmaXF1ixLIUrbNBL
bo1hzHen5j0Qt48q5/9CwiuTE/s421+kxi2RvmkwdulXtWmPOB5JWziQGL/QIjOKqfMoUvzjHeXc
Cz8kgQhjMBdqmzmL64zNlx9Gc21sy1ksTc+OY4mf68QJLqUdkx5l/5Z9ACTX/XW1CBprkTfO+OjH
gxEEsBV5X8tyDQ4/qS4d1dwW9ftzt1y9WCz27/6q9zLNFurRGtEABYzIAsUkRoBB5ZdS0ZNqBtVS
ImtloUFFy7B/gegEUggv2Oc/EaMBr5Y9yKdEnhdy8r6de5zTWQtpr1h3ezKZWszNI0/XiuJk5zi/
V9rSL+ShThxcGoZdehuVfz8cPQo36Z/3ytBp6miKbRB+viFpF+fKITSc6sSolBMPpgkX+8Ln4dk3
/Uzsz52/iCnaniJ/aH6e7Cmpy+qwJuL18rv9xXYmJiRwEu7M/yyCzjU20I3Nt86Ttbl0p0Gimi/L
/dB4t096i9NZcjuOm6SFugBxKWZB64QYLunSyC775Gvx6cCmey6tFmg4M37Fq/E8hdedWZ/zpCNn
OsEsOjP/nN+W3HfRf9r7Tqf/N2AyJq6f/9SjFN4sX0fq1aLrtZobWvuHveIEd5K2mctNZ5S71JBT
zgSDq9P2oA768AD51w2O107TL+gPlO28w7dvcNDprjBvTPshB1vEr4ptSf21tD4GOKz6ZSKTUYDL
Uf4Exsj/j3GzuFlz/uIUBpIGP682g/Oa4J5XDzJNICRgeOsvtxso0vT/dePNxIgenuiDWm7yf/sX
pvH6mzLmSQoylFncIvQztQCVMcbbkRReNJik+fS1P1RNh0gkD0EuCxnbbir99bRX8YD+6cRmNWW7
j1hILUXXOaL/r5We3ABknntdVhuTyqd/f+u9SPXetqwv/WTy0ubbul3Oai8utEo1jwSkFr/2Stni
0CkglwX7s51L1uNKNQ6gWomPoJpB8Slmvf0L3k2GTkrPbvN9KyJyhVeoxL0yw841v2fNVCqzEWh+
FlCraFOoIqNluwCUlCb4PkO6hdeUPLv9W/a8emkFPjiVXZWnm+Y9UoN58hLxqmkrbOLoJ1q1tIWa
fX5akKV1oWPff9lCMvS7jFKUQbW/5YwPk5gcGp4aylTuL8c9XsdWHn8SU+DGWf1wYiOHL9Vk1zPV
DBXgHoGjJB6D88yOo9gvN3IQSI2eyLlgE/uYaYQVeCY6Ry1q7puZtr3b8MK2eAmI2MPB7v2dIfFR
8w91yRxBhKxzx+a3l98xiCGyepQhixh9nPhjO95VKubiCAZGdSMPFUrTskBvddckyvU/6pPvEbSn
lqnTyuklmULz+SBjNw+pXKAQdBJLAHORKhJr8oOZmZtLyNcJUOpYpKE4xFKMCTe3eno7a/MwiZof
osy7fxqfHB4APyJS8o2eorih1vzk+B1/436r0v99QznUZBowxjtJVFvJMhP8U12X4YA/cA0ShZQr
/TUv0+MOXhYwtsdSVI81IBG94zKtT1SOoA8+lm9onbPWehczZOeF4JYcJQCigMTlMwlQVupugEo4
hg2DXm48Hk4l0wamogl26j3QsZ2ZZS9INMGKyNqFCl/pKQgQcvLEvr09ZTIeLRcaR7psZG7iotkP
CeDVlqwp8jMV47fCXJxs+3dWx2cg5CGmol7mDO+r6oMOOFIuYLTD5IhLnoDbzN4SzmiLHNDycNmF
vDvRhFylPNo5NMO8rhnL0GwR0LhXN+dv2JYL7I/9QSROQunrmYc55gwuq2h/Ai0KnPm/S1EwdR2M
9VVGw8HocoAYjXOrRcohI9iwVAKNH7GaMvaiqthPZrWIMwCR0mr4+dFvfXL4Fl9A//8fk9uK9bpJ
ukWpktZqgpoJPIKffYOqeQJNLnZ1HMuB4+IdYQAXkvVHtNDOBfcfDvowXEZjvFeaVTGe6IDS7Cu6
IQi0kwm4RtexLDDOX4E9XaUwnAPZk5TJ/3EhxzXuDNXVduWXz7fqRCKVeKcfj8Q9/pYDagCvH8Hl
MS9NgHk26Cp8J/V8xG06K+A9USMbk8LmvJTlbIr0wVboYnSoN+3BGCj/rHWJZ3Ad5GbQZowVRFvf
syHBE640qGgAZzdIsf2XRujM2G0TlP4E//j9zu9QcSTazWj3SpFN/I9NagXCDVqh2MqyDgkTGTkR
74HFuCd/Eja4i7zrDBz60J0N3jlbWvgPwvqUB/ZRbt4W9f1ODUENaHs/FHXe0IrovZCuNu/VXR1U
brYF9FUK+C86xn0CfvQrhnxSD8E0OzEhno+7N1D3p+NtejwpdWXu4c6HdcV+SpmMFk8dwIGIqb8w
yksC1wBSYCaREzPfoL9+Xut/JDUTZRywnHm34eDgpMXrZxdpB+xHtUlN8kQGAWb9bq7qC/odxdDm
V6L4iRYzdIKVE26cS6cTGBx+1Pjn+L//qtADssfPfL160PbO/oLYhUDdJ7wfVC7Lg6cMXus7ztAz
qSKpJEBHovMzAkFlFGKWiaP7aRAd+xlUQ8EaK5vyyHICdpAxWdWMOqHamv/MMP0Cbknu8z4/STfE
LbZI810uOkZ54GjB2lzkwqPNbfCT8o6mRIA5EK3Bd7+WkUjLxDLWDeEQS68NGF1YAJN3bfcvbuJl
zyf/v5nIwjYG6O2jZg/T+hfEfC0DPVEo07TcWbrXHkzskgfFYIVyrQotXieDxskebuJEy6FOJB8p
IeVvCR9mOgC68p1fJctSx5jvQ42slj/Ovpi+hsAs4y/tLujKvvubyCwyOBK4RXuVKk2tPaJOqIzx
JR1NsSG56fsFTpMjVa7yAUksgjJWSQXamELEw+riNC4I/ytiHzZacbKq/JCUX4UGtpYM5VJctd4n
p189V8lm1EBeET/vw6GT5nAU4flYtxD6/FBv4PaYRUDrF1rUAeOFff5hwdSwH2yNTWQ/5sIybBTR
Pibqifb1yxawKHdzAjj1YrSYVEZo3gItFk1avItl7EFPmVFXZNa4K3+vrXpzPZmCZ218yVtJq4g2
yG7j3WYx6X5pny3FHcSz4BTiAqVf5lR2ZiloU/bSvYTwPT40Ghgu+pKv8njJzuaBSMK9tQ8YQIUy
tTJbilHiU+6K+Wbt3qCtg8VTX6zmoSlD/65RArvYwmggAmOtMTexrw19VNwkfJRFO2ZqNhbaQF2e
NmieGKtlJV+mgpEtBLqhyOzqrqiO3I8B6UQIE56vtF5F0Br4pXwWMwo1FWSI41RjQDrzok8/jffW
7MFQDeMnK5LbPaZIrIZt0m9cyfYiKhkjVHZNPP1NgE2hVyHXbQRAUxv2tMoNWxiLSXhj1M57kL9e
wL7SSl4oz8yxF86tAEnOnZYtgpPn9snrfIjPjHrdHbh5Ns16YyO0sanj+dIZcZ3ycEB9Em3+3OmI
2ZR2xM2PFp7SIMb5n6+k6joUeBnGtde3FBYOBlM18WlV9rrt2sqwUx0BcvBjMEKvtg8MlFNYJO8v
qVOM2WhW1XVL5uX4HCaV1NCrfIfspf8YE5WgH/tSylFlKgVAOyzLHqgUe/R5fq6Z20XyPLDAw+wV
tpBZob4Y8oBvFP99UnQ3vWdq/CMpbGZvS1MaxyGYx9NmfxOiP4VrqQA/kM1xbdLVcpQrjLbIu4Y9
pWqzA8aGIIMWVcqNKBbJltdOLl5HDJF23K19cuDVmjFBcdA/P+Ighk1ye/QvL6geH8TlGY3jHRGL
8tILdTcWsxHimLChRWG3Fo7KwTm49G1xVMY6ugg6FjxwYr1MzSAyK9bnBQcl61pC5oXuUJJ30K6d
GL3LWhOxut/Zs8zeoLtBa7ywR4SITsw5BXZyPAU6jTeypgS2MND4xrtJpatToVegTs5Pul2ipl4E
Da2D5PEgYMRbl3uy4+5//1nOOlSZV7Ds4/Rh+hF10KCC9siOk5mqTgIETk1ulkhLnVT7f2aeMarH
tR1hRQKojjwtDe37twvvOpg0akv+2DpNC4SQWl4Bijov9bCi4FR7Nbtb4l31tAnz+iKJiogXJtu9
9H3wp33iX4ZAR7bqaxfILNwhS4QEwIMHfGVg9uLHzIbfNEkBPx55vU51PgRHal1m9BGrwdJYfY/l
oDgaRwFDU1yX1P07WRQ/f84ijbOad8oIo7aya/Dv/N6CRiunz0leRiJS86cpKwximYYM+PQbOb7i
c9Uc0NCxNYduR/6IXrIeIdazVsTlR4V834rRC2SHWRXIXsck1oDkeNPqMhU0fOT46n3YmGYnG1Hb
4KNVjE/4s8UQeJFkjpCXEFmaWhf7Cyj9fTEY0m97/ZNsMPYtkaSVK5NT9uZSCDYyA76Wd9Sx2jpx
99mzuczGKa16mDZ//4vcuU5BomIz+cQek9tuU6qkmLstdMajiMPeszCV6aqeejykz5CwLdJ36cR8
kfyG251v9QWH0nUMz3RV/sarCabKaphtCig5ifmVMJWbaB1ZY8e5dBfoWpeD6gYunYF7sbmyVEcD
PpmeK5NIEopdSXbSMBzTOZ4+A1Vg/4Jc0m+ysvdv9SMVZGew6rl9MavHHTuujqnXjjMdOfG2zDGm
pJORV8D5hGxI9fkunGH0cr9sQ/z7+InKFROloUh+EdnqX11OAtzGCPIG3Wgu6fnQnm9bbbyLrErg
4f7roGS3Ongs5z2LafcwyIP3Tatg5aMUOv+sgH6U0Ytyso3xCQvAxutuyhfhizenmtz66N45I5JS
zR7fiug44bCFXoxWk3z0xTm09IX1/7PGUE4RTrJGIFUubu/fJ881f/I1CGlU+X/gUH1Vwji/xe/g
MEIStFBjR6GdPQnBIDBEmdzuY66m9kVAw+xVh5+CfBhCQ4I4viwxvZEz72y1Qym+w1D8skhm0vqp
VkfN0xescrp85ee+nwDajoAgSnl4XcP5CKw36Fq67UIETzW3l8G7PEwcNDg2o1152+jnUI0f18ax
VQjkfaJbOa//VgxwpJpdIFLOM+BxOJ9BSlCdc0ZzNruqAOfiJ6chfWBzOToP7Dv6op6T1+/Mixpn
kCNH//eagDNwTnum4HPcaPNqu9TnSItmC7+ZY/1ul//tch385iVsPIsWpGJZU5GkWndRQUPElGCW
OjqscI5yjY0waBnnNVrz9QmA4yxUtwiq+zfWqrkS8dfjivcziVQqkL2FhL3GEvt6RQORsVla1+/E
oiw2UClD1uzbTyZKQo09X6UKau6xWoaC9C6XPi1OPT5QyHpHsuhSnlpnNJrnn82B6yShxLQQ4QGB
WdRW1yY1L8dCxhp9QFEPRoMBCIjltt4PiyCMyESMyVmj2o++xbHM9gs6tmbwrrEzcnyGPyySWdvk
8w2jC56jr/hrAOK4BQO7cxbaeYlcW1nVpK19QItQq74fjH2jQil1YX2gLAOLpyb5cz9wWsuFv37U
TGYYZd7W1RmscSD9a6SBBgWeOHqFzdh7ptdzzuEXeD6WlSm6+t2tVIJGnKhfq02A6fKUKbhrk4Yf
3tGykePbr7IK4WHT9zBzwQkOMmObUP2xGtocFVnFRtKu16AGZYBuwJIlFNJTlX0A0oT5siI7bzQU
2eMYKYoWkMx6IFkQMeVrvxbNgTgzMs+aHj60bLGbQgKl5x64zappSn1lrAfHov9UOrVlsAt5SUNb
n2+LbuIZ5MfaYapWh9aIhi9zNy+PMvf+E2L9Zf8emWiBlhbkqa1uBzOLqM5waGeLkeuoXEqbtfd0
kGXjsOxhGoaMkh9eYbDF2Uqjg86+F5NP7M2GwctANf5j42qEH1CndQ3K4pFGn0awwwlXqpQg0UMi
XhHesu+JYMlwP3wSbyzhHbnmWcsaJoRto7m03kSAFyH9a28w3PBCJ8CYLMjhIHAkWCZA3yOwICT/
F/KlgzonccCDNXNDvBoJ7C+FYNgM/VPgmQy5gHtMBY1sLoNvKnX7gQ9j7k7Z3W4qlyp4YEoaSs/s
YXOlow7Y1xZYn2mo5lAYXtGlwoUhr7ZPeIOZopZ2wlvnkCrRQRoct4UnzkRcrO5QDRXmNTyQ1lHa
Kv/Rm9VP1lYhWgBbPOu7u2PvebRcTxBvqm73ZysP6IM0XmmQ5NmgbIfD2V9DLhG9ViKd2IkI7StH
FfJXUpSwGby1ENtPkKdoMemNFWqyJBfMHg89zyWbN22UcSMuBSSM5nxAcLKVpJnXJNdgOHnj5Oay
LsIabu7fg3pMrNEgudhrAvG5ujYZUoLm2oQu0CnGc3nxZWgDQkmtu3xuDUk49kyf8JUm7+iUj1ot
+e5FQUlIaqKhdgKJiY7jl+6F3ABR7txXtapWSH0y3p7wjg4xbfMqIK94SZ1TxXJKSrcIWvBCBWFG
0o3NLpArmIjPGzFRgNVzVQrCkwpmgfzocGikJ08nDrmS/E5iK0oZb+Qpe6Ly2s0Q4FUSW48xp80z
e8Rs88/h0Fq7sBZVuI3tOIAefcZ5bGaMkFfAKz1AlSAC7EWcVFqZAq1DwYAs66mXWo8uyzlZumqZ
qrGKeu7o0xHFka+3ioIyN28TarntpMxEcXRuXNggqaHyn7MkPFnguoZKVp7CK2WdjSm71AD5/GyO
zNJtZa9zPqTN2S0pFeAwlMi6muhWxCvxY/l4pmb9zaIPBVUvKgiaWZgpflxsdpM+WGDHltWNn7Sc
PyteLdWDI0VYPcty2euWAQjT3Ym+EOKepfuEmj+szwziRDXOglnfJKyIXlRYVWoYcb3hz2hP0PQh
5KYgng7dOOunqGcVBS4876M1KdsYA1aqEyGbAt4h5tsVi7czqqFEEpFXAqjLdvMa2gVcCRRUT7fj
cjrZYI+2xmtC3DMYvc3XShowf1shO+uzTWDiU3WkFYkAStgo9lf/3FJgwgOCboyvCc+CBY2OOJXs
1r2t/BGbKdhAEmPg8ihMt7sDePnGQPRPyPLssZG1AyCAoWaZRMmAbg8f7YK9YXdau5RTL3N5kUBM
3uNKDwTDHkyeTotgHxIcwdDuz//3K8kqSRp7N4JIwM0dfjiGtwSEv6dEsBrG/IjszisaU8Xe4Yul
5CLp2S51/yEXq6QTAgKsolsWNcO6VcytuUMGJxOfArlkIJbpHAnbfQvzsKMmNmAiR2MUY7gvyGTE
8a5I1TeVTil6lb/l2F/ewkjzJWwitS1561ahxeV5arhnrA4dGEjo2uoQ78ptEMTnpNU31rDyMeC2
yZFz0YsrIPJoW4qk9jYrPa0MKCPxYstj1FrLuAM+YqK4dr5ppa6VDs07EnCEjjAZtwfGF10GeLhq
xkaxpKorRp1JWVyx9J9ls/9v0KaWu3IuV5XabAhX5X0xy78DdYVTB2NP2L6+eBtYZlb5bODrWcKM
8IXS+VUZav2pJuj2yoL/GbWRtOL0wbaVmsWLZwfZtzB8ihmgqu7ZveYwtAbIhOsLQ2hOkilhZn72
R5RtfSVG3VE4pcVKMVopET2+rAFvGnr5HmPoh+AYAYMXTLIehaQVAyRaJejNJAFS6aXmRsGVz5eR
dDLjZRS/vdRuTYFIpMM4WnBFDwjeuC9b8+IEI7SaqjpG0AfN6s4WIAptGC3ykVRbC11ScXyNDMWn
Y+mIcBmWxpeAzddl1lzzo9Dasu7BbERVCmKF+2vpESxyfpXcHpl/tFKl2jzuBHaeNMkRRNy0O2Tx
N2WEdOMm0GJILrvqvHLAapPP5Lq7ks7nqCeHR+fmCox1Wll72qvkbq794mTHXFad40yn5kg/fOx/
aH3vzYMZCn6XzyawAbMC4mWapI/qrZo0GBOKlLsFMHh6mggaMd6W7cU7aUWc5hNbCUS5o7wy+8Fl
7wAsD+Rz7mI5keRxCmCFtUkU2RLpDbGGAWIGgeWMSFzLKdbUwtLSM11EgiB62dq2VG9jEHB2N2Y+
ug6c77vexrmD+yYK09hvskp+qv01wXxbd82Y8OnMHMYhAdc441Xvkx1YPng11qNqXSteGFBcwiaV
gMsNppYZ2Dz9JiXQDx8roeJdNt6QRsfyf7BL38gkOtQZbid9D3oizcUl6TQ5Dj2YqNy22QDjTFq2
1KnLR4J5tUUIhZO2xVpPdyAumOY1YxCII5cCxnh6QSuf21PVgQB+ivUw6msgJRNGyNFxIw4BGGa8
WOOsVPvB7MfdNBj1mHPUVhJ7AJgk4UvunG6Hv5/5pGSvqlw8ITiEG8RSNRyao4KsYBQYhT7U3Sxw
ftjRURXCXcHwa3XTKegbyeBdQghjMC79YnQOIZOOvODPCWp/YqtuocANZFmwSImqiW2rUWEzGqJG
1mUknksOZdNZxPxbYurBUoYT2aV/WN0/mDx//9ChXNLzslSPaXsojQYNXOWl5YCJ0WTDbzftMfWv
I952TM3jAj9SewsgSwSBccZiRTIFYjtnejMLrNJfzQZrlqUhZnyn4rniquZpZKvkNheJm1igN+IN
GMX5Uel+1sViccJ9GQFdTjjWBVmzCHgzuz4R3iHuGO2xHywsSFyRBn/XcZ3Cjer68R4pDsOUab6n
Pv4ZSsykqL+kSCtqW6V50pBcVMY/ratCHdwFrY+QxzpM9pweDv9X093YRpgRymcnMHyslAJR0Ns/
6JSq7H/l+05JmLBKFRJyXr+tniu3lQ8jhTtFuLKGCIzYfXBQy3JPOn4j3tzqzR4PU5XdQB/byHa6
JKm9QYZauW8kQ6x+lo9VM48t7y0rC5woh4OGCQRPB5+qm60EcEJO0eDCsgxBxTM4cN1qtpOtFDcG
Cq7czaLE3rFe828QSawWVh8diratqxMnfhyC0eQ2sM+HPekm5vN2DlejqyUWR9Gq/pPBS7sL0wpc
dVu/mJqVM6yoduvymK4dH5rzBf/VJk2HrHQEzdrKziu7A4bAM6xoccCnJc4wIhMxwpCb9DGS7ZPB
CEPpHa8ChdY4ocBlRemlgQJMVl4hLSVSp2595DOZTjgwUqDUl4dSZ47KF3kf4m+XRmY/nrsm8ObJ
5S0dFy+7fQDRQZLxdmxRkHwlrhiWYU1qOfc13KQIjxotS5UyaMAuMvvy48hfaa/CzWocMcPra7jQ
PfEMjZQ40sarULb4pk49YskjD/D/SEW/LzHJ4gLmFFRfjRkW4CluSV9C0F5JpxLaWKnfe90bMQeA
PBRCppH1tXhUfsYPiI1PyiPaJ7Xf5Ho+T4SH2nd+rdCIxmyQEWadB/OGUcHXWURlQPWWOvWyqpjV
6xMAsrOJIx0HUS2dAkWhiiPwIggxbKcyIK1u96MGC1ki6Iw35ZzhSkcf9UmGc3HvX3Yu+JOO3xxA
yNcMchJwpWYEquTDPNcod+FLDuDAfxlXVSPOrcjP6bmmCPOSzyl96ZEUvFR2vhTWOPwoj7smaDxb
0dPvueQbXGMZkLkA11FU7KKFQ0r1e/7BnoH8scf531vVMpnrxse/g+v9nvZoxYmlM/F1nmM+yZav
PY4WL/KYQRfAD2qHUFEAmqfZpP/eHbdPWFcD7C8LqWmUjHSFDgqzPdXIOeGqwANH7Gep3YIAQd8r
DYviXBy6ZiEWdWYctocmqGf95icnGTeX2BlceFZmdBdhO3w4inbjE/RWJyUaXlzZ7kNTJZMq9riF
w9Ul+VDdvwskW+4iIpZRbwVPbxrLLsLjXZvwJ28El0eXIQlUl2UnBo9ann9mp9eFrtXrNaIeEMMy
1cXH2QdgSWynmKDmyS/+AXv/06NkgzCGjRrAIpnhKAfRuOkydIKMuHybKKH7tFQx2e9r1lhsI1XD
E9TnXEGMXQZ4AXjAXgss4MQ/FZpLbaw1D8HVce2puI+FpvRyutEVlXB/KqSszyttVw8+wponI77z
Udy8G5IPxLhXDzGM4NpMJnQPnIhUyTlWorGvtqc58FkdR/XVnBNGFy3lXpYGPugu9lGrE3emN4W0
o2qgDGuIwrhzbmO59NOIZyJ9LZKLiXw1Iic/ECJlcWnIriEkTzEW3YO+GTT0ffdCrQwzBCrTaZUe
1fuM97SRa0X6NfM2n0RPzZTrWl0z0SziF8Sp7eeFZs4NrgPmEEVrA5C4T5EpW4tt/0dx0MrrtJKw
W3RyhP6uBueRwGbaiApa/gwG77h2ZEFSoA5uFaKPEqj10d3P2rZhdgsunx/BrKvWTlQrIh3oc8w4
0rpLl+DjtM9J51zJdpjdbbm0ez4bFBw5X5LH4D8LE31lSd4H9E+OwAcG8PHvIjGbdCjXxMscKK/A
K0XEVmGDURgzVhXSxhK48n0aGYX89dJ7pGMjV1ZDatnHfeVAYlZgNsrn1Mg+aiX6d7bZNKx1WPk5
OtMoPkPqqeStu1zVp6gokfJtL8Asd0H3p0Dh5guF3QgOD9+WeT1oltlb7PCRdDkrwVkWlmObpzFe
920jLqxHfgqB+a3EwIdtytpFclxZWhYp1KhRbPw1E2u1SNzoM9cg/4uS/pCCaorhm7GwRR+fdUUf
7jTNfZhAucFA6jB+5dgG1t1hxZw/rNZbdlZSfp7qRYO/q/3N29z2Vb+LhkiDGmEMI7H9c5gAPVa1
o3P5nC09u5yuyXn7Rh8pwd/Nr8sVecpynoLiU3dSq/5elQvw4bdmJtmYyGCmneY41ktPwkmV1Dft
c7xS6XGiqGqHJBpDGzNeP3PkYlaSMPX7gASU/qtQVaZb0CzU6JBEwPxSgo9V/+5ywk7c0MIYP4jM
aZCUKJpSsnp42sdqtj7a78HITP4u79dLDsCweELPr14n98fFp97yqk5R5nzDevZhdlqHF7BPmLr+
BhyOm77Ir8Sq9ziXBiUOKP05sn3WTgm4S8n+V12+qtIwkXXFPf8WNSD9avoeNMUkdAxqeSBQkgCm
IqwFDpc9MhMNsMWT8tcw5+udc7NN9PeAwEA+4uFQ77cNSTnTrtxRgokEW/6RHwYP28eZkEe+tJ5c
Rq8YGbHYyFkluiw1IxsjCE/Gx1ash6jc8DQu1/FtbuJxjaHjThTStwwQ26EaNaCyJEkCfn9wWFq3
zW+Ao6Ltri1GWdmqccoGbO2hBrpirwW0o2388dNTpBoC8lEDVhEOwEhCr9Q5PEB4oVhb1fqohGni
WI2nknqyeMQle2W/aAFYCWQ/zMCPOTDNjxFsX3/Y2J9TaknpGIWZEqQu6+E8FNMYQJy2G5xVPXu/
6xh545UKGWtY15FjPyizWul9alvLTJoEn4xWOtRgSNSBZUwwyHXOauURDxXJkmR5gYvmGIEzviMR
sxWA4EyDlHSH5+Dp8JUlmvyIofHf9z77oysu0wsvvmUJ3V6/8GyRa107tDyjPU4TAnUCdqc1apXr
K5G2ObR98/UjxzHmfs1jxvlHG6GmAyrJ7XLw/+8QQh3A0Y0Ipz4SlSK35GIxGoAovwENznLV1uc9
OHwXxxWepu6cIFseMpHQ06vZIGk9eTk7xpX1FgCzd6VEaJ5BRgAZOQ1oagZEcxySNU47eJcBiAZ3
CAuAPmYaQIXWr8PPCfHXV8EUU5FvlFOSsOeDhcpabjBVnJjCXIv2oYWpTUlHoJqixNuhykGi2dmS
RpPk6VHr/ugh8i7OIKjySB8V2N/sVOZ9amyBAlD08qDi058za6IH1a7rQTSxkGNwjggtSFih38vl
+1WT2vRTXdv+nYZKUONvfFcxR0bqvrxvp890X0B8G1lhdbZMy12EKqR9FMbx5OZ0XruPc+ot9vOh
4YgrWmrHeOhHmgf6M+VZoyQHi3r8YY5pL9vOhTwQussLWhxia2qefcDW6TFlSQLlRfJiB1qlJjsG
omHxgiR8IGDJTICpVBMZa0hy+l4ED4qXLjeDGYDN52CZGsI5iSzssj0Rge8PiCgaV9lO9D8gyqog
0eoMuMM8wCTPqwTcx2V+M5jAxMckT0R1+25alAHmuKfivT2yLUC27U8ijmXssa7iFyBvWo2LBJkN
dSqYc2qnHRKGX2/yHadbF/saCKlXYLVOrt1tfkwyjuD/IIKMyEpwEU4Pepoyil6SaGML+ndkDF0K
LB5isxoQXDfVWOoezWIUZh/f083+h66A235wjNE7IYOTdXNTe4k+rhrzEFha7DFlt4NyT+tP7j3B
v6vzIAsnhovHkXPOPXDuMdoXp+0NGD+6stzSFoEI2pzVjdqdIJzZLIxn0Cdkf3Ho/ZUC6PgrGu8o
3D5B5v30SFSN+hiitu/C1KAB2Il0cnNssEOHa1YI0V1s8mVqobTwy+bSmrCsJnEQyH/ZZH4O/f+G
nE1XEAoSWRM4m4vxNBbK9JkWeXMdHOARFA+UQGYJFdjje78ykRBPYyYKQ0p9HhgmZUF0h5iy1lS9
JRNNam5ZA0t1775P747KS/DzPmsIgNAWXc4Ro1AEXf/ZpqBaffcl460t7pGsGzGL34ck/5EXRMYU
fPapPQmtEZIQ7cBWvyd/V4eH3ipKqeRLeY6rjfHEE2C70umaRMbAZviQC3jggjpHVcCgWxpObjf8
3bKjYnw73/yhYk52iiKN6cSDwuJDvLgxg3BZjcpMDaQJqwVE5368sXb6jovWbXd7gGyLILKqqNQl
RWrOKdGm0BIMiZ1JpWcekjLOqC1l7Z8ckPTwtwW+lo55hSeC2LjHoKyz12I0BDC1yFF3p4lervaV
tqdopL0LKHRZle1bFzrBJvsMFLed1ajT5sMlkXSUcni3looJQVGCEvGvFccIw0v9C0WjJPFK2cqq
cXK1adDcfGd+GsRDxvY3zWIhX0F0sgFSXj72rojFzrxn+KFCi16298vbN4FyWVbM3/s24CMx+dJ/
4qJnDf61g6cadl/e4nQT+ojeln9G3QUfwHaisLET2sLu1a0hS6nI7toDNellwW6Mu1cAqS1LUPd9
gJQJB7FqK0R782E3JIytU4JsFIH8imjfUsjYgNNUJb0V1zUGac3AxQVuv+EZWW5vx+9KJFO1kmKZ
OvEpUP8u5imo9ukoOJiYplMCL5cvuVACAJr0LGZXLh4a31I3wNLEG5wPQMNwc2cFcxK8H61GSGAn
WOaDmfsh2YCsPNzWREsIglX1u1reZBOAr8LZh8EO/cL9I/2Oo+jMMMUN4iXztfOc6hOdAjZJsb7L
XS9gEctScNcrpwLKxdtGdts0mdC30G2+ns5QceA1ipwOxnm9c2l+Yxp5U88YoHzm9ayxxCuvw5ra
hylEvz+OSLnv7k4pvDamyWCQEtHkaofOsnX5fQdfv4YbPXa94/8mmA5kzm9hoqyTbrZiR+RVGN7N
THH1HpizHHANQZ3x4GJa3O5253k1BmN8oQxwda9wLchf/9l3x/jOZxEb0u6E2vu7PwrKuxuNPS50
2Y7GuIi8gCBa6lBtbEn8x8L0ObpwIPSY4lXgZqmi01rFHXLjcWNc9Kpt2KqvLsxaOLywTojR/lMr
YufK/Cukjclyi1bjGcEGbYUgHAslBLtZVCZq1sov0F2h4/EkhXddWiHmTpfaqtn55wy8ZhopSDvS
Toyle3VY48eEc/awVy+lqWT8sXIlb6t/7yKVKuvIJMApK66EhJXvHqHXiB2gKMY5WYn96aO7tmdT
nifmhXlLHT3UbYWB9XFzTvs0kEUL9SmTQRYdGhEpfLJSoSQ6vH0OYc4IOTdfAa6CDl60W1dEMpdp
0cyEYPIcBFnCr4QsD6SSxW/5EvEyyggvSyvTkIwNAZdN003dDVb+UYWdc8nlLXyZVB8OOKzNwqHw
zwSaN+z+90CyWm/Pp2w2jSgJoE9C8lfxvrJu62ihC1zfrB/B6OC6PuibrW9OQ7J36YMfurn27yZT
bUBRqS0skoO2it8f49STzSYzL4QXfZX46xOYkTsJdS6osUkEIb0GE1YK4XEYo/MqhP21qDh5q0dy
ilV2YEl9tMuH+gfEPrzLApKk/hTdJIq+nRa/hvajsiA0D7Bu7jlfBmk/4Wpc0ePORE6OHCMtLcPD
mBgdTo+9bwGHjtAPPtkWeZPn8uHuE3HTtyFLcgp4U2xgUws6Lu9WVq4Hfmf9H7PkjQMlPuxhqaDU
aDVRt8Y9dHocJBEb0o9GfJ5BBtLBIAIMzZ8dsDmwwPoHw/zD/7crnSS9doWm6rDP+x5Gy/x6K0c+
Ea0hMEhpf+QaLWxlgWkIgSvEyx0HJpmTq79ZyTQnsocAyoYJEPGTYBLzqMR7FBE2Q0lEUaGW4J53
pIzsuQTUovdSc6Icoamg1vo8tv/3umzSYFa6WCvZxseIzJguYnTcXTVnoPFv2SO5VS0ekWbH/tJk
Zgxb1q9HcTd+n1kJsXNxlnrrMXRG7P+g5wZ05D4EuCnsdoFS2eiLGUmYDUj8ydAyjx6xOd/S2EzX
ftV0uKB5kl8EuvM1zJF8D0sJIuwoOfb7ql+fmacjSY2/YCOLpPG13ZNmpTxOHU3s4vu395b9Wjhv
6tMvId77UGBegu3QqqzSClkMC0GnAVh3+S/xYVjln7luJglpYy8BLmjQsBOjQaZMwdkJhOwAgwpE
SDmOydz+rwJeSx1XecQR58Fthp2U8uSDC3Ww0tHOgSBcW481rDDsETg8P6XAKB5kHDWdmMc+n/EV
KFq0MFab+jNgJktJ8HJ99HmCmeaXZmycy91ZJOyF/Ylzy+9m993OCCuD6Jhy4+3TwpMnS5it/mZ6
/TRgtGR8+r4y0q+EELnuoEO95235awSguOsaV5wEElQtdU3ZBBCMDj/6dXyg+i1ZsiUXIjUM6/qX
G0ePltzGmffpcwX9vy6miK8CUzm4TKxQ8cjXVvUN+M5nQlSOBh+97csXCnvIAWECnYF9TVprt8HX
J7y33XmZK+28XJ6KYsQ7N5j8eGY2uX5ghxc1r+QS7mFOugvIE+63gapfgRUsolqWIJ5DuyGDHbG2
ZhHiGRFdtGFxGWHKXeOAEY/13/UfNTphu5g+UC83S6/vPb7Fo9KhE3EqJ8wtXqvDQBodDCLi/gVU
1Dwd0KYNu2Ugkz4Ywc84MhSIbuB0nbE2BtquMiKCOb251Jk49vpETXQC0jjwkn8HbqkC+mq72V4m
pujZOZTnggbtb62QSO8I0X2rGNGVYH30uDOl+7OKxpZzfr4CpCpkPejCejy8ZGikQEzVSoH2HGAC
MrAlQeI81Ke0r8D0VAjIGVT9ELrWs/saF8yOCD2TOuIxePmTkn9w2YG4sJZHuakDwCQnAT/m3yvq
BCsku/VL9iGulPwXJKKhkA3QSL797lVx38oBxBapMrvr0AnfJE30JSAI+sZ1wljd7Cq2rfYO0Zbf
33v7AKz13/7a9RzWymJzk6weudd/gvipWpxtSi83rWlrnS5QGDGqvt5MH5uNd2lqGAr/ZkBfWvI3
URb6Q2rI+veIEJnOiy9sPj1VeAigFFRkr2O2BGHGkg3LKNcIzxZEoM1u423CZLgcPf0RnXpt6XsR
qORz6VgiKHGtphYGtxiQwxZN+G8npXxB3sIo9syz3dtldbM3ULkWd/GHxpz68vrRe2kToWVC4ash
Mff2/KpMAe4MiFiA5OPvXEbo5GTA51aizG54934ri6vspcE66FXm5BPVwTCaJM8CTlTvEzb3Onlv
bj0dSkMjpHT1PkmKU78iG4owbPD7skpV4SVV5mQLfgoNEBS/6MvU8W4xK9rqdk6NMGsdDf13dwgP
LEMpR1WEhMVanLT7Tq5Rw5FyRw8uN+qHDEYX8og7ZhWtPWEj6D3AtNw5XU2A57cBSSgA7OeekZqp
SMKZg7it1uhTY1X3sObOgGM6vhEh6N+WWwdG6yaMi+Bsdh/DgQ/uXAX/Zp5MFucEiXpyUFDH3Nnf
1bZ9oP1Xlk6pOJOy9wfXT5jbiXRAsribfEVjH88QKXmpVuwX7KAp/RNMEAO0GxI41nQ3wKRPcZ8z
Eh35SWfGeOVImKp8yK8OTVU7Blqeq5d5hhjQFhECgURwkPHk1Z22vfMGs2cXpuRnL4RAVE/lZlmI
KMJLm9fX0IU9zYUiY108mOYJDbyx6uEYDUq+T3eHRPxAzxYruyI1UybxfdA6+hDG7ePXw33QeCQc
c+4yhziN9MrmTX+VVemPv1ESWpgxGrm2xGBL9wcWBIoTpAE9gRu7oCj0ZPwaXq1nIUYG3LC6892c
UVPlIioiQNRyZFLwFp92ZC/DO5n2pB6Vh0CewFdrDKEIpeZ0L2CtSV3bgnl+LylN+8L/z/h574Vz
jMVnAEh7vGkk/sWwu7yExGahQ/ZL6/a4ifhKL/x9hP7hFY0vXz7yACTXrSrdps89rBjB0FdPfeAS
2PVTvnfNXONVLD3N8ch0tTjLsLnJ6JyltIFz24HSMmxu9fhtsG4i11qj48Ge5STHCGJl7iPA8Dfd
UU82UyPsVKUbSE/KTFi05ZslkjTv+FjnGMcEkF5AH2/WhF1BrUYA7wq9Um1UMrFWrGPgM/NojaR1
8j/1NIOcouveT3IYe76Tk2dBhqrhe++C28uVpIN95yBk39he0Uyv5ttB98vaRE4Z0paRg6fQIDOL
XFMbc/v6KG5YtEiVPP6wRsNY5yzkZ6nSWCmlh+1Am23qU6iEDaUPMfsYZVCljLI56eO9L815v4ZD
224XCRb6vcRF6VqaMrYlNE7AtSlCnYUN0BXUp/quU+qzzbZlWZRW3tbzt3Jr9vik/K0S0uFfOLl4
CSYZpIJJ4CHLFRDy6m16slVxwGpT9RHQqP6KslxpC1ZbAUb3q4WOkWvrFbZ0neUcYFHHv7pxEVbf
h+hwrCHvKLSin2qNgmpKLZDuMm8rBSmG+ymvNPQ0GjZWXGUiG+y5h3EEfcAihQxy/1jpuevbz3mB
wpHRR4OzV2S9eaQ37UCZfmB+Y/9sOeTTHllx1MiHgXdzTt49ARez9MCu0yKV5hNfIhUNSun3Jf1Q
nq5p68dedqi0FVG4naPX/tlUFG+h57Eo1EuEJ3REW8HPrCkPEjENSXsI8UizzZw39XoZwRP/ygSe
jMXeBqvQSilpp10cidYv+0s6d0eIiGN3G8YCybMu0FcLCd55LpKL+t6YJ9ryo8vhPX1gNCGiAS2T
KNv+2yK1stTLgJTIP2T8BMUdx0TwWauMHmz3WeamglPXcn5kK8/SjvjwohkUx5nplRWc2TcI0uwY
nSRKv/m9DojHCl3nda5B/ypjP4ppX4DSnA8Ld2dQ+zPwDm6mwHt56HmvrpUlBJ8fggYofIfz4Pug
O8fCYEBkNfXnEB3NuHGj45PZ7dCMw1NxTjiomjC2irOnw899E8KfiUP7TKNSTRel78Ox0AYqk45I
YP5ILUJIvlnIlGg7NzeVmGRSt2C2STAiUwy98WopkLRpyAvanSvuxV0VZ884Jdzf09/I8PZoUyFZ
WmdZoI462qY3Yg22KtRoVrew/iSNMuLiTQy/jEVwpOKSFP88xQwlCDdIfQ64AKzOu8N+4wwJ3Pg5
1dkTZ7GIuaEeYPk3szWpEfYCTURAfv2hNK2aOp9ig1u5kGF04s04fyzFUKRENtT2FicJRlfYYOSd
qYsTCkjzuAFQtck2WR3SUXgXCpDFV5xC1BFYFJ2NxpNLVz3yRoUqnEZb5djhcTxh/uGamzuVJfvO
0RRh3hvsRZZGHZYQ2pFePQ/FRNFlHY50DO/RHP0n2eMpts2OT40NRBKz4XUYmH4H5OclY49OJDtB
58A77TD6B0uUtYN0ECR4RMcg8nguW6M4Nfh5eU4bvIb4QuXQqG8/nCDgf296PpavdXkIYLG7S2NG
OeB3/5BpSyrvfQSDaW792bQdRypFzPHMa1zEBYKpZfC2znJbzkyt4wm3wcu0/6mqQDYzs3FXkxrT
pYWfXJEf8TIk4NBfaP1mkuJb6czH45Osbu9tQOB5/4daMfk1Md085o7e/dD+EdeiJPEzahLQLgZM
0uBrsMNxG7gQBgERK9UWtxQOcuT2cSHke3WuMB+QpVcxlEma+hvp+oM8oL4bw6WLs6DCLmU5O0qb
fa5vB2KxLYBuHCCPXOZWuGYW1lMtf3Wfh5Xhd3UiMVRxS9QlcsoxEwEToYv/E5xMUd3+wNIdGudj
qQ6gqjJlOlSLcVnzemVd/ra0++bP0KFaywZYnoIOf/jbTtU+gKSDCxTuwv2YT9mJZGj5bSksZYUW
uotXXqZU0WhZBthpJawUSYjjhyqOk0l6xa6nN8kpOhDptXkaBGvx/lfNZtJFWB+hEMm0AsW++pDZ
TVEaXocc2M5DgDcuaF2fC7hWQglxpdUg9D8KnGbLkHFJTokBXdJuzKFhovrfiQDqWCyPhDBSj5Vw
iDMFEO3RGReJ45vtDB11a3xeXKnGHD/8PxlI4jYZRgSp06KnPpZ0TEALDqne/sqlp2raQfCFgKB3
egl4A8QFtC7DGcaVApO7Mzk5adSRUG3oEurp7yOAk6ABetY0Ph8YUiOUQ8YjxemNNqNkz1Hz6xvr
p4zVk/5r0k9ZgNdXo28vUy0Re4biXZ2LGqwRwkcucHVQCWM56knPbyWWrjJD/n0OhrKJ4N42jp8k
PiP7YCKBfG3nB3YfzIMJgODZywpiT7iBMqJyFCIsCVnB9FpA5Gm4hhnnnFmG3KVr5JCOxhYLd1k7
iEnhbB26UunwN16wzHUIAee3aSkRP4rci3peTDBm+RR/vOP1Z7oMUYWaadiThWndPEG6FNlo6xAt
138YhvIeAoJqn0T/qDO1c1VfmCFv4OD9mcIb8mmOYj5WT2uOaiBrwVDAhdx0towZHKXH2bw7jrEZ
/LP6EpLy4Omdt13RnAsIdN13VdWNg8m3YisQX3kV718CMy+Q2Ne7VKjBnZ8PKpjZeQJBlDMjUFJi
ssa6Il1UXFDZ4gIRWWo0sJLVYMttJ0bI7NhyvCgRV22uV6tmDl6nbibPAmdrs2ot8mttVxLSWt2M
8xIakUhnpm0acM4gEd4kWN9OQQNicvdcfwFWb7DtZCKMuhurhbnRwr+2uXx/ieM5o3o66mf46WI6
XwtCEgUAL+8ZYFp4NeDvstRgdEm/5VscounlyNjuk2Cjb7FYbFfIAaWYZ5QJnYetKMaOLxDFD5kW
uwm6XS5oKEsG7EGA7ah6CCMOqHdJOGHkfGh4HO9zyxvuYDj3bWBCGlycMrueNx68fh0CQf8bsGNs
Br3P6xyht49jK9JjG8BxTucBk8AJe2UXth0bEj0TwhzqjwrhUPDmbJ8Y9if1lPlNEqHdMn5wCaJR
Iywg7CJ6FVHstqluxyINvKnKNEazzg22onu4komapfub3DIbiZ8FegU5hW79nz6OI7eTEGp3gbZi
gEXD6fI1PR1FDv774gK4Y2NZ8FHvXVOtfnKokOGQfrCRLyCO1xCPZzOL5ri1w/X25VnVqrcvkaPK
slpklXI3S/gIvQhR+zAEgW57CEfkuxBZZIOkKXLGUG4+1VAqVyVqLoOtTSu6rsXV7oJFAIhmitHE
QGMX/S9yvxBuMIggmxsxxE8HK/rhtZW7phuPaqzQgzbzNclKnMFx17LH0b9+lx7YukfALeiUAvre
Q3HGcLptH+0yQMgjd0BhhabzYRWGAb+pEbp9Ccf2/OC+VeUwZ2F/tZzssveVdgtEhEPqTqFYQ5yR
HqZlzND4/9otgjvqYRyY3qMZVQh9s3kjYNHK8w5bPg93XfaHDQPTCfhp2fDgJcBIQWjg0UhK8l8e
STE8reQI+aXqPxeDgaPwJ49gAucRrSVIBXi5GILWNTLpzPfpRQTF5ffb79dNBZ1fvTpLTjr6FiGS
bYEnAF9wSeGXwy/MWnYTPkjgHjHALBV0N1fFndFjC6xLetPfCgQa0o/Y5siRU27GdHXOw2iiw1z7
47qVO+G0L45Qyilmest5EIzcryaztpHeX1b/HL9NSgpaX5Hm1NwhWF/WJkJSCbidn3MYVDRm3LYe
etjPr7tapXxFqL9l+N+c5lEnDaVXdVBlVEXbbMdRMGz2MYPvOFIT6yB3Cl39MST8LIiqFgdmPWMx
6bZOklcLvtVJ41pSoT9hxDlJaxj+MKGSPpMuQgTK1vUUr7+fx0itTVLV3cEKjej/qmtRHR97dh/N
AFsUdBJco2/FReExXWMhpXjnp4bJs5P76iXh7wAQfxqCT6KXJugUsz5CW0sZ9XC6Xcj93T+WwmmQ
voqRzyouUId4cAK48bny2Cqc4wh9K/neMDnIVuttnrEcCov2ryukG8MfmBH6d6dQFfQY6xyAgP+Q
IGeIPW5koH1lCo7AVNucBgnTIitXAFouoPpytTWSzp3J6PIxEDGtjr1zwhSIpyW8A7mT8J7rra+7
3VVfIN5Pbo+dPN8SIIYnLfg+hSKesYS8+0jNjyssjyuJzARTRwgaJXE9pomLB4p9/AYWz8dWif6c
5i2b/W3jnfq/W2YXPbkUEXifMxTHTz8E+PlBHXAgJbcCLQ7zXIg/MQmIXiNKujwBxDrkP2iuIF5q
zzf21QfYSpnUg2kzYeRPY+v02lAi9d767phNKMDHOtbOGtZvlpoJVk85wUweIaieCfIWcX3mkqUc
eee3Wk5veYI0nBvPnxdlL5QM9NCIAEEH1GuMOWHsYOVfoXXWve2VlWu+U/R2tAxhTw0Ctu7VPZPz
p87b3mRljEMOzs/vGYyxwy1gS1tHd7H7IxJ6rcSF1mQKfPlGM7SZU6msktKLvqWR1b8GmDg4AbzO
BnUF2RcdQj/Gr1lzqsR1RQEmf0qKytbevSj+ptqR6AVV3PPIaqX2r/FHO8mVSEid+N60L/cknWSS
JsjfnGsYssxk8p26f6oCceME9lEfCKEkhLhO9m5jbcKa3q+kSQ9gwQs2NpE2P5uYoGUYEioGvRXC
mUkUlE5BaoTrZJKtc7qGip6jTiyNyDPvQgkug9O7cRHpnwvXCsTWWCYY4zpQQ5m/nP8IGYPbEmw0
xT4t829NdORC2TWzvZo0IxtRji+sUkYmtvIxdOsa2RC4ErpEVWtVlxdKK1yIbU03O2/fNnIyMoqf
je6JD5lCEZymznAy8cBbg101llp+a3JZNpoTMwHgk8lYFrCsHhksPugT+TocIZkesuaGfWr1Tk0W
6ENG6isDgAD8hNhaPIkclTe6RGH9uHrczbx7/CONPwTtZaMl08i6k3JxvtPSDY0N+f7dIjxQG7Fg
4zMI1TE0qXAIZu6jkld/N9ZAWTF/X7BUH3/DDLTDvTTjIXXzfot+tDt085e/bibxZAmVqLghvQci
XFAK7VpfIjxlG7pyjUUWjYFx/miIC4bD2Ld7rDr2yiyMHgBjb8d1W/qR13doBHzSbeZ/CyThQOAZ
6+V1/UAlAbdrmwM+zoV3WSrBd5iy9xzLMfAhfgf78PD/IK1ScbAW9fDNNpLaaKX0EHJiQ7/sJBV5
8Aa9X9W3XWZFgiarJh6FurMSEFC/VHzN1zuP/Pxlj05CQivnFizy0A75+MERPgil+L1sSNLLnnBO
M7zkRoBY2kVuU9w4O2VyiimuBJD8kcRHpXCO8G5/wCoC2WVFcNUCTg0VT7S6pKOGcaeYWhKb231J
sxEShilSYtKTBdP2J1Kk1MHhIPJmqm3BwyJYm63QXxqrr9kEgcHujvjBcYSiQKUN/G0pS9rlBnuH
Q7J8sAVn9D7sfWyNd3YLnMNdNWtOjwOvf3nLSLJnRjxRiUHW5ZJTE3CtEzY/9ybcRSU2zzhyYJ8J
YX6z0vXp1sCxBJskxCZVcfbHHu3AJ2N8odKvPcIaZ+8XZ3VEd0/ApA8sULnLZASBhW8YbL9I5SNA
JmvDcjx7zO7UPx3OyQwvU0lrOUnHOWqWoTP9//t/ThwEBsL2ZC/2TXwxHVYPLw7T+VPqkDs3t5pp
TV21BPTHmwv7J8CcNA7xc2UGHmFwClAshQ5sB2S/mnnagnF7hWRgPV51ikRfwGMGcdgROx4sfoaz
QL5p2Wt3n8EKE0y8FcvUsu2r5nnT3U+FTxyT9MQF7qyIXq5GSvcl4ibPPwvuV/OfdNQX1a6sEogJ
aEzjxuS/E83L0msX22ILD9trTr8H2GCee+D6elIFY+AiMApxdwM18y0BwiVUfiB/pqaku21lLKqu
XbYBRItvhD7JZotXGZsORvpqUpBgDvdHoSFlEo+R4zUbZTj2cCJqZkhlXc8d7DbqHp/inQQCD8kk
DSUT1smvQ8EHDDtmhMt8JyuQK6KfSzr2devIfEdVh/c4rDStp63BDEj+502RjGDl6zIGj3Bvw479
hfjpQYyCwz/OQK5lYTc0XJveDAz5IkrNfr3TSoAKnYn3Z81m35K/qva1m2QxYGjhe0opmngAebx6
SCMC8tyrz0gs71Mg+GVSIb5fk88rAPxhESAORhqGNSpsX7bhoH8Tnp+47UlE0GtcJjGwQ/O9De4D
opwJ7rAcMIuOZWR80tZxon2T5wfYOFbwCNP5AbCzQFDOmdQWDWnbxiS0EQPnK4tuaEWsWzFcVrC+
8GwOpksghHr7/dbMZl9AK/9Ew+5g24Aq3MuMQrE4fJIBu+RLxxjCcdCojjN3c/n33Tn1cic4ctfk
yBsGuw3fyuDppHtnmb8Ft/4+7yKaIzCN69SJTRe7zbT6GOonzhirvK2ZkYNgS4ZcML/dEZbZipF+
35eD3zVUtvGJ8pTtNrs1UhxdW4LKxvqxnJ7HiM0b9XRgZIp3tMX3hG06QS1l/PR6QxApkeguw6jd
AVSJgVlEsN3N76j8PF6CUeS94+hSwWq4PzPEJ7RVu5VRVNVPQtRq+pSAi9tuYD7nTHpq3ZCKd3xy
iTg0LDO/2hE5c0sXmWbMhJiS97VHiUDmv+NDb6Ni8zi1E+3AOT4JfGFywT+JFbU15GjE7c7XyzUi
QJQE/E+gLfYu73cw7XR50KrO0h6EyyTHWPUmrjPg8nLu9mWoThtXWD1MXCZVWZ69EIXBEktLdn0A
/OE5NrYifcAF8/+1fMCN19ny/RlKexSxHo3NfJAn3S7h79EPqnW7d3OaNaebyLTr4T4WriQvFp4n
U5zUSmCinIAtDJ9sQ+5kbRKunf1xdja79LEu+A8iYnorR28k/zp4QM6fJT6steS06cJXgRivbu8P
OtaiBwyCGxItpIyLih1RrJVkllE/blH6Yia+re10h/PLREqseAt27UVTMA9y7ENhM2OTEGrMyHEh
l7T4diDblMh5gGp+oN2kMK9ruJeMHzYWE3UESCH6RcKR03Q2XZ0ZGvMZYj59x/bo77AiS02Nw6Wa
56DuRNR58T7jNpiEiWr9FJZLZrd+nXuWO0Su8ukAXAw9p0MM9eXUHBjLIzcgPTC7PkoR7/lFCoha
y5UG9T2da48PIbdBu6mps3bvQSPBJuQ5os5mjIcTqJGSPJx5q/yDw39oY0wHm5VkYLOiqkz6Fu5d
8kRw1YsFblr3oOwg2Kcm5fSfPWso2FBTrSbMnclJUNSJFC22V1Erbq9mFFoouum6jyvz+ekC4hV4
cRO/fW7CfeLa9zWXU3eKL/wTh70QjbaP118lmTWkRucIe7lCI7poLlxcL+J8f3Q/WOm1pdxiCPP8
Ci6Og6Y3zgWugTMCs8V4NakXCA8UlMIHVeCidgYDLRQeVKZD3PwTIjAmTCI//25ElLoYsk3eZijJ
BEL3GmN+uuZZ2E0NNGBcBlYVCFiDHal5kVO7ih/QL9obVnmztfJ6FSV7VaN9claRjVnmNUhp1o+L
mc/cE3yuIdQl5WGAynzWergkvJyXDvMcCD5zrl7LFc5zamd1LckLT3p+EGs9oPm2CcOnTvTB12Z0
RItM4aZGNIUPF0enihnxWCW45rrEr7VcL92z2S85TJkhWWKxCNbOV1i0cwdZd4nhM+7jOY0u5hWG
uXDdapxzNI2oRp8pPociXaOZKjvGUwCmco8/sOUP9PS7zon0nMEv+sU/jEawCCH7keqr4OWgnYvT
RNnNY8KQFLZ/umWNMmiIY6QC7zDy9ViIS+Gnc2Jg+B4rLSguHLEigVZvXD1RI/ZrWWE7eUfZdNlo
KU0wi3nPqLuTMyTuGyQ6x2ZtJD/2bJuUM56l6LzVRPYMOmWn5JAp9iycZ7TiutfaJb+xFUAorG31
yuwQeDFNp5DvaD6kneZg1eUXry0DaaGD2dxC5iHeDBcA5ZE+FN5gGp48ooyUhmuoXs3OWRbHlCu7
86XGx0rkGJ27NIIdl0xAKL4fUGN4D4G2PXanlBBpxoSfqkgdaQFCFlbz0sIxRKVX2KsjCNI8t+6U
ForXlfPNZ7MhFYL1TQZl/LGIU3WNFWXD5LLjb6+JJUaVGcVBFu8g5mHWFH/Q1VZevNCkMO2mo85C
95D3YZWdUakpQ5694R9rhVr1LV54R7LCA3zhiES6JvflVBo9HDJxFVKG0L9kbK1/tS+MHcYcvz/C
PU+zY2WH1K0VoRSsbhX65GxeMPKx0I59PucfCBqiaBSj44WfiOUReBsjzFzYGrLBj6N6zBmk6MAF
cXdmwvaM1JzxII3PD5ad3cu1bQf7fBmnts3oTTtYRIP8nhGogSNw2y/J68YbVzxrscGTmFkIkSBy
F5WfQw6GvSrkYprpgGEMzxkPgYoQI2nGUxUE9qCkJMCYxY2ULtv30mdA/Wu72hM4yRSUBhoWCWzv
BReZiy3XW+4u7kRuM28Svcq+QNKDpk0gLlr00bna6WVLAqSpsCCpQkCCN4pUBcQkuSpfO/iHmlOK
/aSL5fWYBYEfDtSuagTsygc0GOcD8mBKhZNqFsu9FDJWR7p5VHNNi92Qx/s/SP91TAwKdhQ4fvUV
T2OrfgBqaLCNX5Qes3PRESchOfV6MEDQ3aRwZWxejYlJZApH5Ewn51Cro85JZJINTwaLy7CnbE/a
H5tLfRlNddRAF2NXpxEYMOt2f2yeajQcfiLRiQ4kXYiNu9zcNo+mb9l2CuwENKg3el9pL51rm2XW
RKHd+a9DWewa/8iy/7YrJ9YlNlUS1kx82iZjKpHphjD9rAZ83ETFtVDoBi//shNFmAKCaZdx3ngn
2BFs1i0tIvl4bNrL1Wal1TPb061xwHhuSzFmkpKAQdB8eWETgSBaAL89K3qVt5ewqShZSDyzWRtr
Nw6+TNqnMGise02F7x6TeTo9ZHgjHRH8wfKZubVvbuWLnF0lCKA6ibJK4s/o/rShkUz/X4bTo+H1
1c2xaly/PPDvhymRPpu6hswbxGr6DfmpUHt2ZmMRRAsLGpAoLb0sSS4XWcJvSwxA5DCVtuiSxj/V
lBmHR700hbYfxpJiwnu8xcbXo9Mi+GX6yot0geWie2zPXYV9ypbgTZQmfcA2r26UladBD68AStdl
9MZ3FdkQAwjRmjPt4/LgKJEZ6eoNJrBQnzp5jEP63GO3szppYCprkzKaRJlBYIQx/TaNI2AbhgkV
uBaXfvhmVYrrvh4oHqCLKnBvkoWaFCRNmlfWjZEayBWLUB/Wa8DLihJ7+a0Zd4YquEmbWm5zjwS7
3i/dgrWyoAXIOWEdVeCyKSQcWJmt5I+dTvN+7EQc8SYOiPo8p92vFU1fG4i0SeJq7EiwAXZXBiR2
1leDM/UYYAF74aw8uyePoiwwrknex8tPAPggaYp/l9NRg2ytaJ2Z05vkdPzzhHfqJd77MIbogaZZ
Cz+VBEluP85akP24oBHbLRwgC8EyboKzxZq3hacwBdpHx1nw5JrSDFSb64VH5YtpUBmysCibSkSa
Az9qskK0sDNowBsHKbkTBDb6s+y4x/OjsObY6/sIp/IaaYAd0gQkkkV08lkIDVFtCKI2UQz9npsy
Qc2dzv4ij14er5SWHWx8OFgcYe89IeMp2YWp6f57rNmC0t5ZZgmPwL+Dgv4y/VPRHQLYl6Pu3nP1
Q9eM7VqYl7USi9Z5oFkCNsSFX4C64bptXj7R0TYRs463wv4tz8Rwcx4PFoPHy36hmoYjZpe4lyrg
IW0QIQ7mDVpRw5Kap+UFubMgRlipSV4KNEriULEt/W/4AYsLsNoQXhwQ5mR0BqsNLG2MTcgHCurP
IWDnAU59ln8jDylLeFg9ll6aPzAeVHdzuEKU2MZmJRr8qCxa5BXse8E+Ah2cUwUtz+t92KUi+LYf
6cqsF03X714tLtxLfdcDqnNPsa2aRM3foYoYqRwXu4MPA4vAFuh8Im+GSjohBwPU34yAm0uWGfAY
zi/seT/ACxtTsHmQEwxGetNorX28Idd5H3Mt6myqoFZb0vZ3jwKBVP73TONsWTZL39aofJCaT1GK
Jstc+/OISjceZGy9e6socEGFJfEv85l9lTsh7/MkC3vTsfr1wYzy3+wSle/UKmxeghix3E4PNjNg
SxmpmEx5fZ9oY6DOrRVGD1gVOqdpJD75qzFg2HqCbkN29gYURZhqvlqeZ4NJ2Jl291Gcr1UuGr+y
9MyJoYtKlpwkH4Hl3CVbDamtQY3UxWd7VxGHl9sYEmkDFD1npmS4DYx5dvsW3amph3Tf4tYIYBfq
Kplr343NTDbSUMm7gXveyYZnFlP+TCQeGCbTvw7DFXzcCh1XdYbNCh+spO/0emgeltWEl62pz4v1
TwCBlxIdSqjXZdSjDQQNVkS0No0H+nBzYrZT8czzp7a7Ji749YJ6/0w+mwJBJ11jeZ8aDd8Vlnez
9ndVUEoY+awyYZy1GZ+FIKtwoKQfORhBsof0lbP8928lnDKU0GNpCM2GfTA5mE2YaWBRN8zCiTgM
+TUeI7TQ62610ybzAmCpklqb2/1bq3mzBoOkEQfaWcUcgDiwlfAdB/cIip3A4BT/fvo7cpIklWa7
fy1GS+zkPFVnYzRhlyS9nS5CUNw5U2r1NhRQZ84sM4OWxU/I72a2bl7AhSrSUa8Tewf0d00jiZmL
1DAbRBptlcbV1hs8X9QiDK+8rJTksQy3PFRvcOmu4+w4WQ4UyNhhLlRq+OjpEKIkrGK2d/IA//Nt
VPX0MOTGpUI6Bt7RU5yvTtYuNMXvlPsvSoXOmF2ckzRR7W3H4VFXhkCmBsAZObcNITYP9RRGuait
uXz9pcqEzkru23DwGulR0sar/H3QJKpFoeFz1rrSxtor35Toz5lQL5cC/qV0CwIfbPEV0TI3eHXo
1H+sdi6OUdjFjd1Rxo/thQtCX14JUT4U5kKHUYQOBUYCNop4iQstq6Pf+Hf0gp6PPw065hrRd5Wr
UVZg101uFAif+T8QRsKwltOAVb5/U88pOt6i3QIis67SO6526NEu0oVv331iqnN9L0ozFiKf3deN
IN2Iu3tx2MO1E20A5REKaj6YbdW5wV4cdjEqWjbYJiGD01EbmcOhYw5dPYmtRMiJwMpWvYbSKvx1
G7P0gPi1FYdGkzXyWb3Bxktu8oDSC7cdigEMc5GHGp8NlH5lKJzvvLwDNAykVqvVrW+xIRRGZlxs
IZ0gBS5Zvd+lnkQa808l8Y84Dcy28sK8qa+5rZJtqDShiSFnZ6Y8SKlFbLodKYNTRppB1D9+yHtt
SA8ykgIiioTNO1XpCAgZ62ccK94LsZgiMeyC40+q15xzmFvaPaQUl+ei4R5j/uROgFIBvHVPar37
ko753Qxpa3k1X0d9kAnXYgsz05SrshgwY8Ue1ldUzr4ubPdoy556nrM5zvvcSo2zbMEd6gbNHJ2D
gF67xfsm72Y+JIfiSL0W5e3CKbqW4lMVrCJaNXlDciUJZ5ck9IOMW4ebEHDn3amr3HMhLZt4DBQd
XN/Xg0AahbvOZD1lqOfCXxF2Bxc9x8MRXqUhrLksMEh6rbZQgY5O/mCvWX8dgB4dlfbcjSacjZtq
xPgzREv7L5iYrQBXLXDWtbcdgpW/lnHWaHwXUUXT/LCOltDbFzhYcKekfLHIb4P6XFym4reKiSij
OOYokOdCD5FLnaN0rH8qHlQWOdSal/wCA7kFnM/+f4LfOl3QlMyjFv6zEhtKUl5YNmBlTq80vgyN
t+LTi2gltfZ/IjAnqRSKGwmmcvuisctid2ZDTQsd7C9BDWVR1CsJVtICPv3uuFBYhXPDCCcjGK1f
c0DO/253hDUsXnqGbX4hSoxWVxXgKjC1LCU3C9k4cuB5mRhV0CBx+yCZuDGbWb18zbAC8moMUKG5
y3b7Vm91Z2ejTER8HrxqeqmSIVbwsX82rCFoo7Dh7XBvGPsrMgEOq9ysfbmK9aAtFxncUI9YzlqY
zzKv0Sp/MKy82HJXJ+cGx7vtn+koKyDtNU0yI2ZMCtFmf381C75Ob2rJ56WQ2/ThTOCzpYjhAsXl
2Fb/g5gyD7SOQJMqMW+LYxRNrPlniU8shi2sMVQp+zEcI3PafvaBX1ufhwp4fbdrsC4zFJvgej4z
An17jo7r96w7aZSSTJRlPokjlJcgCvFRxKEdq+yw3xDD958X1GB3rUsyN7GOneIyE+GyTKKfnUvK
ZtZj1pdDAKIbdeQlnfK9j5Kd42pKoaYgQVhEha/5fxp/P6RoWzk5Oyf+tivqVqkYj2wvbagsDHs4
sSsnbZffo9uciY1uGXgcLt4dIZvgBlfbrjjX9TGgC6QnD9G51GIHud3iH8ginjBU/PT9Mm8wqC6r
9u2Iq1Vg0XU041T/f6rtiilhQ2yWt+WeGlmbIr3VltlnQWjU63zPQj9XI8GU4WX0oOPAwCZiTVo2
RqSA/CQ0rO0x1Ic0rCl3Ruf4bpHWHXl55f2zYmTlTrAac7tZRSa4lzlsXZg8J/HU45QzhOqCr6WG
N39s0Cj3R671LXGl7w6vP+Y0gootXIdSzGqclYIKK4B9+GXSbsguiIi4D/hqn9DdNi5umw9gCrpp
iZG2H4LsIWzTCrPXlpBTKTX4FTks36J5Jwz7UtTnaAICWuxUw1jQfdVM27KG8/u7N8nyAqbARn6B
uay+gM80KJjmGQY1QzVz21MhTLipUMj0MFNdhLq9FKhxKJsqzYkFFsCeQ5OvhLVebapxPnXn4gMs
B3K3tLUtSc567V2aUfgyPzX++ICJGAEam/uXb3/yPSE/YsIfvdyOzr5qlTut2AuFbMJndHMQ8cPz
9JGkkuosVneGXuL8bGQnjw506z+ASJ45R2y66ZgPWxEYr3FB76uUsOUgFei4fdCe5gJq4ptSGeut
ExOLhYckpITvQFgZkGV7CGNs9oLLLQZRVrpiYPjNB2i5zZnWBCPFTXx6LWg7Uqi4U4nwkFthS235
37bGFgAVm7/TtXDY+TIbfvzn4O40deigrqQUhf5uG4lzY/MZC9P/tXUP9GthCFlGX4hFY2K+/wX1
DK11cSf7fdS9DvAI+n1XRiyXloBsZAn4PjS+qkn0eYDNQ75bcG5cAq8ukzDQsO/s23V+NwGexDuP
6ld97anYtC/H3VNg8ZCsgM8T9BuKOf/q4zffF0f65ywsAjGHT/wN0hct41K77pS7lveGiasXgxO7
MMXK9LSnQkfQvCsWNfroldHSx53h1acH3FMkGkwjlhrTfsw10V4jeOlPnZHqPiLE2eD1MTcRv0m7
lxYdIJgHh1YnaiZ2W1+ZSXn3VBAAPrDZ4Rfjq6P/Hz3z6+vZ+lvNuip2dE4S6jRHwFNL73E488+L
NWTXv1xrajCyf2gOYacEaldqUjXR7QkyhvQWwBFX4rB3iUJyv/uGSbtOiLZnYdNhbYHxKEnH9gEx
DTEepvedXlrRojgRHW8oDFsJQ3IIfh3INzrTXgBov1lUwIR04NbtZhxursJ05F+Jc4hpBzXrVK08
zDuAYKJwBnYyIY7vAX1o0W2U1LgNbvEug3FSobxqMTKKPiEHmv2nvm/jij/9QJGfSK2A1D0qnOlr
e4M/bR5K5PG77zJiZk8UtUl54QXyb5jkZof9uvkuWalZgWXIfLjM0mXwf7nqv1X0jOw0oAkMkQOa
tedmFMGgrdRi2z31J6e4j+lKoH6OullYaDo9FPzjUYGnxO8L18Xi8JNDkkW1d3IPRUAb98zCz6Vm
a3f/+4FDFZKYPc+l6qqOFKLR0MyBHLqb3zq2ykcRir1kea0BvayDe/injOmtoVmNNtTkSuTIQ7Ce
wOjhpoY/wycByDePd22NRUh7ui7zuNly2fDKkFidBhuOdpEwAW0R4E9o21VTnLbU9E9TkMTMOfnK
0MGUnKhDg1wC/rRj1xcsEV5+NCJ1t21CJZcEVs3KeaFUN63NlhwFih7iBZbMjmnXKxnXN50mIN2T
eX1g6P0X7eF4VjYBdTWuLL4ZWgDHe1mrifDIUzd/sMh3gC1Qpk1mhQhQXx3ARxIihjFjBTFVNtAi
71q18mWlRx6ie0zKptO8imsV0Hn+EBnMM5LIMpKrcrR2Nare2A6PfmHExz+4QnC18lUPNJb1QgUr
SLUn0czNFLhs1sZ83p7nbHgF7uN/jUgZZZfP38GuhFz8J1XOTOjaHVeokjllMUW6zkJlM0+bHJ2g
wgszlXVVGRU8b4VF5gJtjfxKtX8nHcCwBnrBbxyM271wgsIL49cJb8vpj4gOmOl2FiGshha8+AGT
/eNRuBUFUWHu50cr1H45hO4lwIYM9kQyGBzcMC5ScPkk+mfOxivVnCT4rWA7pCZki2nkIPvr4X2v
EGJNYdniEbaz6Iooj9byL8ydRIVmEhLO+JqcshPZdEgpzQy+04ksa8/G7ww8tmAQA3oPQm5TUZnC
MxRlG35i2YgwIFYGoNsdBQna7/6dlCt1Td5glDg5KsAlC8Ze5muldbbShMfWSBqhPnF9tO+jplnr
bCGWZ3RbtQGbNMwuTv4L/7K5VkfTWvDG8cqdVYurifhXR/tb/pCt/9VfFivdJe36O0ramH0PNmaV
jRStCsD/E3NsnPTL/4ibsHhoT535MDuSvvf2y7jdOwAAqIhQjpjtJtvepx8zP5bnKNDYZF/CPT1V
IY8y+RVJUiy5J7N8W16qK2vOhxB4TK5bJXkeLJpGMiRyf5gd0lZR1nzggJ+Vy0bHS1XrTN1bFCie
JzrelUH8cN2BGCFbqU3l9smgZodf7U2NMNIoS3oSVle+4snPmktdrsrhDKk2xlCLSATAX94StB4a
jpZ6/ciyY0NHyHFrVkThk7Yt18misLrhYaNnAp0gjGjJupJNX2E3sims7SY6EyCU6zgXcjNnP/sh
rqqKGJfub8KIEoRfspjM8MmoQieE1qzpcsEVUlQOJb4icGoJ5tduzJ3lPiIP3CWPSEW4+L/kSfmw
JEwd/KGOjLjKu5ck8LujNVRF9kIuCZGmL1NScZeojU8frb8XDc1Wiq0I9A3ExbwygSiUv7PteMyF
kgqZtiYau70IYXbzBKyTahRRCN7/nxNOW1B1BAEO5cdOW0AjqzKMblLO5msXTfB9rQFEXym9iDSU
2X1rIRnekVnTdoeN5XVWsxAvQPyWyJIXwSMLA3mfYZknUuJ+j2138dt3+OxHXXkGzrztdbOv75wW
KhwTpuNs+xi+kZKAxcYuIqr1BSRCcJJXAc29F4k8bLr1BdEmcifmJagfVq/F3SOrAys7+d0h+Lyb
xRtr7Lkror6bzvIZBciDXrG6PD4zEvS+q+8vAeJX/GtjwYFffJ2bnBA7hl50DilPknUcPRbaJZF9
xDUXdM49XCuVU7dAf9Ta4zy9DzteZEfGV2OktRY7D/4zLk2yI03eUiBWx+6sSYrXVFNtVVhHbphV
GUfz+aNWDAoTbVlNk/fkBMcRiWJZLMR8szzjrxq5Xg9xqdUrrM00OJQPYIJGajNmlgvnpjbutqQy
VlfPk7AuTFlRv+4ueztzUOnek64sUDqAz2NJPimBJQS7KJ9avzOEt42LhP5DvOqtBFSJIUxT6WUE
dk6cylvXR4nR1pdPDHF1ISS361M6UCLQMNnOiwXpjvbEPHln8h3Zlh0KJcDZt6HHnLhriv3Sh8UL
8hcKEjXD6JSpJ1pdP/G2KQ1A2u/pzH4FWLOf6NkQhnIM6em3iNCxEM7U7ftNeTudjylNvX5PTSWj
cAP2c3mo1ZZ2Iq3Fm6JdiHlq0ZrTRrrVgEJTqtqWGwMKT1KtdwJmtUEz57tpfiSLwyn83T7hyH5n
b7gI3Dr8OOo37IfgruFIQ0GMli+O/heSRU7/5rbvj1f40i3FqUwMr/C2XQPW2jEgtF1ZamTqN3O5
ymqi8dLxYC2BF1uWoJmNbHs8tAx4Bkk1p0t2R0rB1T3hRolpDzuMlch5ySWxij8mTFS9LwvAZpTR
oNKOlW0UCY4WXtFtN0sNARcniSS47379RGn4x9gxAribbThM+0bq3QD3ds4Q0GGi6jUo3qs/Jr6U
Ik1U+WPpZE0H5UTyy/U5vahoeD7laBp+aaU3/zt3CL2JBovLoxh0bpEY65x4JrdVFKa5eOEJWUlz
5U5Z07unyZedkCZQOr87B2lLYLK+x/w0fBR+6c0L+fRK3lmWYTYEjcqni2w4J6Y0ZXzPzi1Rwy3K
pkc4XUk/sfrH2RRbLVsRfeauFOQHYx4/sBJ6P4SerWATap1aCxYVW2/11nyJdZX2yFYcRmEmKhnE
Kfz4Y51PSysKYY6k/2lA45qGvH4GnsWdCpdcoCo70HOpm+fNpXgr/8l/lwbe6Ka7ynF3FU294dOS
GMlWzo14egkgCsKricBAxjbrazqwSJi9LSjHXErOW4/0cMVjwNogA3ObAn+Xs2IkWcqqaLt0vUHc
ptelKEJYc9HLV9s8EAghUdvCfq9BheeNXYd2zYG6pBLPUvfQHrpqj428QptNR9komvPSJsye1B3l
Vd6yP4+9uw7ScYFIrr+P3JQkpRJhNxmtEXoWH717NK//uztb7TS8J2J0UUHyc8XTffiehr3i7YtL
54CgbeL+Fnhzc7QdkoNc9aLwkcB9ZTH8W9jXBoXaZxpXfIRnC2mJADNc3JeDagrvJlhzEst2c9uK
ZhtI8y0WAb7h/IAZG6Z1EbI986pqLjI3Lu0opC8DWylo4lxqZ5kXiqtj3z+llrYpbR31SJUg2Ie/
d8iaE3NE8PCTy8R4WYCjfFfY8Kn9aZFosYqrPGdlXkEfPX9ElotQYiAL3V3Z1+EE11Qesnb5lnP6
IOn1lZtZ3/C8Y80MmWPMr0AQT5c1MfkTdtjkvfaJYT0CrksaDOgVlcZbQ2loDUxeq3TDqHOhSaxu
2+SqSX6tk/I0MPRVpFfSGXQTKWmUcgnrkMrtE7rbJWcm2oMkO9Z2AgccSyqKx1nxiOFrkdc1IVVQ
LmYnYOAGhgxVQFTT0xTwUYRp45mcnFy3yUimEDAZQx1us9kdesgctugnd+jjDmZlgZSBbKasDCBO
JqlTLZ3EtcED3RvVJ0LAWoevwFZZ+Z4yw+73QqfPMulMgyRAwYVu5TOqciH/uHjZLdqDBpaFQTjw
qgke/qHRIZZ84zTgxBWqwrlhNeLAaV4clFlPG6AnPd7RZB4vgmp5dTicD46AL18seOwvco6BCkdm
TKfkwB5GBPef6MEfy0iUC/dGCu5NWBq/Wvhi/jiXa9+RrE7XrZxOUEvhyE1fQejx2E/e3mWwRu7B
sVEFR/v0WqwGdZkwOOXyhCI8hqZv1v3xFuUan4KkkxDYiwCQurCwmaTvWbj/fkkttA6M+9Muu0nF
GM+foxZwXQDRwjG0LSBlqq/8SxFTOoiLKSygZR9PS8T659/Zo3jg9WB5xGjK3U6tji6+KQ8GlknS
dQOWLFHmXDFVefxgnoJ/TSPT6cUbAAYb5FaU5uH6kzcra8TPIKackbvp+fN2pSCa896cOt+bzfnW
H1VqL91GoQ2weq7EPI8k87T68eaCPUNf4q/cuqmeO/qc743REVh5Gzgn/pheh7vLS+bXmEC8I+KN
violQkHrlXGsudxeTIjmIoM2GV+PEf7lLhlh2A2Ps5r4yMTy5NQQxlWJDODcWbH88/uuokw31l1U
XLvJQFXFfhEW2ftfFraoPha7PSb2xlAbppplUfS3+YZv/MsdR+voqicxvQnxzG/BELcFhnT6+sxU
p+nb65rQhyAhNx9POsUHVJqn0l5CpZtfZf/HcBbeXsJBAdSrxtUQ6iCVZCFepyhSNEwCB9ufZkLB
9Dt0sSTly4OgHWvKZkm45RkRS71Kc83W4MhexAymcdN5m8TGdMGufGdACGV1K1mGRcFrItwuTDRv
yv8dvAdt7+H9vDrH/xjBubEOtJ5K60OTg+DUyakdDR1Q6mX0WbuAy7ULPdn/M08Di19k2DdWn1q1
Zq0c0aOZkD2XqRFao0728d7wgT+SFQcSLEwhOd6JEGsAyld/+bfaBr5XCfpJPqKKrdf4r6CPXz02
uWCLcrCE6ppd2wCultAFMIBMkvhYnYTqGJ4TFs38BoPR4v8MqeQflpze3Aj2SbOWv89eL48e9i/9
DLXBFikLYVcC42Ko/icvBljgU6Qa9/WyFxKTfZQGVU0KuO7MXUvTiUVq7xbWu1uw2lPYTywvMfaA
/BLeQjOZE7KPSfvir8sKMmzWBJuYGjzERAku2LJqmKkZbnGIogKo6rIPZxL+riXeFZvRXKbPMWqr
TFxbcZQ1jdhonPn19ZmsjdSeGmZTyLMICPF2vzIaImLTqBU64SVNY/MXO3t3SGoMgPa7hrwqAnUK
gtRcvPCIbZ1bsSZwekyxEWCKdE9Tm1xsdFXwWt/vDSdSpIWy+6A5vLCUR1mvHU2F+ZalzUbVySrN
gCBLt2Wfd9hbH/lSZp8kqhHHYR7aFdu+3EpKbKLw2AAOVxhw7WDuVFgRF0MVO6yWIpUZZfAOLOdO
ViyCLVPyy161MB6hrQT3A5wyF1aD08ucTrP0TrsiKRILstCX/J2sXWN69QvARFpINs9G4KhxEvJ2
UyqAKaQozErhLEdUma9IdaGLIK6kcN7XMj2PhFOYAMUQb7vq7UxmSG6G1afJZUYIxn2OrZWsgX0b
VutxDIWXrQCDkh7DK5M+hMJnfV6tdKHh+K3282KOWvG49NHthoj58ovSCMZ6DKHklfuMaZvMqW0s
DiMAZZKJJmjgch2+u37bqdyhit0ilNhJd1idA5bHYeylnHyMkae3qI8zoo+XJdBH8lLyNSrzln3F
WoQeSgkB4r6l928DkDc+QDX/Um3onGLGAZi5GacpdwBjR3joWZmErsfHHq8Mc567s13NYhfiE9+E
SPtDQo3v3yvnxWkmal6XOckh9kp8gxfu8+1gF/iVRa0QpLXbLLlExZthvOpQf3+AICLXQG4eD0q3
T5LxpX4zoFzJHMvLJd82WFlEehVyWeBo8CW/qP0ITnkdkjkpJFrGORfUGoZAb9VUEAWhaeiUScpQ
bMxxTyzHqnBjFjEs4eesgreOZmJK4aiXGHr4zEFEoSBbtyBMUomMnvCgGQhgk19x1viJ809dKVAl
cxwjGsBjb2ZSzMMrPfCErb8pCKOJ5cHtuobjpPfKhMTChQfHYvBC1GpDhoGHeowMRIWDNN/K9zkk
ZCZcWAG2SPw2HwckSPSQAqQ8WZU4GHdHWk6A5Ie9AGzBOdeiaoa5COVbdzSji1IFKt4h5t7sbAQg
mSUWLydoSKCjxzKv9VB0X2/hM+d61qzKaWdGxpyIVrP1IosmbCi7c5fhgo+2VEHGpfoQQWm+EGur
GKwlY5tPRCPdchRvAUc55WODFe6LN6cSFtfEX/7YZEF9BJGYo68rfq8Ve5ECaP5LcXWA6E4tNNgL
x/Bik3cSw75i8eyjsD4G2m8bB+BvKiZp5aFGDiUJmQyZYafoUitgZpzlegNsro3QhLpIuUUrsQsd
/2ecZTfs45W3T77eRi3iYcHK3xBoOrrlbBu59mp8qEGaKVvvlqOresLkKtoCy++qtX2Hzb/OK35H
sTGBQmechpF92l7O2frV6LWR2jWzmhIvjZxJqbmnRq2NjFgr/5NZizRQ4zJdKS/Mmh7nM9vws3e/
AmigBjqmK5YBypOF4+EoYyLRDinBtfRCSNcGFbESOZOlS9AblTla4jO+cmhWovOLLQURbyeGkL1R
c97utrRheZI1QucrVvUV07hN7UJbjDr7tI6yjuWrH5cW6hm42kXaAm+qp/2rbTUG8+oA5AZ1zqvF
jGYhQMzveFK6SMfsWYC5ENJu/VvUYwO4HF7D3MxikZ6LrNQaYufZPmavnVn0STcFIjKl8Jf/pzoP
ie3drBCoZBfkSAo64TxgdfJ2NNVC9lqT1x8vdhqEnMzlVlPi5tYrNbK0nrHp1iWWquoglUZm8l1T
CFunBfDMmXq61GdbhNe/9gFfMOn/rc6w02HDDWqEf1hJvhhxBtsSGOtZ77D6lz4oGAhHSuLyK/7l
GvQ0unQXmWl52c+BRDJM2uVeKvFCavrBTu0RdzakFHFDr2KN6m1aORO3004u8RrFhCE32y3ey6l1
i49NFsP7eoXDkSk62qEtHRIlGjE5Qywffc4YPfkAEMsevyqsZTY39tG2LcZGyceW38KfmTgOr3sH
zA2s7KwKbkMUF7sfb2BRXyaMZsR1tSPRYbFyS+Z/ENtc4mFr+BcdpmXO4tr0JxtEidnX07LhPRMI
0lbVRLFHcenCidk0EVStblSFV3+ZRUKC+xGzlwulVhJGjOlaMOOFHPugrg4fS/m8SLgkFN21SZb/
COvrMsvCYMH/UkJHNchAueOZ7CmT9s9fsjexz07qToER/FHaRVxyxXmXj/Je3s6Z4TP1EsrkSkCa
hElYh7BJwigTtrYB6bQ6gH6omwcW2sI2N8qny8X0GhLwXR48xwoy0imsK8JNOS+M3liNYczxlHqy
BfTm97sWySPn08GFRPcy2zGcvdLtVscTrWlQDOJAy++mEI2hJOrN1IOJ0iy9UibUeLV1901ZRQVC
GyklFFK4kX/FmyrE0P5P01Wy1XZb77FUpj0kTBwouFAYBip54LRf4fBAyT1xf8GUu6Y0F+yymwXq
PnyOZwDEjnxEtCxYSPC+hgiFaiQUG3LMVB1qTgCmYaThvJqRniIttm1OUGuIXnNh97rNts7ySeoS
zN2WiRDT3gbZApJ+p444V1AgbIFhxvzu51SuzTMt6i8KUHv4JAsgvGXTZ984KViAyCs42OfK28Ym
Q4CWGmOIxNS76Ah9bnARyZWRtdRlbV04MBQFxtMMWh0382F9Orx//ZdmY4Fz+Gn3MZ3452YTc8Om
1piPehIqEslFC2yRBsXsyQz26kO1N7O/FJze23SknOr1uZYRzagdjRIv5hoVy9pGNb6PaMFcf6bj
+c4lmJApOP6IgMqlioXYOzVuILKPJsp0EKIgP90ytBI5n6CffUJYvzVWDOFxN7todxPlIszubB1J
/DElM+aTvvMMr6v9tvtiEKRLBp6zWXYZaCO2/7IOgf2zGEjbpePs6NADtPXQY/FcGhG6/QR8p6ZR
eO787oqUENxIuT2JWatoeWx+1qCXOVmGtMlQrm7J4ln9HUN/QTiBTjE7e9ywwwgtoKscKN6XoOa5
z/J+mJQcMj/FlaEE9IA3YaOAk9ZpwMs42hWRFaNu0jJUFiD1CxxP6xCyIV9YHLDb4ZpardhuxfI2
PmUxwiop2TGIEwwXuTNZ3CULx6cBuQWrKaa3+nG37pRBBLmOEZzb3Jup65/8JvTuS9AtEvYqH5VR
vvdFwISbnYHLSGnBKft66J1yOVdCL9H4BYj9y1CVyddS0EHQo/T9/2p0is3wcg8fx+tR7EdLQym6
5Yr+kL/TVbyaiSh5DNc9gpC1nGuThMtJMAS28KKWufniEuHl/QZDNokPW8kX2GcdTxNe52t0oGTP
V6p8naAlTc5Om0UKW4kNDyjKoB7J5mUOBrBAPCifS2DLPEUZ3XyNXJOPBqFHVnShbtqexupUyzkW
09nAeTl2NaB0C1jcdDzj1OPeN8Spv5pNaOpkenqZWUzxiV9j25O/BuNKkQJzXT3lwK1qwzU5oV0I
6uqKrAf7WkVCzWDEUQ/YlFgr8n13QJjABtprymPZA1csIH9lsYeg/lbMPGXMRB0DKXCpQrKe56OQ
zllzc8NuEt3s8dISpRfuw3EQDx3YmpY0eb2T+7lyPxY07WyKMhGpovx7kwDO2bUjpf0+XN3mnNWM
RsZ86RskE5IbsuR5I8gK45cN0Y3dykIb6ismvOnNJjfRQy3yP485X2/JrBJAiAZBF9gecHk+YxJs
L1JxqcY7fFaQTbYaA0vHgHUKvQnDMOcKGWez/+F2H4yuID8WT5IJXm6LKs+DlsN+vEHX+DM0b4s/
aUvNIRsiuidZ33gyOpKT2HqkL5fsCaR4AuABHiU8ROTyZoLFFZw70FvMS0kfQmXDykCJV7TZ4xUd
/JlmY+x2NMOoTz/xKJ7kFW80poybqlr3xTXozMbIGCND3BxNuKSALu0fRae/YtpRx9iwykAbzU54
9Eg+nGhy/VztCJlgEdheg3BQug0/cRuiZb8ExFR3i7fds7xKWKHGheNT3l72bUBBqeF3/EqcHZD5
nGbXUOKAxEWWtZvZEFa7RWIQLdxIxtUbjTP1U0HzvMYdFV5AmhiA2I1hlWgS3WRVYrQ3WR8I1OzA
UnVxPSG5AdzCSS/IuN5duzvEtLG85tJjurDrotm7fO+RI+wzvy0xsf7WuRLEU4B+YYGTdaxsYsqD
KeYGMKZTdfR56T3leLB9cZn9Jq5e203jAb+PpKKLMqn+8pKAJCJ6HmJNfgQT+SOaMBxg7kD/DV6/
sEjzxtJeWfoMeP9IElLGBACisC5BmKTU9Pv0CpEkb+RI02GPITOYbsLsTQL2C77rF2IokxeniU6c
uvnIVkbd7bezFtyBz5vebi76VcUsAIUp0AyOB9Nu6V0IV5O/qt95VhIBY0d+eCr/IpaCpJZfZexQ
jZ7UimUgrFVZDSWo4Oi5QpCfjPKPo5LjPT79do2rpizqQjwhfwAOj8yPrfLdyL0cnUAy4rPUa10X
ETV9SoIxQAqbLpTwX7Au0InfEDYnRXyzXkfuvBUuGJNJJiBdszwYwFo5LFyX2aa115iXl/uQibmT
K/V4Owqs39E2ZvMBzc3WXVD/CgBNaLkskWiSIVMCvOArNg51Iysm5UZoBi3hNDgLD2v88ddr9S91
rEefTaB6dsI/qvV0vQSRAvMqdWj/pPrn/KmQSCiHAxAGPM34ec0KDPuyTl3PULQPtwJjFL/KERD/
rWI6E+u+WxvU9yBAoxjI6c4M+JbPXdVCkZBp6THfaKvrQ75FCpoyqnIUsdvtBNQ57D3cNW3hsuFR
fk8lxw3BY9HnP9B1gw56gG2bkYBJBltdCN1mhs/sXVnz4JG93cI+/VflhtEPXJ7u++R66p9ZYMUF
8FLH+j601mZzSFFLyiFOYpj1GmJFpHMkY4vnM3WkXgvK7tPSm8fgxPKYaSvtEyg5VVRBfbApFE/a
LLUv6g2qn6K4Nj8FUfDg5HIosZmZcWlkYjzdb1pwNpQgrUGCPMp32raY7ND+7B1jrF/6UOko3Wn1
rc7zQ9sp/Bif0buWeb7YsECN5jeJdMXeMUJIX4dLrOH9eFAeil+IJThQCOaFgWoN7bEu7XaQxFcp
6N6tUFquSygrlrcsKHjSSzn/f+Rhc2ScmW7WLjqJK5n5qMDyju11Ssn7SGgat0BZD4ISgnA5gtfr
KX6jTKc8W2/K8tDSTxDtyePQ5KyzF4TexDbJASd/LEtxs6WFYFtoofJDQUy/Natn2O2hcuNni1pA
71iuCICQMIgGc9RpotlthR62StL3+UNwh3vIvTlywWfMAvF7C2VGs+TEIbBg82cI686Xy1GRFRmy
MhaWPM/v41sxWs3Q82vl/v2Vi0+81VeV0zHqecYjCkplqgLGwWrn9Taa8J43xtL1ZMXXOriA5ZjS
6eEFZY99+RzINly7nhm1IIhF+yOC3ULubj1KTabjoy5wKeZjARBXSOMmpS2Y1A/JvKRxBZLpgWWp
3s2XMuyuvFkvLK2bsxyTzmZPAmTeXwv8oVvqdzOCxdJza/z00kID155XEKjqdu2/zQC6R8Yt00Mq
k3uNzk9tfGCuDhEs3gf51H1P7jAHPbDBU9mJHTHgyWF2OyyzFtbpxHS+KNxwcEBhSJPCbRmh/g/t
HuUffwjjaNVGmlZ18hvnw/lrMG8XibQPHEWq3ytRDehsPFyE7ZByLFa7mKLDPlrsT+mFQso4F2J6
uRpzLiDFfa1GtkzHu9JjXmJh5L5V1ZsZskAZcMTd17/qKsGzUXe6Hji1n8Db07n/lArUFpiSkVdo
QukIt+VybmkG0Qgj7DFGHlgqmntGdk10W5AX6AF79QgXcPzHXp4yhZdaINyp8ClagKo/Z/VxjV2h
kQZv/hw5DHy66DR88ugAnmhauviduCKLxiqtAgjcuWxv98Wvtr8KbD+JxkZsFgROhSqZ2TzEjYYY
EPWRXZulddZyMpINrZBP69MzpiYKbGDFEb+J4l56bnjvyee9DXY4oDXtL/khub61D2Oqtv30S8Z2
epwSVzh5IaRtpSMTTAle41ATB1Nf00ZYxpqeBLqg67CXWPLvJQrEoRJwrhW163vdBQLUGdAQRwfb
U36FahIuUeMz8BAhpeZON6g9zvVDGJfbQAcHKEn1UcHJFT7sH9rVG8sE1etaRavalKk26H0MGRhh
msSrNcoR8gR4/WpLmJ4LU/DrhFUgpv2beNEF/4Ph9ibwbOriTRbGsviLc7Qdg4LKvzYPcahLMCy4
G7aj0Y/FJN+N698v6vCqYhHB4jqigZ2Gpt16k0rrDEBRwmlIwluvF5/4nWQilHJ+cse8fm5TFcBx
r7KnQG5AWh7lXm4UbfOcHmOfit/i3r6c41f48QuaTN+Sd1akofdT5FtXsUl0TqO1Ar6lIrD20kwM
jZSW+7gmJD+Bt3O0kSgm11ZHeci+oJ53+k4JPD4hQtt/sMWn7rSwN+pF7VK7sr+S4+nsVvVy2V/8
Cr2lD/DGUMBGGo9PGxkXSTmkPFlBPsveGZNlPQjbYN4pyfUjk1kUvPgokI4CAW5Nx4jeV9/Hky2W
Xb8YVVvKFAGfEjSg3QKWvj5MnFRlIrD2g9aQlsAiD0aeASDgDKLya0i99QSqooikvzPTD5vpluFS
mq/QMDdtgr2gZxLolcbV9R6uu64y9DF9MYX3Izpxxvr2wC9/GyW3sdgwTLZhKdP7eMZxNyQqHuzL
Ci9z/q7OB5b2LMvUX35IARXtQrOPm6G2ut7fft0qGklCmaLb5uJJ0P78u7r7ZpcU2dhfzNL9Ol6W
ZqfZ94tsT/gYkf6YYYPQDSM0z0wfFoubKUF5jpZPmGj62Y0fWltlr0aayqvPyaMwa20G5kvYo/c2
OIesCH4lp/sPNKFllXTvldbIEe39d5lalSL+YaYZOU1vGeoWj1uzLFK1YZ0bmtSLyG2QfZiVcqtQ
6lYzZXrlK8/q8HwmsSnhe+29/Zn7wnMCdavvXNs4Y7WTS6fsu1hadh3PGztgGy48mZ8tINqxN9RZ
f8HDp4pcOuxgKBwr4E3GgUISDNfHY4kcJKIWXg/zwa7ArNvmfzGu07I03Llsj/0V2Yt7SYTytsAl
jtXst2Dia83ghGGZVgc6oUUMi4e+x6dYfN4P45jXgkdG9yVfBLR/00oKqsIF0VtYUD46Ut7lJc28
MTJCxRk/3hKqmUu/6XLUW0ghdOFh8r3p/yX58MDxd7mfBnDlTXcDwHCAUmHqf55VzxoqiKhdkV4D
KNg63WtFE/o1cuu7Bl3CcmifT68D9caVAkl/+vM2ndz+se7qTpv/LDrZo13fZmWs3gwuXoClWo2T
gvi25a9tyLGvGEarfJO49DYwgmRlaUfkC8ooMuCj2TrhI8bJqU3tSF56MuftEDtTCEqIRqksInCM
lES8u/9eSWGan+Moi4Ozyv5L+8SbHeIv8rYvKm/fu0UEbiwABq3Ai9FGyPeVWf66Vk/0JP/ZEQMW
CjJYLlzAslY7TO/chhy9anoEMrIhy2ZIVMHlW7Fxukv8IsdDU+fBD+1T7geNymdBdvHD/SDnx5me
LIGMsjvD/wKzL9NtAePfM1exY5a0WMRraSJHIGPukQVCW8zhh2UPCYnaCkSghWgdTj9gkPcmFO4v
Lw7zxkwVJNZU4omusgUrjPzLfpxyyJxoGf/8pr4IbxomVRr3XeNZN9qewuw4nGC6z8Mw3weX04un
y9vmyeualx+o4H4eIN+tovh6BJqkgCBCmy+ar6ZgWXrtJvcSPzSKFJAtY6dCPQpRFxsTCH7VHdBp
2Lq8DBZkxHS/N8d9TNCPRT7+NLzJldP35APzKzOjqSG7g7X3CY9qY+LBx1G0qWmGi1QNZL0UN8B7
y/wJrhyNiqKVT6D7PjJyDDn3GWwSWLfvk/Zdt+9gZpCkgcNRmr9+f9SM69yWmBvGNGiSjhklWQaX
YVyTzEGPTmv61OQUvMP0yjjwHCKKMSCogyeb3t059pjMiz9j07a+mRNyyLbMUsYv1a2MGjBxBNDq
nlee+vXUpCgm32yl3jaegqRI4XlpZsStMaZAg0i2sOU8HD2YRnYdOXO6P45+W+B0Ejtqna4zW5iM
gfGg0pXnrmeH1RBAfhMN/IXZZcJa9zcoIj73nxJ/rzsQUxT+B1qaLYJGKxy5sXhoTRhutuwE+fsc
qjirGDxSKJs+T2BdqEJ5wJ1qYcZ44Nz0f2JdTsBvbhQDlxj4c4HoEO9dNhkvQWhpbThpqfZ5jQBY
1g3W3I67IRtDXMC1/J0917vVhBmLXw/qDfPw40A/tOUA9yZqiAHibzsivBdypLk+yiBOVYPwDGyt
D84ofPU+vaFVvyx9HXP0On6gtFCD9pZB/rljkkbn6DGusyUusEgPLhiT2Ml7q4ZPH8bPahyxTrRm
QA99ppW0gJhWzRbWAlTV217q7atoRuqDq4taDX1xCEPD97+jglXqjB4tvQ/gkEY3+yZfoYlbs3n8
nMclObtOFuF/IRFNBe3vEBYefkqZVEe7/v40H57U9IzhwmrazwNdiD+B70hJja/oETQUyVH/JJzL
xDU2eapR6ZZBgwLKSjtcU4e7T2d0lyTPZkX32+usDe/0m/xu65TeEApmUm9ykx565SLlLFCzoXC4
G2CFGzsApa5mKWUnvp8pLfzw1uUBIVDFw3zdpLyEohwVULKxvvjDF3dqvuv+4v86Zny0e3OeIpsa
G4QLzTdd4atZ4rln6IuaYAMcC+X+j5Y3yjxithi1JFqoyCeYEsplUtwWHReMmLEHYkTveIK2oKra
5X+6tBW6z/iSg1EB2ib8x59wn/gpaI0zje5noZlhg91xFLCyMmNZ9FpsuayuQK05frEVKQtFOvy7
/bZ/6hLWlcRjs2/YvYdq1lwWyOz3ITnLswonvbUOPsPfPpqd9p9rzdMC4XwoSTfsak5UyXzbW+qT
LeE1bcgAUxWC/3hPP1r+PcjWIZgVmm2ETiSWE/nN8P3vKg/kxWq1Ar29OVlPaPokjxg+9ACaZ+x4
xoXRs2atEagokkfg6su4xaRVSo5XOpEmQiaTdybFI9eGXJvJLFeZVT1i4NfqiJBNURiFB/WjWb0h
qZD84Je0/0cff3Pi9v1UdrGUnoewhD30oP+WHotXbLViozU23UOIdvHHDefi0RlXTYFgiGooaanC
KKqAcNcRf+qsQ5X2vQ7fC22NcWxnNDvOw3zbq4eH1RvgdYbBOtCshDMjdp8u6+gAxHtp98aOhiMr
V/IrGv3RXhitWc+yttC+lI1Kpx6x2LuLLVxelMaKmG5W2TOuXebhsABEg3ukVuD+cEdWsuTjZ3YN
U9waqtyom+BQnKh2AhMJ6mj2qCvuNPU2cQLXFio2aMOINkyLUj+1CQVfa5+lpep2Qb0MjDXNZq/i
avobWIT6r0Aqkun2f1b6umYq55IFvzRxcgPAVG0kRHb5yqt94Ta279EGPCzVXI0P/OeVvLXWKgM4
TYiZxFzrWpnchz1ZMOr7Rtn9uP+o9Ei+jkjTe5ZuZIZYYYxnlp1HvgSyq9cIKbYRJqUobz0jr4Z4
lYpnx6j3MpZELUN9MQzrdtl0RArvnUiJ2em6E7SBrQByaCHzNUB7lxiOOKxsz8FM4n4dVe0Aw4Pk
Kt3ys8a/yXrDBjZ0voz3ajKXHYlN8Our3SEKQOt90+H78nghI/AdSYayCpMEmXo9X1YSKhWzJERt
VJInlP9sEZq2nKupLDSEpL2BNsdoNGhW302LLkuyviS9SIvzJqMsbi8vLm8ihv5gzehHdjJKRn5K
fp/Qhe1uWFMCcKpTax5BC1C6ZKGhWYq8DN28sjuQTTryqQogepCDmzQV2ztTmFJ2X9BZui7A2y0v
RB76dKgXqJc/54e9szBRfGbRFJUixEoYw3oGPRpguz65cDTViEZm5QzAm9rvUY9gjwD2y9vRhcA7
COdmH1M/qb+OqFg0KZzCv1WjvjgOcW+1e9J1aPFXGdAAVe4RP9vdDAaUt5oa4MgUCHA4zzTvpNMY
HvtYwTBLYtl98LgU4Uq+prNqA2SEItmzHc0z2eWjebpEsNTy04EB7zlTNySVWXOZdQTnvBhdhSXX
TMUtQEC86gnW5IzgyeQEnD63elPwISn75xTyo55V6DB0r9RWo5KZYiC6kNyIx0jMhU70o+x1DWDg
1BM8HR6HCyzYOMpJmZtClqE0de3yqlijZWELYjyHBXsr8vyogDrPA6329QKZfSAkE7tz5P4hAV3/
25Gea8CIceEGyzg5e4BVR00m3yS5IKO6Z6YANQwP7+dBtWOULnNGqUKkTQKWBYfdDms08nJdVp1Q
8z7Nd28nBQMLqGNfsFKE67XXQuS3xk3LWR9BCZAxagmYO2iZtdnp9+KTDkbCBOMproRsJctkE7eL
T5VMyXS9Lu1RGiOfbX9s5fsxKFL7OcqgV+NWndFb+dcIL0Fd/rmwwBPu4kv/0e77NJuOe+I8M1vL
1WtveDMvV7yjG5asWaD1CIEgLxyaNxXpS4Q4oQNeWtpMnePLMm9htnf0kbC7W9xsISFCwJHqhxme
M6fIa8iYyvd7OgVRWQzuKxma5Ppc8Vr/8XG+dT7+VFbgrt4usKOWOXnmheVA6J/NAJ33XaJ20sYd
7eUIDO9Hvno0egJPas/ut1YtzfyQjpIW3ZtxhIMQGgnr/IBNkNp+KjHINg0QC3UO96PcMKOjFDyp
7z2tALq2JasYpn9YorPNjN/KNX/dwiaT3RRKVbxTwieuO3m+/D1Vl4ATMZADLvlC42KXL1BDU9iN
6ozQeVbHsylsvBgvLPyCs+3AXyUjzTsvwNr9AVGdiPFdqkZrOGK/S+m24sQ5VG8XiKaKVj6XdfUi
0M0urFhv/sXc2eLhghRYSwPEk+/MQnZBG8/kJ9rjTNuj4a3WtcWM/l3atyBcyzMZCL/a327TpgqP
PftwWuHP6+paS/XWwy1UCHXy4hEs7leESqN5iLQgGMbdD18UK05L4xsNv2AUY1oRvHUQNGeI7dXk
0ooRXJ70+BGn4sIaLEyVBR4yYleIcD/tSrr8JOCaODxRL00DQt3WNc3dezSICcDYE9f0tTALgUvQ
40j8+mlFlE3pNJNtWQdakLqSydlqE4aTznJhvlGYkNHzxy4YXtc+/nBOSQHAs4fmg/jPDM4PAT7r
WKr1EzDhY152q1FKuqGJ2steH3pzVQbhFP5auyfqXh8f9pgDchFNHxwx4+DEx72MxonQ8g2DCXZO
WnILIl2d9HNFB5GKTuDUGfN1bo6SnazXd6zJD0VdMirE35NitL3+tP3vxukM+WVHCXaMCM+LCHnX
8SLo7G2cFFDa89NmVdlBZpK/OoYFoTpV1Gb9KGZG5kKlGCQU9TF9FQHziFeFUJk/fgu9TDLDm6O2
WPJtG+FYnqj/hmoWfNKY1S9fhvlIWrYnj7KFZ87JJC+bUbW83/qfR+/fIXeSPS90vmlRVYrWJvwN
SjjCUXHSwDG1OVK8vse0zuwe4kj3UIDC0WclRNM/Q+bn3b6mY/aHl5phplH5SrYDYFtrGMMwaH73
VaxdFvBLYB7MwODfACwe1pZol/scpGOWi0oHBCfD3YkETWxCwQfqcKjlmIZlXTJ0S0Zqco4luFC1
2U5EonxKv59VvcTDbjXtI2XFKBTDA8hOpxWZ0wMMRJg9REcb3B9Q81vgJ+DWau9KHzoEQaa1tgA7
oj/Yd8i7Fa8lP5XTdTrRfRh3wGq+gUnWtVeD/2coaOI8GTRzpxR8Lg8wB6VvjogHS15/NJmYMDHG
PHrSo/a7hLA29hFozKEEZQxv9EiF3Bh4SUD5qf3IW8KH5vWMkIi2rZDnJrPbme385b60s8MtblLd
ZNTJkhMiQvDIbljp8Bc4rTvqKylWKHI5kmFO5OUp3FJhAu2XfpZsRSgGyeCVQtCwm2ihP/jH5lGE
OSCq/jtseg87qjXbTAdc/DHE6VsMsJnsFTM97ADmzK+BUqFDvmCKac869HCWXUjz+fbcND5X3qx8
rgE3vPr/cxRoM+wkP1oeQfyI2NYivPuGwz2umIcmJTNtPdF9Nf/iXrUTexwpaEr2av5mOIuYMzkb
HEkHipNkNo5eq01o7eoO4LmB0OkqaWbOWeLqfPbV5fBwvLQeM4Vl/ZKuyY1JUqBxuRrklvWdvD2R
tHPTog0ZwKw3Ng4D+X37lKyer3zugvaSM82Z5KTUXcDqBfAbckrBgwVvWtXI4Kx0hY0LMXRLD53g
JsOqPSDDAJsvAcxOUDtzHBIQl9oI7CY6obHhM/0Rsvvkf0nYMKCYb4xflczbKbJXRWAt5vTP25Iv
bklE8wGCXpQ35bNUrCzpdFDwiHtJCx+t7BHjLBxAxqhciIEblu4eUz9MAfSdT5YLFb3y6JfPyUlZ
Rz2e6HjJI16PJdh0FJvmcIO+MFTQgiB417Sm5hRzf3Qza6KhINDacYdnsaH4zBBXpUgkWicusWEI
EuRb9Mi/cPK5ILzFVDdOxSSMSXAEQbevwB3a1kDAW2Zk9cZL7f67ShFVmrNpgu83e4xUA924Bvjm
21vNMlkpKIOV2mCB2VT/OUSQGENHLtK81RhL4QlRRK3s9y9TOTuQPv8hdm+hZgsrTHHdXsxmADuf
gBjcX5Oid/AQkB4CigQ6vxAxQnzw95u2+Ha72CW84YLEGRL1Jay9rTQtKCUU1LB8X5lElFLiuAJ6
GkuLCP8IwkTw4iFtenACH+v87MUl6QPfSY+3hwk2U3OmFpVgesF31DE2NZrQ3CbRHDXYgJ12Ukfx
5eMG+wIDOQXKnlhRIYLmfipKuvhVEO8k+QoLoYCQ3TJr6LRrHjd5idNnGY2d4NBA/MnGWG77A8kD
D2RHbYQgGTbf0B9uKkIkBxghxv5CzsVgdPigthhAdB5KMzZMiXoGe9UFxFgRMYbnQK9M/wa7bp/L
MBwMB65+awgpALKQtZ6jIbCYyqU2vojGR+wO5AjIBH2mT8h+UvEnIY0eT519bUBC9aDfqA5iScT+
+Wudldm7iVbAz8i5UQu23TxViilwrFjp/+ML8WUQIm+/fDsmr0xCtPPgvaTiIcMh/Oa1eHB+n3yM
iBgVym682YsnXjkEUnET395c1+URALN+HTjMFwIUjTuGxtV5yJjevTYqZlRnPGd2p6RzNGRyScNi
WQdh20fUO/9/JuFB26pZo1tuiK41NWjXh0HS0cpUBP/rwzNgMHRNXNRambFAncP9aiwEe9xmk32d
aopuSxguDt8xuHBraoBJJBKuqlB+6fii4Mc1u2VbLSWEcecuWvtMuaB3MzLTDCStnHBxf1JOxhLP
0oRNMji2tNIvD7H38C0mmVOsHZFN/q2B6zrcy6OyeNBeQr31ef1SCS4XisxCrKiNPQIPYD6VgX+o
6I8RJJLVF4xTi+F0lJF3IiecWLRmsSCBSvi1KBJhnDM2Uwm6DTRvB+OxMsuwpX/1jYKKZ7Am/gPR
60KkyMEQ7rNzuGrmH69X5u/OFtZm9LW3PHJD2XhltEv91EHI2fI1/M9LUyN9V0ktsgPK6+8y0RzT
lcCLLF7Yz8ZTR0If6XpJEDNJnXejYybzUQZyA94I5x1Lm4S0Zwh3c/oY4r0u9N6qF1zLPgW37DdR
dohspf0ZL1neJuEMSghmDw4PIx7hL+2ZYTs3qEcZs472lrkzBD79SsaxpGZZgMQT3Fy4aFqc+NzB
H9bsnPlUXwwx6RgRP07r8XTFl5wePqxmuJ6qM+7guvT4ZZVZRhM9pMOuowNhFpkHU2ljGFHVPZuk
iHhC199bWXsP9Km1Dhr2rNqjhF/nRh1fS8jIR558BMtTgUxcv4jGEppRh6n0hsP4QSg+P/95SqLg
sPqRNsRzGuS3YfWANFCn+MJS15eGwQ10e9Icx6BOy0ur5QvUL5uMqPo3vv+/RIQwnIAGuh+7HM3J
vnlFmWjGWR/ww4Cin2qzPU0zjmORjSci/FG58A4hi8o+/OMpAv31DefiW3/JF++28E5nJjqmmnk5
//LKslPWHUicih55XiYMF+J4Rh0bKWfnz3pDjdrq/rl5gC/sMjpxd/m6xTSomGLeE1FJ0cnJs03k
B+U18pFG3KzVCEzq3+8nDUV1T+ey+3WM254NFJeeVfvz0MJdRB11XyI0gk/Egmym+dxksrjpxZdQ
bhiWp4fWBcwAT2aMqJKiHA/iSelUxi/KU17r7Gibnmrqj3LENWaymPYUt8nHPjl9pmcZJupVOxGE
ZKd/PuCpGqsaME9WHLYf42s1m6HlO05jQKq6ekN7YMw3/ChPIvtNK8vr6BD8/r3zVW2CMrvt+Ttf
U7J2NBvjXJgOMdkyTOPJcnicgNk6NmUZRgsw+rZRSEDshnF2wUwpWcX2GTx1qUIZ5zTcstgvIWR1
SNASWWDbccj/0cTJYuZY9WXxWsE1Sz4Fb807GItZDOUA7Q2poDxcGbpLBG5CNrxUJ+LCNOxe8U6N
J39Vv/+JbcA0CTsZAe/UP6gQBsGuhQpXH6+kVWFFuBmk7vLO4wE2dMveBzlCWjDSNgUreETe5S47
Mqa+n/9hDlAY78oTTtYr2p6zTSmngRkMUohs0JU8D0KN5r9WDgeobXodt/Qm2wR35HC02lem7GF4
lybZWSSuaZan1c0dyMLpByA7EZtjBqcZVrVlWpZLUlBvOgNKIWi7Q8ENSETFY6Uf89jjfnIVvtXM
AimROBTXck3iXfTrbhlA2o1JGbxioTshoAVAVD+Vop59XUyRjZwQl5C40GagwicZokIaSe5P7gAu
ex2V9l7QrNc+VdpDI5UVvP1yJOZ6waC4aWFeiP3Ee0mJEQ7/4fx4IyE9LXfNcEwB9Qgd/a3W6cyE
3Tqd/cYwpfvKobA0/QBjYYy8zzk7NyJ4de5zvVHDUYDzmeuVJmUWlffqsE/8I+ES+IWliC83Wuny
QRXZHcz7zy+Blzm+WYtGai9aWI2Y7b8duzQPr5NTQqF7cDkUBDfpwI58h5vgWg1rMiAMMeBEMvS5
yuFnumIFKqw0lhx9i8r/I5793kx8KL3auyJkovdMoLp3HUWMLMBPfJoZIeSk3m7l7RM+bx+nha8z
MAyzyFbH5biSdb6jlRzAVsvvT/2WElmwMafiJbd6Z8c/Xn14Mt0Y3mJIYbee3akUvW+qaB12K2J1
ZoIRvf5OmKkEZurcc1+rs31EVHjp84MQmR1hlGzLJxon14JgNXY3y1sZwndq3aTFvM6C31w9xhBS
MsXLLQ6qowxE3V7xbvaL9J9a2If0B2TqBW7dA7pcNcD74R1YJ5j8pZAKiHp+SpAKQsL6y5tveCCP
ZTMgNZsUybsAwroCwcrffNOcyupd+gHOKw7mwv+tpIr5HGcCCOJ/rPB6Ur7yYqzhBHtMfE/4+Qvt
l6qpG3yph5QXvy2hIcRMLyfLAYpDfUvHtQ+DYd5dOQHYK1CneViX8wVMbzWyhHAELfcgFrK/HXsW
S/uM8Qmr2s0CbOsJFlSY4KoFlSRX1U0JRjz1CKyqQTTM5obBUeuP5yCSosNSs2zXhsK+enym4Zl+
uE8CB2KRalMfQBiZAykY8V0NLHx0KPdHS8OE6rBN8UEXUd4wO7Ou+yl4l7K6LeUr6+vMpIHvD3JU
JVC6QH1uCKGfiiApsIG9Dr7mdDtedX4nQOG5GseE7xmCVk96IwaKtIJ/S5nTrvb6if5VgXKl28lQ
Sa95h/XVjze/Tj7ZZ4mb0I3wPDg03BH15ZLzlqxN7RsgWmQFBEslIsbDe+aSHr6isZjjFl7c8Zqz
P8Wi4ERIBtjYzeMnQfxoKolPbtcuc9UXaFQpSIfwQzKgVnXWE9y40rlVMgIXt9pJole8ekTYnJsN
3ojV0pzmcLUyA/oQK12Q8yvBNHR8iy+ZdQJh2i/vWuYboWxfOItgJ45KfNMwvNNT8TEKvx80912H
6AElDeQcv97U6qA7I5bqCIoeLD3zvupP2smvuxIESk10/XZ1+ZU/NR+/menKdwiGrcXl5i+U9WFx
QLkH+3FqtMHHvxWVeJFc1XFZUUAzuETkX8Wqp17nboono46h2dAkUiWtA9tCpns9dISJE/L7sSPD
HjX9vD9HPv/YfMXfishxYCk31hwUchVCj3kCgi/qCLoICCe3OXKKqZ/n5n1ezABBDAn19vYDulo+
k6J4qm74mPlAMjn6IMIHKXYfa6lHubyC9SF6JwQ4R5t7034G9yfB/3z51JqRr/kwzDHVWw8u1Qi0
9N8OWH9HJNquPYKKWm+VJdWz4pCtaoE6lANXtPi0yVy+8zRyDHnnDtgR/x1s4vGtCZkQBAcDOjiL
WVY5sTi2Hza73UQ+F+4r117fs16xAftMO7j+gw6cJBfwGZD9CX/aB5AhIXAvP+PE5Bn4ZVXlTjgs
bNhug6mpG6F9KuCUdfPF2LjtiEX/WYgZ/v87E2ocJyz2fNOgBz4lfirqMBlRt7JyRuu/docX3ztb
7MEtaelEHUQzPcHUe/jyZvyh64psOK8IJ9Cs2aigJEnAmYFN/zJjLA42iEp7k4wWgzL3Aak/1rNr
nhX6mnV8QXcV1b8fv9DrTWCvXJswYJnd8TC2LjYKQ20j2Hpt4xrrdhITrVG7omTILvwf9ZS0RSBt
YxzF+eqw9VrcETfJE/z/6GlofMQCj+Go4H6Kxd3k8zpxr26rT9IlSded4wU+o6PBxYNp2D6WfupG
4MfyaKaSeYXcBk/4CdniZ1d4U9G8XWTs0zQeMSYh3UmhhkPYTHQQUZg9fkc5GcHZIdDu3ot6E2ZE
ws6+sOmF1OhTAqoLo6wufUZDF5Mep0wQYDeA08zV/aGw1l5CNqyVsPcAhsdKXjcSYtyw/XUbcQOQ
wduy+mw/XJ5lmMdlHcVeQ0go7opFCs02Va+VMOAysu0wKjKnte0WLQihDx5rpA5sCGmz7S0h0zil
lGPX7LCkonyQY7Ynb9XW3/JcobagiSEkG0hP176v+8itLQJCp8S3OnWfvotiYoM3zK+a4Gmo4wxc
MNO7CJqbxIAydbTTIbo2qjO6ZuawSVZLwE19z4wzU5GlZZAZNFwnXjDauWiTZ+XwYwAfFklJ43kb
F86r6Cu2R94NMB/of/6gKnhAR5jEQMEYWC9cNbYPfPr4HQn3CT33rogoXnehVgUaz4RMhJo0cmP6
K3Kpv8o46f+8kU7U56da8JPhFVF7bw07ij/THX5lu3vnW9ZyFrlryCqkYk4Zn9z6vn7V9J99Zu0f
M7RlP2ELvgcjlsIbKCaN+xTUS5K0e/Xl0OxSs1pdvvYKxymJuiGGpyOnORdlYMuPgCb5tj1NKDtf
7gzasaDI6zn0MgPysAwo/E14MGlJJGaOgShce+l0PJ41urxNS8wKrRizh1lMIlyYV8Y2BSKx0Im3
ieMI09qkw/RLLrO5Z1cH2N5KaJeNUCkFHzxzbjA9vzR+XCk3PV4Rm6l9/qadl0xf5W0A5ihvXZoM
tHgZkG4AaRiziicfQFjwCVran2QaU0hpLaPv8K/HHAb/Drkmoa0mg0r3EkNnUeeYWwg+zis/y9tT
vS/PQq7mNCM8fSeR7Atnxdix8HzCa6m4nA1FAWffufYQud0X8l52HIbpmhJc6JaYQEOL1/67umjZ
0GAyI1JT3uvtbo7+6e94vYh2213pGnTuZib8u3I6cl0uvVjBuJHuENowWsG32sZxvEzjMpQl/u3f
KgDfBABNq4LXadKFBmv3dZvDBBuk5OHCgrIujb0HedUsASUosXgZh0Kc/0PmKipR0jIfG2t6WqPr
sRDWZZ9y+OnpWYIoHq8HLlzaOlqP4VMh52H33sYAL4zaPQN7r2VhFNnjVafdzPdxqAv0z9AaPVpU
UfUrMXVwM+JrImCMhHOUZYsBBFjewctUrMrkDQUoPpm7SnPGkoSeQlEwiif/J6ww/3vJ5nzaf+ta
BKolsd1M4U2v7FWxpFtGwG60+pfC4yvrprc09DVn8p1hMAKCzg38DGao7CYw18HxxzfYnNQI7qkK
XCL8vavHo8kqdzBMQXXkpJUQJlIMd0sGQ1uqmmpkZJQm4/n/TSsj1EJIsXVSWnlXLoKUa8oU4PyZ
zbljCcvtgleP/H+Yk7hAguLYJvD+uRjWAJlgmvyx0jlAxfZBjREBxzzS7g3zOLIsl62WIWhYCCgi
dW2IdI6pFh+++AwOm7dHAh2hwDroWQQACkXNaFFplB+3LpDNQbglD24ftNnmpienNWKpSzP3dxns
DsCIAt2M8iMuMDTaj5YFYUkxgSfit6hok6VZ66R8m8INC+MV6tdN29EMEhAy5SSvSskMbugLdlQC
KMrdn1Xt7HMBcezeqDIQSRInNHVErTnhbbhDYFTatLieabxig7AgKWybMpJxm2SKJkAv33bGmp3c
HuM5c5KtPNey7XwA1rC2CjQhckp2x0uKwfw8qWuSp6ayEF5Q9PmZkQL4+B3jOpCWWRpej9hS3x/Q
4QyHICWfsa9BH41yvdPxU73OG+8WSmxMIj7qZqu5V4px3z+b866TlkADiiq+I17nyQVInb+ayt47
XHeO3jjfYUwQ1JKTHTCe0VXPC8JPeqoFsNckhlNKMQm33EnUApgYCVCezyVyBpXtxjIo4tSIX6+A
m1AIwaTi2A0Arbc9NxjCc6zY458TczfpJPVgVA21Y+fNqF12sdIdaVss/JXml0y/Fw9KyVyE8t8j
FG3GyaFp5J16SyU8TtPBXVamaVQbF3Js0D8aIoAXw0QoMHMFH8qs735AnJi4ArMr+sBt3iDxHwRX
AZxoB+oRoO071Z9ZrZImfmGBHjaEh5DO8cw+k7diap9v/R33X8ETMW2i84gs5n+stBurf2YFwNNi
iXupt8CHQ896ZgVZUEE7TyZmv0UGSUMpForODFPiB4s+n6L0BFJZVUzc1YbKdgXBvuSufrwl4RZJ
J/qrAAZhfXadKakAnY0WplEGag4hbInL6Zf+RrXUsEjMHrHiKz/wc27Qn/KbWeEVbPZNjJ6nqWYU
wvZzm5gPcShwS5x5UdTwVkBuUfhH4XrZWSD/FhC44MyPvKv7Aw+8dHni4xrI8s381o1carhAMPfC
9oMrBhhwmSzoTvKUQG+2JvYS3P3uGceqXCSyjOtn3cGMX0wFgXZB7r2jW2l6HnPn//VypDsRsPT9
mSMq3JtG+OAZ+FczM4Eix9exvJrG4ceiMsJUnel+Y6esFRjdYHODk2rTi6ZEnJV3zhoS3ql4wmA8
WXJ0zRwZKUU/N3YSyOXBCrompTrP3gc5YuEtxUBydrPEA6EMmfdMmcXeu1cbe2CRX5Cg3SsGKJem
MSlUctunZdpT4Ce2lN8KjmqJfFx0BFs0yE3vV6rUmn95C7thjIE7L29Zf6jd9UlhL8Ljvb7jQqYV
alKQyaZ7xAWEah0SOt1DYaRU/SzsE2GYWtROaNGJp12x6C2Vo4oQoWQDCPH1GF0RUQHpx1b36mMd
RYnc3Du0zRzSbqgWCzP/PRuZ7r5YsyrKsRaGrKuD8Na3hRC2AElKXsimiJTRug45wDcAmnbjzxAo
MxMKmWH5WUtbRVmRzABwA43SpmGZhPATGF/c8bw8kpdztYZ6topuZ8IEd30X6yf20ZYOD7VfDkik
VbUQwp2DpaLw5JlQCUSeoKSeRPMeSEOsKKVR0jM6V1YgrVDpkBWfm7XEOjkK75HynncZIwoBJstF
lfQokzG1QAQA/n8ycu5PUPTri4mWhyroSJWuUPhgCZx1RwynlofYcDrvTM6MgpjIps0Bok4n3HNF
tgORE2fQi30lixOYDc59TVrwVmjkBgWAVV5dADxFTztUrqH2XrOzQHjUUrHlqRx+l+RMW9RWuX0D
1Nw2z0bjVSjG0PryVsb1HalE1d/G8CuXd06WK4OppkaZs9DxrlAhwJ8tMpPj3T7IlPSZMFwHle6/
MuTg671iytK/uO60llA0dzelBCEDz8SDLE3CfJUb3hros61B/fS4PLr6IudfLrvSXH/C6HchF4pV
roL1Lrc6Wn8ygIHC62EAr55ZFcp885mhSvKagIZHhuVoV9PJyRub40EcwmZl9y/zzFsqM7MbXhdz
jXhChs6VscybSlKnWq9f6EWSAS9H8o0u6aVje7zAjUfKj1HWT9UkDDm5AXriO/DZtt3B9eKcX1VH
5M9SB8+fPgSpZScUbM0XsmQZ2W1iFgCQGZ4/gpEsYebKDLJPvorJ8joWIPOkzvyZ5zbpoJtN95pO
2/5i79DDzD+vNgCONyZxwivwLdjxeIvuMytjq1lw3aOzj8x+ZlInItVTY7lyXxvlkgio4gUNzXnM
CsHlZ+dVzG1Y+bJhKmA26eg22fpnzqDax38ZRROmN5BQR/ap0WB8FM/uoIZK74Lvtl+UoO2cZsl4
mGuMtDRe/SNY15wZneCm3E1KgEoHlMCZalym2wXJe3pKwmh33xdx+EhvS3QxUZvFbKUyXP0kEg27
xV59GsHgMOPOSQLdg3RtjkAIH6hFfT4JRtPnFCRl+nk/2HZMSgk+rhnEyAT88oOJm+2+BtJnVXZ6
/9gT3UA9/d1uh91vCfB/BB/nVsNVjilCHJJcdH92oPaoBeFHBhI4VKsRlo++KIG/bTxY1iXEW3dU
nevWh9LNk6LqE903uK7hUgT1j/kpJySzJmDALCRFxGSlPXib7WctJyC784oFjS7ac+TrdCtCz2nh
rbui7Go15HTN2v1uDGfhfaNlXiGVgTpcM0hhwxinlevnRfPAVnLxz0C+urMvhaCg9Yrcxbfauc2E
pUHJ/rgVwjAxkSXd2XJGzkIHr5okfU433fBDah8UXVnYs9JWrZAPVJA+ayCm0ftO0ZXUc4p/ORtR
BZv2XrCUb+Pa9zbqUuWy4SeDTPo5OJmch62vdMqaOWAniMGp2lOPef0LU417lcp0xf4FgaLefmhf
bDqz5w1ibAQFMTpdZRj8uMkWTJncmICg351oDGvWbTOpArrVfi0Q3WKQ1uQwQ/le4EJv5x20ZgwP
odQ/jLjulHzdXDaFQDLaFnYX+yZo50nB9ns8ridNPOVZqnwGsjuCIDlYK8UshB94xTj+A4D0I4H1
XIw5CFksg6HbknWDy4GqpxrEfeE1e3+iEpqe5b7DzyqXW3ZRRY7HDVNlZYzZK4+sfWrkpdb5LsbG
n4BWkBAvI5bSpOmPMX0B+xepWTNTUVv2zS/OeFIHlMMhhZuLVh0aUKBqFSN0NkjMiZwMGsOTaLso
XZOF925+12ZMxeOsbkdFjLCxgnwDATYiUcVs2o/VTwS3ztI0lmPDiBP/ua9hjqwOEuYe/UB3JakC
0LOiaNhlh8+q4ubz/IdDD/i5DTHcKdmzWRU7TC75SLMxZkC5wPlSlytFt5LZ6FL8uRkplGku2ADS
Wvz4F9NOZ+FDjQcwvwLnj/ZJAjJeKFpHSLK18Y6Tt1i60vR3zuHpknE+zsCUKCyDifAyUGm6eXwG
PFLNfKboNNSTAQ/eu8E2JOcn+50fhBGoEBp4PwbFDfcSxgb7bWcCxFbOJ5MfbaIBz+rvES7THWWr
S3UsS3M0g6SfpoI6fkM8C3A1TaxEeN5O/YJNs+eFLwWOFn8CXsT/IgOlnZRyqash8GaiwbJuNrLO
C/ZLwAec1wv3mUvz9eoqUI5sC2CnT+yNmtsst20LXKodHx2Ghw0crmS2APqcVcApOyoXrlL+HvUo
+Y6a4yxqhBTaDpPNlXDRpIVWjPXP/5NzHufBTlZsNs8QFnv+bdApQeo7Ze+PZ865YwMaAADjAdDS
DFwI6w23CBvMR5RfZVjKQnK7sszPjFvK8OFgk4Brhre7BQGpxldJiWe373EmOydm/FWw1zHhxA8W
iVLsGc1NjEq+MEm4fY9j3StwUPWsz9ejDgLSqu88sXyFlTWsf6Acm3YYVojtD9DepELwIXw/CkEn
0OiBa9V16QeWYQDbimI2Yr+m1ekabqNqpWytp/79z2t0i2pj+weKLl5qtkoHj2aGGwo0i7r38m/5
Jp/RKhOw5bHZyBjbez6FlIHEGOWTKkjejazYa4QyF/s9T9sYb/jlYyBgnD70xxniPvDgE8bMDaMO
OpWnxv8jcwMRp4s73UX2hjT6OoOklinQ0TPj87LpiWhX9mcYDiCu8sAS5UZzL8xaG1dcG7pef0kz
2BJdOPmwuPVnhgru4IpCHv7Z1KGYY+n7D/7a5HaZnBBSqOhap3cyogjVFURl7JcE6bD8mbRc6ak6
un2x1+e0YnTMABYeOicsJSrlZJySe491akRrDGIw4fuNQ5AET2MccwjagqyeiJSU06xZ7u2denKz
fV8D0rJl1jm06JwO5E4X7kKy3y61p+KbNfVqElhiO1/yuq2x9WFVX3hcMzrzGlyiMZ4LBI1e3tVG
B/xZkZ/cb9gr1ynIDOUggNNxYvQnvC1DmPBJJrMcdGtILaSDb1/jR7fbOI2h2hbbfg/SnqQXtBvJ
QuWuGmPY2QHrwKy59SPM6b4tXmip0cleSfyQ0MQr/vGh/YtsL54psXPlujqZMtX6qc3RoJPA3c7n
vspfE5GFqE1nRMXDkcxDG9NlTgVNiNsCrInMlZmn8rLlkUtwQME/yQNTTGUjKWbN7nHWa9253HaB
45DMwAJAB81RcENeJ3OjeOjrkOWdi9MXzRk6bpzd/OX/eDJjtKo2/L4eeGKRtw9wDU/lpVkE6V0U
iymDTNMWCt183huQMiwkSe1n34F3JYXAonwJaQmdyp2hwU2T49R/wrwXqGfKzgQ+7u3mgeDyajVi
BnvUrTLHuYFii1CMd6wrSqFml/mLw7DOa6HjZ63SF5g2PZ5cTCGx2Ln3jh9Jbh/tq4cM0XvGer2Q
W/UJ7Ve3Ct8ThU1yOp9dvq2xxnB7fV8ulzkbOqIYHlffWt/9T1mJGSDnpn8ijKjmQ+QlRke64zR2
9mFsiv5eBVtAcxqijFNsVpufFQyycIIFB1DYKLOiJ+r6JfqvC1yz9LiTGWr+uzaafrrWRRT8MwIS
snTkDvfTTpoS+QCAzH8hu1/JZ3yff6iM/We0138Ql6LqInIDUEpMzxLl1L9zhQXW7vmZxXbStDIw
uwZdfPIrvMgijOc/Tysf+nW/E0QPqz3Vk0fDJy+8csDIGcEj05G+L+QB1r0KEMNwB7ckKoVwNR75
SbRFt1QwQE+DAdLLxsC129KVv2COfJPr9TtFcqjBMPvpWj07Hsn9RkHzEmkRIO1rkIkhtWHcD8/y
poxjXZoRuWJGXjkIHE7xxRke6UZsBNIVx7yV8VjCqgDEsA1S3fixl6Bs7ZiogGQ/XMv/yZ7CPnBB
Cgb7BlvFXkiplL/j2M4GVvjvevmJGQpqoBRU9BwxOIqAfp8wKcdKHtup3X1jfpIBFsVcc7hISwc8
t4TlGnGugf28WxqlrNj50CdbXCTAnOrYOCROHv4LP474OQlbJZlUo07VTGTfR3+fHcx/DsU/92hS
YRZFLucbMVvVnQUkfMA3AE1R18tPbHolT72hLS7gDorFcDBWYHRFf287rM2222+XGu7vOrcAMulz
CFkq+b7lH+RxJHD8rovekXy4fH9vunXnhktn+oCbrjoZbVJQaRaE8pjx51WPYVM9vnPw0GKmtyq6
EAxVOHhd5Bl8XaedJN2h8JXnp9dNiEaQ9AfBO/vt6snS7XUVloGDUIP2hbmDUB16Kv2arXitwNQz
PFxH81QOHggBuNs9tx/J4Lb7YEpBP1+9kswwRsGdEf9Sm0Jw8PQ9TFS0wYf850DusqBitoHZmrDt
rJMj2miGI6amhhWoC4ksYL8tCORx0bLUG+5z2imPtJV9F/Q/rLeBjXPiJTZlk3nhk+Lpj3CKFZEM
mdnDLeE8ppCAWqOc0C1SzYRLAJ84EMBktCKIb2MwCQGZFSZHsCqgzPBHZkh9mZxRYaZFv4KtvzrB
qX0WZPAKrpvL1pw5UTbbLzNJmFyytEDb5cnvx1+C0aPC13DkYuPOs2ghHxAzx0o9AirNTG5jVWCH
OiarKJN3snTsIMHd13yLiWHBejh/85aE4uw7BtldAPexlOZp+nGwba/dN3/QMhODW6FyVpoxUZBG
Zb7erBqRqCePQxJ4znNU4mTfbu0Tv5oIHCnayABNFVXHJhcS5KW+abIFH9BaGmOTgkfH+rSbp19N
uj55a0ZyOL4KL/VYUPKj9i4ZmZIX5vHx9ArzzEZFJ8KRAT2oT2d0DLrwVR/6NVbbdYShxGgNltRd
J8cBZfMjxF44/33idQRRV2jq37Qhws6l0PD77WKah3O2UGVeLF8YhDfWICh70J9cNYQ7DwP3kWe+
mFE3ujAgIQWkZzYY0yUiSu6NP13e8Tk+j/U8Xer36X94TQe1npHMnetaXRWl+hHOnDIHk/5f+69t
4WOkP3qGgO6gxdu01X5M4W2JuWD2AN/Nm4HS6IdyMvN7riAljr6lfznljyMUd/OKTiuPPUHPSBeg
Oe9hs5RNl+rRLaxJlEsSEPV9z9AemSrzn9BR2bOMzKHg1yeWzvqiXlrapsv/voujiv5C1S0u9625
rfeSs/saj6L6D1u/cJd+ANTf73BA5BjYlFhbekvjkIsg826LB1DnorNsU/10X0jDwcC6ldLJyiQ4
Oakn1GHCDrY/Wfcm+Wil1zf7J+L+4UIxU2It9FzeRsLG8KRcs7HGB/BUeehVAyyTzYnLDDgOABBI
fbO3LuBUYeArKI4Tt3U6Dc5h0FUU6wxOJ4CfNcUE+133wtCU+nllrY0JKsxq0b3c+vXsPLpQ3nux
Ew3NkOslIivceBrczIo54eYcs17na06Rg9AegATWzYLqqAWiNVGXTuHDpFZjfSQlcMjrWErFFYq5
Qh/x6ONNMzrXFO9nbf5lL3zhgngRcZAU1P6aG8CFcmea/OaP3U51wsBBAuYpncX8DMrPjq+zA1Gx
IvQGZmTL7n0meuOQrZ0iHzIXiGT4bwUKvxLnPurv44dD8nZWAo1Z0TqEHVCfAK7NmVhPQ1slhoq4
fjnM9IGYqDVvaWL2Aju3x4FmZe53qrbm6zHvh/1NVgYgtY+giGQdLkBjRU8jPSEDXorYHsM2cHDJ
5FKNEKdxc75zAZTUtIg0dH8xhsCmh+BpibKlCfw0gRoGoOsdFMT7a31hesyJGbmaZkQ3e24RnrqI
EAByV13lvtnuyXXVKDo5pKZIrxsirQ9xGKSoFtept3P21wrExM5vY+2I75ptFkvEZbFXvamuXPPT
VM1g/3ygvKakRS/jGsSRTyLE+RcUJqr/BCoUTw4rD2aeV7Fr2N/2HPFul4qtMBQrmtmj2tjOGj5p
Xzo+KldMX3+oR+BblU/AIWWvQ4fvoJhciNXzysynzcSgvU4XWeuV6bqW/RGO33y2HAtHymWnJq68
IQbrJPyceJn4DRsWLpPjjfH/T4sYXH5MehOLwRUwI1Ich8LbfAM41a9NSYBfGrlsNCMgQa7yUIiU
H3ndhrr5IePklZdklOZkElB4HzPCQ0fW4Uy9wTaW/0hz8K8P9vWhNLr9ahZdDbqm7Og8cS3aiROJ
6Ln30qWgDkeQ2fPej6FreIkD61p4Zowv4weyY541nrL5EgZIo0g2qwU6b9nznHa0QbUaiznz77LH
mq+O+yN0eec/WABzJze3PoVeBBeFBmP2kgrdct2jxsk4GPzRzGs5SIyxTV8o7zsspX6t0ZZPIBGS
tpAOhD4WMHLW0OHghJJyykGOyVcXgwStjCRN0sc99pmif8WEDZDx7lq36tKTy+HVN397pReZtTgi
i+TkaaP6b0HH4bJNKKcedrMUn58HqbBHtn3/rRsjqV3eX/920tj4qzaIGvO1zTax/4+Egq2DaWln
H6AKO3Pw+l5L4VV6NMhLgj1plvodn28OpzPrFGc+IpJX+dEQdlf0rm9imuYziLKMe8JJdgw4QXO3
hG0bvwThBjPaOWh4EBMy4eunZtUn83xwG0MjgFKisCK4Zdk73xX/vHqMklbbCBuTQsX7f/q7Q4pF
SwM+Jj0icEVog/Q/+0bJ3x2W58Z7GnmQHCctEQn0F87QkrILQG1aIzYFWVyFQ7BinlJnCkGmcg40
Hjkp6qDGqfInWKhVFbE6G5xTg8PceLDSc+doQFCU2pQXirNQKAtXgo7THm8D8eh4kcama1SlvjDF
LX7PaQ6orJJbSIktfHJOMrZ7Po7gtvqjLbNS24NfrqYeb8ufeJ9fGCd1Y56iV71mubKrJ5UYbzsb
Pk/MJ45eVMFG37woPwsyRxsN/9mc3qgcnn93Ylg+EcV3klKg227qW4VX5DC1lXLatBFj87aOT5Ux
hs5RxaMFZT1LDXCncfr7g0KsbzQs9Dz5gbItFScYpsG0HG16gkAp+btSqKrXDuCHF02JQMsjc58l
e3lRL4+68B6xXAldJxZJ9FT0J99XjTKZeZuMdjKdvIA0o8zqpRS0rJfAmWZoZ1AIGqFVRlCQeL/l
KuhCKGMdSlM/SVhHRKnrFoFJFBmviEolY08v13Aqb/50JkoOgBLhycNSLk/LSaBUtokZGbiG8Hdz
7QPFmuip5enzjHXUoNs+qFQCTh/lo7H2unZL9DVBSBXD+RZhU643lnHz5PERoYaeuFXNClEOEVc7
bEiPRv6OmryRX45JCiNoMmn5mBvvnczYuvpF5snSDWOigJ0CD4u62QoFqN5BwH4vp/Q1kv/0xpyV
PNJeiGITCmCEDHlj6+nr/WkJTzIutUkX8Z/IKH7lGp6S0oArUzGVlLldIlVIhYGLvIJMOReaXzQ4
s1d42pVOL9VE8HcX7yCw8o/YG6KEVoh2DzF5X5vogeJl2hcSZTtGsAZtNE39QfZFWc3NwMyH9QAC
+D0QxSXBEyG9K3BSo+hFi8uqzAp6RC88qOOpzFEnit9IkD6Dl4JoVQJtVXodScwDS0JuDFhY2qMx
pYqA9qHd+JZCndPSYRLFCIxbOZT2trP1nC8EPVYxNFZr/z/EnhJrtikqnqH88oHZwz8+yJesS+tI
Py2PXeADSqoqzKbh6NnP6E76hCau20yMWPLVuwqN65iMhu54iBqConHXFXyclJzQ/96aMIoctaNv
IOYPbGZdVbOTXuES6IyUyCxRgg8xCZCuJhvCijoNl1Vm+tTZjtPaiQLLvsAUz/bxDUhWaAWEKEZA
9Wn8qGbG/LPPmZ5ut2hDv38Kos7QYAqkBAn/NmxELyO6uOceDv0hWbRfXZD6fKkoTmLvdKvEAauO
MTLkCnxLlbpCxND+lcTbAxHO2s1SropIclev4F3vJuT0aVyLrQGzf/ZCfmfyvPFIRG3SO3unmI0O
WtKVoU/M57PhxSw5/fbSxK48zerHJv8JleWyeghh/EmgFs9SqAKwi80Qy0NbSfX03JmnQ60EJiDE
UVotQ1vwHKQGMlbDkcSLUv/rDLyg3A5pZGdsV0LqL5yC9XX1Rsq2X6WjxxspJXuqbTpCkLmieZHI
KqhekLJZtZEyNikQy1sjatcHQA7issuhVB5TaqX4yMHE7XBUNM6GMDJ5IetN9aRi3GvGiDTGZpJR
1wxJevSTviosjZV76uyV4KS3A6pC4u6hFo8OQRW80dB9B8BBQlg4k9sc7t+ix7nC8gBc4q6wRT83
PpdpclxwhAfAAGXRW98v5ktAqxhjICmQBRpMzlymwbgj69PmiaZKClpjDT7DnkXvVP9ikhNgeV9D
cdhEt/vZknlHZb9uvJEdeQ3nLeUFvv4OfwTlsjD4R/pRb/78A3fEcrv1p6qsYgd4KcGcT8CFL/YI
ALl6k3in+qnvEEf/8NF/nrhPN5cWhuhRY0zuBRhehxQJezCVOtoX0AcjJwe69uKGBUtMyievMAju
/GA50wRyiLX39pANiPO3BjA+/nidg2jq9SBxXIXHWyk0ZbMPCtCXZAvafDeEXDoRY6t4vEbIGR6C
ZMgPwe+5HzY9FHGOyQ7uMkeHzTaS3WFZFEICUtba0WsPcYuylwZ4ZxecDZTfxUDXLbh3xX16OpZm
iEm+CN7r0Okgops140tHl8di1F3o6ddxODApShrPHPPwYFjxGOF+AgrLz75fLBCCmkhvrkQWWyGA
OSQZQZIlut95acEPn+bV6SKOCfg5mCQsa2j0rhVr3h/AQulv/hu1qQCUNSeqTIm8qlb9O6jW0FEh
+k5itsx1aDV/uIeZEPFG86lKFC4H1KfpCyCVapx4eqzGtWlOiQ9GbqLDI7gm90quVXuyPnlTXXD4
Y07EAHztLiEsHMmqiIjb1qsCjsOVHO2pPOKNHYtgqNdsTSFeUPFbykGRTAqZ1VOpmS5X/iuY9TgI
MhKcxGqFW8kCgNYWjUW+c9vUxb5e3LQsbHRmVHnvXoQLsT4DDZU2D6sdesvbUGSUghVNd4oqlh5H
NSVviF16JDxo9uMGlobJ2byhRjE5UXfZvJyZ8B9B+iqqL5uFzhcLjrs2YoDYQe0yLg88KunIF1uk
fS4tprzBUlGKt6PG1J91qfM+40Fj49d0MwQlfhCFKaIIzBaw7BPN1JzdsuYFJSqAGwwctBJF4krx
0dqBjwa3HqJPUCZvctyeyIvD1maQ2BkgYHiR4qjJ8imhjYS6s8iMpqMo4Ym3Y+6QMWST3hUl3O2g
pe24A1DEpW+Pynm5qHaHOA3Lys9jEZk3JLeTxqv0nnnCcvfGM+gzMkaPt2jfihbnMpn6WQps4PlN
+zGE9p0Y3GmVbVyX4dmOcQbycjvNWfMHgJ/FBr8RcQzdC/2bGLUS+9+QeD/lOWJFP4GoDJoD70Lw
cBQH1k3ePSvvl/MqJS3GAYjIAXQvZyvJKm0Q4/thfmtBzKJDOy3d7wq1nQGJSNg+mdlDzYYRN0OK
p3xHrAbkkemoWo9W1J4govRDhLGskGojTAWSmWhMJoGu7NWLtpBdLgpfa0ejYoM100538v1N4pii
7pb8+DUUmuHOM0JC2qQy9hTmTX/NVKbXRuS5bsPv5wfy8sGckPxR3C8xY/PoGMu5bos1IGfU3AjW
x3w3naHMRtjg+jYy0QpRyIcefZmeghhMTISN7B39M9iMjOm4GUuJ/VzuwWR2yrtoCAblk2cncjT1
YbjyL0Z8KTFAS6eqs2WoxHi3RT9PmuQ+GSYmP0fRAzwUITe00i8D4U+Ir4hIU8D5h+SxL2m7b1Az
ZLTW2aRzm3SNbCmNgCFN4mPzSNYfOwSMpS7LxGC2mY41ZEadZWnEYp7OXVyIOOJdfu5G8RQeVfiQ
hVsikDFIqwCxbuvTKOFXuiMB+6CTrzpz+EgY87V0q9gzEeKRfIXAxzoOgwNB7hzY+HNDMeyMgVG6
bIAIWN11bXvfTjj9HEsxHJNcp/4Gfv1mNkJPHTcCZGOvhdVuq16lobCuRHUbXAhhUtTOJ8oNYtVa
HBYW+qIdJQJaLO9Q8vej0vxV2H648G6BTneV7qpoVWBxLXYB179W6sI0wfuFmrUyIPovQmwOcKEn
54RLVtOyDViMe5/xfZNlLg+TDMAdon+deRCg/sOfZ6VpGR3CpmrBZAR9n05HCsC/BjBNpA6YKr65
JvZNsdGX+EU1CjL9Gz21PNK9mzvCucaJZgKT399u9DkFZEFk771CgPOw1WDJEoPvtZeeodl3z885
nVVsdPlegy7lc7rBVwvcK6r0i74I41BlEGkSMXO2Z55b/tmMJwOucKurgHuhqghnJe+wK5wLaerH
2yDA1VqgvtwNtM3zK57PSyV55C9MBXWBYODsrPt5gzPNXhW49cPYuJMx96XbKPgqHovhkIcdAEeO
KAo6QMVsQfrAp9walqNh69eA39WjriqiUniYRyvyX/H1HLmk/q7gnVACWQMQvp/S2tsiTZdnM6dk
w8ff7SCrMkEaMLxDl1qsgQeXINRW+0ybIEPb8zyqyksoF0iat4Adbs/3BFqaSPHaT+4wQ5MpB9lR
1KDI3ooietRTuNIyku0LOWhdEMLXpjUaOfSRW6RMO1RAEwUZ5ECIelP+IwYHF3S5dz8ZoWPy2g+n
9og94hz60+RQh2h5Kzkg04NG3DN41wqaLejrYehIitsliCCMuwmMuAaNIr7DH3mVQ/WhJpwH5jM7
jT+NpuLdtKFD6xNpdB2a1fBr0XChLEg2Pmd8Jyolq/NHICIFnWFTl0jXP/hxDUjy8KQhYc0wFM4P
Y1RDxUHn5n0fVCT5QnZ4aDEYjAtLBvYWlYJvNdAbMgOVNIUWN3o+QwZAtUs4qE3Nhs/m0uZQfp6X
f0CV/fdpo0GS6iIAYEmwzGppNLTSbUOeFdgjX4iT/JK0jg3gE630QrT+vo8p68fOU7qtal8c9GZ8
ZXZJHPwGHu1P+94n3R1ph5MwNWNoKfcb1vl/AXjp4ya/54AzzzZ8e+/irGGxEDih8Ojn2MDPD2Yw
WlUK4jVqhKrn7GFZZFjgrGls72vwJpv8+07f5k1/vraQMNWQ3u8Whv9RF4FTHow4kf7f84vqbVpk
R1zERk+xgypLtPJlh7AITCsZErlyC53Dj1qqePDGSQ1Mi8RVQjx1ThjLRzMEHabgQvnKB7gKxh8k
rUZ+I+dWsi4GaVUJYqMDsAXpSSg1Nhzt2JLiPUfSop+ucz9wpsNodKMg1gUjayBqIUINheTCPe6M
AAhVIPninsziiNQwlxw81H6nc8qD+wBB1nAgz5P29EyheU0IJhKN1s4Ro1ybcATzOp2f2+AGpM9E
pHlV6IEAaN0LCvTgb61UyAa4zneWKaPi8mDoeQYZClrGHWbDqs4Jc1JP5omuXqnpi9YNpzxXF9n8
5sw/zABKmgWlv1yZp+zzq6F913zwlyONGJogaUl5i16Nm2kHsb24WSBM5DlS3d/TBeu7rCOsNcU+
n5FFaXPjb9q1B+UlDQsPdq8lu2UN4W6BYe2UF+BviESrC13AgPCDdzKDApu97DeevAg0ly3tx8yK
7aVO347V+j3+O+q2cDcs5kQspzCp/KYRhdduvc3wpV9WSSTYOOxTaKNAHCzpcgn4K0uzBcESJufW
i1Dxhe525AI75rAn8bGWFwzheXj/mkRAl5I6VF3aZ+ScaeU4ud0Ydj2RPfujTs3WqSwq7V7jYfY7
1G+dNh8QVfvIhs49cXTsvs0yLzvp+uwP1WRkZ78FEnM35EoqAPnU4Y/Iw2c9tL6TPB9at7rproBU
1zw7589fcR/LSl7GdVFd9Ok3jqUVDAtPxOgptGER8oRkwlZDJqlpYVRGZ5Ibm7SmaJTmjl//2DLP
ReG1iG7ENGW7ITcicXYcAPYnwG00INs7ymCdjai049Q9jsLmw6rAjjAp6ayE61xHCUmJHr5vIUGq
h1mMLyqyJJZL3upCJMWM9M78ZudQ1t+SLWyKBtYsj/f39qy0jcKFjc+yPDgJHVfINuNTcwZ9QN/i
3q4ZX0gS1srukjaLBSln2CQXqqpRsFewnjZD1lE94McISyf6h0xi8BY2X6lAD3IWxe0yIIPyoPmK
mA0gmBEsNt05Dqj80NOzTpD8NDWnQSqf8BTY0Lkx1dKT5w2AVwdShebpLwLw6aQ8fQe+nI0p3T+P
3e4xY96b/wh3vdGOxiJkUtxwk9hrUFBxMVV/oLR3JB1Zl2CV0kXb8zkJ/uTV/X2/Iqxi5V8BXgB5
f17Qm8V1OVMfryvqw0B1gDFdei3T5aiVKGOczJD8/waXc30GcclrL+OnHRtkelCy5iJWeI8XOwrl
DUH6S9uWAZMp0EpSvzHIIQrFwzUcAxCpM1lRKATi5Fh/u5bQpCXiVcWd0sMLbfdPFLSUBFdq3XFn
oq4VN3ddwSqBv9ViDSANx1hyBAqkyZ4kGDH4A0YUFA2N1q3A7wK7t8j3+twj8o/mHXQPdwUjeIn3
vKUuSxbIb2vonZmvjuAUt3jdx4lXk0RWQp3IIw3Q/u9lEnazXN0cdiBJCqGZK2qxXjJRljt6eoeX
n5KMEw0XVcIUV3uVnXc7vHuvNVI2Sz/jYkKo2RQWITnfhKm8LLaXzpbCY48EbHTm512xfsvoZSR4
nAxozQPxD3rWIQwtCtwfXilgklE4/HuQYmeUlrXOO3hvxor89d8Q1tTqWF5H2XNHB4dzhkWMn2fv
7eDwFFP+dpJwqzZnEoQp3Byz0NF/qzoEfSd2lvUiGRACobdIpGOobJ5KXFq8uh4V/RzSz213faAN
EIrPItSM/76hHapR7sKo0jKqlhrXLnKnRMFBlDNc7nc5oNSudM8WYmHg2U0y1oYUFyGdPwIdcGrP
lquRSpPXSYngb7CEdUw/X+GBBeypT4rkH1ReF8Dik8LPL2D/GRgUme1hLpMxI8ygLeTys6X/xUET
9Ry5CmkwVlVmr6g14uCYBelekduLQc7aZecB1Y3fNEsZXbltEjh1ivqQK6l3UKIlu449tkoahvq9
Jh2N70qJbws7uoM5zdpAil6ayMFDdUTo73uEaDrmmD0+S1gOP2M87FFvT6YfYpiBqQPIhGrNtWFD
dai1lLmoi9QrR7rpFpr2cqFBKMeFfxg26j9FdXDiBvKyVeMLitVxlta/zYkZ7Gkjj+5MbMYnl1ch
nnKTT4F5bdZzKvaIL+wPDUrHTkWOxg4i8wIjMQMWajVPacVeKttshazFbaA9iT8qUDL6sWkIlTor
dhLvHJ1hjsTlldO0xoTR5eYtZx3iwf+kzIAUg2iqsF6oJAf3dx03/Sh+h2tSBe4WMhNgfvY0KsEs
BC/S5TchPzVAk2+o/hw561x3f7LVJfWY1XErTp0DiWyycqFJb2t+bvpR4qs/6+muJpxw8LlF+oA+
FkQbO7wb4ca3AV1xxvfoFOJy2Osi/S/Vzm5vXkSH2n4m9zW1b/0S9uLQvxZP+xGVDEF495gp0XzT
s2cFe30DuKg3lR2gDUEdql8p5DFeA2pUl//iUlpNWMtGbvNpuPvEPSOXrB5cRPSo+S6f7bYihnlx
IbJEiHC9mmQ9A+fHzveqHr0dZYmXhPHO0KmjwrpVK4OVifAImt3PJ9XxQBX0ZhmaVsUGAXQzsuNS
GNzug2ny4hpkuWB2DFiGmgX+PQcZ4VzulKj+8OD2C0xwthF8kUNwUGvWAMCCKnZRTnlYKE7rVnOr
oO7YjAFSYwM4ibBATwxjO/imfRubGuJziCWGlLUiU34tRqZpZWm9PtlVlCr/r3I++UXbh18hd30p
XdvG2w6GN9luzrFiFRe6wRrtijFheMU5D4adhipMY3CCAKEqorJbsr4UmqQbHta5vOIF2bXZ5H0y
IdJrkDVkWu0Qnbx6gHPLEX9UH9hiLV9GbHd3X61hlnm5H1QmSXqS4N+f5b3vWfaKU4ROPAxNQyAX
YfK3/tVVOW9DVjonJbjkqLb7PEviF4Jn46xQ+N6y/EEVtHBu5IdIXRxXeqDTGrUij8SA4g6+ffjh
iCXastIsGofGbzQT4UpMacp20RmwrdEvOc6rQoZLvykOPfXcTguFzOyK9jgT3qpB5I6lqCGoJQD6
GoJtnQ6j6Fqmr38NFiOf+jfwN56GzojrQfMbiOOFZaEpixwdbJ/X8o8PvOdpjE5ntnj8eXADjAwj
ZgPDPGpXRfEonyEDNHBDoFr+m/48IzkouI1g1bymAReILHpkBFL88TQW8kTPN0xBAqsRIvuYzL31
bElIvaSkd3HOPraFozA2XIkioLqi+VlF+2wdGREAmCApAO0e7eLr5smp7nUJZNNbuKDjuGCdgfW5
B1c7DNmyArxCFQ+OgSCbbYvMHcXaR75ukAz/T0sqGIccErYod4kNfscckI8L4tD3VEpcz7eF7YFS
yxifzW79a9rUmVet32hD9u6EnhUp7KnBY41J5TbZstdEUVngjSFJxQ8pCTsc4Ct2UQgOj57VWzHR
sm1pmHxh7EYHJEU11rMGZDRPhlo5Zj8bt5xTm3o5tzg9sg7gagtFUzbIoyYllm50DjTOVYEZQkiK
oGhgCHg5SLMI3lvzbklfQvidyWzARcUqRbxQQ7G2rfqEt+1/Sc1uXFmDNg/18X+qp9tpAsnwO9FB
0M3G8/eD1tavvV+UWMOY0WMzYrhgt7LIYD55+9S8FZByISWpnu5QdUISVq/JD3mFGcJpO5xXs+iv
ylvPLA62sIpFqRVDEGTHXnO5/1G+HpMHKNCUvnEuZi/WERHgFb+CMEWeJoQZ3FD97TuRJlbwk1CI
bh8CMuwr99OzB9JO0QFay/Pi6mz5mKN7jvHY9oHmYeuO5eIDr0eSlycjkswHN9VXL2AAVUUmoDeX
q7TsLTLONSfYoqpQUFT00JjMrg+Ht3mgWP1ta7FUFLOIV1Wu+aDvVEDCV6HBIoVwbT4uyUV2YaIi
/HwC6/7c5CO3iGAtNoF2RdFwmLNSe30GSSrL7eHGdMPLi5z3Vul+IwPvsFTZDK51bD3jzSkF/kt8
j0/z+UnXsDvbIBdMghoQ372EtbEIBDfsMI/uCgBohIolptvNlqz+p8SzmcLNCCy9/s8RRON1+e+5
ts2jI74R6KAEE0UJNsWYvmWnVl7zPO2edJkn77A0gBDXz8eBtf053pe6rOPvT55A6DbaEMVxOi/I
k8lgvTwtAC8O+c6CdJ31sG3wgCxQXXK4TCSKXHBvDIMg2x0JB8f4eZLZaHCXYmx8GiniUe+rkW95
YlRvjF/7RYnBx1vqr+lVfInGb2ntwCqZ9eCs+vyBdXePwzi7G0Eh8T8B1ornj5FCgR0HoPKwP5/4
wdovxff5xwALfbQz2U02cNlj5l4FReveLlw1wly7g2zndXER6/5MvVmZ5thPGO0ogdEQVvWdV39c
UrSOngeoBOweg+HdTDw2xcsVU4fdHUcqGeH7IfKkABHHFrrIpxlRHUHLWO1tqImAEEKy+Mi32m9x
mAp2e/O+u11ZPyNgVFXw7kTDr9KW74vzlxXy4KOQ2jNC0lL8v+oDpFD8gzhKM67ka0xih99w8b61
iuo18wa9PGYWwGtjvWzvF6Ik2QZck9ybity0EYmnmXvJuZdRyhaluOjjdXxK7MhxWJ/lg36k+apz
+qdstSOEd6sVRfxJjc7weiPLKIzYFxZ4pHAestByjbtkL6fRgEi7mCj6oT8UBJQdv11lHYziVbei
PctTeby2otu1ExHLzQEpc8aul4cZ2AIIir65qlBpVw5zP8im8D3gMIVLRs9D9AfBSt9okjdgnLpb
kdKDzq9h+6/EZa7XVK8Z8wNXn8MnPUOGcUEhOPglI6q8SbuVPhS5yLteK1uv0ChM2MrXK/u2AXH9
lNJdS+EguVh5ZNY59n5aryiQWBUlrZiej8fIagHfcr+JGtlILge0s1Z547Jn8+JAUL31fFmuWSj8
VCwy/3Q/C2ZQkWRwwX0m0Ca3vsI0MCzHzeAl3PavA0EsjOIuXZG3FSGjkXbd9HdQpfadX9w+EZfx
2It1Jc13mez7Df96z0lPS6xhWKIVzSyCWRc1KGKNyjjGUA7oyT2tmxo9esUwrg4JpVyNg/VMSJMA
a8RMjq8bwgg+iUE81zzk5t15sg6cuVFJjHyx1L9uzkha4sUztI3NdkWLDYpkuqx1RIG5hNTlaTcI
atPrtkMzxXL92DEx2h3h8eLDRGzlRHIuJ4jyXMLrRRFt2OmLSwC5pXuIyRyyhVpTaFdDjQlSUQsJ
WzjwN6PMOun0r5had1wcJFhid15oANJjD/Frl2ufBvfRTNwDkXUrlteYSjSKpcrGkHItajo5fXYY
IcMNGZyJ0j+r3ulEIn/K9klbWJvWg+hpH0AUBtg5hxaHXKk/ENCezqPSNlMrxhFM3GyBNkMExmGO
bjBW++uobfO+vHytDCrVrRWpWBk751eNjpQpYijXrwrOw/7TMKlaMAZaHlLRBHgpwXkjhKM8ufKS
2hvh35/E+rumq2VBwcuyWtZO7WV8iIetromfllYyk7gOqk238+WMgv3UZKdk2SBZKlfuCPDYe54f
1khyfts/86Tt4ekUg7RizaucKU9r9OgmqdI6Ted0LaqMMNyCaQ1y/gUU4uxQlNN697nC5uD5d+yb
D9QS25oXfb0P8oQO/o8GlQR6HWdgClfq31F1Cytmvv2XBeapbWjdk99TeL9ww8+/gBnqOTBaBDZ+
s+6mRLBejF1SUUJ5jOK6pNNgB7eIelAZHTgRQ3X47Q8l/dQJ2RFg7YLQva0BiqTATxItCfmPJKmi
7K02cO8e7xZVUNeBMPdWkFEFYmmklMvDGu+Tf3faMhSJF22FxmgyXpAm6IoQb/UCd8mYQ/Z04vOv
36/FuRjqWATAdHvaHFUL49emOSaQ8IjEBWIyk+XQnxCd0JiemPaFwDhvUvQ0L/hKl/pkvXzHBnKz
kwUEayRSDps8BgsZEkrctw/kHlRYUU28Api6SbRCRnMERoN0aQgdSg/QXfSpG3PHb8MhdT7peNft
m8AM3co9IDrCEdXetg5AAHF8+jMS0ELvH8utc1nzSZz+kYGhSixYCvmV721yHje8JcDYYJ5ynCTp
GIuN7G3ZEXTmoKg2bCAysVX6yAFvSkL0alyE6h1lKxdL8ZvAfzD/W6e+TVYWzvJ8D8s4WOntsBxd
s5z7sCueAJkutefFEvzHV+sOX3IogD189ZlQN3O+ioj7BbgvisbQUS+s2bws4zuKelFZur7f2Akv
iSpsu1R6P/LG1N0JmJidSD5UlVdNfxweJLQXB1P6Of/ILdwBDb3Xki2Oro6ifQ9CbuCYKrhR7ViP
fzRt9d2usi3wePN1nnafvk1/oDYsUkpkAwHb+nCNN4kHV3q77zo3WS4taWXiDEZidl+m6xdp5WjI
YhEtGzxVmSaFv9Qdrm9CahiFseYTxne8OWEZZf9NFWjU4OYyHlba+IW+3uO44uFTiyMuqYfubhBw
n2oooT9Jq6Sb4Af288XdouRzv5fL8DTysFy7m78Y7jvIqtx6yzZFfJvEEGzKv/Ji/AJvcNxD27F2
PRsackFQTyc3Fmre0/2ROCAWYOD1pc3WjodMRuptqwvfE/0YsYKk6ZJXSHm25iY/2rxCKVVR95II
H2LfDZQoty57LDv4CFeeN7QjgpLy4prIX/356EjyywLGMmZXGasM4jlAduzWieFeUUSjxPXmuhwY
0RvBzZ3QfEy+QzgLEsoN0xFG94bB+MHaFt/ZCnjQ3vOX0YEtjmAFjxeFpqvP8usC8M5A1gideaLp
CiwOwG178Ei90FlphXcsDl9Di/SN3BNA36+LDoGAXrKDKUpg/r1x+yOh4Rl8q6cSPNEm5uYX6c6M
qIaB8uEmB41eO3pkonWNHNNyMKl8pAhYRTMd0ZoA9Qq+07BjkCDDQbI97PDHXvmd3cS0vWUWnepH
yJyxgJpaXBhsGXEjYcRchucUGTSjmjvYOTqoee8kn1FCa0CZVgcImcAWQA9UrzmuIFQIjLrrY4PG
8df2V3YilzYv2UwJcNZUYUgZSlLlS+zosJtNgVvpl8jAK/1XRqlrjdPRKAv/uLgHkfMvNsVEfFNl
eW4vg2wOMZDCpLvPM8Sq/Mk+AYqlpPEXVq6vReSM4RdJ2IG4/Zeft+ZyOlB5C8itHRRXCHcRGbZu
W4o+hNVnzJJYsi9d35X6x4RDc2RUtOH2Soutv5secQ3XUJsfc8Kjz/XWzjfZCQJuDbOJJMksOI+i
S9IZwy+i5d3+typluI4y8nnYjwkt73ytZCzDCvl0pjWsGsuNim0nW+wNV3+yAa7XlVyyf54jB1pA
Na38cuGl8CiuJE/VaEVoEWKa3+F2yRlC0ICv+8W1IiQ7ZMXDkxkVjlVa3lFsF6jFVOZgfam8TNt5
Juv11TIyvfWRPrmmwMxRDApSBAcjKr9Ab9fDqOs8Jce18eOq9pueNo/HxADcMomYJWE69z3YjZ6l
b5wC7n42/yHpHKh5w6GPtZUOSewwpxbAJwkil1x60kxqZqtdhu4HY0E0bO4ogJDkJcUSZMxWXtxQ
0J8pGYfcIo6W/3NZt780Ue0eWMqrnGoTVPo5VnS87omY/tJspjZykDLjiWlBlpfPlGXeHBDP5ly1
c5ib3y/U0ncYGje6zYiyalrJblnr1EkNSeRnIbYvkSreRp43Okl109A95XcmpY6UYvsQwMz3/9Sv
N4UsexmHDvY8YTQAVHOip8fhGNK/Gc37X2KePMsOMuSkoTd5PtKKXjBPfmREziV3snWtKUd+iorP
r8z8NS/EmulLUaYw4NehQoOgtpPPxZJxcNTQgUHD9yOvCiI7jRx2Bd1IKLevB3LVCM8vcPE4phHO
YFzsGUZmJlu++hKTkj2MnoKDTE0/mKZLzyBiAnsAECoA3PQE0pRI7mL4NPAmGY0qfutaVR9ZRHUp
6CQzvMY4J/DJjG933yczMcJbJt9uOT+jeDoctIh5Ns9Yy/++cnuzL4mcBTVRgdIBBaJB71E1NujN
Xkqy1OgEOkgqdHoEx1ss790R1wXUwsWbfpT3vMzAuXDCwrOK9vgU/1FLlNZl9lf5OSvmKlzT+0RW
hHqJvTUzYJn5OqjYWGDL5yOTTUcp7AOjTNzlCQD2MSQz/fnH+biFsYSRCnyozOTpy2g2zay99YxM
Qie5o29TLfLj5mKOevNO68eqTbhHPUhhWIFP2B8pUaugjlEvRVCU3aKqrmnhQ/LdbARKC7RRIthp
9aenrjwreY3TBegi/OLM473sdggQ3+B+weHYYBavM3QP9DOWQKehwg3F8nP6DvYDSIakt4/tiVrO
XVhxiEFk9lCIDwmEg1EcHgh9a6TFR15I5w61ZtUE15Do5dkUJ+FviWs+Xm57e2LosIMOFTROKfkX
R39t+WHrKmWDaeWt0/uqIlBxSTbH40RFxEAlj4q/s0N9uKZRkx+1J1WpmsOCnGcHhscY8wu11+uj
gGXag5X0gdtBAwEWh0AIyrbppfU47RJVBe7vgJCxEFKK6QlR9Je62+oL0ovK3Ej3Bsi3wmdmDB2Y
Oc/W3dK35zbJ6mHrMlMZjzQqAPSiUxUaKQJYupqjw4oEf5ASOR32aGY5hCs70YvCjI0Hq661VniR
xj+EQ0dVxofeJF+hG74xL8GCqpicpo2qhB2SGkaddt7Z6iKa4tMB0Zet6Jh24RQoQLNpl46NT9/r
sJkEuMmP4JJJopdOdQ3eraOe/Qq4fGJATT93Ze8iw7zjl+MwOSiHUdqay3Y7HGqBDlDM0UrmqvwV
I+2OZAKto6asVA2yjhCPnei9wNrakFlxCkDzfooIc6uEi8yhctJME5/Wq9GlUSa6Qpd3n+RBJMPR
bneqYR0taFq9XX4z3ZXA2BepC78a1vQ8O4yMbd/VlTxz6iPNgzjq7NXXSuDj7QIlFm7OUfPUDwvO
3PM0UbMzK6Bow+seOST8PrL6Xx/ZC2mJfx7hQZGAtBBDoXX8n9ys0YGmI2G+OSs7Vb749JrXSuHE
cVnoPsAD+XRBLsK/zmGXmEJuFxcTxDGWH6LrFb0tQpcTIBPly10icqDNY1NDLvht+nF1sO8sDMlo
+Ro/S9AGLGrn7t94unxC7UWo/fUeCtd4TCIFnovS5SxqSgjUXo3dZFyd7pMzavmgVL4a9Ov9FRGa
tXWHHu3i2nvguIxMBCWuM9aEcucM4TDJJ7cSE6mZtkdNo4AXqBVkcgxD+bZLJN694J7ge+MxmvCf
s3WRQuCMxTMR1txXVvbtL3XWllSBw8YXMCNzBcyIr//mp03ZvbxIbNmtH3WCxuIByiu0XjgjQJMV
/spXdQGbkZBV/gAlmywgGtWVp0Eu3Chy4dPR2YqeJMZuJppRk3PkgpmVPBZ2qCEVy6uttNS2o7HW
wiFBc0a0r2Z91S/yAe3c+DvgrX163uNg/xD0FQnp2fBj6jtsfjSgZj/rn6PbJXM3GSo0/xGiD4JQ
ZNPgnpCdUjjWHrGH4PLBgWaQbeXrYICrz6FrarHH/Hd2pTkpY1MfBMzxRgQjjI/C29imLwELLpPZ
3OO0uSfqWfTItWOwLNJnZ3hu+4PUC6quYzd+Sl84X8YBkAnT+3hAMP80HVSIHLT4SHI4fuLaYwh2
qQnLBtsnTLJwHeNZDn0zaqNztxvqXxCFTQV0pAi69z35j3615/02Pp9pfwQ0SyED90BXvHjJRzrp
1Zse9C1KcTqDY45UyBxnzpQeP5mHVHTm8JSHDY65pnn6UR0a3UvwXhaZ17vz86D9BTX+inux4ftA
FJvh9ksSBftbfRg527L8p4FmYviYz5OLjEzN3Z4ORTSEA2jhvUHRQSIjZDXG74QEdP7Qnivjtr1Q
NF573Y9nrGI20UMQumXaj08QIoO+uS7vrs9G3rk5VDrPu+jso3gPxE6LjBAd+nVOgnGfAoZvw+rl
6lVK4jLMNtThKUEjHbp0G2wg/6pdx+gP79KT3dvlqAK3tahGL8z1T08eTZyR3tgsb90XZFziq9Uj
uuyU5Uv7yYOqTdO+yDyx5XQLE4O9oh61TOIvJIWDA3S7JkdwjR8ZFqzWf7ovyJzjGAzD0qzijukP
mWowYkEydGaDQiGQOCu12HadcjMdhCFk2cNmX9eBV5ahDjMIz6QGCpmCGxREOotDKqB+Boa1ePVG
2MhesJHQWjJSgDWnEEuF6qDrnwiqBsCmlGGm8zjstnY8ot1EMM9cBZyenVUsa7Nwum2bkfbDhNWG
MsbDkjOgCLEcJdudiHaUFAFvtZRC3O+vPhXDtCguJSOblKprGCPEqFQVXqWoOerUPUGCjKbi6BM9
AiyWn8GzgZrFCmjHAHpHKfwYm/IFRRtYzHpe/xmdgYn6fdaZEIY0/DAW4ZhVcnCnz2iyU07VcNWy
sQ6C1Q8L/1lcTlYEDuP4LqiupADzKV2SZ5n70x5o+DtlubsuxRnNwjPUofXx8lnq3BWc7l4lk3Bc
QRdidVdl3/ulGLwgLNu5GzPsOxZI1B3rQjau8J7C79lfpEGRhBk9APGxNc3LwcprppqMxtNr1Sa3
vRyYoVhFVXW7vPv1FYlbBhXKePcfzhkxv0TfvMSu1W4TAfe4UfMoJThd9EzQlcKU11AaUlnqxumT
s0968VLV3/9lSjKRF/99eeBeoRDXRZjC/XZAPaJ56cln0FGYFVSGVbyT7Ai73/3ub2wYM6Jkza6L
hkDXLYFkjVhHjZ6CiPjuaF9IhDHBsggbffOGMOs6neUBegYC0SSfhKhfPTfNPeciARLiNgmBeU8h
B3Rz3wMAmgmVaaHKstMh7wdFPxPDX1IcnYfR06bs2+sSHlMIrXBFfcbecpcTjmhJEo4Z/YlSDeLt
zoexnNLmndNdMOGopYQqa+zYZ648kC5XN67ljXB4ObW9ff9QmRCdBW74HZxQ/HToPrdbBjLlL05q
QO+ZaXGnsU1gWEbGl8ytY3OzEhrJPeRIIzLoy0fs0LLUPVCpvYOFmv45mGe4p7JRWxYoopwLZXPl
076tI5ilU6OBZ9ddMduI12bb3ovQjtM9IklrOCLeb8eD2mWWsvFTz7RrfsJYKP54SCqSjXvfpj3A
wSewKiC3wgo23B+gBvNz6bktc9Q+C437nma2uWk++kZL0krprsuIybETjKEcLTdF8u8q3BxaUBOK
cBIVsf955drtBJA0L672ppbOD+tcbdHglfQpRZtqAGm2+L/tRbaOZ9zqPhYzKr8p12jyhPPzMSef
qhc0qr7g1tfZhwcYwGu9Xy7hfdNSCT3N/AzcG7GG8w48RSfO37P8VInGS3/YuRjkfHxnWkxgSheT
kFoHXQbapfikSnyRyt6PVpKjlBoQSmsI+EDHB5987f7rfxSGHNilEXOTXnMuGqmwMUyxa0rcmLLK
aoZOxxAiVzfJwzZLwU37tH/AMBaFI9o24Cd+Qo/R7HnAKYgA8RV89E/ow7X4UYENFFhgqjys1jac
2N9JmIQoTGecn9bHxDJr/LZIHS/nut1zV9uW+pSsNCGp0EsyoVGRqjBnaZ0+b6RDdm+yAsNB1RDU
0KIOlhhvVJw+nsfN+hknWS9sjjmsk3VKHO6XfyCVSWBnEcKIVjDlkO3R7lAEUS3S2SiRVjOCMu8j
kptKIHOYM683LUedeY2KnvNp2ISbmeEQ2sC6S+w7EsbpyPriZ8G30C3shA/uRus5F/jkm4mbg7jO
5mobMIYshAloM3Slmz6uCaEFIInpHFgTJ+/ZyWiHDleFIOMMDaV0frN0ggps13kC/SwAebcayreR
pmn7WIYoL5/gqDGBUoWbIz3UCV4imLZeHXghA+BLjYemPqoaF5jkEyuRqQP9pNTMd8KG0sOhW8Sq
kVA0CtzMXMzFDYTgxipv/gcbyMVWFRS/LsJBNLObjWNK+r0hSc7KGmkkhIwROReeC7jnVLen6z+Y
VGbcAgzUdA+78V3SkXzodRfXfm6o7KmfNc/ADBsIVDr46riEK5IUmwkQWR8mpxRGEsKtVnIQrIpB
K+oCk9AaxZFyqvFvclTVzi3RHLkjyzSvEI6kmZVNZblDc1P+SMvq4SCy4YxurD5+8sm8JYGXZF/X
IUQCFbfgC1xNxcr/Jox8JtZfrY+fHDx+fHzQIKn0BnCjaCe4KlnJo8YyL8ZRR6GUIKccqEs7C8yp
dNVggfkZSIO7SWliFJ/jcOfYzS4SZWrC3AzkMyQqfxDViTyn2vvw91Al+hMWo7HiF/IcSTBzJSuE
COw7HrwcdAwwA0mZFfgntYVUzBhau8ImEGWhXhzPmYoRhs1tW4kmwcqGGm+fzCV5JlTamkD4+7Iq
tIszjxF2zCRYXPwxuwBg5UEm+B968/599mj/9pzB3EkBBGMRPs01SC+5tfaG7SJIhIOsNGk3B2ER
+oS7r47K3lNOi9Xc7SClp+EimZwE52RUebqVP6MgHy++xC3YWh5WYYhgoejoFe2WH3MF4SObtNkQ
yaeMNGXQGmH6WfdDQxqtyrmLMr2lwX0aMV6QxiiPoirmWKgz+rP/ASj8MAgKEknApIVU090Zr7dc
YppxLV3g9aGtKJ/P4NEJbA5xUpEU18sv/cvfF5YCKJlJ6T01/S6WGb3pIMTBlwxw4tHhkRkGZXHl
MpqKWsoIUKal0vyfeGKK+uC9L2jySEUr8V1RT5EfYtEy0FAtFMo/5aNT31wW8pp0SqzJe4RUKpmB
zX09c2g9qRF/yqB57DIB6lQIDa4+H4gxvWmKGV4GViRwtjWw6pm/zQBgYV1EVr6Nz3yjSZpE9xl+
9l3pKvp8e5L3JuSwLdZdSWdd3QwbOOVsx+d8RAVDgWE7KwAQe1wlTWrOAHGglbBcZrL/ItZ3gGlz
3ky/Ki9ORjg+LjlPDfJ/7VauhlX/FCb1bjIWJN5UWFXRKuwYfKbwIeJjlZ5uxQ193IE9D2pQ6Gwo
ZQsZhHPcIe6g9E8CLq5/Seyi55/0Eykm98goYO+19wSvLhV4h/4vfHLS6PI8IsUm7g2WAy4Mglx3
rrUrxoTvP69B7qf75fYDouuhj1zFYn+l2MLN7iA2wBVH7rig+223bvSZZFyQ0eyNzt7pBAFHcEy9
dLz9JW2lbSuk2spX2kAcvNcppgsAnW6Ixz0Hu3oqTzr/WX7SS4RVeiroBAkn7KQtsjXDJr1hcgui
VaA2zX3L7SeEozY1CjPBW3kn6q9SC/fV49MTWu37LRvB1UB/1a4Ysey5sIdjHoMkRSHNIcOl0vbK
UqmW+0pF909k/9RPnpLW2S5r5glKa/LWD5CBzl4QG3pVhj4wrnBPC1DsMKc/ZVkUFk3N+B5wTCpU
t6SXmxlSrEGVmDExLQOBynGQXKakFkko4Kc07s3GyTMoHOrlMrtkMoBr68tnnwXiOkpQAvTDAp6x
tz7g3vTK+yR//MZ/1DJRhuh7waYg8GGziMCDLtyGN7FiqEbDYMEef/SS+dC/7NpmJ7zN21heAa9T
kUhk0SJH1ajavlzrogFaqfdkV9PLvPWIFImSl9EUjBvsEPT5Ju/aWwOoMTrUHN/Ou2Cl6WqrKQVI
B5LfU7Y/U3haMR558RCmJf3dWvncmoMP2CqnQb6CAd+4WLUZuUl97nKGn02AmzbCBndQnf7zO9RY
wRlC5mIHrtBZh6TvfyLZCDmJ+oqfsNaG/AE8LVmtJ6cZnB7yUxpV8LRWzbHgNyuvm+F55qqm/1hC
4oKabLo2wjlPygE6Q55jJBLtUde5TNgYvGtLdK/qK5OF2y+n2NrDbS4mPeMUIEMjKmE2jGJFnakM
sB5ju+v/3jx3V3zQrAZsddTVsfJHLnzbFU3dP3DGk095/vRfP7+KB8k5YBm40YE1jzeIKELGVgUp
T4wvQ+ajVpW+i2z2B61cDCHon7YufFuMVZTbMDGw0PEvMe00jJNZQnScwp2Ywomy1h7poAwidwWr
7m4cNKBt+Pfg7w/kseOLTXec27UgWnfjoN5XzAXkDHQCXvuc7JGku3GN8eFE7vlrTp7ufppiJbpi
XYX1PAMtWtVk4523Wy0UtPG5/evBcs9ZNYysaakINv0eB947DMo6tGguqC3TmsRgl3cCEfxi1bC/
I6y5WuH9DNeqXDjJFGTvtLykpN++NFWtpYTBA77hA1ymIIhVsuO+NhP4Bi1IOY7bNdXH70goa/hB
b4Lj4c3+i2Rmxy0zRYR/9DtiuopFkTnjkdvKJC5c+IoZIRPIKHIorcw6yKeupIGo6B+ktllOtPk1
2OC2CxioEsm3iNPZZDujQhisRyw4ZSYy2Zn22l1iRmCwFjk3hlKbiWqYcm2Tlb867JZpYmyxbeQ4
+eGE4sMvbEBLVdXr1u0mOFK2CwW+gm3QJQofmpCen0lauw/bYj3WNFW1o9a1HZPvslwShOn0UEPx
4+aQ0760LqKVltHEupZtMXPyDiCTSlxAAtqdXgRsRrw69Elpxjy3l6aB6DGyRaWZT8YSbeOpqFMk
F0vjMY675ZeGlO9sS2dSqLCzMMH/eLNvKXohZxiCJpiwKU4NR10AHo3WXy1XlujdvpoBwn8L3YCl
omtgZXfMqOIsdoXnGM5Aysxw6XzlphHuoIXLR59cownVtBc4A7JNTlJHYQB56RmsQWbGjCUje+NV
BxNFgzJRCZf9IxQm6Qmwzoae61hcx5ZIQldrKI8wOomJIpT1NQ7kFuBxc5jYGePXfFzgOxnkuRI2
G3CGy0gv/R0lcpAt7d4cb8TDuIQzVWbYmFlqXczqC8o2K+llekV05eQqiZRFZlY7+jEyNK0Pe0yn
MkR25T0jEfZfPlmYSnVQpx5UC3mSHQO9daP08lPcHFEMG5jhF9duyF/svCKge4DBcyWI0Zt9uRUI
jpyhIP83AsCCh6KJwDaYvlLwHufeiEiKHwin91hqheXaJE20IInmMGTAbovNTshKEVwK8pkzWc9L
r2VmK00AM1sZz2awxe8w1RITjoHnTZUe3S3eo53OX2307L1euAm8sWXz2+6wOu8zE3k0JbHGrkir
2cxy2NCQhb/N7cZ18TdyVOJuoYTvnA3S4pUulCuEEBKUMq72YcjFeoybBbujhauP/4Mlv65hpL3c
+tqwTJY2CT7DD8ZfNf4FknfX3ju2TXSD65uayZgDmdn2urKxxT/l7jtS7rfWphMmL6buo/hsv/Ee
yUP2oQ8w5bvWsHPn2vs0VYFdxaLprmINvlAawtYI7Iz/1XbNPt3aURylfBW9WtbQjJWzCGNwCjdd
8upfWutLOuB4/7AaRQv9+pfhZJaVSxXe/vnPBbLxIwjrPw8elc+PdI7L6Gws2KDL6V4OxTEzp5I+
/tx4LufDpJL+nX5yb3+aHHQdXfJPkc7Dwa+I9CRAA2N2fho7Qnp6kIhXCtFH74w49aNlnDXjwdq9
w1yGOYq78xD0M2lfOrJ8HGtkLr84UBNBOjyZfoCr9nIy+93GVvzAP0Jj8omhEhxCKih1niKWJvAi
34e9eMMTyCv6J4rSeePk0/ZM2lO1c7McS4wVrOipId/e5x67KqtmQ2iIi4yvOHWaHBSG+nklcBJB
7VfSCqyuwD5oslJrnxBWic4ZZnzETGrmpBGiGYje7C6XhQOvuuYef1MJSHa3aQ+Ol62vGBYaWIkE
nVeQJ4tCHKBb8JmogtCWlGNdyFqQAKy1AWulkFkicCawbpiaHW9xXVRO1paklkmLPVQtFBM5AA+9
tw1y9ykp3msIO3HWsFh08fK1WfVNZb1gzr/adAcvC8/peGazI9sVYskbU//2yVZlntEl0POG4mER
miBpkd1miuUP5Ucx55jnfqD5EoSlcHjbvD0mWljBU8N45MrkrNHP2zdl5j+hMLkyILJl7vH7tXAg
ZacOrCPXkPj0xG3qRQJZJfg/8NvI6y3kVU4OYp0QyAgSckkftpUT2H2w2sTMXvywMIllCRiizGQe
W9V9l2LamClEjP4L1LFOhdJR0zJjoGMM+lZwz6bS9D4JOuAeevbuALVowEjhG125ocAVfTkJzkUp
Pii3CsnIPFa/MisuvIP0JXObTubns2dBhjIjvBXd+XdiliHIxmkecUvdQpWSpC27v65f7y+odjVA
bDz3V4VvYIQWq1sRdxk7i7DnchojES3dGX9a79sggZ5aqekeEdw8RMF7Afa5Un+iSoDZK3/1mH74
7QxBz/Ohuz2K4Ki7fik4QmL8Y9kpvr2S8Dt27G/PI6rgn6YuHTxPv9jxKRzBOSFyieur2cqydWOU
LwkeHAmIyWUOpwhGsReLEAAJfQUCSjf4IVo64ivSeyY+MhFbtu1f+0lduL0Ses/CZV/5g1nbrsEG
eIeLW6VjisBRyHj66vUoQ+JBhFO/gv/rcMgYS8IEIIX/E1HLkZGxY5BPAsYmQd3M/yDj/S58mTbM
AWe2SB0RPNBfMukJpTs5jop/dfrxmDCaKkp59e9YVizVgUdPVVktj5DQUyu+J4N0cpYKdTdLWJ7Z
XRJhurJfCJdjlEaYso5fkQ5qWg7FVa1EON0NtinBkyUCB7qNtLYBa2fZ6t0e9KLB0AltXk0KdMFd
NB9htfxTw2IQ2KkLMuPdHUOwmNUaw0nmCj45Ne57aFhhkeFqvnLsQZSzCrxcpw07UjlDDxZuTWwQ
9EVYQr/dEVjUGNSwCcjN+xYoFeB0m24fXjXE7gJapw2mZ1w4bw58gWSn1oM/lvmwRss99AvTHHBP
N2PcBqN6MXoP+y5kyX7moxByh/EOiiGz6ZoN4K6jV9ZywbofbY7bgpid0Zy6V9QxnYHB84EiO5rM
xTODkyMxhcJA6CMKLkYmsY1ct4XSeXTm2qMamZZR8Yd/7Fdtl2EfdAvY25bickmM0RcOnu9heEJv
koS/3MXZlhtqf0Omqvz6G70Y7EmPFP7j9EE3bQK8L2O6YOzW6a06QEJ6awBZU2RHhlKvwit0gk0k
43Z61hlTvbwxp2JH+gKTGcfkRLGbLmcLZ+N+NCPtjaCAFEwYPcX/7uTpspP1heOUZ4tnkbcQpZWR
92xEaHsYakdBdkCCrBlN8bP5shmxjb7s3gbkHWEhxaXi3vUVHoYUPlMpBQHs00FYlFp8ggHsWH5q
vZ3bIDkmJJ8VeZaiL/1Mu9vgbEDLIA7NnFp6kUiDpUGH8Axx5fn/F0N/iET4V50y5qfEP0+LT7IF
0cC9EGGTZ6cFMd5w2uG+VbXTlWytOQ+fVvc82hoWRK0UQBquvg4xtM7IdeaKUam4QFFr4OVOEhln
7N+5AGESg2eR3VrhiZfSd5d5BrXG5ViD5K/BCmEMwHIqWKRAeWk7Y6OIMqAi2Rn/EatGHm0GU7/X
j+5FXVvYaj3ZBPJ2FYYqHJt7WlN96S2hkYBQekoyKWrlnF5V9vTLDMtmLyB3GyMXT2L1HUDyGlKl
eEroeKbqEuyKN5q0O4RYu2RkvUpMPdixVDeHMiGzuQ9cR2kasYDV6f+7UpU/VpOFwkJbqeG4lI4s
pdx9xhVm/TEox0Uz0EtJ6Kwedp3zxEwtoicZobe/XTJOLz/Zs0frI60eiVZaUUmpnUPBg9SsjlFe
VM6FL+UXeQ6JdzeJVFUjPPNYDDgTBB2lpMnA4l7ZJAB/4UdGC67FwAOcGBC7XPXXhPTkXnVvrgRX
WHh1CnH0rfQcmLH6fJHkroian7UbVN+HWHUQii8hQx8a7Nhnq3jKOcuImXcqK+PyYFqvP/a5reh0
2hf9++E7umwtYcnwHyiUg9adp8IOS7bTlSTmD+AEazCKOBw+BCeyWN1qKJH53QiAilssHMqcflDN
TF3bWHSLASQqF0jJEiiGQ4gGP1j6+mHOTg8RLR0CO38vtqLHyrujBFW59aU4Z1M5GiHRBzk3G0Rv
l97yArDN/oNsA6aOqnZmMXka/7MMoIMDSCnDjc4Xz/hfNo7h9V6dI0vQ42ehBYTGlg/vm0AEXtDf
R+GL5NZMsApw05LoTCE+PNYajnJx9nyVc51KzqGfPLRCV+ndBD/EOIcRF9FOXMjoyKak6Lw7ocKc
QXW0eLrtQlIovBI7jLFBSf4FjXcBTE25xFDJVVlDS3E4HP98Ciqpd+UcfxVE1xF20KyELlAigtCc
3j/YTQ+BUUKOlZZizoKffmyXEs8Ugg7mMGXGaNDWJAKDkbTIHH4mIrfxgEkdCleb3XSd9P+h3XU4
t7CRIvMeYXrqBt2AmbBM2pKkezVilMVjLrDR7rvJz8HIbk1wuHQc+lwDCNOtKTbFx4WN6XSeXMJI
4bWGTNtHMEl7injtLnR0klH9GXdYKfdCbXAWHkwgqXrl+d9/UoULHluS51YMBmlziVqOzYBTZa3J
ReIVnamR60PXKN9ut7kF3+Ke9smhGivXe37M6D5KAlkElWKhx2CRW5/ix/Q4yRsCo6N4PrRYjnt7
777TzfWKA8WMtGbxWwFGUhdsTIG/5BxukFJ/VYtv/R+fUYrigs0v1FzjfyEmQ0JB4POhQ+cNmvV1
DwJ0uxV4bjrybBYIwhNnSkjY7Iq9aOTqoPrRUcn6uRiSC/ahwk3GkrBwSS6fQ0dMWtXorkZX/QCJ
G18b0/UaNPDOFPztpGyGEvYimpjLW/Sd5OylqC+XUupDIryl7MTc8OxZnKTmOYt5s4QUDd9fPH7J
OLpZEmGp6pr1bbo/OoM3Q3RM+y4OzdmeyRX+mA4KUyvlHDVkwz7bDAb1YENtGmWBeFlAYeg/EJ7G
1pVH8Z9MnJzQnxtGKbOVLoCVkxZrS8TzfpvkGIs7kfGajXnQ9ObsmaZ+2KEZgEa8c9rTAK/B2XNx
6Zc25dPVmo0MbzvHHTvV8LWRFexPlLs/s/tvEXI7roBF5XN76dahOWWqa9KraphqmuavQQzGFqmH
1bSCJGrO47heEtWYr6PeROOKEEhugC5SbIufvAOCRKmO+UoH7GEklLvD2JJVHKEc+E0aFia/lHNN
FVb72X9uiBfVmsjFkp60tr9PKLRyrFDdpaQC5ClTqkJxiKviHDF2TKeeW/MTz1/Sw+VYenCIm8Yj
2JDGYjLu02wnItwGbxABKLQcz4M/AYwM4nBzXC5OxSoX4kXe1KQivOyuyvrrUjwkLMyUzONWWmIg
dXYBDwBNO8fmnPIKedAlxCeqRKzsW2GEFQhouuSxlmjnkZ7K646WjpQpYgAe/uEnP6h8yHnqL9xK
hZ94Als9rQfzM7NUTD+zc7Dclk5fczaft4+nbeZDVxNnbecBbf6j+8I9VvrpE0PBy0R5X1NZQvct
jwrmwmlkDc+TPrPcN0VCVDLr8aUqGvIr6By2ck8CS4OERPq7hLJdWyFKSpe1CoTEGLT6wUZ/a9qu
ClWs6ehFGQs2tJrmSY2J2qJBVr72q9+WvfEOJ/WTFpxNOWkCB6WQc1vtod/kqXYC0Zx24/P3TRZu
OQTeV5f+OO/zCgTuRuYdUD7viDiq39+u117xwtAF0eTuoz14WCXponpMuJIOBUx5w6Phr0vgtd0t
NsvLXGfBEK+BWkLQVGiCdg/o98h9UkAXtuB+pL6oT8oBn/NT16k5XCoEcAW+5oT2C4zSqfpeSfyc
tlUrSiF1+ksC/HeitXQESqN6G2tnS7/g/tUV8XXmxRkYiUN9ag7oSeBMJPEMyQfRwiQ/maIAgkjT
vrw7+1S7QJ9CRukSJ2MzJX/IleeAv2bYPnjtSLfs1RktC5YpCEADzODjzo5EcspF7VDxRGoI8d0y
45qXb7Qo3wfcV8b3mijUf6old0OqFrdxxlrKLaXUizcLHkU6SLZxMqMsL3wAlZG2QX91HwQIWOYM
d36ZWXCz4e19TfCl4/aTBJfLiqSNrVMbogZUVOdmVxoJMs69ooYplNVyFSVZTKPRsoYCEzBJ6Ji/
wO/0Yo6yzoDBfhjdr+Q6R2uHqna5uby2ooZWSu56aRlCAmYb0g2Ygj+bA0amytq9h56s0SNHRiSZ
5TU1acTZI4PTFsUQEJ+imdhaduvVZTVk9CggfWJpJAJ5Dfdf1SXlilOkUGKRSGbvuuQ9pKPp2qCd
L2R39kxqx27Ej0p5ZexkSK1KGC2/IXPbIWuwPKd+plodZCm+lH7+SgZzF92M/HdN5G5pYXh6FEKV
KtwWHLTukeNVf8etalgKqCZ0GA9g4CKvySEaXh1R2JgdM0objeMjMDVIW+ehEPJkuKBzr1RycIWx
ZGZ+Q931bTCJlxXWrZMfoLTZYnnWNvrijXJegZyiePCwV5HrBGIEoUOR5B+WkMzENEh5+UFqSLlQ
62WfiQq1ZFL2TREEsuEGzEvjOn2fjl0vi52bD28d6VczoeZxbSgyRqMXCME6qAi6mKnz2ofuOig0
K+r4uV2V96fkCOuqY+3eyl6OITsh94xOD33RqJhAhaBO4UGlaSwOsMOpEPkYnH5WksWbDy/VnTN0
vDFZYgXr1VLHpud9omLz1DMBfWu2UNZFCOyifF1gNWTRd3uvKA2sljgk3qkL1GffEpbD2ko356yA
WuZ3owND76XaKAxZKXvh7zQDg1+LSWiSdGwexDfRdaEZTK7tEDUS7o0qQ4JSMR/SWhCu9C4OUidR
OLy1n3O6+btl2cQSMFK5tt3hMOX2+gLeWUo1N3uZGHY7TauXp4rV6un8PNLGWz89itSPlz8l2+IH
QYJaHQ2LFAZYGMKRE6mJUTF7Dld0ruwVdmt7J05uJW6CTvgktagIr3fzflXT3yyx3D6yGHlfQQN2
4LFObOihJCir+tU1gAdD4BuDF4Yhy3iABlABDV5apz/wlOFQ0XBXZM6HAICzJC+6hPlNkUhv5oPg
HvHXCW7Z3WR655mnyWWZWIx3ds0Y7rqt9+OsQ+bglLwX6qy+OHNYgwqKlepPCiod0XXqP8VbSlz3
KI/5IuDZjINDy3YK/V+sw254hKh+aOnjE/jQGuTl+Y8ARGlxwy4Yn1sQY9011AgPuc0RQdaHmOza
BsmFmcTqI/5yfOvYrtXTaCZHDnKYcuFzTB/HaXOQPLutlmVhKuA5YvodPGjBi4djwQc8ZaIdeVvu
lixBTYHXc8idf9rpmodVA9FeouWzGTF8EHTHtuJZewO8pTz9iPpo9AMF08e0CvJfx4GgPHKjNnWP
q3IM+QSvyCxDmH1taqSmZ00Teo9Po8DKlMlulu8NCGFn+Wm8DhL2XWsDY5rHkH0KpVRGkmd2S5PF
gS/u1YDAR/6gHIA/3ZuivDjjvtq9Hgp9AUkSaiNjRB6STS/xiqqdwNrgHL4p23SiwzKWHD3UDKgw
4bz4GZTaKpmRrhNg3Tvw1XqvfNb+5U665xiBzExGj+uosVAIu8TRmAIWvyGqZ3oWTkIQqYWUcEu3
aom0/96o15NKstNrkZMA6D9LKuRcMoN41H9wvzE9EOIAqyUmgnHJFzw5XpO/paDaYmUw66vqDlJW
WpIFwXXqwfgGcP3TeNLAzsPCfmnqVZfoqacvllBuhwaviDfckKVI6fV+s+5upZ4QK9ATjNHstMS6
gw3To1+bThPqr1VmprXjfIoXUDnkcE7QN4hlYGYg4xiO/kLw0tZISqBiHuG14ZHlC6Slwi/LOjkO
HrrybKIxCpgsJbnYYUs0SsVjT/UkfKMsWWhwjByW/9MhWGHJr8rgfGy7KSHOvIyJFrIdxQ0a3zsr
wHmKl4eaY0fqUwkr4zqs66OufCPQJ6I14saWbXt/o5AvB2eBEnpZsZD+CC2qL9AlaGsRXbljrEfc
Oc+4/MwU9kCyn5gign6o1Zbzzh7XLGPY36gsS98PmmiPltVSXTVYZ7AJtUdM+b5DmhuBqRuVlnj1
nbn+8HLzi1pBzjE2tJsEpVA+Vb0SIbzryCJhe14lEtHw2rGi8+pmLqgJOaapNqKkuZnX3Y5M8tgW
YxzcSCQfboERFYz+DuRX0oGbVgSwye7ervYIwl0X1iovmIjKOyccsIPxZk9nyrR473Ld8QiYT2uV
ttWrxwQ4JId7ieKE4Ft9UhS73r44K4+pmCGcllB1LLCNKu5eQyEMys+AvM0iOSU8k02CZS7JrZ0W
6xkF4sGbAlk8oeR5ZdgV6fg/jiQMIOKhlDGAzLfE2Q1q4qqRpa1o0lg6QDujJq4AftvZ18cYR+ak
0vnoMNhTpoMfMwzppYPONVD30fTYGgOAXXWFiHB6B0qtIKxRFxu9z7rQbXDdswvA4HI1mcNIejvA
AecjQBG5q3zLDOYVfg9owaCPHarAth9fyeINJXyGFMJK5Eaz6lakWxGwyd7kj1SeU9QC3wxHihIb
KyGakTnEAmELAn9zSTTDWAI3m3M8ceqwMIW6b4xRIF7HPYa2RF7ggkZ+I5A/N1ZoJFIqydh4Vj15
ab0URB+lKDtRE0B+rd6iTKB8ofEMZKCNNxMHS1rcN5ABfHXal46VDMDqZ9z+Br5Np5ka8qcmnmv8
8zICsBKIQ8/iRI9fGDsXfYBI3OjxxR5WIMyyVEirW6/eQPYL4vE0sJRayXBPBrWtO+jXQJJE78Bl
so0JTFoc/6wgyFqk4iKD12ZbatiIzcBw6IRHIc5nGpoC+LHNktSMlFmJM+KtYpFTavPX3QIEkhMA
TTrGCGd3nn7m0K2wFt2k4U/XZ9hh4QHsJusgn12/E1qXfTvutv6h/TYjSoVUdBG2saxhISlqYxmO
1bGSVe4EHTcEPH5swxXsQkWxK8/h3rV0DZV8gNXQo38+Yc7Lty8zOhtyF4zdVO3muJzrH+zR7cmZ
9Q7W4u6RYYq7O5B//2rMB/X5MJXzDizYLN/Zg4Y4WA+4hsmJLdvcUintu6YQY5mSLG2NZUFPYQ1q
tUEaxEMD2UYBD7KVQW3anwQhfqqhmfOw38m5SC0Uv3QRDzFejFL+zewiftc6AJnniif74r1PBNCd
opj+tVG4aX5Wy4x7k4mSvxFRKUXe6gyBKCBNjX9lVBl0WaGh8/nyJ1PmbQvXN2A6kyUpHRvRlO/C
ViLq/wAoyOwbnkN48rl6HtwFefVUfFOQn5jtDcToyW5M6kFgxQxN63h3e97EntHhwx/OdICWGphU
aoi2bm7OblDieXU45k/OcA3MIN+yev/lj9XDCiQ0wvvoAxaB91gDpE0wnVOKLI1Ubb0giWkDExal
vsEftq2HPZx450w2I/05bFbSgc5djCOTFB1GDF1FQgZ5zPwtbYx2Rpl61C8GIKG5ZwbmrT8qyThM
1JlYcTopcrohj+2/Yn9ymhO7tz1FS89DXYlnLJPBcYEnQn5ePH3qCpZ8M+EluMthUEXsA/7dysT/
e6xJe629hYe4jdJ4SgOgNvYOEtePeCZYKvFvU02jyeete48VlDDxMKeScfCLSNoTkg9SpXeVwolE
v7/E3qMthezoP2PtiWH/KDACnKJakViKKvjH+AZdL/2SEaxYMCKpESRNx+2oAq+00WlPITYaAVIt
Tloxj94QhKDJbgcZGHUCFMtfZHWoFESINEB9CMdpwTtVeOuamhMHl7xmtuVEQVI8QF2BYS7DZMP0
qBb7uJn6MNPpQ29g7Xtpm7dcPsxSQMAfM8aGQ3EJZt9OhbT2ADkVSgPfn1K3p3hWqalcDOce3vc5
HBwn0scR+VQ7kwrLfsxKrGSeMpzxWOG7TSmo3bpQOsiHjOk5x7dC+FeZ6W2Lwa2AgYnBEG0etya8
J1xnaYiwwL+rCXNHAC9+Lqx4nwLmRJFtnfvCkuZpKxDBO8+H/UP9g649C5lZipOTOiyBhUkXLNpI
B0ntOhuMGWnVtdm0pzcfghAb3ZcjSx7kUwiZD2AkbUVWdhoy89axTWEMvhPgS+AXBF81KPAYqFH6
1qQw6L7tvRp1urBFMdSWInd2YNwBPQ0psaQRFNW+sUGwa9YTFhQK3zFWroKEpaCqsvgDB55AW3kA
Q1I/RAgBboRCAS6Xmdsl4ncB2bLi7Keoy5WvRGVuL+TBKfvakDLixiAAmFjKJt2LsFjKXbYkTlPI
jgHLmXJALH5f6WMcuk5y8GJZ3ai5fVjwljXoML3+qL142fv2QNtS3AGJn/1MIpGiDhmSB2jvzAZ4
IenL0nUjT8s8V1/t5p6lZbyctJ2dsjDrER3iIiMrrRRmIEQLIB0Za3jYaDMKWUF4ReB8HHmoqU2I
BinkM8ornzSYol+RMthlIWhKaKACiv1qMTYy+xBr7ePkgiCfQ4jRUZretu7O2D1aH1nT4894QG0r
LLE7YnEXksllzD29qyJVnLlepe9rNC/pXeLPCUXuiv8RgMPPf9VCN5zxhvS5pgWxQhO+srUTspjb
JSMnK/H/jTcMkFd0Gm1CU6Qt/eYS3gFmBkbDduOfUArE3naGC4SSYdfCswmX8KvIq+wIdGG+CrNo
EvM98QFBy1hZ/PwlCM1AupcQGAFEyQQKcton5SntxGQxmoAJFVVzvlh36Sw0raKOXNoi3MXjHiIX
qboYUzXJWXvG5+rKNUYY9QB2m2DzoM/nAq6kvdC4C8vPUx1UxXrNDWt80rjssIeoKR3yrLtmXsrN
02jtkeMUikbh5HEW/Qs+X20zFa3GS0Q9mIuKr3gbuw5n5o5GhMrnGB6WZHfKNQ3civx/f/lEVvjJ
NRwGfPsyJv2zA6fQck+54OJCuNAvNmcKi5PV7DFLPxodiDwmcWMv6XDXGTLj3o1ocuStI0wUhb+Y
wLHpa88tsGwZyJ5w6upjAD+hAVb3smtuoA4fDameVikxQ6YT7NiMM500ocNjIebXwt4f3MXQC2eM
H+kjLoyzueGEZ/uG79bDc8B5g0eQRVHRpd3cmDIKFO03HQ8bJdWHhsshzYi9iesOU4Au574mskTk
S964SvsnXCP2OIroybSokwyk4ZoDahF0HgaNzIPAQ2oPDXgnciwcUJczPJNELoKdMNjaIYpcL/zE
6Ye/qTV5A9w+FcpeVyyRWDWOn9KKxkDeGkdZE/HtsnrKoZJAWJLu34WH/9v+Qtjmr3BS8axqvqAS
IVCDnqsqblVE1RNZ8J3rVEL2qcayFcAF9VihqaDEco1RtYREwvA3/lka54KaUrjLXITQ36Uy4hnO
h9s0rWQIXcNuVqO+gojoSIcQaUWZ4UgsDQ547o9lz1zjdt/r7UfznNZWgzndH8HVhK5UpROPtXf3
K/fgWsIOstpIULqD/8aJ65aIDfzUrPBdPsaRBkKemZmbQBgRlg0/VeBB8OcSKY/YShxF5VYLyBXs
UmlBB9lvPegz4mmwDgZoGdanNQPyxr1qoPSwbJsV9kK9Qmavi0aaPIOqnKdB2VXW5DDhl1dFYTIs
EQpR4EK5z9nAhhNtqpXaZZyfCrOoHxFpMI0g5VmLMHZyLmBIGdY8s03oaH9dWev3NOxb8jmXbIeq
AouPhph5xIzxrueWUIjjVNWZ3DLOR+/c9vmECxSvFoaVWQQISSO6LXrbKaGM3hvc0NJrg8pOzDS7
ZExB5N+t+kXiRs5riI3tMMPa+UzZuAfUk+PUDjgHQyknpkpTYuk1UuLdT2T71gcWNcad2tQ1HeTb
Wr42IayNJD0xEDmE2Yd6ITnU+WPiEXWEAh0koGN7ddLms4HPRXjwa4MeBvXd72qrC4+T6RKbBZbz
1PR+zfJBDtvtQ22tCZGtF80FVQyOTNot9ilKikf+3a6b3lOtgQkY/S7xeONYAUNbmKtCOaTyKE2Q
V+BuiVexBmv8bHJ9aFDIVEq/ax5YsSTmqLL2R7vpCn5ZKQwiOnUarR5QWNXSmGMZU9MW4MNWfDOH
tw/ZbmHy3/5tmkiTNLGEU218Ua2MejlqM8U5JlBttRggI8MQBt9Wy3ADZFfwE3zaNwA0yRX/+bVN
lKoYgGunoaYYb22/Ow1FQgx5L/NZJr64zaalHP+ePcU6QxB0LR8qUNoYx2inMwiQbAClu52rHqtf
UUOlc+zsNtbHn+krYpa1DK5VD8eFcpPg7AwNWZ4shu2FXTNlZtAau15SZTtjtRFx5asCpHqy2d2O
mvQo7ppuBInVbe2NGRdCjc9qnIS+9lfylwOqZpQC97pCEp7yKP3aViypdlylmx01IZA4c1f0RVWq
aHdG2ew4bC12EbAC138HBAp1YFGB5N81nfQ59vFoV1BWWNOXILP9mKZ1Sjq3DGVBSwKYWm2cyorM
tTLh0I/faOFOLpeb16cmxCC3aIn2h/M5J6Q72jDRo+IwT5pqjCWuSwhIzuIV4L0EwREfZKEQJXLN
zoHnhHZtDgdB6F/DNq7JVYpz9orBcb6GNM9byz7QEOPxufJrIY4VRXVbyr8XSym2COkngdrF3kNa
h+EWBUUc7Eq6KOWrj0Urb3eHpAiofLPaJ8tb3xHl6+6PJZQtaZw+831S5mWzc8Shr4I5tc2q5b6Y
eJI0MCWva4E0Za/2Zq9qeNwERJ0la8iRTgYohneY5IyqosBescjtDeKjIvIkiOxTTXvYLAhTWEQH
909VxajAHd02Q/PMFQD6yaotBnoyru4vlnXuuh/S3RD801UQMpxBc9fCpgLrK/yeqWHC5DXzXg9N
pPT4E+TSJj6y/3Y84LfmzbArPjjQuprD64LisB/9b6MOypA3hvqewWplkJnbFU13fEeQDlsGzzmf
XKGdCeVZQQGRXbUVqfcP516DNZtg/0iqnagmJba4lWBZizZPdCWB3wvFXxBJsvd6Tq5flNKweckF
yB4cvG/RH1rphBn/KitcbWgb1KPjjxuBUe+0SZ9PEZ8lIn6VIhZCmh5gemuibRvSvxi3+vcd5biW
Vh1RwBu6CZXxyVcnp2zI/3qXLtZxmMeNlFkOunpz3j6OMw0JrCYsY2KkOKvOEgYIRStcXC8V/Ama
qDDGBZ5b9pMTK/HFdCTdUk9tw9nHswqVGpmqKnSNMQPo+1kt2zcNEMd0L6DzUq4/kLnE02oSA9XC
lzvLUXuFH64AzOVNIA1nq08r36fOF42wnHPnZWOyZfXMB2zTOb+qXNmq0NoGUEGlOwazB/CmAPXj
Qx77k3HlXEfqHefHFMNIqSjvuqKSBOERW/BeANflr7hmp638uv2RT/1DA+hu77nls8+vlIfFjwLb
ASZ/FvKYRL4LLIe9/gmZZYAduTpIIa6d/m3gSqkD7iKSS+RMv+q/uIolKdiuS+BS4vBt4xlLd5ft
nfvwbHeHlAi7R7R7oxYyAkRDMhw8ctHhlhvJIsEpSa0V8cwtrazt4cBYPzF0V8Asy8n9NK18Zrz7
SzOTpogD+HHj7j/CaTxf5OjcMct5MK2ZK6b3gPkuHU4A+0rQy74Jsm1xdbS8YuqlpAHhiDWMV62A
ZGTDLgOefVPVIjSIz2Cbh0kx5eZNkP2KnGGv7+blnBGWVxx+cSrTT10HgXsV0mD3FUNvLqMD9eER
HdFt0tJF5SpHvLsDQQ87mj/0kUN6tfXPSH8C9RZByD7yP2utobhj2FbZsN+C0Kwsmoe5yRrg2SLg
X3xH4ezpCyCCO36qUZOzXa0oQOJqVUufCm4vGX6ot1rLtlTJ2QhILbm3gQLx24FJrt1IHRfhDmaj
M0ZcALIO7KXUmEO05L42LY8hb9DR0EJk3ZLF/v1+HprBdnG5t6Er+fF3vikR8MQx1aSkuSwz/iO5
Vc7eSmEho/38wrAsmz6LUmFjA3NiCD8dB/5vccLpEaCgP/9QUJsDPQRydeK/0E4prDK+f8e78KYi
DXtGcNUKGlrYkI9ak6GmRtOUjQ0CZiO7fK5sIzDRAC37+VvJ1S16sUT6uwNk7BDRoc+fQNqfhcSS
YlOnKHPOANb1mC/ev8s6JcNoGHRR/2zLMo05mA2eUSVoFhwQlIJuL4Z7IGJo16iMgy8GwAd1zMNs
79uXepiCrHY2q4CsYoQ2H5wyTUeyPjB8Yyl4+Nj0/r58+FQ3Qob3YrIiFhH0KI1QIG/h/P63sxwa
w1bDZm8VTYUN/n31qqvKc6oH1bNxQ2SwrLGpMAO1frKoUwDQ04JM0GjvZnvxexx9397Xyb/5QP3y
aLTYewhP453V3LfwryMvOZ99XklE7/iu5B7LSE9oF8z1mrFw+I3OWyTiVTbWVgD7+06yLPJCU52R
SWEXMpDWQ+rONmSBrHkoUhgBPH8UYFT0pn6/R6bcZ2q+7BW8Anx5nddJoL6jCPoYd4nFRFycJccu
j8LDbqB93FlKCFTun0GnmxYAVoylHNfMuSHUS31Uw6Aty/9p8hb8H/F1NkKL2d4uCHHnX3trCZm3
d00YaqbmAPyptrm/vfxo8K7DBq63BPNAupO6ro2cXXQuGSci35CPIbZ6ZePL37T7U7B43UweZNtZ
oR1oF5dmNIcmQjgxnHCthjN2vw4njcee/3IZgiy6XXiWJ+gjE5bsdUypv4quorztDZctE38sSibq
8yyzmSjvK8dW3fnNqN0W0UhjwGmXCwQ+JOMBYT80wLYKAm4y8YCnTPYJ19Ek5fCWhIIx6omzN1RV
0vIrSEaDrPobfTf5FQTwf2R+NpR6Ayar5oxK33dMjCBxlm6wzwCN4KRpsdbRNVT91KaCu3iLf10W
9e4KvVtp5GhW5pKa+GGRwfIrcdA3j20EPgYrK6Uo4f15chPVY3z1kaf5cEZhJJWH7Z88nTaZ6o4D
WgPl+YwbY0K/f778MBruTXzgZ6Dje2KDggogiDqxTlrqQDaXlV89xYImC1eg2iA3n4PDQW3EvszC
NVApXR8P6k4sZQmUFL6L2HuADGbmwpCIhJBA981hgW7cVb8BCQznR1g+5sJpN1TE0StJ2NpCkjfb
JX4MR4oMe3TyRx1T5ree/zOVX/JnFDomO3G98awx5WiwMShYRAB8jVmdefIKk7abtVj1swU4yqe0
PCd8kEeo+6GpG5kmsP+dWutlVK7T+q9aBjR+ddXQV29ETHsnTzZcDznk28G2Shm0sNdYAd/802nR
Lqj6FAoLAtbiq/KeU26E45MfwqwSQRLrKVwKWGQp9zCqcTBws7YLCUaBnA7Z5rX4+37gfdgBzjJq
38DFFGlfM/X4I+Yb02d3veu3yv4m5b4zrr4KufKQZkvI9Y9laR5pq4g0rWy6ueNs/aG9WRiIQR5P
oD6Pw6yDVfFRYpAZ2SX8tgxV96KdCf5kdyt9tvr/JQ/3+djsv/PBXcC6xT6ql/yYST+bfR+Pkk7g
2cgla7Zu71J/2mGAlMX81VAkjErWw1J02oviy5r7vAQdH619qYuVXmekGGoN4KqX3PKGp26N/mN0
WOUFRuxKDclCynIedq7e8/9wqlypALQySX/NSAbMk9JJBcVOfHoEnMlA77d6XBKnb/Sjfdi7K0vB
ENL/Ka/LryxnatS9z7zHTZFydQ1VgRcHr4tVtBUrBA4hkQ738xZPYkym0xomTAm8FDICEHcD94qc
yMr77MfOFskx0MVgkzXLYo4C2ZIJGakLa/ImDdvhizk2OdCoLcPYpKBKCBq+Clmg7V+5qH8oesbz
mamG0GCB71IkEM8X46NpJp84+TP2dhYSiNQM1FGC8+IOr6JxKD/G2whbX6lH52uzl1JJjkZRnVbN
yc13UW45D/eu77LMSL4MyQV1BOWz+IEAozHAKt736LjlJJ5+Sivg/qhBZ/h42AKzh+GzYYB94g3P
3F6gRewf7HMZNpdiy3VYZnPZFiChmug0007mL6v7q5TNbACAZWbA8XkyOzFfYREn2ovu+4qWiDPr
hWcs/TNpd4Nm8prbYdpzON+RZBhlZU0vWG6Wx/B1WeDkAnCxrXnJsooNTh8G5VkqXf2y7lqwkX0m
joBuqaF8LnJRrkMXz/saRCvBzgo7XPlCB+sDl3BlT2AEnzBUh8wiqL4ZRBBpAjefDna70Pf1k6bc
dxE63lrEhvXtGo9wkZWniN+HiiPfsmFfAFVv6hYXcYu3zWhjMU3CTeAUis26P8m6gNnDf02sAaDG
EnpDo3bVi5rmvqiJveB9upEmwhjBHtZRFPNpFyEycjV+YvAjoJo44Q9Wb/1zylKZkEuP8tGBaoy5
36Ev2erLu5G5VO3a3GUSrmi4tbpjPTbrcVtesWd61XQ/HPTp7xHa3SrIKUFN3owDuYdfCqoDc5rC
H4IAzrAj7Ktd/CYosbrGz8KOYE4t5RsbUIujG5cj29C+FSEHnrP24mpYTcP1EnLGfjo5X5YRDnXP
cGRe51M/szrsTurXwOcRRt0xS3IUxJXslwiaAVGAvkpayec0kZ9OYMG2yMWxqzYncnvT9iFZtxCQ
xyMFZHX+zAfjHcB4sJ7MTg3XmYGWF4puzC6KNU7FLzVUtKsD9VtHXDZpbgz0N2ZDWblpJs200Jy0
8nMt6UvOcUJKTWYwBp6dpjLqVTWOYh/cIIj3YkBjvXUI7LbyD1okhyRRJS4CzO52OKf8VjXobarH
pPvlqqzEqIq2X7TsztnC2oyfSwyE9UTWsj5HtDbSF8PutviDdyTMQPnOhoukY2n0ZItGHNGCulsR
PxdrZrYbv8kzKh3NYKMGn5zL5TV5MWEDDFfmFDl7yb/QwNQ0OvInn5kAZ1akYRVWKye2zG4j8PMU
sgUoBaw51KYZKm3/nUAB4M/MaoeazdG1Opskkx2jAVFpWde0QQ2ubVIu1LyGM02scwzCNipLVrhl
d1mo8CR4y1IMANyKVaSKBd9Xk1vtKaCKSHiRdGRK6VKAz57od9zewQNlY7mXtYCoL8KV8VHgYwR/
5RoJhhuj+1zKE09p5ZreozQQRyi59Guf/rKWJyQmXo5VPo+1dYvMV5fqalrmZH/xWhI3c2wh3YsV
VUbXKvcYKQifCzJNNk2PRfGumxkmAWF2Jd1jxY/mdxWft9+AldN1rahOnQmcQOh89g5wm53UK1jJ
X2s+qN+ErN/+bQarUC01K3q/UU2DXiK6mJfVHv88nBvjVMPEm2aSyu1hx22Qx4bj9kbhvggqgU6U
F1GpPNhEIz+eeqvPqjJlbEWX6rDxwgwWyfuauxssXfHzhim6dzKEcSFpP4AK5J1NfoQ4E5iWe/xW
3zc9s7WX5jkD+8YeeBRUxk7SHGj93rIzBI9FtRhW+jYKRL9Xfefz3qw1LC73wkH9IikYG5cje20g
rvPSlgDc88mPrAQBWHKxiHJe25nfGcyHHfQfbUveV6ADBQCGnnG9oxVx/2x4wU/GpzLi2piTRnuZ
ry6gjeWJpvhL1NFww5nMprXF1N4MgS4K46FvpL+VS5XYD/cgIsfMusNDiXYMc4Jgsw7I//TyvpzH
sOdc9LZkKfhSnruFW/Wr8HUjKeTqwjC4zQdhAvBADYj/gqfjEUG07+H98lhkFGPPGChncVxnrm9q
RYBs/AxHeGm+UdiU164EQ/Ufc8hTXXZuARv98l0IOoSdxeOpqK9k/idUfjEvZ0pIKW4Pgp0HNvJd
za/7zlwq03Sne7vWJ3bejbbE/snhj/lK2lSGrik2NVLoHnGAKL5DHLaNkAxwltcfwap1T8S0KPUe
TnKJ+mt/E+2NAOwvBdpmINvRqyfMIPLAOmLQzba9tqPKQCLgqS8sW1R346yS7tPI7oLZbAZsBiQM
YaguFQHNbpEpt3vC4ikwnFfuyY1uU4vyBUkJ7pwNPkpG20nCAotFLkk6kOixAWPaxjmaddLp+YC4
V5rSYbCkglTkInAMKXpsDAAeOhaBeE5bfYSV0ZStCeU8elIKnhQnUYbx33553zlLRqbuzSH346je
relbu85Xprccop8PIwFq3LeD3w0Zb93VHKpyMIT+U8xE8fHP1+9Ey9pjsYCo7XaiHrlB3/01snbF
3nWeoMDSppJlgTkHVA3XwGEPBQSjaBtqSpqgBCg9cwA+4LrM7oGtNWJuFpajBXFb2lspNisxVjrt
W9KPooSfeNQv6uM75ZtWvBYubIk6nLctbFb+iHu6W55cgbotF9xlCJe6H1KrePWgbC/vo9hV9gqf
U0eGZ4jbH0vvih6W6FfeLwlaa+x/p+alnJU1CtZc0yBaWNB5CaIVLOfsO9ZZ9Cpdtq0UpHz6iB0K
Mc7IIheHISl2zg2wSXqZXbiM1RUfF+pS3NLNT/XA+I7Z4WFApHFdcRG5IFyO3jG3hGU3I2RVAB96
BjJ9gqBROh+ykMYgove3TK88py3XQlPBOIQuPMj0coI0e/ym6DFLfMvIhE26caWdpZMBKMLwGB+v
99dbILhza/RKpMoXuOdKMUq95MjQ/lkgOMaR8inhmLn2y7N8vxZSOtfehDD3QHVm1mX+PbCnPmcm
1KSFwmQWksjOdei+EIObvpV53D1WItRNrELiDKJateuf4k4NLhjNtQW47xIcsTODCJJ5o5O779eJ
Au49JvZbKIm7wyVa+Ewbanue6nL76Aiq0LC4PqcTTFRh9ySMwgkJ/In/zjQ/RQKxzypcRdc9Zda7
Fhxy7dK9YQ/7UlhGkY+UokJucObpF6Ccj+n1sIv2PkS8d93Kf3sVHMuOgMOupeyAvxcnenAeSfgc
Vybv1Vq0Zs38xchhHMMSVP9Xbg7NQFc5Tl1RvibPUTLdII2VzVIzwXiK6LL8nA0I592vazf1OktC
MJOOBLIXjQ7o+3GiMbDgi3I6fP4URAARhEcQGrG7Oyzus31IwIY0+HHJ3L4tU08oChE0GD4SDlcH
1/6pqMZdhWxtErJGPGj2ELoUCzOG0oqKcGcGTwbsHUpwOWt43gv4nBr1v0f7J/tzc/0BeCenN463
o4dwkbDMzyUinAiCMB10gSWBknrztOCNPPnIXrrN7WX0n0dUD+cD6aP6ba+Ddea4iGdbFcDm5Hvz
rLJ+ilvLKMRL0VivLy9dpf+EkFsH9ErbOOujX3tgOlG/0xj95zHyATb44wY8Q0GEnQ62trHbW/Vq
EyIfhqL8o1xj0hvF+NOZoSKvqE2100Yyv1T+gQt7AS0UPxSaAJKqcJA0qmTWn3n2IZ9MBJg9lbpR
i/8+HMGGP/93bsNNzCf+3cd1nbmgoxHrXwYyzcdg6TDtszFziiDG9Yo2sp5VNDDpGPjghD6sncoH
LLOMU5pdPigQXf0CMiGDIG6CbpB6PFoKUg13uqWstvk7CN5zmi4bvwHaNj5cx14AlTFDX9V/3c1r
BqLV8GII3bhvVAi2c19KgslyOJjpJ6EOarvBqlciHI7GKakfoSRHFenRD1Erl4H9Rw8pPoY+jME4
3aa5eRvVyBLlFb3/Fcc9xJ/M+1oRUmqm0CSL03ci8mLj6bOPzgEFMERCKLSH7gVPLItiqg3s31BG
5HnNLYGS3QwmYyEgzjWWLQGi2/9JfIO+sBLeRINul/MI/3NxuQzTY5CQwATiUttl2rPWDJc40d/T
gSV/UT9yEfE5tyQ55qEY8Bi9n+kdcOywu0OPaJe/HAAbtJf+1BPtbZ3h7rtf6ZgS4g8P9Ln8w6kA
NRXWjvoYvEgFNNk74/q0kbH3gyn+4Oi5V0s59I8hrZzryRHWNqfeEdoKy3VfuPzaV5dshyCJxUCH
iduXLoGFUaBHmiKW37L4QPjMbGe9VrbqI69YS5wvSfvRYufeHaubTeSbOdMBOATLtjQkl8RZZBvO
pN0nZ+/dwXu7JQw1zmvd6I+BN5hdRub6NXL/j89wwNVFsApIjmpO/EXSYISX/L0SkqsMbqOXqTwr
itYleJkOvwopErnrpnRx5ujGTN+MeFENjLoitFjUkM6jFt3S7UuQ2dh88KpKUiZP9C+8dv4llsIf
KEWhXMbOIR2612v8vK6vqqFgzZjRzzviijbbkzVE0/ucq35E607GH0nHXUHEGwz0JJ0KocXF7sJL
fxzNZVOvV9b+NKsqOMDcMpsGwNR8dmYD8xjkQwvzN5hyzHgKM+xSc8hDN0A8BVuXe3p8nQ9OAI4V
cCl3b0XKZ2i3HXBESgQI3U4z/jBRNF/87VznwLzGTzB5Mo7tLGiodRQY+YdQYETAZlhbk3NeicRW
vslpV4nngBkdryceudIB67MMqDi6wTaBTL+Z+lasSDJ9AmCm5b4ZtNY0g1DV3qzA3P0694nytm9P
XDE3CSXJLrpM8BmMA8B8OiAxDEcW8NXOe3lEuOVoXKijruHDroaK25+o7MLNXRNytFNlGKGKY8yF
NN/kvidXVpCbCTEoePdttJrASlYLyA3PXfpgz3qAOtBYlYu7ndjcA8Kzd0hjXckbr4heS9bef2KE
br0PLbjERLB4BHS3M6Vv1Q4OUZ3cSdNHSrKEGzTX2WU/R0vD7/4uOQ0BnSWW6SV2Zq6orag0Bna8
BL7SXC1q+bYRbtqscbZkiZGfBBpRK8fyKqv+70JSrgPreqgb4CAmlIRQjkQruapGl681+Y13aH7a
R+UohW9K7NjnUDnMMdJo+dgzOD5s1QfTHLV2BEPBZY3ew+HIBjvyphcDU9xnOyPN8LYfInJpEUsQ
ScEhD45kqM5hJ6wiflog+6w0vdktEd44OzPVouZGn1Ru9z+0IAVIDuFTvx/CZU7JbHKSjH2oj+dr
qSKPnw6smUbCmsCxmvq6UTe4vNQp2KSAzM/p7ev6YnHANcOJtY9BaYOX8z0b+odYE6ji0EXGst7Z
aOYMkBaDUHDOh/p+NVO4LKWwN512LyuhkggaheEkM2H0IwOn9ID0bs4FrI54JPHTvgr6kznU0mkT
ecaRoD9Hw/xG2cTeiyi5aUYwbjNpLqAwkoSmFerVXkIgP9wbozWaw6W6BD+a8/04CGRQF8P6hNVi
f1+T/pinHodLR0aAZS5/VjOX/z2r+SmJ3UUKHJRYt/aaj0yowulIcJA1xx5lIVzjSYRWZbG7ztbf
B2xO/mx/TgbpssvRiyWPhhkSXDM2zV6l6Z95KZNHxlRxq4n5ItQ5SxDgit+Jfk8+k3pWDg5YuGU3
qkkkciYyCGtwCBYIt5cXyk70WXJs0S77ueNfeZhUFHZjFN+dQh6uFOrqVsxZIcyGYPDApLl+nbsx
Q2pjoYscXZYagoDxNNQB6t9AzUk5AAz+9CAa2HE7+s7HPQikljOoeUoh240b7o9HVOefz5+3OlPL
UZsN5jDD3j82M/IfcbK2Jy94KSiSKs9uQn57/2nOLVk/mgD8jnO0iYwdT+EBgshWMBI5gTI8/iEl
BiMKGTNyNMcFWDfiZ5TQ2lMzF61kr0HMn7xfdHmMHiUvHk9f9+7mx2RcTbA2Rq3ssUOg3jZmE5Ze
3j66+QdFQ0wnOh1UKt4X/XHSGsbcmNMRUVR51mLfsxYd3JSSYUr0bh04I6ewhFa8iYudp7QYFv78
kZgMhoz8DNCLp5n4n4n/qMIZtThnnqS1J4AeTfDC/hSCv4rk625RIVklwmYqNnDBPRgBNQblesbO
Mph4zJiu8cGGvN1rsati8cqdktxcaq9ncyHoTeW4yVWqCjRY536c12UejItMStoHSPW2PIbdQNLS
lwG5ojpYuVWTVjBVkhn/hI1exNz/5hLMhVoPsu4f1A3tYZJ1wmvYfUf0htQJWAkblczRpLSngEQQ
UKNmk1vTI6UKnPgFPwdWXiSmn6E8Oopn58R+xatKHXtpSQop7ec1PNiGQY03kSk1wrRF69eoS3eF
IS04e2mQTrrEHWbqjPHiFF8uHGIZXYvJDGs4vRG7BtnPR7/Ii2JeWJDUo9ObTjtV6wXFJ84t5Czv
OjPb3i/kvD23cD332SR3gNu6RMnH+LMN0U5Dg+BHbJsRtGY6h7fdlIXOsMYgd2faPio4UGHAS1bT
6GFwbNlUoUcf0nhFUggU47uBqx/s+j5x/WbCRlrLTOmq3EwWz4xwtYkdP6LvNyox+nb+y/ofwFzE
OTGeLHH4jqnQQGT+N4Ad87Jd8RdVLNbIklbqdQo2GbKUQlvIcmgcvn7eOVZ9pmFcUvCDe6nR16Yp
5elLo+Ftm8vqTyCuZH1V6PFPqeO+DwW6FDS0Mr0xavvSduWoe/k22+bnGqWiZOtbRBPQXNnBG4M6
9UofCKW6QvYyV++oC3ZjCXp0wAZhN43taLH6AfjyhY8A73OkG1Al/GfjEcI4lN/cTcmRes8Fe4z5
Dy0FRhasIXbw31Qn1K/MI8hRW2UW6nGsnSkhvuHgITSCsqYT8GcYdT/OdZQro6tzXzyqjnEqb5+k
TNIM0MebvA0+PKQnm5guWs2Yo0V9I8YzP+Suem+L7SQGhipitCigBAMa/KzKLqw18rz0bS81M43+
8to1tMpw+hzDiGxH6Yph59JhvkIQbpSjjK2SRwaE4BKXFNMX3sXlWX7o9wCOOmuzDWCAGdvVqQOj
KVB9+gFE4crGpxjRlpBCLuTkF5RFBUxV0K0lSliHlRIwnGQq6RJ+1vEIWlqQ2qmjHh4uYwE53gnd
GkgrP/udjZL35D7UBs12NHt3xJFhkDUREaJW/E0OZB+oStQ9P4ln+kpvBJlNZX0pO3ZMSRA67fk9
P4Wd+A5HHdD7QoVawKRUn7dOZlFdiw67wMwnsRt246/ont2c5TvTBz5Hv0FdWWkAz+VVNJkFpG3k
u5UewdvJA56IGANxGcsbDajEJ7hT3F0ckP+SXxaEschFQsEpYIuXOBrYDlrYsSqbDQpICIKTz5X6
ZdtixGpyKmmqFSmBA2MhK59UhmA8h+P1YyGXFwJ/0TmEI1mjTFVGETtkK8WghchcjuPi//TR6BA0
qbWs+Fkar99AICX0uTRtFnUSqmRXaoCUGXyacHcZ8GaZwOcKPoMRgoIgWS53VZ2w+sEwWVCubZI0
6e81Ypmsy5014UZGE11JP2meOew16I1So7W8SsMDtzKyDl5cNccDIBjcjKNi8WG7u9NaXnn/vzwE
7hUtB3IHD2f/0tGxk12I81HNYpXQ27yVeZ3bTxJ7jD4tOxsdMM7YTlifm/QAe5iJIOsKJQ9XlShR
EUwIkkSHEydgbgz/B9iJHcz1fqd1L2SOoKci5+1wcHwccS928n5X73OkYsflbWhHqwgZsB3Z5Zxz
G4G1HByr2351eZ/f5aowEuPqtDRB2KdaRt2YxrmyHwYWlZLOtuYmpGSPss6h6Ah8pOT/gsxFES6m
+GW6q36Vdg83CCoyENL1i3PBFkloxcRg+uGXCTyxN2pO6ZLQKqXyLB/KRnRsc41/tpHEhalpPPAc
WiFdFeBsXCF1qy65gsVLVAWUNmgOqoOIRatFDzB9VtuoDfkkZlg7+mxOyMvnfMwnLw1801ZlT4LZ
9u9G1cD8u6JVfwpS6maclEe6DwJhkGccmruLsTx39LYyKf2FZGOEXV1Ge6n/4xGRH9OwaZoWCx/D
h/JV8x8p70QrO0rfp+O0h/zzeqkkCXF5mEYXZo63MYTri2Et+rNTcdBmxlvjYC83kXtMk1DZPSVb
HE2DpkEAlgugMVYgqmLuLL9EimheW51fuQOib92ZgHvEnHHLMBzOUAdqY/Az3YYOpi+BJBsALE/a
F2yWsVLefi0EDt29ZuUvrkDCSAfqMfH50AeFxNNMmdWiLs9f9uM4uL/edgSU/XmRTDSS2YpP09hS
ZnxJ8goSEjeIIPq2dE59hEmwx9Tz0aN8UTVv7dSbOHu+xoX54ou9Ed4Oai9oOea67tGCBwHs1WJs
fCPmns2jRIq0KvRkgMv4gWNQAeXQaV8hajKPjZEFZF3ohxNs8z/KvXTF2ydwnHh+90uoU1/u1VIS
+MgM3qjwoH7BaIxYeYw20MJC+mp8Q7UBbTe3WwaSABpX2QkKt0Pa3F5hD8ID1r0KhfxKALmYnRhB
Rh9nE4R0Edm2lJ/Kz3LU1b42NsBT8/Z26Cjblc5fFaTMdV9csl7fq14WqkglKb7JzMAVqCYsi50q
rfVKNpFJLmUoYjmXxHMYwz0j2h0vVDG/WfaDGe4zT85zgKFJSNweEk7+gMnO1YgX+tdY7imQyzrs
IQNvyNeHZBkosCe81Bb+gnhr+b67x2CPSvfLikkcDzY7YNJcV57g2pvVIQHxL7lIu6zsBoHqtUyd
ykQF4GrtmfDpA05G1qKYkXsnOBqwJN+VpfnOLRT10d5f9E/rKP1ILjAmUyi/vGbaTvuvA/Ydfiy/
UFbOlfuoZ8XljBTG1IU95qKiuOxQz0gWDooj3jZsHEDh+6JaObt60MKeXG2zQxVmPr+dvbgWU4XA
KWqTd6r7W3l893fZQlP8xqJ9RcKmub0Q46/6yKOSu0daf9l6LPTcEi6wn6yzCfFH9/MOLv/WJZP0
4Ni6eevjr6W2eGDw3CCFJ9zdI2UREUifl52yyyTqm6y4Vdr/hHraF5uastFQ63bA0+ENPrFO2Hfj
OsqsTNP+Bel7F1RmD2il2KJLSEObZAet41h/HHOja2C6htuhm1G7MD8eu2mwd2KJMSpwD7o81LgC
Ps2cmMExpdzKnBi0Y2qO50rmaojI6tWrqUY6cilTgPW3JxZgRBX8G/QOpj+xs3aNeBOJmKE0iisa
B9DfVaMEtw5h0NdyysViFVGkzu7J6Be3kSUbcbeV6FB/QfBLR6V+RQzMBc+9nCGNN8HEwogX4Ofv
hsuWgDjHYXGi1CI4Wal9GK8pihaZdTj7TJ1FkqzegbZYK666fpcoZiKPla6K5QPUYA/bmdzBZczj
U+NIqKJtM//HUdG0Y/t/hw9hF/HIiukyaFXEQmrgauZbCeW8sqKD7BQliCui/1suAQeqLqTpOuFN
1gG1SCnA5ikLZdMCbbww3EPLxLssA260WZObYl2kUoNi1s/WEMk095+973uNflgGas1dtqPVrHv1
o8+fDchq+CIP+HoZieqSOgVagyjSu4OKEuz8ditpn7guVe/cepVT7pnAbKVc80WGycKogjIfH4sK
9x0o8b2wu5p2eApSvZUtJ2ZCd55uTE5BuH0+eiksH6qnRqvZpyBhtTyZLmnvbzC3yR/EV/MrCanv
yxRPT7mGlOYKmwEDlv0+33k7UmBl7MBVRITlscu+Qy+hNh0+/PHxSXchWEK0MYFRSZVUFgd8a2dQ
XOd8zIf46TO9S+bcf3mtFRA6awAtiWaojQ2I84/8zWR567hO7m2zeFRvEcwxzWENChpOEu5yG50p
tVD9ZZZiTBdySPNGvMq+ct78W1GntrKO5sDg92ynQVzJ/NmmREJqhaMb0+LwsC3BXlpRVfDJ49G7
fialAMw6XH4ZhFecgxMRXV3uBVd0D6K+mV3DJi/Kb1fz0fAb0k1ki8jWBAlypzVnvi1fI+KwuBli
wo6m1OIJfWbzFjqBVg/Q+jYC2o4fJoZ5ss+OIDia5Jj90pF3ExkWZz1xQ3+24SUgkYH5fuqPX1YS
9yLKeI/2fltqef8K0EnOLz+vHaccu+Js+i3QvT7jGwpebmFsG+kMSOf+WUQ/LGH2h+n8zFbPcto8
FFqK95w0bXDPTXAvuj+OnTRfCFniwZTlT+CJ3zdxChF49G+iV1jY3C9e7k6Qyk15PTYnJQ2JTKrq
fHd6ckBzloPGYTYgmeGCSuMVdz/Thk4cqNL0NPVqhKyMOwQqTSytdukkNptd0tkaE9WwYOsP4yWE
Qd057e4gTXRJ28b4lEzUsw81IF09xjFmeMCwum8Fs/WxrIIQiC+RT0M1YHZj+glR1OkbNTN8xNAy
L/69V9vznOdYZb5K92HzgvxToxh3hPCmOAW/e0a0d0njmsqt7fUehvlwBC+/CqR3qvWBwsZBwJVr
Hh2VtJiNjRhoit5lS5m+JSzg0kJGzJ2+kLH8QQuQ1dLd/2n12OrcBNagwW3yobT7Ad5aUNAu2i65
HPTVJebPCrA/dok65FQdXjy+/GswwV9Dc49aGenju4A+IYlZf/VdJDNGzFWz28yjmFKvGAHYRWGR
76O+3nSwNaEtKgpwKnCsKo4aUuZBygPSlhFw5xrht+klGCclCuLKjKyfnOaqf5WUFa2HGg4XLf8z
RJB/g/dHoEsyhzLOWrHl6LXwDJ44+8x6Gpze/L+DBNZCAdfqBNp06grmNJdgClg2/zDkeAIww0c9
jaUI3QfjpKRo+Hx7rxH0lL6plCfzmjS2Xx++leCzhPiaEkHCDx6pZRC8mcHrfTbdWsV0bPfh/JyN
VDyxFjvh/ZZTy3uzWs81ItrpwQiF7YaNdtSqfpc+QlKDlNW/uq/3DeEPNlwrk+7b2EGF2QnxxeCR
g1VrZiCyLB8pfRdqTkaDBQddZ3LkcyJhXR4pKrRVYh1W5HHyBT0hAHt3COt+sjdUfEfAeKb+/C4y
7whxnb+E8k03IdQCtldXjgQ2qRatejE9GSP6ZHdSN3qjwvaz6ZmJ9UfaFWn0dCjuQN3qM7Rw7NSm
6SeH7P4hBHeknieFJfUfpJsAnXda7Rbact7Xhf7jxBF+3X95mISEoMiO58+K7Sl1y3VN+ui1PSix
/1A4JV1vysRGR3KVFpbIsoHz06psgC3XtR6U/KrKRAjH0D4JIFtJL2M0x5h7pSa3GDGLTXbbeKM2
etQhFQ08i2nG99hlAC69JAU6AjNmrKWOMd8A8R02oWWCVBtHNQbiUDdZaO7+2IJc4/Qxi9hAETLv
1usBvLZ2zRV1x0hQVxxQqBizr4pESyRWErzdR6tYKVCR/8MTHcgchV3Nxm+wTnocZZjVZvl08f8D
CMgqmNwPdnubRmp5o6ZairZg7fQhxtui9XfccTyU0sst+pa10meApqkqmO4FQ+q0upb2oS+8vup0
aaKrRXW6+vz5BPet+ST5f/wLU8sSdoqu04klpWnskdBOIsKiB3So2I4B47a/1WyiOJFJtVYZMbuM
phd3XY7ZcLxTXGkZs9QRMzvvdSUd5yHopdKj3sDIUyYJ3Hr4h96b9ajHa9BBnGhDPhMvmF9laSwb
jlbGShe0qQ3+zbrZsDYbQOSqjBpUR8cgq0rEu8ek8zDyXSrYQtaqt48gkDXzBEEZwulJir4HTFOB
845n35fzwCq76GRXelvucKQ2apLZgMUsMZHFQ6UUgEvkO7wsnUNzfMbaFzkt95vBCMyCNX76HMLH
aeb7b0YjNhM9LO3217u0RLcqqM2cCnFY85vonjI7osBN1lJAvKzIwuyPcHPhuTKcZwa7ENZDFIb8
qTB9KljH+5Q0dphceWqsMD6xLWLGQaQpQbE+eZEmOs1Yp+noKAVrgcMLg+ZHRJp/bsWqt1/4wKXO
rRsukWS0fneyzgvNJPvRfv1R8Ea2txyMvBmMwXuIkUiq/CWJVa4/GNvuWLHVUDc+WzWfTEFaaOlJ
50b4r+rhAOW178/Ps/laOJn97OB8vWe1CHVYl+O8PtDJ3EchjChZEiBlieFUetdQgbWhsdh171Fr
kpQEvFX5aYjsRPay08Jp7oZQW9jYx4itc49fPYsRWruzObbuELw6Z5LZT7tFH7lDsmgsWSJzyqa1
DPB56Jtf10NpY2dknYbbv3PQPtvHveorQuaoA1uyY48rgB1APLwCsIPWh/jbYiREUlBuUq3v8yec
5wkLrjc7VCUjvTvIDKfXTGB/bKa9kn4U4e90LYRsH1jQ1lFeP2DfCjgufm49yopFOjLS1MElkmox
BbKk2zxiIpUB4v1rDaFil8MBuGWVxgR7su4jv89iW3Xl5NbVTYtDZUJpeWsemGzl332PWAf1S5Df
+7zIYQh+CIzlHHWPnz9iRVmovhWNAWKTb+MelnVVwxPzR6zAur2iZEqg1ZyEtTs1zLJA4uIwhX+J
G5fh18O8OQftwzLpCvRzUx39XT6M4t5sHMGRAJZGujgvK3sqi+Sbbxq4uBVkNExEG8ktgtDHfZo2
rWJOg1O5P9P7sqbnb3/L+WhErMMUIBcIWJocF+i1XLDEpoTudPqaWJ76smNO0RP+X48tTIgn89P6
peVSWCeoHgTgoO0X/8kF7KnJ2erDTJm4HKODmaESW7piJqqiJpKINMKxdYdcG8tq6xejhiZ58jf0
KlJr3UVm22feitoXFdcjDyAGIF+NarL2sXV/3h/ivEliPRZBY+Tcvk6pzXLa0IFrsJzsTZ23vrK9
xzMvPdBphhux7H8EsUU6PAY1+ArzqI2QuHL1v7T5OVxToLD04Z9ofVpKFPkOVQ9u2l9TfWi1ZIU3
DFuilPHxoWyGt/LAewS/hf1Pm46pb8JAIqdQGYcTJ8O36E2fy6G/kabT+ypRLywyQ3UGGQz3c3Y6
FDpyEqunyzjx9g+OuR8Hk2Jsj3iOzlZqOsOsf5GrobTy7Nl+ZlT6Mf2GwTOEt0YCX8QYjrHXqTZ/
WBWJ6FR3flFtFHClPLzg+aW2aGCFQ7mveRjEJn2FCVUYMmxod+vyeduwPY+xAXSib90C2v7UFLyv
IBrf+XUkHCnk+VupkPZXZa/BLFF5ko2sfoMDr8YurKfMNhpRgKOzXYgSpZwVhmak75OKooO1OA5v
LOn5WHfSwZ4VI83189SUa9kG1DHO/CwcJun0eVg554VCj1bpt3WksbD3L0b/DzOsCKbxxKDEASlk
s3zs/tSeFUj3Dp/ylWUnk+yO+xai5GodJj0s5sQGugYJKZP65VOFLHvdRKed0bDf9pg7vJZ47d6g
Qp9dJyq9O8saxgZDt4oiZ6C/wUXJT8kktT7IgC1MLxUsOR6/fK0lhu8ho68h2FOHBkYvfjhNKuKX
A7r3ikAEP/SL7WxRTufLYWrg6u83ufGdZXw3KAAN59wcvFpfsd70LXltm6OyN+6miyr7WDUzsvT1
iKtXj+9CfKO5cojRZOjujV21SXYp9KYH2DdhCFkuArGR8fdZC54YqucePp6PSNNDQRpdpiNRm+9N
pwTr81eIIewHMqtX4xAvHsd2L70TBL8WecUgvJQ3cXBGxK8Y8NbNVu7kY445jLyLjqosr15HACws
+ngbd6Kl0ZzlDpPs4UtZS0Ui2QBQ7Q0IafHCr3x6hyrW3iihijkFpwCxwCZ/x41XBwszdb4y1tbx
0zo1UO2JDAhQS0qhcPbZTi6Xm3nimvv1LSKHc3ASfiqsYBIPUWG9MMb/ChGF89OeRrbyZCbLalBS
nTYvHWfyo+6xw5vUhEJb27XG/9W14fbMw7FUKWHTXDV0sUA/K0T8aH8sE4rIhYCYyR/7WeWtzlll
fnqQIJ9JIJexCxUbVJiM6LoselLedkq8mN7UFvof/nxci1miMvygoFhZ6V9dL93KmXzq4q9KRG75
OApSlJf9/1NMNEUiqfsxaH1ucH3bA7qccJQ60egVIi2o4pr1jNYyLgmyiuUIUjeIHhclgUDUTppp
o/CmnlT0J8pwe3zKqrLiGuz9dIFZAZlJfQZz/oWlcGOoHYCd2lFWquJCx/gPnGv737ncch54Trr3
v9jwPM+Te+87a5dhjSfQFgfu27f7nQzpUbSUT6s6WndfcY13jROBn036PgQqZdm7qwIG4iJSIgp8
2ccYx84KFVf4dmvcM0zmTR0bgYd00sqxTJMBlfjplnTd++/dYIb3r2iZ0pZFVIAQtzBH5wbJyFGW
aeJIbbLxn1mphCvtn306CXgKC2JyFvJ+EXhU3pVIVh/G25Z1qZAiL6YmW88eCzMgk3Fhvcdpmqmh
arfqfjY4apwSLsoHBdT/VELW/noxcIfJCDidUjriKCY5mVOmleCn7xYVGk8nMJHDX7SqpEK4jOGa
qL1DGvB6U37e3gUsxwTucvlKlE1ikfHySpC3IGz2Opqab21GdeY9R/AiGvf7umGm1Y0MBWn+63RK
8tTeUhG1UtrbGPMYyH4N2yCF20V0I1aqdhCKvgRglEHqbJ0dkY2dzh9tsFDH23LYOvyUQqPy4RBm
nAJp/QU3Jpy7WvQVbSTMy417yz/fepG2IUWd0le6lilJn4wV0EbRWnnIOBjRGIWNkasSP1emYxQA
3eOyTXUjBFRI6bVo1VYoq2zurrZa7LdwYq6h+HIkP7P5Tg5S6CL4/35bwNnwJEKXPRxre4DL35DN
N97oI2FfgjkW9Xog9Bf5+ugzs2dcMHz9ahnK92Na8UlUP03744kXmI1or0yzicakPQwRaomGozkP
XqIWymTcv2TJcrR9zgb2o3yftgoCXBBKc31yDwBwWjUqcNWYEBb0Yhaia2QsU7Ae7pNiGR8A3+bi
pYRinRbY5C4d4mfHk3eK/aumVPAAZYoEwFPJGx1gno7MNj6x8mAsAlVOPcDT6w8hT9S1Y2D9+Poa
m7Kk2pjGv8Yy8c3Z88G288ieIVu6rSH0HDKWTwRHjeeuxJ49IkAZdA8RhbSoFNAS9KK9o3KXBGcR
qmkFlcZ7iLLYhHNU+rtd+tASKtyi9nWT2w6yI1j2B1NygauyfxdR3Pt1VH83LZJzz9UoyehIzimu
gOSO0zLTzaZQlfv9esGkpe8+0zNUsp6YWovrBa/opreotoTHIaiVZe5cU4OWfi9ScKFJugfLUsxi
QDAWlI5D3vGCie8bZdiXXwSq1TtdiiYalsbWBMzf2vMCQEpmkX4zXInmIHQLqYeCllQgG6aRg34E
Frt4bAc8dKk5hcfP3AQBVuQdgNfQ8zA2WgPJeJubgL+BST+m/wOPTNSS1kMtxjQ9z0wsTtpqnW+l
EaHjdehHQezbAsghZIN5aBk4H0UM60jrFzkm/FdxJq2a5pzQLpGR5FMkB0ebT1uGPENYGQXfDTYk
3HWBdMCHELJun1rbGuI6vKvcbQV1eukIun2ol4bTOuchaMlVcIf4hP7hVSkLiOswaJwKe0nSnJE+
u9BqNGAmuLE68H32SreOA+7214lApa0bWJls4uuQvepzr/LqxytFYzOlmgR+xlzzH5GMSwmrh2kR
MwNrk8aRP6frfcjt/KSKvK67U3HnQ1Kb812q0iEBJiVJ4p5+3cCnqpmsUz082Cqgq5gFrTfCCkfb
5FspvAUlhZiKG31LFPn/rtibS9C0Hyjz0kCxKG5TpCXeKA5moSf20+q1iDmMEKL2TJ/YxIzKo0Yk
VHv/KLtICGHZSUw4METQVw0QeHfe6LnkiYswRgvGNmHKCKB7meRTXSPWaKGqO7cDjIdVMtLrSbXS
wGH/JsMm1dnBzuJtIZI4g7uSCutiBiqw1AopAR/ZxIYkeb2RffsMxJCMA3S62LZqYA4XVtPf0c9M
ARVqXs9oOQIk/o6SnYTv1I9U+kk5R2PXOB/As1MSQqXLSxctrReB3w3f8DKdjEGKt1DcSgL9CAzS
aoFHKFsjT0bHxAntLJP+XHm1HWVQm8XmDubIJi8+7xTkjcYcv8lEyuNhQALdna3eOzj2e4Vnjrai
NMp7YO7hS/aWdpL7G/NIrs6TxIhRZf7Ees+1nkhYvsAUx7TSSgfuarVQdwZ1T8wzMBaPa4l+UbKX
Q6XZUs6rEQBg7YEMl8wikzhq3Zcy/58AsqKGHw5Gg4wN24kL3y3Gk7+VdbZBjbmBC2Y3gwQYWy7b
w76ATeTxDfS/Kl+p5LhR+c2+zWEQHJqJJS4kGNxPXWWY/NHMwEC5k9iTGVPaJXzIp4FhCESmY3HU
8Riurj4cnAHxM5ttp3EiRJQ7fmkLvEliKUahA8B9eWohQq+O/UxLdyZgn2iHxppik8LhPYeONoEh
i6x7t5bP7gYEtkKQufByEwU6LcXIX+ENHfBCX0fiiQe+HCdbKIDswRsj59+d842WdsLw8k8I9Orp
Nl2Q6Tsf1LrquHpYcm4xdy6Rd1qN79P5OVNv830kBT0NMRLILOYt8kx9+CAxzjTaOA/5OrC9q017
zIcJp3SnaQkUP/Nwv49rqCI0K6Bu0kHutouaxN3uwdBZlicRhcWziWwKgwOEWz2AF3U7+zc2ajHY
6R5nrYVE2GDwkcQwrPtsTfY3i3CAXAenlc5eptfRW+7CIiAY8JhGWKF8+XVYuJyuR79tleh0nODM
9oA/N0LNYCYh3X0ecf/JpyT9W7IqK7Zpw7nE/aPd2hemnN09ZWQHRaOCvVFqLkHmzvNFIMlJui3I
XKV5MjyDDrzDwzZEu4O6gkOmX3t6najmtAPjmwbGNTUR5uCKL6S7NJo47VtNlKBhY8S6LW0nUOH0
CIz5qJEhI9bf5F46GlA0hEiMr8sp45w6sU4yM5d0Fm7iKXiMyw+bu3GLrDU7Uh3eiyFFQWdvxdUv
8d8m/mNEPWRYFCBkHwUIqaz2h2Q3sapXkPflFDCLo3QiBI7xj0jPt5cv7t2FaL+J/Vv8A1NpfTB7
FpYtZsNduADK3H9P0EAL4jacB8LzypyyFyUikNs95LSswdP/ZZD8g/+vMU4cyYB4ewLItPoRDgwf
m+4VvBs33wGr5muCm4AXdqnVEwp2q/D4afSlzmeUKz1++X739oG3ZXwb8O6SXFLYYTkBkYlO72FL
3X7nR7rkYFARbB9pqLvZMmFH854OiEdHetBpr+LjVGB2k6NAXjuihviwthwz/8ZBBI32nTeM9w98
Gzissb+wJu8bCuOI0IG44GJVVtn/6npyuN8+VocFRwrjuhewOlWY/d2H8bW/jwBFUApMsNCxxLT/
l/8X1sBHhT96cA5FRZThsSlGkPYby3t53jOvXK81CBeNPbPeYJV2M0RzP7MLsILNu9c2au10oqnl
oXx/eRwNpDrhg09pE+aG6U3pzuvcbX0TrTFNRHvDostQET6l94JPTG8OfumjSFshgDFZIuZb1WbG
3Xaa8Z2+uF+IXOfrC+o6fliS3EJcozTX6ZNOWfoqRg//4oD0dW3ZyvW623K82Czpt+rP3GcEWGjZ
VsVN0+x2eBL/OEchzlafkl2IUaIR/7n9IZBhb+50chr/qmN4xLO9hb0jPka9dGYXkY7HtfZn6GPm
NtsuqzyAwnKVRAuQB2XqFmJ+jcWbYET3fKc7yoTlTFmFWYEfWUoLXDd96MDx4/KKCcBWUELJXNTi
mWX3PsTjv632ZTBB/ofhXZc8kZKsYaEsauYKbRLLd2iA4JVRJgjlwuKhnAF3+zPpBxBnnmlSNqPQ
TPuHVjDB3u5DdpjLHd/m/9BM+dnA4xH1EI6vOewWzoBHUYZBtvKGHgZOy+kfdZw5UcoAbxFYXjLl
mcGBAoEPWktzJjMu7iBEq9uXTNTr38yvaYFV2RJjQfY9Jx1VwI8ayC+qEc8bfy6HgbqGwrS4qCX2
/BDA687Gf0DIiOngcjhNQtgs4nWxsqLjMFcRx8F1uBvfpmRZfJTd0yiiA+l+UdXv5j8HlRK9TS3V
ToT/d+ye/iNPo8Cq717B0b+/CjMEUuaL3s4xQOzLYLHZZd+KmVCz0LNhfgKtoy64v0V+IeiKCTLR
RLj1c9+kxIwh0nNKTfK+8Ycgx7kQp0YikNxiTiivYrzVX8rjYr9pthOIOw7n4FGix00Sn3L9g9oP
hefM2r95DRO23Y6hBshY1kv/qJJjG1qWyGTwysvx7ahU8zYm25juIak923BvMINgAN53dSbwqP3i
HWgJ75G7Q8KZn8hCC70UITu+zbSkT6WtIbPl/IbC34uX+VK0ccM5Am9hjjHx5+iOsWS0T160sQlS
vJ9/lQs5zndxpsyM7nWjoXpkDK0qyXAacylEAvNylCgLFEA+339BgyIWp6U7lKYFZe/9aqsOwX9t
eghDfn842uzgZPsACY9PhGkTVQ2UX5VUNZD7xE7gVpQmskYJ0qDoY+/4OJVaw4jsnvDr+sdM1vc7
yjLU93gwGouxozj62wnehOJT5PkUKy1nVxgbZAk3xgdTdxOUYxcl8LvoOWipKZqgWg7TQgJCIQTn
bue0a8cuzAtAEkEbyieM5d//u4fKjvW+JVz/1nxYtWS3XYdQaMhRC/gV/F2n6NkiookC+NB20eSq
/BtBaxGUPLddSQjZdoWx6jfYW0Phvm4v/64Ut4t1gWHugWIRQsfADZgSJnzIkF0Pf9/qyLgEWIjk
B1JJOKn8HAEacOUDdGV92rg//tl9dCdDcg6eq3PQIM8+Zk1t7LZ8CcGiezzFHrO9wri7GRIFQHZF
vLbkCBoGFWrE/f2WKJ/50Wjgg0zlymqE1v9J40AQJuXdtswjdpKEOtCdB8iYdUo7NmDdxsQueZUD
xxPTgmOhmee2qNyFbooK8p4aezDK2chkXlJrVdgMN7VKM52yW1UOlUggQ5CVXL3rcl52Ct+0QgB6
E6pcTmdGdosf1NFqcI0hn5RXzc7Irs0V90eEyJma8y/ASCHi/HayOPb7mohXhqe7jZZrRhI3lgJo
+XVdsPdZvslXOlMy7XTgq+TiaJMSWAEJeQvjVBFeLFGVYg7lvpXqWsaNlWURPx+Q55wMeQbZfCNj
scxmL6EI4/S8DVtnaELJp2UIzpPc305jzdWJq17Z1kY1M2NqqunsTrrUZ6k075BM5Hh1PWpLkvYT
ok8fxYRGd2T+pP34ESfRXg4ETPUvFY6nVE3LADCPUrHqS1Cwtc91LDibHYYUpMUbv+8qWbRKbcXO
YrUzCCBKtbqYmlOhcl7bHYQz6Ox2Y/yERgSGhsrWKclKxdt/zQ/eJrTMBjUsuPIQq3RAgDgY9g3O
bCmZ8Sd+o5hl15I+lT7lcjuTAsOjOIhAe+A4/DsnbrXOy9637o0ZzA47OC6u0Az54uLEZPycFdEl
3zhVD+zpPpCjkkNgyq3O1dqsRqi7mad1nKEUY92DqgVrFnFwQJzpqoiQlfcFh6UzyGEY8/BxMRE1
xXmqvArAqMzDv6+2pjsPkq2R7kkmPlAI/ek16gYveIM0RTgzdUj68Y10EGSvEZEdn0P92zK+Yr9Z
VNvQ7jHdjtQszTAqBlvtaiylRlQKQyOLS3hgAiYUdIJIaycerishqdxaTv0yK9f4UtDiZwyeT0+q
HsnG7e5V/gj34MRU85jyrm6DDUAhjj0ENfif7lx5m3dy2GLBKGkxnWJXnC96PLsmDzA9gC/fQVD7
BYhULaZinkNBTtMHtvmIpuXu95wn4gJvOEz+U8MXQEg2VsCzUfd1TGGQJqf6jCiyuzVatb+bnvHE
WsFlAz7TKeTYL3EugiNTI/F3i3JyiuHYLN1f3VueczYn30PTCxRxoOjv6Kr8UbJg44QxXQT7PN6q
mZGZLreof1ax8dfULSMqUvl2f/HVjEcJdEyDRbFVaJxJmp60/okQZcPeCj8r0c3sfpGMTrBVYFpM
2gd6eKgvGh21tcy7TPGIA5LIzBWB/FGDHxqGCOSbPVkZW5b8NNmkX7m5jCpRFacJNjOHdSBE6jWi
bObxA7J+ub1KgrS2tBgHs8e0p5YFFR9VnxBNpRU5OqLwvxElKqolzcvB2UeBYpMwZLh5P7ZIlcbV
HMq4GhlOgG5vPi0uUwog6hjTdst4e5G+58UjwzL3GDESoaGCIq+CHG3YC507EybjvKxWQb7WQUa0
E2nA4VgAzmL1QR1rxYp9HR2neyf5EIAbGObpEnXAvjMuUeBimX5JGy9SBJIXDZFZFId4Y57U/W/O
CaH1XipLHSTA+wyh4B3YfJ+yjE1XnUgPg6xXjAHp5WNWcNNcO8lgY/N0RRSSpuUgPG+fahNH+ziE
2OsXkfGZLDVJVbI0STlFBj28NoMZNRR60VAf+6Wmoo9UsTXsobAzG48ksKurEk+tzPey0+M4aIq/
UFRf0G/T50Ua82qrv1GkvL1/0FcynJr2N82Jy9DVF172mvZIRJHH0Hy2sMOtMOjjg9WgL4v+wkcS
CV2vaA4NxeIILgo1mBQkfv+QGDlYmAcVCccIJLr2ozSx0enUDvph1e3YM/fhmyebQUpl3Eb0snhU
Tl9sebaq6FcNzfNKRjV7QQcSxwd2WNpgpDuHqYfFExiHsHpgIRm1PyUhTuCv7osPUvWlDNkD054Y
OiiXL+DfX0zoGPJ4kIRVqiQSlK6Oz8DldLd9Gz7v1rVKC6bq1x7Bmb1YNV7KBXHMfGHlK9hCd/PW
QzlrUBo3un+lDi0U+eQbiPICaQz3QFAfm6x4qZZxJ6UfTOc3UqFu+AyXu6SOVz1sjXtVbIgU25/y
dI0R+VzMbEwxIXUHmeL+KIS8KSgfbATs0McWpBu5W0lV+BPnFgLf3t9CxCajpM6y2Ku3W5IoxKgQ
ktW9WeRxH9UD73XS30xcC+h9peGSSxuGH7sfWo74xO6cK759OOfIAJXKWvqaBdoOMKFabaymsUdP
ZwlgMcPWMInFLVTAb2Ywupv8+lY+msn5cThU0vTXL2yMCLU/VM2jQT0Dy8eQq2lEgT4injHYQLye
cuYVPZqz7dpbY8V/O4KkHU10+o203DB/UZsSoT3bqCiKnLdJFWWL0GQ6hs8k5VgUTTIa1MeJmxT8
nXO9veU1eFJdqfH1OcLSwc2Dik4T0jRp6QB4Ix8fJjcncSHfUbspv4m5VfOD9odPB34kosiIkCUt
OArzD112llJ/H/rauSiCXe2ER07PT5I6MSB1roKPFyGaHOxzgkIUtYc5Wq06frmU7WowrYNVoKBJ
m12TzX13p+lkyRuLwP4vvNAsDLBJmKKRPVyCyp5KWuuD2rk8KJte6Y4/1jexjKqu3Lw3ImzNTxPT
agLaYwac6D96jKSuuo+cj+0f/jVPIU2Esn6fnYl9nOEJIAXdtERfJK35gIk2MuZcDl2lMS5aJGrr
c+qY3CVxkcQUpmKGowDwdDNR7mS7VbMaxnsNOJP+tNbU4/jmYHCh0/pTxNTQQqilsIF0fmC08sAO
22mYxXzLZ8AY3T3JIRe8vt3Sn0EpnC1XkEFxhBlbK/C6xrcfh9ogM8E5t5wPD32eAjbWqM/HOLN1
sSEuhgKiOpP8nlXRuPZYuzUvPln90qZl1toyfQCp69aRjSV2Pf3D9BOqRIGdZGmXsJUt70nw5E9q
J1bmcBq3I5IwqDxARnaPSsMUYHWAJnJ2So+crf+Nx7NAhQetz5GKcQ//jX4iVjHKxIi2KGhRlIeq
0R4JRBIZ2EMmzVVrFsrhzP7fSCxj6+lq+R5KgjdnCP84CNfXXNlWGNqzymG5i7SAOqMrfLjM+725
Q6RInoU4AMUbE3v5BVP+OLm6LNq2vB4tR9fpkymfmI14NXfx80wCIZsl4oDv2v0RYgfqDsZIZUfh
IMYkfnr3t29kOCZ6N2a94nrxCBDwJ+Q5pEtvDJORr5HYSo+oC6ZFsZqZUq/XlTa9ghLq+dvLgeFD
OAOr0/jQRhOWVsgR94CFJ/B374op0Dgz6rML69lzBedS9fMijSRzoPqGtUfehQSunWY6mZeks0vp
qlwy74qP3DNws6B4smEqnB4VeGbEm2cfmjjsDJkWB5L++cGyq4nibx1E/9nMYRVHgNfzOjoIyE/i
KVYEvRayN4ci/GXD2WCydT6cvQeHD4HKQn4kJMqLt4kuk6T/dPl1esHqJgc2gWX7BkYIgwYDJc/D
rT7ZlSlgZylROygWKGqscGW7WZ2lP1A4ryZaILupYO+sm55IKu39nJ2X9V1gRdfGISCSQdDI7uTW
pMaZCCtXJd29/PXWf8rFCTm12ZXVZ2R966mvpu0cybTRPrqxH4Y4lo1rqG+GL6tXdMGUyVBLYnex
XG9XW+s57NQOuAHKoFR+z2kUDZdsuWgzoJfti4qRTbq+MN5eu669CWTNhg6JUojQHaDYRXWe0YaQ
ZDSezevdjI2g9gmMLgQD7FdRs68YTv1LJH46dSwd5K4aPl+hUbhfC7pAtPwuSkiPCPGPiRpqD7/z
Na8dHUefR0xTyTeXB9qr0G7LtAkfj2FGlTz/WG/1FXajVawnd65p94yCIRezwwvszoBA8PaU5vBA
fb75j3LdlADBWks+Znvce/rGKA5eVuAjg4ZXBkBD6jcgiStT1V6f2kNIZmfCotagDixF16jUgj/l
cTtAbxbdDCrZUbOpYYkZT+IzJgoV1l25ia5hGzhQwQmtybMTQdSxozamwblWHCpijmKWUOMkRjnZ
HaoHefXi0IVs3pmPiBaPNq8+gcLzVJB7ugexm4q/0zBmENR61QiEBDy4W7NNESn8s9n25W0WSMyh
y7VSxsuUlZ9CILbj4ovqTzoBV+yuB/5CKbyEUm65AuIZfi9dNBg1KGvXGEMkLasMhfVPK2kIQ94l
IAVIREA+XsfE5WjOsLxj+zDZGbudTEsrteaGQpCqclkVUUbG+/YZn2OXlOi0fDSNN8doMfaomrNV
kxckAm3Ay3+HJpUFA6GqEir2tvCbq76ZPRzfJ+l5prbRd7cNHyFHWQKWQ+2dWKIORFYfxQhT++3d
3jry6dm+C6yPtOkbeMwddxJfCVdr3z1u3Tefp6csT6vwMo2BeJJImFAM+v/rvc+O/A0MOV5MsECW
n/u0KJqlwBeUxLJ/b9LzG/kpf3Pma+n1XbwgYp293pF30sd78yvmE+YQnpWWF1jqWoaITBfjtv6U
S1NijOSBZYKAgVw3n5IVZlzWP6aK9tEXAvUBdlq+xcf4bWjfvoIdfxzeJyMshGkQQ3tr7emK5hOM
QVNYg1jBgKJ21wQWd4MjGxSbR1OfmSIM3I9Pfo3iu6npkdea2EvgiNI7vhQd2nj8fqQ5vMvmTBBx
Mte7GcTfy6j6JUNRY0CUCYbQzlUYjv/TVf3UNQKXFNdSC1iaanasc+YvRpImWjb/nxVmeJSM5ioU
r0OksK0CJosi9CdnW7ALSflOJNK3KtgQ/HGzPpTHgTc6w7DgUynrYNgJo3zmQu/eTU+wsvNz75vV
M4qRzNCn+0BznACV5Bd5n7ogF4Rx7vidpLidLiAYcxTzDq5VWCFPiFUOjankNO8laDEElTgrZ2/0
51T5v7eJCyu+bQWJj700k2wvW2Sxe9Xg/kUeiy+2e88PLHSRpjRkMRrRrnMhTRxf1KTHHjtq1NFV
VZXIhtJy7yu8M7qOAbX1IbJqnnbYFnhzr57roIUjMvsR2lGaH7V+q3Zos7yhyXMHPnj0poEASTAb
mJ4Kj8auSYFFePha2dVI6bCxlZ9TNu5p7BZI8ABOLeF+egQgfImT41RRGL1W/qFAFRvM/KdCFT5P
MFINaFE4OARpvTqzNeNZUbBNs4lD056zf7O1ZBU/gCuwcr1ZeJWqERn82NQ3XBu3hdHC1K+nyPIs
XAP9ZudHTZ0OYopMeOWlWZ0WsqBFYGQJpoCn7XPPiZP4DwmGrAOaKrlegwJz60/z4qWwAwplptMZ
xP2oHwiMRWMSIaIUuGfqQBbqqx7GzXlB656DK7WeCw7/U+nGGd4XA6bErhpllTvzwGZONgbXtX89
DWInzsG/l6Fzc3gN8rw9QQyW7TcVGenL2FtJQD6oWQzHbeM0RFu5xS3iAFgKT6+pRdGzIIHmuMp/
AFlQflknC4unOIX9+OP42fn3Kio/LR3IC3gIymsNd93aqN7KVtbSNcTcvwdt98vA8Ebv6l0N3Sv3
7G7FqaxRMxJSdqsF+dpTN9TW5a3JTcaTkOblyaNWZUl20rNWK51lh9JHSV6jD98dadeIMsgtwZDZ
aA32mfyNIeCbw3r3io1+4P3Yq0JPAtIK7PUENkf0IDhJnYXmoMk64s9rOC5pr5qqpHki/olesUsJ
uAAvdIoR6RmpOZ+dUtkfEVH84XoTA+vgcbug7PebCwjYkJRqjFr6NdiG+fjtAx8ZetWvRRvy1h+a
9t2zxyMysUtmgbR1DeJBuX+X0WjwyBCmRmKEH7MpVykm5U6FIDUaViiAcGUJSDpStTqr3pMhbRx6
1DUTkk/K/6OQg4nOq+D5MLhrIEJge+KbT9M5FJIfMH0O5tZHZjURJxFlIID+eUK8nEccrSB5Fy9Q
SyaFhheeSUeY+/G0OvyT66INVE3DlsBI7QjATuijlhSfGqwL7wH+erxo5P0BfMegADAI26dLt3NG
BjaegrkEXN7jj7TnqbzvQtRDyqLE5KW7/8MzNXbWq+yOYCd8lzNr+RmHJtXiNO4vxEDJbCTfIDO2
JVRXXOvGbRq+K8IGKBFB4gz7Knpt8jdtAeHd5grHGl190LORUHSPKp9OkdaDxYM5BchFaPzSkE0P
iTtZ5YtHI4641quY6M+PDO2Bt/1kci4B0goBKHEe9gCa8WSRjFtLKvQBgip84J0Ats1Nr9uYNb6l
03HgqnRbTV7y+zSQVQDauT4Ox93OVaZm8c2rrZr939zCl79w8pbX9FqNi86NJ8+oouOd97Gz7Ook
pFnNcjjaGfmKKzyfMlxtCElVfUFcc0OSOUfJC72R+05Unj3+x2Sm/ZyFercVCCychrUNJAPuPrmC
ULKaU9/REavXAchUJ+vYm+n7FbKGqqbbpoeXrwlYCwtcmT1oUuZzVoyEcV3MgxHgdgKdY1Z1nCsw
Kil6yABk5JTTQnxOuA/bODbLolBWu59btRoV7SfUrV2oCFIFWuaS6i2pwLq3grdoF5ZI0fqTBYnk
cg6YTKG8fukKAbBwnr4mXN0cEJKrgXbPxPy3fSI9nRxE6p+0gptUUVFJ/tEEY+H+wBDNgKg8XWZW
DeIR4jIBvD+fX4Rnw8a13n8gRlFq3V5WlFT3aiq4z4lD+PFdYF0tCX+ZUtUHjlTOJY3AX06l6Yfl
WUFG/c28p8fwS6AXyy/gp+Wq+o3VJDWrEtrr12DWtrZRkMzrsmALAJbXKER0eebtrIPi19YwKBux
SYNMNQ40BNtrIq2lEXohiQrJAsjdLpNFE91DPr/8u1GCPnWesx2Faoj5dMhKs65rsnrY9MNzTvhi
ovuDDn/X5R/ezjKn4jXXkXY+Hjy76A8uMF4f2knJBhuIY96n07w2oivAhGf0XKuWFff36X8Ffu2s
K56kf4c2TtgYKRDLe7I3+VM7t7rH+Tp93SmHe3+YEozqU5fO6Z8V9pzWbkNQMOL3yGgmCgEX+tlJ
8BbmHbK2kk9e7rEapajXRiuVX0rXz3qF00/MeNb+GmH7mxoASuH92njN6SXbFa/ypu4JoyA1tbcG
lnvq2Gq3zYN3TPLuDBbPN3taIG15j6yE9pEz/4W9MUUWf2fhTJZo49+MEV/ZX8Yky/o33h+fq7JR
OVUhjT/2SRXk1BFXU8daqG/6sOc5TcDmuGPVQ18a4OWrnhtwnyX8X6Fkt2wV0dfCzbvZK5zEGi3b
WC60jZzwlpdOVHhczY45ugH/j4WnXl3pzvGTuqFYFUfJFXwl3UU0pESYsfQXHQYIic/AZ0GAkNrx
9LPMtoXD5bD3vvzR0IF0AzUlk8ZxfCoIZB3zbtDd8jNN+IkMfhnP9B2/8R16MHeUXKoESElNH2Mq
hcxegBGvI5HMyszbwcjQ6Bk7qmto04+Ak8XNukrkYmOZLGwytB5UfAQL9HXdiXNe76URTyVAVy4V
6eBdcPJdqDVIByoX7TcykUn6ji/S5yB8RHTbq5Bqu7L84h3QhMjc+ew2wnpkbrvzHreFrouuy2sD
fZ5646gqg21Q6tXPQwQ45nrXjVbc0LvJd3kuADrXhkV6GDUBDcbuQBJmUvKDqHZhM2VAKsBFwAds
rQa8T99G3epwr1SbeWfS/7GTtme35+/gdUdB7brY8/+crDTd6lEeBABDcKwFPuRXYLxlKqdy53fg
pj6vworG/lzp3QoijI9LurZ2+LuQ0SDwGVJXj9VXwGhuL8BXeyGe9mEvQU46NiW960hu8jfBhK8J
fr/3pwHFXA0E8Kv5R3AJVK4UsgLgA7P86C50c98C22ZbTEA5RsDIZHAYuSLQu8/GJ/pFoG4tnj3B
0i4SSlORgAbTpv9P4PeCLyIRQbyb03J7v7FjOv7bPHyELXjgso5kjX/uPZrvS16VzSdmYXEe+fSk
nHy76HR8Sg1MwgA6gmcq3sVp15bvMNwPThwrdixAjhOqPQhEBbBYR6h6/0e7PXGztKTX1iVCJ+lN
lYcY1YZ+nD1NvAbx/mwmqSwuW0UwRtjzDxtiDkkNkZ9eqPECV9T8+xN0oGzIMY6Fjg7gu+dKc1CX
QKJa89W7XB/pWfCoXtMtJiWd+ibhYO1LkSsiwPl5cnEuq/Iy1NNG1dbQvJli3IL+f5GXobkE7V6g
1GqDMaDPAf0duvJqerQusD3hPZAZFhcg9oXKiDeeZklDw1skyYrOU7Hn8zPi/3+C9aby8oFHDNQt
2LhlxQ51os2YPgjFxxANC5kuttdGtFKkJhwLFH2nj0CHcCXeZn1URYF1N4A0+M/7HI7dGwhHMgD6
pSTIoRL+tWHmc2KCX32wYuSHItahMWGY03X31vcD0zIUt9SexbCr+zgIATXR7RG/Na90lxs6Q0b+
0HuKJfaLTIv5KokTIlr9ls/raAPjeyZeaKSEcAdyBpGX4DsULMc329IkU3+IlJnoYe/gApAcVVx8
0WCCy2nkQPFzbbeiXM8pC2JwUGyj2iwJXsI/LMjXj6JQXP7P+ylB+Euq/OAHkurYP4vWdwUZOysE
STYZByIYjCla2vZmrvwEoOzAxc0O8Vm0r2DjSsPFwF18kIYXFTjAOWk5kemWiMs6VW57C69MO0r/
zik5665FIU/pFFvnJJ/pv/75WdTAzPzkA1FmI+/GhZAiYLWrtLqFau2C3uSViJo9ksmcs41vh5n+
45PhDpxhA2RLk74NOSstCtNhWCLSsOIYu7L4dITVKlSBAZanqRPWVh2wlAYSgETAea3CwZQ3ENjk
5eqJXAY0hs3y++b1J9eYHYTOBDW61euGapczKcqx/rVR2gyh6dcWnG8HQ60DjoESZPqEgfeH7kRl
Z3OBP8C/Hw9CWpoTLCeW7p/riqf6yp3i15PI403aLOHh+4wMYbV0MQK9sWn5vh5hzU/qar+6icqV
9/WRB/Cl/WKWJZ7pUZ/+aGLI9vKiWiitWXxupl2Pc0SBMzdhhkFSF8dhQKK8xOPtEIeGIL0SZuW3
ksd8HJHbjyFR4t9bNF5aIM4AiL2vCvQKdRquwZOLiEJI9Aimnka0sutAACVwRBrnwMcb55iCQpzP
IayqA2BikvPlcWwIzjW3WJZoVzxw8TyDd9Att8pZnxVdPbSmYMCj7gizcXzIpIVI94XPHfDSD2Hl
bFRXx6eeXs99a3zwIJ+3LhcViJVWPzkxKi8WnIkNqlB2J5bMxkNE8XpujiPRRV21XTs2wwgL77Ps
1pDLGH2gZ8yWeF/a2zZjcq2LWfTF2620eXdaAKtsTa/M8qZJeA+q1E95QR7WWW1sUTLOGg5o9lGT
b2SEhnIckiRjDfQ+bjM35ETfFPov58r0UUKl/gHar8WrcJL0yfWsBFAVssGXMl/nBLQwsL/OKw2s
pq7eP/cs5FyalT4liPZdAAl+tVRnCTV2+8KA86oVOL2p22ttCZqyS08r/OhkVYLg2Ow+roGbsGoy
67uY7UvtpGe/2DmScTKjAgizJTtvtZGkxRQahyZ+LhK7QhJyplTqJgNJ/PqYbl5Z6fmNVKKhEd99
xawz7uQlFEzk0/UC1cjMujggyzGN6sfv3aktsFZ1JoqoDq2Dvo/CrAfvKVcK/gBcu14tyaWCJuVb
fQ8tKlfsXHRoOL0HIp3+qwYyXy71LaMQqEfwQts27IUzTBiMan3GYSEOnmpGT9T8J1wLGZ8r0HsJ
WOO39qvl0n/2XHlrGY80SHvx/+lKzH6DuoyfAQl/Ap1ITXegwHm0603VMMtXH8SMK5tLMW/eLQG2
YFbNaHmt8xdKlLG8u7o1SBXgPXYTTaO5pBY0SLjbYY5fb6WF+OTNh5k8AkBwvuiGloyfR7akwwcH
x/QrJcl/cCUG6aX4iY9jV0F1aYdZSQadhm7ZWqXubQ9vvGvWbhc5GgJK+IRSooTbjWecTcOeQ8Zf
OLZLmQw/qw8v8ps2uIcrtK7vMzLp3vguBL5WWf5Gnd2m+iaIVNCO94xg8ymPiczLcKlA4lzyY9Li
Tkv043s93TnWCUbhiPGoIKMCOknEZM46sB/pj50CpYBfDeNCb0FWq6loDTERUWofflMUjqNIT3uu
8mhSc3nqq2rBoZnNaopy7AURFSGOCXzsG/vtNveIH7tRUv5oa0NDn2FRLayKBLbGVa7GY67ecYwn
UHkDAxKc+X52isjIMBWBC23ZiRH9gNSu+h6LjJkicW5PG80JUhxalGgijMt/SbxVH/ARjMOU+bxh
fnduMSElRjc5GHIx6DJERb9GcjxOffEFnjnj4zKz49oOQ5ngfv6JVwGSlzoAMGGN3BdILsevulZT
WIZd7uVyWjBlsITt/65sBF/6sYnxRx9qWPti1EeIrg+qoEMMA37B3HX3x28kpUJc/JNbVUUtMcA3
iRWAWdSANTXJM/TE+z0/1ojEWMuCBcpKwmfHRn8T+P/0XP7eD755+hlOjiVyhat/Ny8MZumELlQY
fyPSEACTzBb2negrnJoEMetzKnxEjIMC5ZiETvL8d4Nztlt+CGMKZjj6o2Y8PeeBA3dWVQfKcHI5
pMCecJV1XiCRdWAW2a/T/rtxMMa72QfylC07QwxUcpLyUeqVYlUldgmsvA9Y7AbbNIdefSrc6Rqp
skDe4BuVSCDt7bx+/JbBhV3DVhOdH/Dp23EOXS1bcFgiE3tuxWX+Y5O3wAQooHAgN9kLu7IY32mW
uDtM0QAXGD4VOCO471/ge8H3vJcgBK9J9fYRG7fAX1+xm+SrPzi8W+2kJNTuNPYvL+v9IwipqyV7
TZNoVN49+2n/BMnM9tMmm7hzTOMu+JcL67wYGwukqsLgRXckPT+PZl7jDuFx2a6eNUaVeXFxcKqd
tXR+Vg+owcUKHzG/1QohUsd7vpE1Whu4LxOWLRUb5DwEMlNN66biJsa0EbvEaN9h20/QxxwEJQNU
5jpzlNg+dOD3nEsyutLtTrpYKfYjHpZqAnTnloyn4bYi1LSvzaKZW6PxtwrkSWAPdDeL5d9jVV5+
xbRT3yzch66xPTTZobtwJhVx3xY/To8NeJ4XQgc/ex3T8TrExKJYJdrolbLcqcz4a2oJcb6LWBvq
rg06LTPAu9XtVMfGlg2sfHSBLA5DeLTTqhB++btbABAJQyVc/K1dANT49jPBZ6WIZ7WciBgl6uSq
TbkshexRL52CjB8sjqPOm+M/cs4ZfqsBtk9R+d5Y4pJd2jhwgi+2I630wRyu5+zT5LkIXjWiFAHb
PJ7aMv91gtiWRsc1+MtM6R5SSt/wlS3pXnVM4rL0c+N8YiQVrM7eTtfMAJI1rjNg8F4TTu8yzEwm
SCeHZln+kb2rpxiRGj4Sm3/zRzxHZrkVUUMBnmXIxl6rofixmgBelcWOYdeW1ajPuFlAxdD49/k7
1QwiGZdFx8uzSWOLK+n1c8mRf93G3Kp6gBnDcTyh/apHTm1NfL+ReUjSTs5Rq9dvY1YtwIKaBE3/
1N+jdtzb9mgmkyMo1JnU9onsHYdDAdjFWcKsOzuV3Z551klSLz/JVERHXxWlmsq2k0nZyBKGyzJS
e5sjBtogwvEjokGbNubvzXH6LhcZoFG+B7C8E3P0scDyOs+IBPSZt0+RpfRw595nsjj6UwBsr9B6
kGAAoFQfEZyMZp0NIxScCUxgpDhINKrs5DiGVs6bRUchg5xnERLi0N7NcksDAAmTBlEwAjaBD1xH
RtpoFZoJ3bkA3+KZ3OyJBC6aVb/aJW2rgKGaQ3VFWXjUjY8ohaVS4q488lgIIyhzBE1zQYPEwbTk
yR5GydtPmoriZnRUByYL5OAcK+5ojQW19vyW5KAezCQ8mXEzNWG48VBmvNxh9rFkuZ+h6esRmYRR
JNPCxrWompX9K/xSws1WwFG7oNiAOfBCtWVt6uqYfpuZ4rcUpmE2vn5BUTzn9nc90aqzadFgRCi+
v5gAAWMFL9MSgs+0Mh0CWPxLsjrfhhanx8eNcxlnPQprgqnvM8srUiQQAbDbdOfpsUGcOfwMF5ww
T8YyWJ8NjJAaEeMOx871DzXa7XMse71KZc7yHsYud/MA21ZxOlePQosknweOqdy36x1+C8qKAp7f
gRfaEssg6Xk0239JmIAKWyWCTcXTSjlgvTAa9wkwYFGz+ulsBLgB8VKQJiWAdeN3k4IMdK1yEOYY
J9fODq+g8HA+Aa8lvef9ybydGoKFVYBjMhnp37bB43AvS5N3fBvF9wGPFDhjDInhTTRXceqfKh19
oTOU+0Egrq8YdQi3HkFdIFuojkj7x+LiCbzl7a5FSXixvGVCvp7CqrR4jkral5hfMPQxhHRdqT8d
VIHFN45ox2DDVyTrnnNjM5nxhe6QW7Wt5D0dqVT9BITdOsfEJPuBp47xPTtQ30W12iSGaxHj1Lk/
Vow3MLp2NXorwURtSDwGcGHmz0Js74tQ1nxWsU2fk56x5ahLYlIAVjglB0woicgqVwODmpIXuwCh
7l+Oad/ycVCv95ncZZXWtAabv7GSRtWYxgJ1bUgaN8DPcngOdhsCQEJGkf3R8djTOpD/aoWY0Dnn
76f4REjD9OSuNiaCbfRDHCmczQgduyI93fexoKaoJV79tgdaD/hc4DcVrMMf3EyIYcgF78Z7o13D
U9zqRQmArsQijvL69lzU2KwpkvAHsDSMsANxaMRj6o8eWOy/jE424HI3sEjlkr0ID0D2C7pQXKx9
QsoKVgz+cmcmgHku4sCHrtFMqid/J/UUiLlP4r1gfCpuTn8MU/w/WIzESrzc2AkoSRJyUv3nyXrg
iYMJ80igQTk68c1cWCmyl3y9gVKtewRKJesgIfprfmOMCHJP39eNovVHLMLXxwwGyvr+1FiyV6ur
1WXedLFOSxuGw/XY57TRGIK61qumiIrqUFEkXRfcE9SgScUVy12w0AEa4wqd5miFasAloPlnYYXl
BUmz4Az3dF/EJFCtH0tIekBz4WfJQhZuMCTfK4nKwwCXTXwvSyeQn7yaldsr6N7GfYJ8AtmLX/Jj
TwyHM6jNc+HQ9OzhCjBcf8YtGrPxV4KgKF9ZwOuRZGa2nTFtlmkf1YLTZObhTt+hU57ZFVyJpf7g
W9ZTIJ7DcJ0gQC/RVApyRYKjAwxxm0Ol4rFBH1bWyPxxhc/dzyRm/LSbxCH5/Pf0Utsyh/LpJ5iH
HBvHwcdwhGtFTIvT7hVdfyQHlPYbOlpGGyZV4Ml/8KMgXkaE86u9ZHlLxlVMoBEqluU/o9gmMUht
yqYvSzSDkw6ysMVPWBtby8y0lEFEJCMIyxhYf2+vNS1Sg3+JVEekguEwVoGRwei7TSrJ35HsU5TK
L8jc1k26iZIwcRbu0moEIEXjri8EskwysctzAkm3N1nivxeLW0siVMUPaonRLk37wyglwQwc2smi
Kls4oRjwLJFcqcbcQOSZRbCm/0QJ78CwX3GSEUadg5P7lNzowTGQlV2eiLynWSluzXDBU6gFAH8A
eM5VrJqdu1Grxf0p521WGes5qOE1e6tZ5FyYQo2986QRGgw32SeNJumpHW/13nDUWgdBC5FdIj8g
tY4d78TfezumLyLmQfWpa77yOzrVNPQJFnJjhvYtDlk2EFFfOcFI6TSyhYnqIlnjHJj8LB+5BCbZ
4XtbVLCROSwNqAL6HEYqACJdlnHRDApy37faBZRP7oB3xBNgRatd/f/3LeWoXakcYL+wx79Q7BF8
+6RT01NlLl43bIaOFstMhRcIqfFf15m4JXseUutKOL6eoWwSnQOmzWQvRXDmkTmGSCnBQv+xyoyJ
RYDVaAQhRzy1eb00VoJk6wMcFerOviwecc0M6mCEKV+6Qir/QbxbN+esamOu0H7ZEjy4wng6vH8g
Aiq1PAgckMEDCVdv2tpaDVkcONmct4KMu1JcOZzbdcE+tOH3lNCZjEFYbg243VrsuxTxRD2HaeFB
D9JcT3U94XFTsART5XQSjv6cml1Rv6ltejVU1qyKvCoaWyKBEZW5pCw/EeM7u7JZ8XNajKrEBcOu
M1r7Vt9EmnB/S08CmRcMmRSBbEEiKnI0e4h6jtLxYGsGbuYfgxZz7oDO9GUnrtN+JJnG5RO6TtQm
j2dAKUCroEATprC/HNrA/P9XiRFBZCTWxdAdlli/BHg2jxGHT5xW+mW9e6cLrgfl4QmoB1j/OwaE
O3L745nS5PA71+hG9LsULKHOC5Sa9oeKVmO/OHJJwv/XvdINdvZd688y3cbaHt9F1VGUusgOTU8Z
B+ds+pYSbbQzQa0jT7vobsWctyptrCPgg4WJKcQfHqB9lu5FLjscvnJMp9+8ia8PZpMLC/JKyaZq
9FXfFNTOnz8Mtyszcwk1eAfzksWBNgws4lENvYoavkKqIDEJsM4SL7AT3hvN/GdauxR2+/WMIa8w
Ok1IY6mq4uRncXeeIPveaLc3BcE7mMCkgfidrzc572bqBMQxUmpZFtf+R9L9oj9UAUQIcfjMa+ED
l2yXZrRgHx6JYZLNobZrW6rovHhfSEMlK8EyFOSTyZc2m9aVkzRu2ywlPgv4s/Fva7swi7QeUZbm
UtU+eQNmArH5nIr8qDfh8KpnzfnQyGUhBgF/l1WIThDsuwDIoTpCdSa4+5qEXIB/+yO6NdKS004B
CBO3awqJkv9vUXNJAs1ZOMcL/QU+aHhxINc02LzBO+6leOOoQsXeWJZPdKUH40H4EIqB2YgBKTA9
XcAyuxjxTrg0+LBtkuP+hRuHAjMA6DZt5UE1qAdLm9vgqMnAwcts/OwawX+SO4ryLjxjbxB8Z78B
aqr//zvY7FYw+vJ22Zm7/E2u210yZr9hbB6a30FoMo9nFDDYxoumA1cOXJoUWeDWbXIdzmGc7Z5H
Lxxd2cu0/dCRN6LWKC5Qp0cOyLrb7W2VZr86heW1OBui7jTpicmqfObR5kotz6Q+H962IHvtbarZ
ipjIU88VslAjn3aWMWMyn7gZSxfUUWDrWmhfimL/lHKcwjR/8gYvaV7wzkFrnye2WDFBcub2wKTY
esMAdbfpiWlTF+M9/G0fu+BtBC41FNnwrFjo98ZAXK9Zhu5MhN6HwtsEOYYOOPLhj2JUYLCnn5GJ
/AIryrAnMzgUBVnUDk4eVhNvZifHDWyANhoGokyPj/D5BAyu/Xk46ZXsHVCkICf9qoHFLFABJoom
qrApcJwqIa3ay/XTNoDWNYitZit4kzJ0CNkB4XITz2TIlqcZVUuJATCp+Os8ZUpJpGiZu0dnP6sT
u6l8WyguHn93HQIMTb7AnKgD3yl6kMbBkctR0AfWk89iDyQKRAVp0iaDefn+Oxii234ILMng12jE
OKbTiYuySaBU9Xnp3DH+Oq+2/yVxrbv04h4GeZwtV7RHtoaj6DcQtt24MmySZAJoKqlc3BneQQ08
MfM8pWLq/uqcsi3pbUgyOGEfY4y+Kl+BvjS7K+iX1aid9aBNCnt83kL5NMLpmHrJFQu6k9KV2ulJ
Eim1KYmwIBr5amdCq40CXHoIUCrQXE9810D0KH/pULM9ipcNb5j7Xgpw/ps79k9Pibznl4JbOOtW
25Y64MHXy34qvViF2gzDdl/JxOWuMyhrJeEn02r9vAoHH9ILNPk1O2UA6CSiWDOacOhjUNtLCKDp
HernIsPtBWKdjCaTAIDjMnLQRQnw85BVh4f8N7AqrNCV0ympz3G6DbtsQ/0IJ1G2cVE4JIRW4gD8
3Jhs5bKsNds9Ki4LNxHAAgaoiSJZrTI6mR6XZcwO1DMm9VY950N6FM8uru4adJLw3FzCYoLfkU0X
jp/PLJ2uMp8SOJZcT8n5ynoRqRY5m3q9kt1pUfEiWlNGCpvg1k5jTtt7BfWJOUhKYta0b/T688YA
e+mJDLfbuaiISyT/rsK7NsAksp9NaCl02ZYBOTMAGH104dkzQMzarB+IzmZtJD0dHwUG/yWMvntI
WVeD956ED6z10mnoUWjAj2+dpt7fYRR1V2Pc8AXWBXWw09XmGRxUjb+HMUgN0AF6/6DZofXUHHKM
JjuK7jYgcFuWqyKtrXab8r46h0+ZyUnwl6ZkzkU2bpUQ2qUUmJzITxG4qWQ/NRWdXGvWnzucydEk
6f4fT8jQ6R8F0YzeG7zXkA/6jgRbMK3XUqRhbQgSZ3rDgNQWIfEN/Zd0h1yYBitOh5W++BBuK3n7
toEv74SavjhGMMTJ+wT+PVJv3XtJizdM9cgLhB1/3ewY4ufNxQoiqauNVfpS9S+yfwTwKtmuaynt
VPUa5x1CaYINoGaDY4ButBCJKpX1WIrx6UuMucDeQ3/PCBXxuxO1zBIWZPZU54O/W3MqLPNQRtta
SOTir8KMvyP/C/q9bXtMWepwcOLJr8eAo20G1N+Zh45JHjDyVO3fQeBKJ8D1HZ9AGMeObRCMTeGS
q1Y7L0eeVYG3yDHiTifXBxe3BR5zWUwn/JW5xQjEtEdB0+0ek4MUrGhXjGq55G9meIwUl4xUmJBY
fH64HDriv4v7BlUywOTojrLVI4sDw2hctcnvfiipU9DOAewEyfOLvlG7mj/aXX2BbD2Pl4d3sOfM
D6tQWfkRmG+zvAqxUMEiffbhCNYGU7Gkzc2ZVStbjYJIW0vpAIDbIU89HR+kPJJ4XfVBU/fbuF8n
sTfyufQZemc9P/MaLQr9valhWQPdtu7asxeUjxXRf7qGQ8W2KuMw08l1Nlbje2EMBEB8HPsmtjYQ
yuGCp2gXwKOqAJPL+ytTuuFR6i+gLdDEkp/xhExo9c94fQKAMfN+mGP89KDuqqJV4JnYc9/eRSEN
VZr9ZWppeVzbdtKK4DTdRXdbu3Ybu6uw0RDptDZCgugr5r0SLWr0/UByF3JnYvlRuhoQUMzavJVg
vTsOPDFyXz8955+yzaPLLjPHu8yKO1/PtIayEoIu1S5K9q0Xc4zaBCaQNAt2Aam+Ead+OE2sKELH
8AA8mKCMuBB3E8JQpjUH6qMNddH3DZ6skgonQYH3ByWnyma3BvvN4pt1PUxbmtOZUKZhCkPQyhGg
QRV2GV62yhenk+v8PcfGWPEtg2X/FtvVv/o2EjrpTVItsJg+/xookxlZTtW2AHnp0zZWLlo17vC3
HLLU3Ae8z0OCYBGr67Fw4PpY0cgUFulGJnfswvGMrnWJzsiBLrI8OJG8pLqZQ5Tj9Rfj1fpSj5jm
EIEQ4M6fTGlqlAsivgcBohHApNalP8EymD829xAjB3uHcXI7fMtH9Y44I7tFMwtg7UvNNuxE8xmi
pujNlofTvArBU6Cz8Jp7hMipm0cDsQH2PfARSJEhyzfO2rpM2erlle+pTNcvErc6Yr3+tiblhbXX
QXWJRTNyRnLtOBqTmOOsx977x+duR4QI/dfN2HT8fSaQGoCJhfg1ltC41Z6fPGuxEjTf3CWyF1d0
9L1KIvKlHEDsGkieo7CEOJJlL12cLz01U2Sv2jQ1rdixA2k8grWY+ALDUVPhLWBtv9/IgpMGR/aq
Qlix2T5SUX2+gN3UDchXfHV1/Lm6vvrIAzdDw7iAGieIgIiF70H2FrnR55Hsj3fS/q8aUqD9qXmw
xJ/BwmC9PY8WD9fhJ9jobyizS2yAof6XrRcFdFODnKRvusNoEfvi94jCS9FBvrfW2+D7grUVwCUE
QH0DNk7eTBJUdQAA1oIPFcb2qEy1tQw9QBD30R2gFEFED6zYS7fHdFq6ROepXcgxPy71gBc8/cdO
9n1Fl8igaGjth3s/NhI9gihmT+PszbtrQxfFz1D7KhKlG8x08Q7WopEnIoGuq7/0qgMgliutacjd
/kDNy8XbiQ+qNjcDn8hsuBk5ODveNs0QS1X3xILLz5n7LRC14a3MbG4eCH9VDDx6WIJpAZukiGA3
YsMMn6iSSvINDkSTrCMld9WenEwNEVh274wmnaA44n1L197qrOLg8b2KU0pw/4FORbwJeoB7kdVA
A8nPs+SnDVysC1Ei/BkoHofwcU/2p0axMZZdBiUlOtl4FzkvvYLFHVsPmmUIDIZZXViXti+QX13d
2DR3TAKcIHGItFSwYl2cGmO7BFaHKH73CLUEkw/2bCXp7o7+mSCP5sEobTHS3R5vtSTcSzgpyWka
jc3dBkqeUPFIyOmpgneDE2zSMabjEAh6moLn6y3guboVWVLNNivsEDens3HHQrt7B8N3Tc1UP4sq
2fm/cEbb5H3e9Cq7chUg2huc+zlKUl+Tm4Z3FqpVhsmRX5voNrZg8RanblDqFJIM7ASfZykuy65r
LTNP6rcUmBQVn1j9fkxeBi/KyQYXJNGg9RDM6QzCM2FLavaHVT2VRgIVYiRtkGj6fLVtBXS8PWGd
y7zE/5zcvPKclbx0fpISioAeQ22koyx2iPPqC2XDVBQj/WLj0hH2mq79QUKN8F7GKMSFhFPZbGzn
lO6bN1nd5i0TP8OiyzqZsM5UYuHx3ziuRx/RR8jfrBH8njq3twEMskxONiL3YXOKdg29NxtvfzFb
RsaNgOlwrohwXD3Twq1y5A1f07AxsKoNQAfH+mlYiLT/cNgKYnqHvI1gIgQgr9+CgQj6GsBApZvP
BNaKU4yssGP2ZZtK+Wu29N7IqZ4oR41O21cemERlmBS6rce2fiatzsFYAEgnNzYS4N9rbXsYr8pe
jGFMyv1ur07Hrv6rNma53PmUqo9/WRy3iSp+7VLXfJRmN2xSnRZiFeT1PSc6T80oN3wgQHWEg4iE
zT0Ah5GwtY/O/02yG9tZC1ThybJxkLXZNYj1Jz1+xh7SEm/RIzORxM4wMQC0luTfY+F8xuNxtFcq
PuDi08szGuHZh/dYmxvZ/dBT6psho59QYZ5rziVxnBrbgHKUjtHyvtWbX7D9XautSjJzhjbZ/KZn
/dOqm6fnbUOC9ca2DAvA5RU7eBeQ3hSuaQTUO7FJiqB0dSAsWIrsnPO/uCdk8W754luFk7Fu4iG2
rvAr8MAhlCzJP8N5qO7OabPuw20EQpFjnrUfMrUTHnL4UTNi0dUc4NhMPHCCIklqU/Bkov+o6A+e
FDXlux/nskOULvK3zj+Y9JUjhxWWGaaAkgM3VggVjY4lMUf8ie+fsCO0KbWdgWBD68tdJhB3hNEk
anUEEpT3LOk86aRQmmLyrOy3POq3PI39q8VHSn49/2HryCl/kW2PNIMgu3HIGAbLeVyfx8Tpa4nv
6z8LtUVnbX6KhaaqPP9vmPn5UhYBmkAsgwdg/z6UlDPpXqL1TK76km8Vm+ksE1/GkbtqIzHw6R9N
QwJhVmJNesixLdsQndtJ3rCv5FXLqtvnFKF70toKrWnqcaXPkWU25nP98lMlxSjyNofBbdb08kg7
wtEmO1xKTvZC36njVstRQXi5DSRwTTnHt7KV/mXF0CZHg7aNYx1YT87v550vaVqduWm+TfPaqGQY
fW0veV5c3eItljBL69w2mVEHTHfKwq5S/nYb2nM4kbR0hdPGKvI0pYP35Syk49Ys1wfC1rs4/g7Z
TOKCaz+A0XHetKu3FdDbKLvrfsLvs3oY+7e1jCKWQgL7a0B138ob+v5KJMq7+C0witB5rLvdmBmo
9xnXW4pd/uwXl/HYchY9aE6b1Dvxcu4z9lsGwvmI8h+xTS5D4wCDxgBBvu/EcKsL16nVaPa6dyqD
UkVJe0bIpzx8RMvljT6Tiss8TkcLWKXjEZ2ZiXJWxSlvzbcFHQys/c/E5XoByuubuCITb4JJrJgP
pppJopQG0rMotEtqbjmlMLgnShnyAtQg9ieXT+aRahyYQRy4tDUwFGYzlnZ9b4uS/snFOnlQ9OmP
Kq6bC4dBrqlxMOU58/8w8/K9zEZk39ZtgLmxOOwIdxsydovyQ2JQHahM74UPxAhetmZpHncjdl0c
h5lgTO7OIslhw5JQnIz7h+ZDQxIPde6Y9cAdYQgiHoRM0iDsD3DjlmfUTpK3S3N3UTvJufGVmm4b
11r/Ue+XJUWPEPlCjz2hW0r6OftHxTIxjVtr9gfG4fY7+8LpJhwSWtKJNrDXl5ZfB5i3SaT22JDa
wJ5XCzBg9GfAha0l8uFizOqowxklRaep3dDSTsNzF8PAdW+xrQm7w2pkl5lk9xehFqlWW2eqzt6H
CkUqzVLVYIwFuwHQKQ1Ud0Spd3w2giE56A2WR1vUvMEcizEhrdLlbyac7dR4cSgP9no44wQcOttm
2biDdmPdooTMPn5iuvEGB52irK7XQ550ALifUz8RquloURo+nbl10JCCv/i/zt20aw8qVrZUZuNd
5Sok5Toa6ac6r8VbmVz+q3ZMCoIUc2nVuoTZAgKufANdwDDdZ6lvLUITR0TxoZLn22MdXdK4rdBX
2mywMofzyMtlo02kkWW7UptS/KMYw5ooH4VfJMIhNbyrA4El2mKfyHUhnrlD7S7bDNqmKIs5IghL
tq3wIvF/z3+n77Eit9//5NPwiaHIelkxy3w3cK0cuMiGSmtSueYmnh93iIIEDul3HiT2Y5CM4v9E
kia0kKu6tuGRnhTl1rciPPgUVz8GAUWA3zR0CLptEHb6dV3CfcmFOapIx1OncjQH1sG9miIp6EGJ
fTJx2a1JNi3NLXQ6uyIF3Br5UG1zchHXEg9gc9JXF2DiwwHCvkMFWXK6fUIHZO2y14Y0c2Gb1HHB
AS0ScnZpXRQeYlPEo31vAp9RsSdagpfg2yhaTrNC1uFMcVfYqIZ5RsCEJmQa57WtAaKt+zMqV8UN
DqijkQ4U2QDe2upqP8/XOvAvjrf0GnIPJ3O0AA9pIxC2ai9jtY3OT4FTLLSYCcJN7T8WFYQqS0Pv
tYbC41c7X9aD9aHPRm/vMgea4NiGxoBckgZeg98R6G6zMRKdHjITalhCpsULfdbxtpkEofMQ4onV
TXb6yWHSiVh/d7AdoI2PUU5NJff6MGvbpiffW6EhZIKmBxxJkuRwg/sbeFbeunoLCJj5rxBLrGzU
dIu7Zoqs++9Ogx8Qbyk05FgJ6edFdTebSM83xzu5kUSTNok51vIYkJNzok6+9VwFQ8rMyjOSZSMe
4WdW8GIY2jdxmemRDdRNkw3V9e/XhdK2oqFj0f5+sZZWReYzHOFxzkvshL2DEnn1Hdv8C/h+Avfs
vGpX/eTvM30n1ONpo9d5ZWsZ/gqYtp6HYNNlq40cERQzH9Pi4AQqr38kWevRb9WR2UhlgfrPaupB
WjNYdz3Qu+DGa9whAxq4HpgE6Tr7+jbB8pHn88Z8cv7TibtwowZya3gDEYw93XkSg0noy2N7o3k/
0kCY4eDLIzioHHYVU1UO+el9zRBkKh571G3drpCqmqPF/BZbi48MO/vXTXeDdZNopNbWINMDJ0hG
X6VEZsOanEeqNYq3uoVbQchm9XhUdIfvvd45RkVQQZlIE2/Wa6LlS8Kot/50EZGpZ9MHeNsQUVWa
frKrkLYm4PVi6Fjr8r5F2xqUA2zO189N3E6Dn+wpSd1lKORooNsFJngyj8DUKM3/gvq+hDIBC6bO
aw/6YYnKDxSTjKQz5/mOgfMJKpszojYppLGmQo4h8HTAPoYVwtELDWmQHpW5roUQ5RudbOyaX3ed
23O6IAhY+kRy2EQaUJQR6mIsLzRpwxW+8/MIWRwxBeOh76hXXbP6wV+o24SeZ376VVHsll5tBpKZ
5Szm7IlbK2FOnNSRHNpEsbOlFh086Lf0yF8wGMf+n/X4RAn5RaYNW3hAnqBvO8A8pXhLDUk5ug95
iz8FdtA4ZiHcgwlCuFkO8bhuwaWRk8MfavV14omjggGsaJi/m0JoX0gulxWmkpTp8/38MPyTy4tI
G7i3JaHsJodpG+HDGiboCYqF0hKgtav6Se7kqzahvLE45jPKnM4b1FYmOtA0uSEsFsIHig9lVahN
HU7rmFK1rAOVSxM8eXSRbJ2ccxI5D7PFz0OtISD4NrUj8Q81Ad9/xNBGbraNstctzYNodZCfyXLS
zd5G0fRcForxorSzKMb7kl65GzuNzi397A6H5/z8FY/0L/ZZW1AdA8p/izUu53bPI9kvx5GmnSvI
VxN2w2IgJ+bJSipqqTmlWbEA20WhCs2HoY4NtLJhcb7P7pfFg44b69BniHlj6AX/SPfQOWbBg3EH
1OSws1Ay6APnw5yhpVupF/bquhI7QetYsppAhqVLY9VwOu3Fhy4YYKMcbcXjfSkSeC+EK/bBgYYT
CSNhgFWrx9UMhJ3mGWoUM+jEbzJRAZ7gC7VwsZZLzjN4uRTPY4h5q7IjpH6X0ljTt1/VkOY3LoL8
Yt85OqZ6k8N3y1AFS/d7kBqpDD8Hi4lho+8Bs989OXDG4EqUn/Boi7pzmg9pPpTwoB9Ntkt466LN
wBL2ukQDANVLmtrK9mWPYoiWfp5zJcOYfilt7zWJruFal9hgAUdAzbpwaJKfeChtWbOfuhr/b3aV
wWFngp9xnim/l1WOfGGoC8tZKWy1gh4SJRmjB7i96lBzKkVUS1B1IP3ouLYHwbvUIsN77x0Dpr1N
7Q79yrLJ0VxISVQU8VB1oElpV3c8ZvGl0Ld1CumfYdysV4CsJlpj6dNLh0FNoftfljq/AMQLwHaz
iGPYt7abCZ2MdOYIza948xe893xxjN0lE38zDV5m1jhcK+QTf9vzhVOq1TwctjdC+GyXhMGqEFGQ
YzQbV8pcwZVbNz//k2zEUBaSWAzoRKszNkqNXNx3aapATvdqS+dyNy4INUlQCeABgC6brEkkPEfS
t/pKKjdJVGmGfEBZe49ejdeCxSwfWFGK6GUBg+7W2ne4HonUii9GLHWD0eYkCKciuSb6pnVoIFm7
exXIM564gqIO0FCIcGCmrfpm6rRitvHSB4ASJuxmMVDNHR+R2Mt9wKDBhiNZE7BTECT4QWh7GPa6
K5Glvp49rFD5/dihRdgwcn5DU6JbP1tX37B5A7GdnyYhkNkEPxWjCm/J8z5cRKONT3rv5xxh+Anx
HMEl/EK/7DULBKC5tZBZtVpJdhgNz/g460LQSWhfPtmp6cLtdrYRD3EWzdc8AiqVycNTiF5eOFzu
dvvVWXucEEYp8dbmehXsld+s2cVa9niJ88dD84y3vayZXh23pXKwjJHN8kHTBVtrZGyHvXCglws7
7FbhfJKF57gkb3cevI0Is806dDAxHHEacu+IadXr5JwsRWRbGs9jtr6HXyK3gvNedjmbAwN4aiUO
1N7d/+4k2qNt5WX4UMZlxCsIaTi1hLJ2T5KFPThZVM9gtVnwCICiwvuP5ydHmGyFCLoELO5Y/kiF
yO6rAfTUJenkl1cwIuBZPuyi1ZpaIDZnTR11hEm83sXzAZ25ZPJ44iz3X/hwoKBlAHIzy6Fr0JDY
x2fXmWYmzZ/bODL7okmCWFe3Lcy6e+clixRVy/SUC2SK9Qmz3bBl0Yofn5bwjfz+hUnivOgCfQGb
UYyYqeKFXnsr/1SzynXdL/7stmJ8zjCgpdwRlUopch3IJIQjWIEreiEGx1eUdqN+7LMZlLWbqDwb
7BweLxzu/dnx8TBVBGlGMt+rhkhyPTzAyD3+O5NWB89tLROH7Ryx3qFNsKbLuqbP8yQlFb02Aecn
J8mnX8idLQH5toTeipooYiwmHlbt3go+V+3+gbs1KUXfbWNGJsZA5LNAIUuMAUs0/lvOSXvhJ1+P
vPWUl7uFgFESVa07iTuj7j506scmBFEaeciR9wO9qC6hJ+2RezoZYxyUT2zu0/cirOgMvUOAE7p4
UktXDpgdQaGTc+5vQyj/5luIFT/MInvjJHe/RqIzMqZIaGWEaJSOnoNhVq4eQY2P+ouBaP9OxVQG
yY44W0Mbk3AHM9TrIhO1P3a/Ilrbi/UT/BYWi/2etUPWveJ+S4n8V4N/5BnjymPUHoPO0VSmTG0d
N1uMluGW2HBptXbVnJnRZia8fEZY21y3uW4lhiTAkCAEkM5xTwNpwPhwZBUFBfmb96mZE+xIIwUB
LYIY0+a05t06jJj3iM1tSCbFeVia7lVtQHUFAMJLRzeJ9DO3HAX3GvwxyLHPQU3hItAkGBdJlAgb
Cfd3FaV25ifG4IEMku5qOPatXanPadUPcL6FPYdYCaro13qdyZR6E6vlE+13meFh9CHghGuDV/bC
rguYXEhiAmzMDD/80nGXQA1zENm3L+ivQy+19U8snOMObKz6ykjgqjBymj5yu1u0CycNaDlCiBIo
sHp6XjbMmKTYgFUUqN9u+LVTimkUj0WmPBDnXrEcXLh//gee+WkKqhZ54Q+a3A0IlGC4s0xXwr3L
ODfW7gwDymLaT99MDfXm86v5L0BUADwWe62s0OqMCtOsJX5OTZL2dlbT4qe2/KQ010iHlq1M8cD9
qE7ASSIIuGNhGhVWFHOD8u/fExBF2ctwiGuXDxu15UIFkMjL7cX3FhMcH29xcaeXa/vf+lewEYI+
GuT8Y2BbOWhN20hR8qjZZjb0b58WR97eUGJ9qHdjRroNCD6nuAw3Fbz7vVf+CSK0L9HZ7MVrPfba
juZJCqzwWMLowo+bvDRJ+NfZRagautRsTnHOETeeMxtJ6psDuJpW0IMtGvBpTckY7MGg43lZxCft
/60ET75+MjDNVzvNkGy4BxhMTw8doxV/VCqI96jYTFneJggj24Yg62CbQEjOlKBeeOOGxqK/feGb
QToeJF+3k8Z2uXaaYb2YhDsAOtnwF7evrW45yn5Lpkn2mSSgzr6AVKxJgAPFbG00FpmXMi+ua75M
7rYE2BPXKlnicY8vWGlTMI4+SLUTZqHStyHtIpoJ0aqbF8pO2umn8gU72zu+ynf5CSaCCZsy2HLc
P1hm0S563dBux/O/c9Ty59nk//ko8Bays+e92Morw0b8tCuGHdFpQ78tBIQILw8j6CC5W0em617F
OAxUj1L9MEM5+bRpSL35ZXcdIe4cbeZqSOYgthxOsczYSGMhFazDGl2MNosXZYL6kdIbRCmPh0h7
69Ufjye21UqDxZmr7rSbJY4jIY+lXg1Ol6G6qYOYsSKpbZmVrHb/wjucNtK05+Cz97fQOtlkzzEb
ax7t13sz7ta9nNdbvgcUAt3aizpd7u7YsrgYhLRZvwlb0xrworT/EhkvxIdzYVWKjVgpyvl2AIb8
ZtB0aVr8LZerLS2G9TBr989Y10RzrM3f1/mTjVq+y+5Z1VNaItaVk9yO519AWynVzo1/TGrX2Y7A
ADFbhxl4/d7nSKwj6l1WX1GXMeSrI+D2xzOa/5By2QezeEC1tzsxOXilXaLPLUcTZNWNqj1HEtIK
Zw8gyA97WnJg/CooE0cYzcdM1jS94xvWOl5XijRdILNcH751Kx8bPpTAlWITZ6LaIIbSimK/Gj2d
D6sgDazGnEAwXIGyPzHUV5Y5X5YAdyXmfOjvcr8OqDTvgHzt0EugFZWMB9KbLtVEbe/2NgF0Qwny
atUKYGNQJ8LUp64xMORb5gChgY/VTYr4RXw6yCHB1H039TrkCm7XLYgOZF0lkdQeHhad2PQ7wGt/
Pvh+IllvkHr6NGG2u+RU33dHzJal9cwavfIbgBJiIKVu6fgWCqmloJzg8o8rSZQdA4e6FJuVpGs5
4RwEk+30Wt7gUZwktycNYWiMphCxebxtnJ6qVabHwcKg/ZQJpsZJRDuC+lr5MqHCt6DwbfPnTPCE
TeikVHqSsHKk/5LCDbBi7VZeWECs4/KGu5MpZBGJNoBmk71AFJt0v3uiIkUxkUU9fhi6Ou8j2C9y
sTM9bjrhIY5g5v2zDrhmQ17eUH7WffTANVmOf1aBZ+6/tBXfqg4ul3j75MlOaZTAbgCwe1qAb8cJ
9sIGy3Qr0rywi2YsOAzcDqTnjTVUPZAQD9yHJWGPy4CcnhXfdzEt3j1jUJL3xm7TNaPKffO4A7OH
PX7t1QQeV55/HsDJBiAHBNikDSR7aP/7yJXdiD3b9fp5tNp7mcg2tZO18MkjdM6bIZQRVzYznWVP
X6IiLiYKJZiDWHj4+TPndwd/bFabJkpOCXQaDown+s0VJsDT2UHlZThvcV/JyM3aEoeLqBxsnSaB
Cxegkt8zfZyUUGOKo2ERYKz0hctrG32IPF8El8vFKfHy8UDudZ12rgAGlnRTJcENm+vUvXNj51uL
Z3KBETkcTQcZd3uebdfZ+0kPOm6z1FzMnE/DNo4IX+C/Gn7AiYWFLPj7KwJduc02a5l6BaJOn2Ga
XnBNgVZgiaygh+9h1I818oDOBJD7Asnq1WuydTrmCrtD0aTWkHdwJnsPa4zrXAPgTodV4GuCQfJZ
C/6PjF0nLFXFhGeIkogiNycXdbuyP5KYSRVP8tIcXhwkYtAAahkbddS4jkAZlV9WDDDlYYaNYv5j
rfi0PDX5oJ88tg0+xtBR7A84d1AP/8uy2d5DfblFcXNNOa2u7e0YTzIDUpQzX+D/JF4Q8q6DTvTw
AhKeirJdIi7DGNkFk+LS4bTwQ57sGWVP080L6Jt7lH5TLeqIoTh6d4HFgGvcq+IBqxqDKP3MDlli
V19wGWEYX34LaZ7V1030+qFdGa8YSdcgxlGPkmQByr310U4+j41lAVT6+9Do9KSnP9EErc1b1R+8
+VY/l2kRkLzLNO0CpKPn/JbrKJVwEjOVG4WiNHPGZkT/uC9cJjnmg8TDZdspX602N8anxv12c/Cm
s4FDVqJsdS04l2PDxc7HHINiI5lo+n/1h6TmYOHnw+8kDvK72ypgzYCZmXRl9GTrFtfqfRiktDaT
SXGrf/pxLlDjSdtocTLFRCM8jI32VqR9dEhg1Z6tTVhdTnGlVAQGYT4gM+wlJqijLvXG1bCMayd/
fMUIBTD52V8/kZ8mGg0Esc4nd049kjPSvNFSaDNynjkzcynAqIJub0Pud03R4rl1aWJ3Dxs1a+qH
EUzOqsLtRkWH+w4xQFEkWKMMdoGNjFRhkBDOMk7wuAzlk0iBNGUoHsTv8nLigecMowy2tRnJqYm3
N8tJZhW+uPh1wvOR4ZW8XBTj6Pwzci7IPYnk1PSGUK1gO+eqOVV+w16n0ExVYkfKWhs5U9HCWCIs
gAUuIo/Cqb3GTvg0On7NKdzgnF5QR88F53PdGn6oMQ9MoJF7Z2Eh417JXPpfPOUYO+xX8HmhGmuu
FbGy2YpFFlnyRrzJNYuKDI2DKSuuaJA7OLxm5jMNhENE9O7sF+mio9NJCKeuTpjpYI2R9ATfOKD8
/SLzAOwOPWTRqXbG7ndxwfmeZRCDMsz03Lkc4nJg8t4UqA3ZOXrNChTJptV1n5inm0wlhlfeDYj+
smGeGbdMX1ht+W65eE4IYbB8omQh6pUv/xG5xsEceshxtrhIrtTRmX94sOHHbHzU2Oq+o6XKAgM1
V0WXSOnL7Y0BQ9Xik1M1qC2uXJwkBBGQpgz7sd92b/GpVBaGol5/zXeGTa1n+GHs2r09LEcXLltI
jVdZd/3ESJSgMiAVSHOtVR0GDEe9UkV5x5lCe9fLyvOq+Lp0dmbzlZYCxCHKePlyOfDeXJNmokml
Iv2CVOQIUXtwCHEUviCFvQmppW2vOmDUOwGNz7S4II+WCdl5FVfqBUmSXpY3KBvqCk2jMldVLuJG
SlCDGBmDEk9syywLXun8D4e41ckFa+SYsqfOTP5ymMQq2SmQtCQ/hzoUjnbh7GFZYbofqB45beXz
ZK78mZfDhGhtazrvElDRuJZMi6DTBdckp/yfCp42iYpbkZrbdy2SdZBucuUgumMRAwVwgTmTFnbG
IBfmYKJmSpj7Nt/KViXy34qjCdnrWwWzCGq1Q3AVX4tpqHEZgBluGEj8tO15BkORsDbLoV5NRd3r
+av0GviY4rfvVE22iyjCgdZHYABeOCXAhPDg2N2RMR1BuLz+3g356UHHQAEplxw4eyBnkSzzFMLQ
hZTriiaaDDEd/io7SUqKR1pQ6YRrzPi+cScYuEoJXKn2i3mqp4NfgJ0qzwXi2/PfRfqO+o2yuB7M
0dMZtyWwYIqhph335KMDBWl0X6Z6/Xd4uEy9rul87nEmNnZzaxq/djOltRa2B/ArOEOwJKiQTlI+
gQy1+UUbhvInm8zoTgriwwX2KuCwe2UwxfvjrGxPuZT2Y2EgUjZBVWluDq1Z2Wq4GMNokjna2RcA
ZdX7RCyX8l2SKC1hmkxK2Hb9kDu0TJcPTBilOIFyJY1xcH5slGbwmMceMbnOxTeEn/ikfwLNT6te
3r8eKE6IZSY8csb9dIC8zBzVWsY809edFj1BMjpVNamLlOnmLxrPdRbUNNseDoH2cBT4mifllGGm
DWwwuNUUXSiIWYYUNT/Q17T9jt+aLq2QcEi4o4Q8V1gy5CfUZwvKud/kxVMJTD6sgFSDIKy9FoHL
w5oXY+oS7CK9s/WLe9hQR6w/DwZXdSZDEBewHYn3P03NJgp5o0TSNvASHoA+7J4ipdvKbS0291OH
hmGJb2wL/00P2BQI9SSbZfIRMMBuPuO7h/CC1V2os8LgL5RxDd0O7Ju9e388bp3OKcAYg12KFnMr
ppr6nkLHGDUBk7v1kNHVqJ+NTsz0oRbRBANDNw/XgvrDEcvE86jggryQCUSndiiZp7AVuWDfRKz6
0SaM2AwGW1xGqxa1bTlWpfeneWuRSnlwTONqX6LHFdQTz+7DdL1s7zKF+pmqk0k35OAOEF7h0k8s
RgVF1LXiYt08AR1XUsXT+aCPBVGuf4zCYNptlO3/oUMwCn5u9m1tBE+QuhZQj577WOan1OeAbeP3
D+yBnXPhuy06pV/sn82zpHsYfDQYUBi71ZXQMbKjPLHttcY05ZDQXsxfjHuNRBA7QltOVwMw3uIV
XT9+PUVExkjOBrqw4M6uoc2EOKHsKzBsw5YttfpYw/RUBIJ2cltt3XkgsKshj/JzvoNuNze5Al/6
4x1k+2xAeixrI+PbEWffSbNq9qX4K9TWWJGp+QRhtRBvvLbQluRmblhgC1duIyonKumzp/yduHh1
dMTA3p9zLJLM4dySB4NH8CL73MtHFRrUovCzvsn4v8nQmUWan1i0JLd3I0AbvIAb+fOIGLe6yM98
/DDT4Ig41lX74zmjoDSL9/u7WaSAVDy8jxjiPRjxL1YS8sGqfqyg0wzl3aKnv32JdboqWSjvdKdA
FoIjC8cNfnKHNoRdfSOWzevOk2ZSfuoDpJ8zDq0WOzma5TPeGaYycH9MYzUmAQl8vhaBt1EIq/sj
JSCkb1IpH+4lR846Xko9lR2E+QV4Pj3SNpQ4bK1cEuef2x7HAtLoN8fBtFPRxADTTv8FZIjRTm1V
B9mIVyOm4JBvn8SPDqDRfnOSHQHARh+/4D5LRUUsyM8uiN1YKVHqRrLADf2qY+gcmMCOwjOiNvNq
jbsUahZQBQBBPv5Ggaa90md1mXgJgiQzgS0bDJRrsTy8FUcjUgZhIOCBAmQAPwOe5lXZYOv7FTbn
Ag5mt1pqPVk6BCvu+tVlfCoh00jKD7KeE6HK9g9ii3E4U/w+V3fw/WcM5rd/l1cjsdipXs9QP0kV
I3ufPdnTWaHnxZkKH7icGAiKPcl+wKQLqgCAUQMeCkwAB/o0RQImfgbL6frAgr0jeCixNwOO9KbK
cmJx8/sg9EF8b0WDWlB0tElMojiBjDh0YCMRRqCsMxKWufChZGXGtCRt4vY2a57HYV0/H5bwyaa2
rqjPlhf5q19W7uDxxBUfpJ64VA7CC0RB5RtnsUNr1CyLcsKz5tZDnhbIzCZbx/ddMO9ptjYyAc95
nVkSgVOJfaSDWsafyLggCC6ZDWYnUYfcc7VkYlk1dMMfVF621VHvZnzd/pdYamKE4iCceIgRYjzP
2EYj4h3D4uCs1ql0RPKiew5EyGDjfuYstpU9xt6sLsD6QEbdI3UOmqMEP1jLJcV5bQtVANZyup3q
ifF2KIl6cPyD8m1i2mz0ZgC+CkytDNDqCePZc+CQytZ+a8KaDw33FyFTIDgFvvb3UDD2OIbfwQLC
axdGUv53ZkbI1nx5+MXWWAwnSTo0zHXuQvnZXks8M4nO1ULgarEy5nO0e8EFD4/plzxQwDAZYe/Z
pvNLDCOZ6T0qLLEHHPIjFYzsCBC13oc3LDMMAizZl4RagztsCfBMuRY6RHec7ZOdUqr7vpdbnJw1
CHwJTwnkEM8oqo9OrKWN4VO5Ugz6c9TPOvOWmpx9Wb+gY6x2iOuGweNOD7AQtsOcBGTWXJZ7bUyb
ZchB0e0O3r0e51U2dzzmBvX7JqxjlS2njc+HP1T7CMEP7spvZQhCbVs+cJ9Krmr4/QoKDWxJVuB4
XqsHnaODH2TGlDPKN6efCcFHyjVDOJKssRaWkfZkUAf18Zyzgf0Fzta8/YInTAw6L0Nq4fHiKpEl
gHuWo39aB1SAE95zfBk9t9w8Y/V7L/PYDsYO6JBCD6II/30DvaMuMCZVAzdak//4BvMzYEiO4eRB
JLmCJjC6spC/NuTZg6q+LS/QcuJOiBdb/yES3wMegL/KW+6V9Ozmu1YsSI3+6siEGkNcIQf83ysW
4X0t7EztOsApZLiJQDURdSw56VPYbeSubrDnLbPZ3W3QtY6DBgZIJhu+ctpj3Uf3vRf7A1y/5vuv
jsNl+D9zEPicMN5oyd7QSr+KHa/o/ZHc6MVC60OJwnBTh7YUq61nb2DRsqhidI5585UxA1SLDAXW
coNCsKTfMrXoSuVDcMzRTmoQfwU2pdekVJyPdLd23Aw4bbpXrwZw7IO61d4n8VDp3x5Usk7FlPHM
y6r1W0V9lX3nb73DKnJjFUlEJwxL7OUlITAtOHiZ1RGKwa12gm30NYDlrMX75rbK8zx9HZeBifx/
XuFu7VwuvhR8AQUW3cT202p1n8JTQuuua9IWf716LdVUmhW1GyOsNe3ny68V93eMUTCtxxRm7pI8
7SRV5qqLE265BhKh0fwvU76bazuPrSqHjD6PeB5JMMArVhnojkG+U3SYFpj8wJMB7PyvlIlNv3AI
fRFHeZcvR5PvssIJYi3QC4sHp8uNFFU6nFQ5sI65U6tLUKNGCCG9XTWHIYs7azMe25N0FmejgcVa
UkJ50+uLBEWu5vrEwKxwjy1RoqQWcIsofPBccZQrf+P352dPZpVJ4U0sNxd/Cm0V2l8CTeEljDG3
+r3nJtygE4ce4vlYhFopZylHEUNUx0yhgybRu6LzSjSVA1jTFPep0FrmPU6kE4HvYcS39T+sPlzV
wreRHAejFBWOe2gdJ4wmzRKgyP/y4oruKWMYny/bQCAuFmUrfHfH49sskOvEBdJCY76aWQtP7tmv
9LbSCq97oN4y5/6w2/K9dFiWpHAKb7FsPIWvmm/IfIb2JmzFIkYtRpsinn/0pnyeImtlJY66aVD3
kXdsbf1Czay5mtAdOtt7B+1fux90iF5eWEhC5bQ9inNSuYTMp/b2AO5L40FEnISymEv6yRBlOkz4
IMyyEl175yeglX+XtBW7+l7/XjKe7IqiK3jh3mSyCDZ9kpWTkuu+AXSW2L5LPQY5NO6+7W42TQCX
A9uGL8W2NS3zA+sqmRL/bkh3oLdH0nj5dSDAHj+MXCHnPdkxMPFyOKO+mzqaW0yBKRryZQB0yAmC
cRCiHcuiMCiWerWAm6xvzp60+xNtZfB8Dzg9qMqnNpVOIj2gnzuHJi8vK4llTiAD7RVC0GL/8ms1
+8enEhtCO64Rj+uqDx/7bsvS4i21y5gX8fUH3kO5s7MfCrpy/tNBL3roDlGFLA3Db2MpnNToEflF
ZcyliRJDcCM7xphkymW4yC5659nuzxaGjuxCcLKl/ZOqJRLbrvbSSuZ0O7HJXDa3y1+mj0Qp+p26
AnBbh1XXkrWjeODF9xZBxYHekhAtYXmsK40lrc/zk4KLum8GTj8YfzUpWZqhf5Pf6mCItiES6lMS
267r99Zz2f0auvHI6cuqSGVYP+7kKkFpN3ZkvrwrT88ZIZBkXqX+U7LCCex5t1c+unScKe3jlwjO
l3++xiYzhKKRpTZJVWiFhCea217MK2QeZcufANCwGEy9wnUdo2xPtqysY5UYP3b4pE5gXf/uYRah
gpjnJqeHslMxtnnjQD9mH949fijJxajK53w4GCXL/NSCF6E1jwFt2Uxds91yc8P9/nVDMqesE8w+
OF4qlASi9m/zsAGAdzjEV/rRsG6HjmbbLJJdAFiT00QndzSocy8sGY04FmQxkjmhW4yaj25PyVaf
LZrf3dnDMvz2jT4VZurMpM4VkANcgPUby7nLdjMpqWYzlZsiX/buSdOF+viVOqmm7QX7Q6Nysfwg
in0MDL0t+Fm9n3CNHLKVf2bb7SHRVdI7Rbz4fbtDW1JlCQMrvh3b1Tlg/V5RNo+zYj65QxOcK/Zy
1Et9/4n8PdUWymgShJj5ScmaQ9ANVWw17Md+aiCd8rO1S2R6YbUDiHyLMnsFWXud3rK5u2AphPjb
SJN8WnlepMTGWvVL5DNqVV2N/DITaGBkZmSuAvO7MgnVwsox+RohyFvFTaa/O3Wn9ONiJeQEozGL
A3HuNscjGzoHju5zPLw2YrIUQdQt1c3doZRVc7Z0P57//2fcmR6mKp4VMrIUqUnTxYew8G2+IxDQ
HcdGRRzzQ1D5A5PCHBIC/8GbiA43eNsYhZ4kbuyruR8U3Vmi2ZbSSK4TztOPBY50M2zIdGM61UPY
hv1ZZd/ETxMEy/ryhPd1yVxHwzALJVPejZDLNFfHWEKvPorUd4mkNNYPHQbz3r10unQEOXvZFQyi
aK0UP+KdmV5X0vJrJpEanLvUqEi9Txp64Ikj3LU/0vUFZJQgdMsmQ8vNIxJ+VpM0dmX0aDCcta83
TtPQJazafsfb0S4ikheHIe168LGEMujdqOJHyorAefyBVWELHl8UY0MabkqQLpOrJzj8hP5suadd
O4OaRGnzlxtTAMc1+9i/QT/ezLsxDGA0mBi0PRVTHfLy1HZNFg4JT086flrkQ0Rd/p/nTWHFYMI6
rCqIqR5LXRcgmufx4fn5yBclb/nqSva4eimlqIlU5JCz7nYGedNETJ1F44/kiTzkYQk+K+zg7z+z
dvGkBlKBhTKdF0ESQxGVbeMcDs6BwvpthZDjL3gtG5jXy+XTgjPQYnar4xW7zO0LsSDhhEMiEBnr
2s6p7kGbQc9oyJaPi/uVyW0eWnmZj3tJU2bVcFAdJUm0hcQGQhabaFEsOFac49VeF83qy64itfc2
N9I36/WU8/jIT9EEqUnCc6uLZVYp6IubLe+WV8bJaX4KiKZvDrmT1q44QA11omcwv8sDSyqFaep/
PBKSqxylQ1jxdStl8HiXMk90WB6A3RnpDfGz3cem/qnLhjbjABbB37nm9Cw96Mt3L3GVwA6nNGC8
ll+bEYVr6ReDV7+pTlRQtDl6FV0xd/GGMK/1zaHvDz+XVE4+HrSATUkrDPpg0nP9HO5vC+y/85hm
Pp9ORBFCAFyINZ0nS3QafqSeUQZ3ac5dndIr9AWX8A0zDtNwBgt+EmHqQnuVbJDL42uX7IQhPeKL
W4BH5lw0RFR3AhiaExjuD3Ebly1MYuA1wJu9s0Bylv8FB3zBD0Q18XKU+ad/AwFbmYPdfvCOTyyK
+sviNSOdUeunpcOHlkQVIFRZpkPcRHvqZsucvABENQmjtPrKflz5rug5dSNrJZLOHuU0e9rofaZY
k///5xhc0tOvMCpxB0pQrq2fTZJ8VYa+06K8lc/UaMm2hJTq8fma4kADsjb2oIqACmDmKJ1IUdCw
qDt8rRapFTjMOoasBWFlIk79xxx6pWVuyVh4cwmBIiXAuiak2bucJaqtXe1MyeuX1D25FbqQyB3T
i5f3eLMAwmCCgu+CXZlt1d2ua2xEktbuCJFWzwOO8LqB0djm1+nhr1x9/6WAPPbEmmoD7j3G8csl
IO+PCCxbl+gsK7j3CEi6mTVFx/Iu77qnmFLYzxoygv/epi3cqTFzubiW8fF4pVFZ4GvVzEpz8/e2
K1xaZq9jNHRRqrozqEgqJFKQobvnHQltgdyPT0rla31uKrCoBkuglf8T68B7MeZyBUDhZY5jjQB0
/YgE9pOdVbfJHo/WSNoOHkftnTH6O8UT5in/p/k4wKbmZerN55Ot/bAiBXY1Ws0wEo/3i1tSV4Dt
3OVqNblVlHqzKeqoHFF9wG46GCviRJ6v43Sb/LdV5gxRST4qI4skA5YC5k2LxzK4185r2WNRxArD
74/9whZP1uI1p60QL7Hz1fTlCAhyfsa7lUmcd3NhbghxX5u9umoHa48WTcbiDLtKMFEh3eAk1Lsb
fz32jVgsTfysOHIU1uWZfU6g+kbQUrzfZfFcWwRUkWKmpn0/3emOYkzFIe5y/btUYUtxUSk7c7D4
EWVHYBN30yKJ3t68Fzs48UKTJ2K9UL1q2ZUiz9tjfHhuhynzOO3D7ghcntClA0WXfEo/h3mtDP8y
gIWCeRUhF59NJY8s/HsbKKGf29Kzw2Rw4/gbEmflg1IQldZyc9yU+Ffk40h0BSm7iI4IOnpkIJht
WDXkwAtBRM3Tc8w3qkUGCvPcv5UX/Sw/LeWLEajptLqay9j5nKVc882DHedHvfboXJkx9LlIA/JY
u5dleokA6Tc2DJQirSKIo9HjqjbwNJdYX65+0iCrbybLGS8v9/hRE46VavVN2tUrh3ADpmVshoxc
Hw1bPZ67t+XOVAwjlEVXEMAxofMQ2i0GNJoVAxWRzFuf0GlqYI3aYyifRzHMYcg9Tq5N7Z/xyo9t
YQqUy+OpINmvkEXYlgu9CPjqWTuHsD3bb1FP4XQG6TXdm21/bbVkm/x+RPOcEhwD6EpnETaeQEbn
M1f9OdBvsByiaUXN3YGdx2wFSULnmh1BTxZ1k/117kiVfKzZ5R+pFe2OciN7H9kC9PVlvZbRHEAw
7nTbgxK+tX4X/LNuKs1TGdWs6dTXg1ZKkAm9UdDp/YZ5eAm8+lrvuHJdtKLdsi4viEjUUxArMNKy
Lt3JE0+WHXw3G+FdHXWlGckxd9HdkEVFWxk/V2e1OohqhW5ZNp/MQl8HbGAOT1YX5xlaXvx1fqpp
schreb1yH79KXNc8K9bEVs0X2TuoBKHmeljspx0qezqw0Dx/25Yg6rhV/hQVBDfFMo7Lf5vynWWY
ysFFdOOo5pcQ980YXAwY940ADXe//BuxfPGerMPv+jJuqMPadRGt9iMWV66Wm8KLPN/qlOD/20wi
0a08vY4+G/L/Kx/vB07gH0tFAkDJhKE1hVRaAEOCCoKHX6GNRzqYaaa84Pr7CtpqNEGNxOxsn8c0
sNmGdq04RFgY1QMicv31IGRUo4G4luoxlJMlUOLALor4AlWBamkmDHizPdSHPBNQ63eIgQmyzzpV
Eu4pVcgAXws88Vpq+6VkD09TOUVUk3SusrDuhTCr26E9HLGblQzZATR9+RGFC9645hlud13TmQzr
agD3lwYl9pd9HiKK/vGKj7V9FX4KYnbvxHXVY3gGxxoGvJnEyrmAeIKA5JU8gZvTtjoZFb3cI/XB
vEQaogtYXZoR5nEOBXesQRZ/vXZH7tyiQsFuDOaOy+PLHA9Ki/CRyyDCJmItYBx7A73rLgsUY6ya
AtBg5MuNQfZDkf+crkWjBacAa/tbuDIuplf7SQ8eHplKRAIU6OdVQZyIpDmTJzU7eNiGIxkmIkJb
xpg7j5Cwy4BFv9zfBA89GYDMcvrb2kRA8kyfeNfjqs5C0lWs9CaW5emivP/ycfz9k7sN21zdNlk1
IAUtOaR4c1t4WL7a70rhJS3EOcP9+s639EJ0jzGNgebxSfuX508afdo2N6Si0hQN2iVIIQbidcPZ
G8Lpqj0wXxUoQPFmpvSFkRlREZV1WLbrWgi34FYTP7ua3SZQ5Qa4A61XYJcPmvIc9dS0pNQTVjix
4MAbajvvwQOFB2/omepjVVrW+Rk0hs5KzJTyBnpHVvwtKQ2O/1CHOrs4Sava9hz3tRchZ4J+bO+3
Af0xSbcLfVmGPPcLvQoSs55JoQHHcgI9cxh9hWlsijnqlf9wtrMozF2sXs54dvYrY4BSXe0NUpTf
SRXF87jFJdE0H8Q1OLjpRjH5d4J73HjyhVUjeIwnVsAy007+TndFtzJNEYqv/37BOs9gwoLyFVQC
f8+Cto2Gv3Nf9qK80cLVkbunTAtHLuDsRfw4EHiHGCpKKGYxe5XdvKCRK0nvm8ux6DK+NxcnYxUf
MwzOVwf0A4byZK+yjuBVKdMtCwpKI9HK0jU0tJ+M3Vw2V292R0noFMVKqngMyy8dIM+0ckC/Up38
TAeW12+d4LT9N/cHOB73WNQVdk8GhSLUXGEYYAxBWiIOupSVBqsE9n33I02SfIsuXIIlrJWG6ukB
sx6YhHyYO+vmZtdEqGLlmOEBpO8zLNPVZnfUcI6DkGHMgPNMH8bzZVteyZ5nt7OzN4535X/CD4pr
DHcU/mjuAvbhds+SkSJMw44/mVJVtmMRISsgsHK1xsYel0RWiIGfliWdTv+x15HF/+p21wiBcrg1
5Vq5f0nJrZjL/yTUV7cKBkb9T6XLif6cBgN2BMuS6WLynFU23AkLy8yl6EaWn+Bvj7cP99inuza9
TNyPyrP3AKTMmo179zJHmtx2Ex7hmGw4njCQrdM3phzVeUK0u9AfhHYYGpQxpSNiJQE2dkm3YWG/
H4GuC+PpASltR+eF4RmBVBCjvDa3NBfGarLRFipDjGj23taican4n9q97R7U8uGWGQOriAbZRU2Y
GXYmiF/JVWQzWzWySZX9KqGHrMyaJ2xV6sTc9uTCzT2H4c3OEbQhgcb595q91i1seyRaAfNI8K3c
77aAxEnpAvNNqPpl0mdG4YZRek17efs861qIQighhLdpm4wDxWZIvctiL0u9dI85Oo8tjYCyQhNk
scZW9z/ey48yBMg2rUwCGLQJKKF1xYUhXcJDJW+8fU90eEC5DWA8P/sjuyZCWemIGvm35vo0g+eN
ggTp5NPuYT6UBl7W8jyyzjzzvU0h6GwnBXW36izrkUIWxpyyU9E61HS4M3NTFYNkE6CqnDgoxpSn
OfuQDzojFsBAYQRLkAeMztO/OtbHuL8bbSAHtqEzm5Q3FlagxGdCRxZUQ3uE3cWBOpFnDeABv7+S
s6Atpb7VWeDtmHCqS0z2IV1729zwaNXKo7HUGs4flWmgcmfukaDmMsMfmcNzLEoHaFdQu7Jma1qi
hoTXKgtAe1GIwYy7ZxCxQJ2CKI4GJ0cpDT8KHxC4DoNjEcS9yTuqJKlf8QoUE3JLhnFJqc1l255S
0mB+hx97IYKA1TzJ/JSby7QZoh1/Nkq1Z+x0GnIdeG4dfcE1vMI7Mv+4x1o+/Hw/qVgZSEbSZ2MW
ucpG5yLWSP0qKeNybBvJh+7RA2S2CRFTW6HVzy6vbQMTOU86VuYiC/j94agMcVbWEHoCaszmGN8k
jbnd4M4+FJ6s39HroUDj1B9OGuUKdZQKfd16zkxKEMbKksKWtgwxDj78DqYWDPp6ESEe+2xXn2yV
kC1ndnv+a3881wwlgeXV827kBPNZMa4l8U+tr5AwhH2PwZNxb/piLybRF/D7gXGQ1YsjRMsB6wH4
SDSV/0vwciCGJILhtPoSeJtmmDGg8uJyEbbqybztmXpn/Et9JopquOYV9Hy0bqXR5R0NmY+y2irC
TROIsgoInvbaD7BUQQBrRWWMMF+r9zSMKZD61HRdt+r2O5TYdPDbclFHLvvNq4YroZfQqvwiUrpT
tDpzt9xPNPHsqevNFZ4Wup9MeFrhRGkWRnSi4l4H7IF49QWU3PTq3pmQX8y0bUQBZD6XdIV+W8gL
oJzL23tljPz3GH7Vosd+o3+93Zo/fjblMSnDzva1oTDYtOciEjGkP4tRUrL3g7yO9W3vG3HGrSe9
7sDtlj/fg2Id3cawjXRXrNzdxIKrJzRNHATw71SWOJIwea6pCfIcjeZUgJEd6Ulm7Qxs/jF32bwq
180lXTODea7xGhpH3sGjzxd75inHE/boReloi/l8VeFuzpV1LW3sviwYQLk3xX8hDpiAAcfeNrY8
bK7siiYLEkEwTEsj2UB94IUKIKDRAQv2P6aAhvOH6XShnlmeLsQq2RSDTUhSd+GVJh7vTDIXPlVC
FYo4V0RaXh+UWdsGpRwtFesu7kEzZmfrnpLnhfZOgS0m+J8dIZZU+qrh/dlQiyCbnGdh5aDEI9Bd
mjbujPxqPH3o7+N70/6jppxlBHlmoOcas09h5VYE67Eb18FC1UcuCLL4IWSPF6vkKJMRBz/6/jM3
lBrDY4P9f755ZsCsssm88ccidXEJbVdrEaY2H7nM2ImdIn+QkpcZRn1zztFIskwXHSfDSWxZld3u
qmxnsLDTaFh7FsjncWgcI0ypb43j+6DqlxqKcUUw3z+C3pb5G4DoZIx6k3g8MW5oi/RYqFlRrrlH
NNekdmUOJzZUixghmPeBROrkeT54PzaaFOw2sr2UKQ0rsunvMHX9il7GWUVrXktFbRE198UJao43
GNGL9qWY852D6G5jxExcrAjh5SZ+Zezlm2VCDu2CTFf/Em/v0FfZeDqisZxAvz4IhoiSfK1KdQr9
9YYVL0PSino4wJcjO+CYttoLszlETF0pJAE/ondsYQbFUAULwxng5Yzv0sM93HrI6kWAePICOuzN
W8vlGgR9mdkxAx2hZMQD3ecz3Uq0wHtavCukma10Ik8bjF5CFKIf7IDxx2GIEU8srnZ+mevPImM+
2NGvyhYjXKGEpX8ZZmqCvLVun9vsdZ/WxYDyW3OQkfDvUhxF2iHlkTg8Iski7D6/xYLrx41dFJEp
3YNsYRp1Jw0i3Zqe8A124RfquK99W/y37ihCGTmUQ/8phirtQL3E8aJA4YejGC/nqvMI+NvPSvKT
uwEdkgN/kRBVRCHY5CsRb14S1lHlQmwWH5hjZZbOvY31a7DisVyviRJNYQk6ONNyxoDvQQKzUxor
WMKvoyc+0PHAuN9r/WbvEB6+4MHRVjZBAlcgRoMXgq005uvnYoIEtm0kJeiTN8C7HXPMcc439o4I
hiLP7QyS0e4fXzh2Yru3za6GC8H/ZzZzczcN4cBZ4lETVeNsJBvWpGwihA57T+cOa0Vv0LWmxcV7
NEqwkymIMOxRp7dTHtzfBjdk7nMQeFyCoyVFDCYjUXlN8HrkfuKB2UoW+ODqIfFLCkddfBgQFhhW
a/jjOeOArJnJmoYHMjrVWo7JYLR3aTBfut057iOHaOKKuHxeyTy8HRmUefv+8kT8vWRzBYaJnjYJ
ucmJrzQujKrQBVDdnitW/fey5dq04n+Bn0dFs5ZKjn3JllCjs8J0NO/lmyuN+mhVVP0XMsv4wBtQ
sCpRUbzmPMce8Wh+2r06TF4EVeTCwsbS1WyTsMvD2UxC54haPhwXjr753+GP5Nk0rUtI+MqLDhvF
eQtZLW7sW+ZfEjQof3+D78MriKeZTVDjacNa6WjwZsXCdlUuKvV9Aa+o/9fD9Xe4C0+mTPaXYvLu
l6EUFF3rvBQLkSBGSBzoGQV4izUWKCSA0S/OJ9wC7L057IDuvx2O7iXmgRuJMVxncognVPFeAlrM
P+x7aPgimf0pSkFUyEVFFPqQU6LvGcPReNvscsXenQ3w9RxcqsASQ0QbEsYWsKeVeQ7p+aOF54nM
4Vucq4f1LuHxlGeTWMfgmm7HMDud4I2XKVTrmamZZugNX6Sr2otlQE6w5x/3kWox92GnTBpmAbPU
v4z2MoIyFjcpdfni8ipeUgm4jhvxdfwUlZM44r1gNUhDaI7ldOBiIXgRtZ8RcedF6triuhyokbO8
SnDdjSdqBVfULTyT6GAsRKmPGwpq474LuRACJ5lbYlacEcQKFtiavIzDd7qpPKVWq2rsvOYvA7rB
6hQ0Di2sa1gZfghjZLU0PhtJ9nqAgwfePFrHWWDwVBCyPFl/odKynEdhu1u0EuyxrmuciO9NXuum
iC9mxNM+AsyeBbb/qPR0uZq+iIaDzMI7Iyz6CTp/cR0WtCXbFaFb7yOrNT3oyyCNybOoIbcQRyBx
vvZLn5CW2tNAXYHr4RWYhVp4XvUTO6R0WzUnewet+mEh3r83q7d1D2K75TTO0vtljH/n9RrnPEtW
TK5a+KKEZJAqaD/BksWqYKKRepEVv9KCv5/8+/oid9dzFtIocsn+tBGp2ormXhZRvvF39X/5vunj
8tdDqScYyFLSvfEoE+iWMGBjSWvkXcg3DSEdrXx0v5n1lLOEIW6fOeLjZQIWDhsMr4hwbAuiNqtf
onZF7lyfVib1PNFzo0ULylwHmA4AJTgdSZPNZTisLuwekmBZFPWRnuHSI86HSFEQ5o+UoRTZVsEU
Sh2658+DoxMDg5tR3kBW8x80F5Ts8MjgaPrDzxD56yk8jRWrm1y6lra7DXu8cW8EgkNkrDfDFDTI
J4LSha0I/5pt0PBbhxwWs+4p//JP67jvumTWMMaRXEYwQ2AYW128zE5+edRzMpm+uI8+DC4NS7ee
U8BSn/r2hkltb3NycvI9tVL6VrOniyKMRSI4Mnyc53XmL/p6bEyL8cgIvZ3JP30daagl4LaBWKAS
2BAtCc2thiP5Mk4/fCsHl4YHauKVR+SugAQiVDN8jlzxsh2Ag1WTcYzDfaExX/h6l6QkVGm+bSvQ
VWWaSBCxiC3SHPJsZlucp2VqH4AgDVS4/2Hd+eAb7S6aR6m3LgoteYzpDvy4WUcnLIVStcgzwwpB
EO2omfTpXOS07/J0ASiqwWCs/jQ3hF46XquPsWhIJ+MShY/+69ln7BixnVSnoXxsdIJfpLGMjahS
UMg59ZtE5rAph7sqGgADvlA0Za5MjmbdNEJbFPaNrd1EuFT8d8YapiKJdHvmH+syMil11LMiYS5y
qcDZA7VS4gLTgc3YL4kfLpFace7JyGRAPVqPFW8ymBHBOxwFgEcLj8ScDSEUYwyMTuUGnfRXBqo3
Lk3HFr4sDXp2nBhVHy8fBllUYE62hsPOZZ4lToZ73yUikoqL0PnY/dZB7srEczlvaMfRbxXsC5D2
a0pOs8E3LZXI+GA7BNnFWZo9q9++d84UWNMIx/JrJImKbsptZTPE96Dzu7CXyVLNZwpXA4G+dMPO
WpWjH9U7S5oLhVohUOwMIu9yRTG0NqhpY7ynnHnkbvvECqMiguj3k8RMMi0yUibsCKyzKO8D0cAg
MtcV8vQ1XYtfz3mwkANL437LSojWfa5Gsx49NWgHxWd5KuHxk9zeQouZIR4Zv7msDuBhp6jIOMnW
Euo9QORtEBkqc2QF6o+q3JcF/xr78m4elhm4P+fAPY9l/sgS/H9u4godx+eFFiOM9YEH2aQJtinx
oFFzMF0JtcPOFALl+rtDlWt7n+lQQmYENw+syUxNxoIxtqDsNxl/6t8cdDqRrUuGGRcYEfIkzBSV
2FOPtMeKKh4wckOxd3CAHLrP+TWfqiK3VFwWSXQFU1+wYP9YCZKnRtXKooetixhoEIIvH9vN/EKK
Sb3AsKhN5p08mHFC91EkKlVf26dlUd1VEH6nENeNutoHXfLmiJfYVwQCf6zFUgLF7N48fBhpL3aR
1zVjbe/74S5n4UVGKJWpQXa3Uys9ELzDhDmpJ58o37C3cTTfAP0gIh5f4wKlEtp2c2Lf4NGd6fJh
s8Hy9PRuyPRL+vjIA+9qFaYaUYrlKANv1oV54z5MWtXIOF6WgIarky7r5itbLleoVHOYRZ+jzpgI
l9U+QSAgg6h4Ceby7Se6izj2oY8DL73edfby5OXXy/cyCPVnqljHHMALURka/6dhHWa+fJ9mdlwS
6G015rZ+LesnpDBNFtafTZudtGHVc78ihPAG6f81KY17MXacPQ5k5QJ1ycbKsD0VSvNlM6MznstV
JbxeHrjrqskGErC9iwbZvVcaSBfuPwQjTETHvQYeXUXic7VTbVddgMJZc12dXCUHVJaEXhiDueQ7
eiO1TPOTMDVSd7vP8bT7EoUnkA1bxXxvn7YLq7ycvNkEHy1x98HNnvwxvgEukPkW1RxJ8f4cJW0V
6TQkynv1sPFgX0eR+f65grll84NyTY3O4AREcBCZpJPyhRT4ZEYVgGn7m0qCnttvNhJH42MeOkHF
yMR2EzpwY2G2CQuNwD90ucftMl2F2f5tfLnRRdeVgNmC9uwSbkpdyKHHXCPg8JkGl57/srMOWkQa
7XjiBPFVmr5o5R8BN3qloODgRHZ6fggqGhHpblk2b8WkX8uk5DBLYrLsAgh15u6J1heQugwH4ziW
aWnJAQ9f+SEnZvavg3RrV7B2W9gsBD5VG5FY/GnRKCe1IAZdhiEr1jsPbBulRflxZJ68wi9lGrIG
ZU56HM8XPCYZI6qwqusgIeNlo35gxEJo1iRSbDT8gbGorkWAc01ADEsyoWgHtyGEpJ7KJsDFsOwL
5XQx5YrBLRjprPljcwgBDrFTG2nqWszHEk+AKe1JD33XpJvyD8Z8M7yFDgkOeDysDnspqtUw6E4W
TFjXLAfruwQsigMlZ7LXUFTe3Ujz3/eyh7lOJ7ZUuY4dxtSMxhb/4Kwn+BFD04fWBK5myj87AEJ5
A7MZsB6Cbwz1YOhzjgiaysbazQs/oMamcrGHrim6yp7XwL1E6yLlbKKEjaXi24vYhIRftNY0vdgx
w4ivE+jIXlEYfvuc+2i5VofoH9I9RZk3cxA3Jt4FOTHUCveJdStMQo7n/iw6V8VzaS4Wdte0DXK7
h02QggmFFQeiwV1L0UAxBBzT4QkqYD4Q6zspcstQ7Gp5yeCHCKSQhzMvq3015nk/c4nnF2iOWVj9
XKXtSgjTJsJKPGO8A5rx3gFQrb1VNxqTCQQ1MY/06FcBRsmjIh9kX/Fd2HBzEljx+n8KrJuJPekJ
dE0TQ6e9j1cSy2XLLW9efALfi8UBKm6hN3F7YZHrNK5wRr8+dtv+zx+9t2ru9Q91bVKzV36aj+vX
a3rak8gQR3HNVIlpS6W1okUQ2ylCg1fd6dU/5d4O7UgTXP0jzBk+qkSas844gie3BgmJXr4WUdQJ
yDOzVCJMuHeAfLISaiVTVIXePTq5KM6OfzdAecju4ac7RYpnAwfa6e50kHntENBTYEspvkZcPEjk
KPPE30LwBabz0ULLvnZ4JiKDj69uCRSkt4FURAEgiYTPKrnLlY6Ge9KxiCSnz2HsJ8VJJSC+aBFM
G8M0HdlCu+riyEAIN3H3IcOsXus5aocwDul+uaU5MKVjZENAKWx3oG50Cp7pAHRZ3qhstcxod/f+
pSHAjJuSMh7OqKeCigNPo9EUMZwqGpbqh+RZ46mzP0x/s/F1cqOR9pJmmN9T0JBySo3xuApT4rUH
csGZzCdCfQdw6Wdg5R+1bBVywFlWUPlMb1izy8erOsPVuCH2Hd7mMUWHMqtJ3srqbLKblijWn/D+
HC/NMLP2LTyLbLpi/C/FeehpvWMApAwznvUNDYfG82kRVbY3fGU8FnbdPDS/Gkn0EYlDOdUr+gNT
XYIQGwQAN4bRxguccGahnREJNzuKQ95YORXGCCzJopm4fs/UGhUjaFKP92Gf68uCy+LTMLb2H77h
KOVxHFBhKtj3t7zErWtVljAjU5f4wqM+ueEr4NTCdgzIM5PBvzBNgsbqsdUDB4r2rrld5LRQIDsP
Tv7JKtv3YE38d1IADUVMQ5HBaJkTuzgvtoSdA+OHeAxunJOmt6EQMxdKp7Gc7kSTlb4jKjoi7lbP
pl0wl5z5Rr6c/5XB1EEhk1Xu7LUrwNYvGxOSxhi079YyEeF8HeDvyCDHTkyUrZx1nzRTtToMG/9y
FyFDt7mnJ8GzQ66xHAC3kBsk6AJUZfy1nSyjR1IuoCyH7D+SGpKEcVfwRvlB71NY4kgnVK8j8jw8
NF4eUufRCUJwGlQPjRSEWwUDDNQCDjy10e3LicMB1nhmuZqyA+2uaBkhTz2l5Jfs2oKPz5TDQmLI
iTykj/JKFr0GR6iNOs2vKciHmhwejBDOagg37jB1jihpswhO9KgL4xo9eSIwEhB+2SrUpnus41eI
kLavoNj2nb2i5vFfze6UXqeZBreDzkPAQlI1C9PhVS209cDJ2uPs2Z2SvHs8iUdMjhx8X3HqO3k7
eIrcF/opOjRsS0IsymcN9BbETmrGkoX1SN62u228V68iKxQB/eo/l5CzPT/6ti/0KHfgGmATWJrf
TsRYlHI8mzIB4IVf8bzfdUAFOPUHIFMTN9HuTY0Nr5l3pgS20QfsOvMV57jjSI5xneKKuDaMWz97
p4ksK2GZBLyh7HzYGId5ArFXBG+PJsdailhN8ISryPvrodbQfWI65dzoT4CE2p5gxM8xhyNjn7I/
cjVhJ8ilANsN5+ggvFqLZFJRvi+k6u6DIT3jSZHJEvD9o+ja/j38Wj2DIfoYa/Bm9PGnZPxATZlf
JZhr5a8vy0sW/Mu6xgd849ZMSMsTOz+4Mv2nkRmdY6w7vyVvBLO3LG9JXGQ4AeGsedepFOhp49LC
rzDkSSrX9Wav4/+hEmryW7vahD8l5mPhvIN7Wrax5PszvfC6jEdMKVxTtoL60LI95IP1uCp+FBFo
B2qTjQNlYqIpAt0XxaTpbaY1PPjAmRdq9w4uxVzUogAa8mOSlKitMNNdG+9dWWV2r7ihLk+RHiAc
z0nz8nNqh/gsaxcVaVhqZ/Qe09xNTptkxTlgvTk6k5M96/xktt/lCDTOxlDFsVZY45vYb1uxP0Pt
fLHsPcxPqgGtrHvTglZCQ7ZvPY1ukmNbaKuLGSQkMiNE1PSztA4zoolL92nMfF1rc0Gi/IowkiYE
sjaa9DgclwFhTMBoIDF6gj71rGRiEc2cwug+49sHy7JD63oy5508vhsDRNFdpn0MDW/o6e+JQW0E
Z/0WjMzxHzwReTbpeEYKxyED2Yh3YpInwmV5N06lX5UTEVJ42daqeAcxRbkNrDX3T/DONdZUMvGN
obOIbd3ozhY3stE8CufHs4XSdOKkwGJeikAOeZ3+65LaaLliZnbgkvl8G9QaAyKI0F99bawT5i4v
ltOVmCi7URMACVK7qHtJQee7TJytsWmYc/CtpwdOR/iU53oSuGh2kVJsaxdmHiW4ATaevX8co8Cs
VsToYJJAdBl08tPDuRgK3sZaBZm/0sJPmSSZ2VQmXrPpAjtpx/TuWeke2ET7nhzK4n51Pas6OAqf
0IctTFtSEbmd9ZQ2mgsw795rOwNkkeotennoyjsxqj2NhH4TSFC9JTWCmlzuHRMWV8wiP+gB9pku
P7VGorDlWIr6qfgpYhWb7OJXk2h5hZjLgkJJrRhN3i0PyXaKo0mKvRiBeWRl3lslUs47ybCEAiwO
n777bPFHZxYFjDo3NfaFgH5lRvgGAosDGZkHl7CFbKfaiDnrnP6RHFp6yYpphYS4hkOo6eKIaq4c
WJO/hHH/6Ze6qrLrj8otmkehdBa2IS3Qi962T28Zlt6TS/hs8aXHWqAcrBTN0Ie3gH//K2akXIi1
rU7eoc4JJAH+NGrjp0Ew8lbJ5DCbY8rhta5fq7B821iq44EIf9+KMKXVx3pgSC42agq/YbEn5LJk
4kPHc4UPTogFecdwVflR07vwCha2fMYHwjsM46gxlVzXWJEeam9gAludFpNW0BKjGX3JvWNaG8LX
mH1j3gFoOR6RqK8KD30efQvK7jpdlEqLKfut7OJTDajnzUfkMW+Cwb8AaDDJWymUh5SAfwdT70Kb
ru87CasyQ9a0Cbg12yTeB5tJNn19KsGLNa09J6ylY1KddUITawvUlHsi5sthWOR0r3I7XjrsLsGm
phjbTI01mZKUXdHaExkI8/+jPQOR1bv6O3gV1pMc+hUfS/rraUSkkRr95dIuf0aRjM7vtadqgtr0
tJnvLKD47ulibkh2Nuz/umruNbP8hhBUisFglVJX6gA4akely296AzhHSWjUE0exGmbM+Kdx/47r
aaHiJbPPxjxVrQofsTWLpP2lwUcOfAvSX/rLP8JcFVn0eGr6q0HfLM0dXHXpjvSFQzVYUMPZjBEJ
tDpAV3CYI4einUZfHDVB9HRDoMUHyOHYtqm29SCW7p1qIxA5y96Dg4GiSg2FvaLF8VIvwT80sbRU
kAynTscIX3+445Zkla1EYJe5Hn7omQMiE29HkQtKLSIuKVfLOxrpGnCpurYvzAB+in0V3AZQ+3S/
tKqh08GQuZxRSu8IFkm3MFZ5k6u6ofU3SPzSVkOQMtKLgpYr75Gn1uWEyt7hyXC6/wN6goD+63do
0IUC6yC8nFdyHA7tUOQmF0eBaDbgxxrBjWCTsRBK8wdhJLHuGJmjAVdpQQXKEMBuFe9QHYcjikYv
JhxP+9AjuEIsSGBTzBEzgnYEwMHrnPjTPWX5krs3viD1060YXc2U24gEHuzwkGx+sWSosbVUOYbb
jbtF++DTcDW6oMq4RMl8CzYTns2NxmxvGl/L9PRWMOqqOQDd8a3yVmf/EeqTs9fL5mG7mkb1zzCq
wwpxdWLUQ2zjvYtdJEWD48wkLTvw/D1QyqCizNnVAE7sEgs5LWhfH6AogyAxq7Cll3zQGIyoQoow
3Rl1Zk2NO7F5i3mi2WqkJ9Q8kEak1mc3kaRPlxZOEF+K39LIkAyoLqLhiVnxa4h+cqx87+6x1l8f
EJxBnj7OqhL5Xps86EOT5VfjMMfrNGGQU7TDpN4mKmYpjgdyuSqPhepE8ksiJRCLFGMotyELlbt3
y7/ZEwUW56GAGYB3/lvWk3gBBfE6rLbc5XA9H24EJtewxSiY0oBMMvn9IT7ynu13JlOvm3Vlcgum
Ei0yNP8mW2lTqICNyDOuzCJA2N93LAqOj7sL6e8fKsgjqoHZjrnLpayk7wrzynyrHB9pCNs2eMiL
naOSV389weLIaTdMxgfSRH38yl8DCLmXOrp+V4miJUyeZGZ2E94WB6VlxS/jsF6ASdZeOM7PB7ds
VD15B0y4KpstETsBNxMYRjncyV4KhqXvww9//HJ/l3xLJh8CWoT7R0HFxW9XXbJ8X6wwqxO01TuP
9v81f1urZn5EEaZPbrSzxtvdFW4vBZ8aeIuAmncx9LtLySmVHCHMomakLDQtHCo+NAPe7JFKHI5f
sxnIvUulRqfG4D5lSWf7avwsbQPHgVs/4JvhuPJyRgxq15tiNqAkWuCqzy4sJw+fNwUjC9GfSrXv
wgbnnZxCXxfx1zZSzB4UJudtUswpGgd2MV6vTRUCnwsHVL9dMDGWUM6jZGDvdaYxKp/PNNc97AU0
wycLhz/6hcPnn9j2sGuOPItd1/sqGPPdfxxWePGjRsnBj0rmMgVp+1K73MIWkN9ZhwcIxjCyQfKG
slzkKbhBT+7bbfCam/+pxSQyjQVIXwMkXGAl9/bhpsdKYt8EbKmJChJ45MVLqXcNEDEDtfY0m7Ev
Aav3eb/IMklXtPasQFr8uRnwYAWggXq6D/UhiZatH/StW5+ar85JMyXOAkqld983k/50Zth8n8Xm
7AALJF3v8lXQbNd6/ZP5n3/ic6qge3rUpjjnyccFgZUSiYq/yVSzyv274kUX4N4whUlkgAFUnooz
GctA9MqV7HPHvj061hyS8LjVWAcIR+QCy4ABmYd48mHb/p1N1PUXdNOsz5M1ELZnxAJm4CFGhLty
Fgqy/f/duEbfRI43wcufgq4Ti60+fgEYKQsbiVKmU9UjWyvhzOGJWnyexRCRCZ9dozSH4/Wh3/sq
1Vtiz5qzh8LsVRPh1WW2BmPcALIq9aVhrE0C+MH+B5q+1IJ0s7ioiR7fEvAx2YxSjHR+q+OiESC4
sU0zPSO+y3sKq09qOcQK9oRKLqU35c8rVrY/FiEqU93/MHW58d6tSi7g9mVxnfn8W6uOzYlMYL4Q
7/LF/GupTTyEf4g7hqy3nVQ48GNsKTyOi4NprWa7mftS+Mmx8+3l5dsLJjZurR6d7SySSShf3rMn
XdaTZFG6tClDdY1J9hkFY5iVdQhYlgozXXqXGRSFKooyY+Cv8PJlaPzVteT7H8RfhGKFsweZP+Xd
6bmPQWNfOoFgdCgTlVIt3GZXfiiwfLumqhPJ+sVm2poAwI8mnF8BAnWf3ydDlT/uy0FFbk1QVTP2
yZpKYTFMEyBbmhfaPj1sEOxyqQfSaxOLV1y+Ti+dKlpGrBaFpylDzVurOLeS6ygEx7WjCTBW6HwS
4Bk3RTI8papfMw11shFV0WWjZ0PyWJpjOWasW5NP+4Dfsb+IzTEEa3sTpgsAV2GoIrLdT4rojN1L
I/FZCwv9pWtdCkchBYrdm4sheRgFK1s22iA2DE/Ncody8+elBT50Yb1BR9QUJCD99EF2TmuIVHPL
uS/O8esG43mxL7UUcoDKSku2GqhH1xtkJ/PPtSzpX73P60P5aqo9psM6eBSFKMSe/4ZCxmy/0pc0
qR1NXSG7mLioPuTh/n/saPP4OVTfSarmhU5Eza/y2s5S0vOGGaBLuwv1EUzna8WjlvBK7+jobN8Z
8uoV8xmkkj7a04pyP3ZEk/vyXK1mxsrjyBsqf2E5R/98P0xI49RCKy2Z1PY5mU2L+rJ9BRJlCn3Q
wb/Ad3YTLjEzMRVEOeas08OGBfYS7YpBIjo0jWFAhaSKYhDQc/o3VfrCV6+u/3Z4ojMWUiTIq7V5
HI0hFIxEPQwCJOjQkAWyKfzd2KZgdcE3nnhLGtd2qnQQtSsuX03jcO9JBm2FzwfyFliH7sJ5K7tg
8BwyFhn8KjCbENnyZYLX7BCzsJV79lV9jpVZdercCLjo9LwLxVpqv3DUESPkTk/fkuuXn5urRjqP
ty/92h1V/N9mBnouYzUmtgdp1pIhKo3aBhA98yKeu18dJiuAAwmfYfqZ69foGogQQHRZPHZW68F4
s37WSsL6OxpEVrqMVsGvGFSth9EgFLhcYvqIYwPKcG8DnoQ2g7OaaXAYdT9m0d834L2Jczs3jpz7
5poA34I9ZciyPoJD9TWnwDdn3wZRr3Lv35djauC9/F1zg5xRN2s6CrgT3oG3lERb0wpagasOQdl0
QvGYhtlMV273m4KFxG9JmsNp6ZkYE4vuJ+xo4q2gJwGtjT/UnAU3chTzXmZoM0t1W93mFCijtyqb
h/qHcsW/QRVHTjv09Bs0keOtNYjpaHSC+MkZd+jBOwas0gHbiK+PWWrtb7SHz2R1jvtC+6c2ekTL
GwrNlZ1JSBRxaBJol77lQkEvTsPwRzIh3d+IK8JTKQbx4ED2Ej1hqmZPZYb5i8Pp6xnpyaTLaVch
cOLrE78W3DWxAo1e6VTKxsCuoSKahdkPh/YFrsea8Q7KQvOge8DPU1jWNjcOvGyYN//GVD/6B/pV
63cSHD9qoPT6ELHBEwat0oLYGbMjp/Lsb6X6vmeeLqBQZLtySlKpKGW0nI2L4xTXchIAeyB2b3yY
hkOMWgB7H6XgkLfnX8W7+8eNoRDmFC/ZyaosVtnrWHWKvYaVz2YmKOoSqVi7UTqYG//enCRnOZE2
tRPsaA1JLrDjPSkUwx6SonUk3gnmtkdcR0UCK4Mfyywdk4B2gVBqJNmDSO89I4S+v6soQNZUqznB
DUR/K3YUs6lFZGn7omtVQwnzTXom5NpkLzPhTjePuWGpQM5FDWjVW5LIcE6Vq0BtLiXR1LGIr01Y
swrcDv2Tvq5NBBoAjLfupvif2vbFhi+lkvQIPCP9D+1zra8/p0DUAVfUokEUQpysaxdusJElpr4T
W0P8MZGzM/kneltNMIwVoU+VsvqxiAv2M9smL6bUqqGTKfFPn01NIV8n08ZCd/zpC8RpaFNOCDPL
6W+cd6jz3DciEZFk0PbH5MY1qvCb3Rs7E0hEVJH4vb87ejp7EChTd5rA/3WfHfrFUDFObb+IrgLd
sHl+ocGYqLJDsIXiD4gH1ZtEvxOpPGklgEYI2EvBecqHuaYeaeI1dpS2gjsKp87PWn5J3JivTtMp
Jq0bkimF64YlYxDyPOnVaQgt3d+deqDgntJK1Gj92FmlxlSJJ2mmYC/kWTiyN7L261Gdg6kheiVy
XiZH0gcWbXmhUZ9VLwrcJTkYZjB7QC0yVR5QihmEsfp3lGUqTrDFj4yjw51ODCgmmSy7nyLDzMZH
qVWHNMs9sOxJck9ApRuTPl4nOQ4KQQeeDFIumUXv2qvuxgsKgfRRuj3UdWfTPa4niPBOTMTFVY0d
EFauPNQXXhkZWYXwIe+yaDZgQ1YaBARiEQzdpXXYtxtNdm+GZjXqIPFEpZmFynoHlAZta5dE+d0P
gDQ0/csSIZZ5dvGSYl6+km1ZxzMJA0BZADkDTxFbiQtIL/Ookosybezdk632DlxdHz5gIUDMcv6G
51hnTIgIlfSYpozpMZhFYzrg9zKtkav4lxw5Yx65v7/x6vmlDf/GgX4Wk+wLUS5EQdSt7RFRNPez
5cV6Jo6SDp+Guar/6gra+Ajz8TxpfNQXS/2AZcJH9RfccCsG+5iC00SU0nkoPdk9U1hqbpzNbhSG
L0i5rpQBp9aWN0vFppEcmxWd+MFsJWPEywto/fboH6dDDV2qWdkhxIE+N7r97s9hxBuhJ/gNfnw/
e1M2ugntwiAttwDVWuZ+FokPg+Ig8Kzn2SUXfzPSZBIBTJwSc7QUaRTbdIp3WIJfoWyxMSVwhdP+
XHeF1PNx5+Z8zd6VzYoT510z/7CRAydFLiihQxwnHP9y8jxcVhtrzCu54MH4HOsBnqXCOjCT++LN
8oEoYHBL94o+HXNj/tzMARIqwt2Y1da1nR+dUr+SYtCLblnHtwgSCub7hys9E5jYvOlDkwx0IEo1
LO1in6vI2nAGh9z4jOWAbwOBs2CtHfcAKsGJgf5x2k6nDE3GYakDW8vtdAOwKjXP1l3sVekz0zrq
C+Ra3TiJEHYcXd+3K8UVzQyX+LFbp7CjCg2K/fQfhw1OJXY12TfrV/ZL1BM54foZwBthIL6ewXUZ
YRN2vPkG/qVVJSoOW2n93gKIBhqbQQHvOk0yDKMRli/6HLZ9DB2Ch8wqf3hyXpZ6TQntn/zsmCLd
/WHqvZAlrU6rOQN2+hgpch4+MO4pyl1giERIpjrmgdASCku1wgeoOKPNk335HqnWfFZbRz9z0qli
cb4WPrEL/xck3u/CyqVmQB622AC/C9LRUUZDOWSmHzqTdanbLzydkalYUxlqiHy4S5clhUSCvlMX
EgROdzqGk5HTz0OLdCywMookoO8ySYpRON7RA0wUq7DK2wfk6Fmb2AinKXHgtVfEy3A175YtbXm6
boYqtoWyLX+pfyOzSnjH84DdE4oIXVamGqg8RNz7kjrTVdoF+ozwaTM4QLkBYYeMmn8jSU3UmPYj
bHQIPP5uc722NneXwOjTULrIkqA0DH7YTwzerO00WzuVge7XDf+CE0jk7/hwPzFg+Qet7kG0smRj
CVxhaAxuEr4akdRrx7cEbLGagIMcIdamKcR0D+/1KyeJM66zXIPqSiPXEUblfHzY08TIalbSLiui
3eLE0AWxKYp/zEt2Z8S7ocME8j2pC3jTmTxif2QW7fexr0YHsjPMuPxveU+x+mwPO3UKGyHwo7Xw
3Ix+ArJEbaV9cRgQ/7OCTlS6zf2JJmRw2JB8J58qFxfER1OTlEW1OYgMI7vpn2jsNQdD3K8GNUda
QVpSuXEK9I6N6b+10sWNFPrxPxkwtBksX8tFG5sIPQwKl4EYn+eDP1RwXMa0bfE90UreyFC8bjDZ
afj0nXuqsCwfR5v0OTWCTcLW0LhfvQhohxlAKrNIXb6WNR8c+JmV+4k6mSp6jug7dfYhzbaR6Lwz
4lCxfbdkAeyqpPBLAWM/85QUNjgCN+U+Zp1Xm2si25QexiS26VmNHIMsZAcOkPPHKyPiDZlvFvhd
j0sDMJgONnLeB/pE36l+4NlwCLSmdqACYGXqzDXgAjlTNDiMn6N5b2WLU32JDf3J1zj2VQ0kMrk+
w8Q/dHLkliOyUFz7jn1lCjXMuxNfv5rFIEYc2llS78nBuJT06etwg7rMJRmhhEfiv2P+NnAzIVcA
E1EkzRrW+FNdb0P3pebzgL99+/bS1mDhgXB2Xtxu74qn2KJd2OWSeFTf4yKP6YTCP/70OWawX3Hb
z5YDX+y4Cpe+upt7p8GS6MC0lCaBzMc5KSLF8xyKz3Fg/jkOsjK5anSduN7umVs6NxcAy4RZKv9R
r/xEKtcusMet75ppCmFellgo9l/DByCZ1w5JlYyI7Wju0jfiOrWOQe8cvnOGNryBaK5rlOCTQs24
RPZQNWPQ1f82YXeuYpAmw1u9cdXeHdJe2csSd7f91b0YtTIh8JW6NiY/aEJl01jNPt+uGee60seH
HqM//oxT9mgH+c5GIa/PHtq0qMwqNjJZpHOahk8jYXDtFzEl1ZdF6TJTACdCZ+0TB4TcJrd0EXDI
/h06L43P3AOi2DlvF/7U4WnqZAPk0OctC9poj2F0QW1VghMbmWAoWx3FpjAQMBwkwfgyFyrvASWc
LWG/3jcU4u++oB9udgvoT0wLz4KJOLqF9XzC37FRPTb/4bOm0LojE1+Wy3wS5ymqWTRD0N4A9ckZ
QnrrW8Lt1FPyzQTzrme67a2fYGEV+IWhsFAETsHlDeag30/ISeJD0oWdEC7YfCU9z5E9dBqZLTET
HcrdoPW/xFz7R1zv7T/Gzfy6m/xDV9Hce84MMDFPdYQX70kRJe75knkbfjBe7GOpeV9mDgk8gwVI
s+3Y15je5P8gXdufVHGJvr1dXHfZkX/ZI6XF0KsmkHrVT5nAdgAud5mTGC8ZWl1gTvw2DvlYxW3I
u3Brmc3z3VVUzh3EzqZ/0kQ3V4lAP8PMOs/3ugl3zB0mSxbNF5Tom4HdmNlHF6jBZly7VSzWVTQp
bT/fMKNB0MUSGezn8yLqocQ+T4yXAZxUDuNSNel+5vQ75vd2TLQ4ax0TRhyWkWEWVXT/tbWHOd5X
i+0me0A+PQVSgysl9h8FXT4ZfOiUvJnqJeJGApVQaC6YVj/LMvU+2c2npmf2xKZZgF0kQ5Qsp2zf
5DqTHnwfQd+xhXpYLpeXlcJ2idzq8TxAqPWSLjK5QQWt4OWbO915KV7r2D2pAaxFgxPWvxiHbCzv
b2dW6Yzlu7DIXZ2qyJGFORX9npHSdhzKcOHIp0UA0wCTIXQNLG/UwJn8eaz7nAjbDkXjdKieaHPt
e9GvcR/ClVqfAvMdm8l3N3XnGUwKqpFSCAEmzvsIgFTI/BVkmh0dWS3AiOl82DrN8jcwv+4l2zjw
1PgbTSkslA10EnBcbSzh8TbLqCFq+TegeV/bZ6U/Ch4JB0suMHLiMRiE0c0wkMyo3gXjaoDYRN62
RpqwxqwrzTl/iDctbkZO96aRT+buZGAy71JRQfUVO4Toh+1oOoW49wtnH25zJf/GPjPhWMoSrl0I
VDBSWDyN0fi6pxoT+Ne6dCDyDZacBK+qoOBnG2RkhTkZ0lgpzbpR1IPK5Phvc4nNpcjwF6SfMU/J
KOPDD/qZpOKpVPcIefvNg2amruQf+hAj2efFXSn3NtEJLs+ibvxZnW5zzPRXVnR1Oe/ilXTzi9En
d3+nvI+zmh7EzaM6t9EgL5YceXfH/Kx/Jgjol1hI5APUxJrlHf1A3Y3/fu5piXsU0Xyf23sDMFu/
FVLzetCxM2Dj3yJOdsL+h58icjfzl+07LNk4USruOWEIP5Yl5UaN387tXq+TDuR2Fy9C3+0bvqN0
R7QiMtzghOavx1yFw9he21pV/SwRTf6nHlsImsOhANZJK4x5DNA3JlSb69wwbN1tMm9zKozuH8+j
iW3cNTHUdFTUipFdh8XcUP940ZvYf3tZxvu5TG9bvLdhAaPxwFU6rXdXLXs00tphFLJ+BcrDXpd9
NyMX18vX8kNdWpOsuuHerEN0l02Gn66bgdI272US8vkFOtt/JDc72ILogiXGKRgq306L4iFBXqVP
7OIwXLAshnIiBfCwkjK/TIUwWjFoDb1LPd3FdY4v3+e6dPcRplMpFSPKKqeg7Y0aIKHiGu0TzJZw
xeKzRHpEBEy7MKXUoGt2f3zj7ppT2pIuaFD+pglwnhD5PjHhccsEPoMp+YO4m65lEkHOFDkKnYyA
Xw+ZPwGrgfSxlD7xNOlY+vN/rbtmgwSh/+ZEm6GeUjpuC7b2xynvBG1eQU7X32THQutTL989UX8p
gLtWbd9VoeVF50V+9Kg5FcA60LvhsmoZwUeXKnPXhmBhNrvtvW6RBVlP+U8hE8d6Tg4+xSi8V7/9
MoswqgHYuslFXK2UVU65d6Bh0A6e72Wln+7u8YaGOYp+CjqM6nhYLSIVqPvZHIAp/uB6/slv5K56
h+6EkYNMhTvvWoqdDpJXQ3cYRtXqvvqTLcgUg/Vu4+frDXxbaHm3D7uyR4AIAIqUzAsSxVhVQNia
+9+A+YpLi8P+n7b/O4PXWOn2PCTF7k7Kl+qjzKqzHIqIzT10B9gGr7mTJiTY8vSjZ8xVtPsEjL8O
xn3f4BKdhSM9U8W31RJND0GrB35volaCOLsT9+HbOjuYCqeyMQPlZncUimgQz0Bv6pExaSefvKuf
x6ISG9X17NRIO+fvPXDTqx9vmLxC5PyktJGKhN73Rdw2fwlHUFnDnsNAQG/HOCbDITAsIH9VZER9
zKRAlnSYrJYjUrsLBPqTRxREMAHNXCGXOj7kTsC74GiAVuNAmjM8O7Jne4gvyozN1FAQGfKyWkSr
iF7Gv4d1UaTy/jw5xvAqNHUtRL+SWbeeGdfqly5FsTf2SFDK2fNhtmfrkNutwGm6IkhfGIYLGL0E
8OqKgUrDiHxm+D+JJVauJ1Tf++KV4W1XenyYDFthCD46bkMn6JaQDH2XH04YdDeyo/TP4BquYqxq
wAc0xpOEyFtKarqIQLqtDYgZdVbcKmyIaQtZwy3H8pBvWPFJZJqve6NSIqb473k4iufSxORAfMJW
gtgzzbIlHpoOG7XonN/B7PxJ5/WgQXpiEMcE+3vuuEoZPgC1W1XC52kJWlqaRlin/8v0V0DYWGXu
HfXj0a0EjkgNyt0SR4NvTxY7ZWfKgqGalV7vAft98OZJmcpxxiPwzomnPMPmv8y5UdmP8w065vbd
D7wnopGbj+MjELpB8dleTzNrfnb29j7bEB/qPUyff0L/aHYHnxwQkp02ZNA4+/Z6SBFyrS5kZYRN
u91TTjq2ticNoA/HPT3U+ApUsmAg5NuvPTG1xejgoxCwy99fzVp4J/DQhGyGlhGk6hFrG76aKDi8
IpGFkp1pmEa3+/XDiH08rzM+wuKTBbGdDqJ8VD2PaaqEEeNUgnY7vMNzrcNCteC2JadtDQZ0nYg+
QPMnE5S8iAcALB2mJMEru3v6MOML8qJJzvu6kkLmU2L4kXu24sNCMjhvwVBxv7N1A7KWR2Epp/r9
zrXj0m4osXAQ0+EN1leCQ2QZPQnjYJrMAE6qCjulnwOOljbGVWaL6EXjGqFqMPyd7gzubENi4BSP
4XrsnhKYSMZplNFPvIw7g9mc1aYAeE9oxGUh3y4snWDUjeRM8R1PSAEkmAeUR4VPiPQOPwvf0nTF
tdp94qbkmOrVjRAHjR7eJJZNUqCt2KcOAS3s1IwwcalzwDi1jmOvjAh+e0og1l1bpJsEH47T5FPI
4nS0XntG4sMkKdS/siJksvz59dexi0ApD/RKGGB1mYR4dn3R0JzWZ/WTK+2S85A4Bnjr8/2FraBG
XdF7UyQIRTrCeOTdB/T44SuRBhOTTLNv7X9H1SA1+eTuKU7WyRgjNHX2gipQZNnjjuqVrfthqmUC
Mt9WmuOfBBqYA8SHiabus7+FT2F5/upTG0fYKwrByAqUnbyYyhiMZ/0Um+h7qZH8GyBLtgI2BOv+
UyxpDoRVlg6EiiDs17gIOz9cJya+oxNkKPSxRb1WGtTkva3MHJlXp5oqXAOiPgU7c0avVIkQah5X
DaEH6J+jpd2xvxS91QTmgYWIMmVMOU633i6RdtoVlzNEqcbd+ysCRCYsrpcOtv8DfTQTtM34s51Z
4CjmR5x13mJwTp5wKSjz3FSA0rQxqUKMfCWiJKFJVxOlyhBZCzcWLPL3pZMB2DFwLft7SYMvh2/O
BVTcq2bSzovQ9XpITPx9LJFdPK/xF1LKYCA1aBJgdvqI9YdoHJuXIYYvItiCQajkhV9vVaIqzMYP
RRDvlP+GbAjx+1iv5BZ6LvMABfGADYJUXpfRB1jTHMyL9HHN7ndCkVgFLn5kKFUyYk911Vrum+a/
dIQ2or0O1GF8Fk8MrWeoMwMoyioihXIRc0YBoyeDLMuxqjve64E4eC98ZURobrGEKprT/dgzynTl
suX521mpVj3nd/O3tedJZq6cTtlgz/JpFwnDWwgJL6aOwgIsLnsiSiXqah3CEKM45jAaVMHZpbQ9
njcvK/bdGLokmV2LH7tCtO6sccVh0vTlyOo4k8iQDoxnqC1u+DJzslth9clffxjljnYmPUkYj1DQ
QD/ZJ2c7V/AWehFzAUK43KKjqQcy1bNZ7K+Qeo6ZTBo55NYq0arYUA8W/pDgYbIEZkwYRArb5AWQ
rwsxbX5Fz9yW2C3oVDGoftS1+REZwA2HMsBMw1HDAVIfV7lzkV2R3lItUQ4cZAwaIMLQBNfisE4q
xns1I/WH0CP+izPeuWCJ2UhgOvTqEBsb4ltSbjZxcvx5rzxXMWZQizKYsElWeIkfc0g02cX6p5/E
OKRcz4e9NgCIt/AxsM4UzVu2YxcLDqXQhcvo9uHrsr+J3h7A6GCXeJJiqgzVhhYuAAm0W1R+Cxvo
/ie1PFdv6Zzy3LpHcuWXdgU6ul7my+SNKbc8te1sDKikQl+lsHXGRKZIYXv+tuK/rZ/21rjGMYzE
9zangLSnA5ksgF0P3Ln8ywBsxjXWbh2jI1hAJ2urdU0dCajeZYPqXrwDUvYTyu2N7SWYi0M9xg+u
jh0sv5JL2QDmswQgzb8poIUVvZZaTjugCK2bVwbl3ygioW80atCEqyOA/pjRmMxyOud5XqYzclv1
pd1Uud9gROhX0VaOUIgLAOTGLR4M/LivoArphZiGqDX5OPVFXwOaZrvzkY1vqe1gGN69OtnFh0sj
worcqqSLBVyvRjNuz8Hjj3PuXKAWf/44zxI9JqiyVs90r0oPy3WO/NjBqybkhqxYdONS0DxsOyE6
cBtxx3FNOsxmWXrYhiCajBKKmgTBazaGKBGR//zaf04CZ0PcBcNDtOe+Aetzrh2815wI6ZutV8pz
MEklLa3+QoekOysYkDA3uSctzvytHyKgJP2vs8v5tHh81lloyXG9QG/+aeecXT98vvyIUDTHFwjL
feM2XzC9MWBYPHnm1v7xAGt+AQbB9y+fw9ZQNIDZPYiP5abqcuzEaIDjyzFBTTcCkI8qtfai22EY
P20P2PF2NjZw0ioYZ3StpWoFg99gWxPC9iwB2rlq7+cWmycGyZ6oxRGrvNI3huXraTtwQ6cWYnLd
v1keT9nlW/P0tb+r4UnHoJ69NkvA3iQgCLXFgna08+LpBks9S7xOcH3ylPgJYz8Fd8HBs9ImQdzt
U+vE+NRbkeNFAIZe03Z3gQE5RFPTTVx9W5GCvWyhMQLXyofDSkQVpSYTXPxlCDh/nEXMIhtuTlLB
hgP5fxkt1x2DpRh1uIBQUwpplrwu3txsIkQTvC3vSxxeWmnGFjuXf1Xhv1lHqC35TRq+DRwMdqs/
xGLUwDNPyCfi3qzuxu5MGI7OnTbhjsYPheefA3vGbrxqonqUZ4bYkTONPZfTBT/YWAWkb1oGykcH
w/W8K6C8brot9ifnCB0jfIYAjjRSldAddWb/tHnvnr8Ypu+Q+fV7iTZwVfZgtgNzkCNAcTXF4jPn
4xsCbyeUQq9u
`pragma protect end_protected
