// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
BLgIvetfK4dSoydIFjmy4z+eZQbHNlVZ0LUX3ApbW4zv3RBS2GjpvyvFNPj1MfWd/Pq0Kz2+JdEG
GyMOvgZggsX9F6CYDUm0Huls6DQXwgeqWJ2k7i5bsmvDeT7g1mJWp1mpL7yFuXq+5eCxQ/4caEIT
VnJ3btPvVEl9RCFfFR4EacrcF5eNdHqIUbuLPxVTfxss2n+e+XlXKoxf6EP6SW03ZCY0gr0eX8MK
otrlEew0dhva+gI8jvTnEwREjqFE4EWdfn6OfAtJdMUWU4GwCoKSQWj0o/6qPAZGSR21YpjdDlh/
y7tDxSWpyi7PJ72cRWGx0bubM1oqizG2D7u6Tg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
/OI/8Ryh0+llm3B/hSWtqEExJRqLmEvhP7tEXl+0LNmL4SlU7m1v3mBSlUK8FgwACBOtpp3wIdY/
Rd3MopX62E4ZXcNlQVSVutYvmq3QMyl87xlO3w/h42NlzGtWem8insRlYpHuvrcjvLKo/v2D9dIL
Wr3LEgMCpfMqlyFks5WuwAhnihYnLBzkXep14jYshNuC5J6SqKOFvRSCgeGWl7AMOlOve/k4mxRj
nxfDMkLhtowDA/T1tJxWIJM2NpILrLZ67hvyYrr59e1/EbimIhcTMEuCgCcqYMslRt1qrtvB6bDE
R9hRdNXvYEgrywIOl8TyHNlOKzBBGhlepc1Qi/qhz5DbnfOtPAytljXkcKfMD15Taw5xOnbU40+N
M7BVFuLFzCNS04Z95HR2ZdZTBDJyPGtFuQIGPMdauAyprOb42y8jpTnKp92VXO+nvInnBjywDaJ0
lnwQtb/ebeIRBi1Eson9bNIp3T1JyFmiDvzwvNMEYWElyMAxlNyysim7iLjMRoIp0oyZYaHY1gtr
IeMs/xYhpcB/8cQaE4sWaHb/8VllKfPUVJe2dZLX/1ciIOmNmbpfEaIs6kso/7PZUIcin2BzNuvB
YpIKDPiNXWKbQ4mnMtg+nSEuOGbvSby9UiExbddTIoCvxKO+F044yKg3B2NJQxF7FPGfitsyXhou
5wVMuTWKz6PkrlfG2l5h0wB/R6ucgWYXdc52YpiGMItFGOoabQhE5D/kN4uV+HUUNHbN6TBklZAJ
iIBUvKsxOiStP+Zo/x+KFHKg17jRjiwFSBS3Mr18J2BwsN0qvyThqEA/DRxbyYivnHCZ2GlkFKOU
ensgHr7KPS0OwYxrkTPMuRduDuaeEYWIRvlSiFNpCZf+hVs+ERLGho1y8iJ3c+nNxi+5pB2xf7J0
1Zn98nmZN+G6Cz1Qf61yTIAySn+KVbz5TEFzYv4nVf3QaxpPJPG4f2y10rCQtYquCvX0S9wao4bm
3KyCToz6c6I5GZwZSSZSxMD8ttE2YzsmRKt/mlsYcxdeiUvqVWX9aEk32ki06Wj+A6AZtvm7+pUa
qFM24kSWk2lrRa3oOZTRa5a6yP9afIXeAb8myor+mKtB5UXJVeoF12sW3gXcNTFhD4I1gFe/pMlg
jALBIZaZZ5IY9M7hJuSvOH+7DdNkWXIPbwCtohDS4191JCMVGvnBePwx1AS4TUGuGWKRpB/rjoWJ
nv7xkcxgbOfuWwehoaGorzwCr4/dEM5lQsW9F/0mOCrX6J8o9yQWa0Mwd+b47o3puVX8dx4RzE7M
JtJu+SWuJTBETS9fClOjO1LfxbiDwtJxesQq1TK+KYDAMP0y6UZ4uXwnugwVYSt+EBTEWOCA+i11
0xQ8iesHXwzmi3ARIQ4rQkTtszyc8GirD0jk9rXVts3/S7Zc9Iq3OJo5/6/+CfqhaTgDIHgDIFT/
awh45D6tyd9pwJvT5+EuA4jeuyb4Dfyl6fJa3SXdLBam3ObaMldFAFRj8v63N1Wa7WhqsONfcd7i
zrKt/5VZiFU9dRV+pooEb/t8YB0ZLRYNin9cpCek0hysH7yvcKUtFVwfrRTyv00Ja8ICtBjpm1K8
QeetIBVXtXLU2AFlY+7R1+vbYRF29ZJZJLB6Fj86fez9+zAr0pD/c6x2YhImENqtNoZ6zsIFaEmE
UYVimsxOe4Fil4cdWse8KsWPnfkKIYnFuPl7nec4BAP803b1tYaXoR7Y8aHGVcZwGlVRrUd3dDLD
/m0DV/Yqx8yYMuhzMlgrypy/KuLwtii6SNbDUZHdEq1XWSiV+P0XzIOMYSvSJ6cUn2kO7IENyoQE
OC0qAiv4uLVyol0g9/3nwjRF/zRZW90xjxIbWd+v8/jfxHHhNmsvdlTzqji0LC07oSV/yN4cHPn6
q4jf06exKtw+pmgIE1aTc/da5vH5a/SsFvrIy+10aLamrXlIAEZR0g0BcdygE9KuRu+G2bJ7r/13
U5hH2QetWNH1OjeOaR30yIWeaqqrJNP1zbjhQKYiD0oRdNDSaBo+fNTeFzSkvzVck8yby3fWaXaz
0gSefPi4zo8E5GG6VEWi65qIqlRVKC6YQ805UIuCSuxZBzG2pKQo4PW4FO2nq7tdPelVAunrmmak
TUeU/ghOMKt/hxNmJbKSIXFK+KxzyyOZj09aDKMLj4T1hVQ83k3q6Kuc1+81Xj0kIG0Ugw68O6Ok
HK26nJgSjcyEWCN3j1cNAE3qSLLVtO95ZMNXE8uAaQHWSSaizRVhBfyXc56ibgsx/SqDKKcOISr+
CwjF5MaUWZgo2LcWx7wz7RPPgPhA+eVfYoXG5xsfUSaAZ8py/b0rxngSttMAbNAdwOo0yGFAzdvO
uh0ep1q+3kl3iBpRRAn5TvrWC6AgS6QhyopQxUg+cJcSt6lHYdVhq6h0s82GsJD9YHr4F3vA9rjj
qhI4xqJJ5YxNX2bc7CVvIW2nIKI8Ucn9DNbjbZkqD2iz2YL0UPCckIbBVMXom/+BZ9SgTFHisgGh
U8gjKAaw2dD2XIG5zAiQAYzqaZws8QTSbbl/MUFu1WDdZ4KqIYZdcblNhBjbsMxir3y9LjTyDwpq
x4XOyGrOfzf9kXjYIkwKERIK81gdDeNUlYkCMEbBVnBoERQUNGQkjfGCN/iMEb9ZPAl7brWUs7iW
X7j/3GjaBxR9Nta51IHggZh1kPAfjWSU2o25+UWgnjzmKfecvTRR4iHsbBvrGBh1EO3TGLfkoFit
N2XbfGU98dPGFJaz82xx1a4WfNbMq0eAGNkf23FN8CEkRWoYr9RhNAX7F8JUOfJze4VS1GxZscdv
bLPgIpNF5yxCClY3cKNBHb232e4nd7qvI0Jmy5QecvPXkx0RCbl+0XRb+GhTToX/gUVxhrWNM6IE
3EJ/TdF8nyJJwlTS3TyA59uJOZbzX5EluuTjtqJ84IBlCFOlIP5FAJa4Tq+BVBKyq4A1nMmNJnkR
Bhz153dNvFpmXrL5NUHxYCHY1FC9oTnO9FgEQY8tqs91XHnMIIj7pRotA3eXJ/GSaJnU7vxuP1RX
8Ym4s45VtQTlZukWL2T3MhUGb51mEN/9KQzbpBumhUA+f/Lc1dPXriB3qdSlIGLZX3aGnVvD4ZhA
ax9G8UsMZZgLCd4Svz67/FsN7r2l37Zm1MWijFm8ipwqMbGNC8glERE6Q7XluZTDIPGtATrCD9gv
oDAY6qaXxocV+Xh+whhASkyMgERm1VsGs+roSTLd5hNma8D/e9pe8dkLGOl7gMSnAUoznZQ5Mij0
hnGGxGwJEgTL/4XfBAqg186rAnJR7hlIMrQlcCRGKL4gaks8Gyh93mvFVqotzfXCyl6HT6MNwp/e
pZyzYsn//QkWa8dI8DAfIT71DTf6XXalReY64FIVvioeOjV+zQHhA297Nt92SPtQtFnWGU+zLYMg
Unt+yS5VYNs0SCqEILtOKyVdRo/7jEwteL7ZProERjt2MMBz78A17LqhB4vBv1wFW4prkdfzo5ZH
ZYPXAOBlykuBd0mL/XSWsaq2de0C3W8qA0f/yWtEnRV61zVZeke06r9u6T+3s/U2cNw8l/V6W54q
7NO510rh61Y9eoA02G1+e8sTklUNkk8NfLPwh5P3PjHfOJPWDVCMS9VSHcO0VBC2gb7Qlcp7ZeY+
bjWqd2zTa7RyZJRSjf9YgYdiCQfY4Pei0xkk1SFY0vbIg/Opt7cHzdTwC7U2l058qPeDE/TazN5Z
0yjS6mqCza8q3aD/hYno/0DfCibhJeK6NrUN1SFNnvHgqqw35wZdKtYr2Nylz+uBM+6g0dkrl2PX
j8W69ZSTJb2RvXxzQ8YTMU4yE7OSQmrwtKzaLa/lPZZBoBosrW9EhC3tfZ4dXoRYgB3K14KCYLQ3
7syuxCbWhZz/51vMFYLo7QufDgpgaF2Ze9q3oyIEIVARqz5H+HbPyEyAuJR2kqqDkUMPkO4cWduM
anYFEgbegklbFUrfWakrnuS0JcDkiedB6pxXLfOQQo2s0mIyqdO8S/yo/iOHsOaMR0v5d9SOoGJx
hJdo8VJ3NWrhoynUActtl1h8cG+OwGgOzBVgT824RdZjF4Nsu/TVV4evbIpRX+dUesRfytv3KFbC
eFsYO8eWcoeKnqEcEvzNhT9UKfJE77hr+tdDbzgz+bZM8Ruk0Wnxu0qeiMydC0rcgUwltrefMX7N
B14Ap9d/kIOYcfMzQcur3vm1X9C7JhocnVud+QMbVXwiLKJNWoooBksZx0l3vJBRpcykXJTAArIZ
a8i/m56wH2JD0bDv0bBkH1IE4QW65F9ds2ujh+58Yd4ah9D3H5OuWYPIPl7nKPRxYO6CMXTWqR4n
KeQmGJtuIvt2fgUcC6Yyh6xgHbjiTgi7nAhT9ole1QSdN5Vyr6uZPJkHC0cbR7H0ZFHsa/Puyfxx
SlWHzr9dhyfJNWLcEhNfgg+f95G7lYsFGIXpM9zEUX/dF9tq5MU+JdWwXwoxTT4yyULfmqyiV+XC
4++N2bPpQRrrjQO4WL+3hZXb9s6TTMzEIZV6ED9BBpNr7cCGEd5ihkXbKoT3DTT/JLvOo3CUiDlj
+1erd6n8FZzfXq+PaC4QgOw1+r8yLqfe2W7kuSNcEFJ3ug01JifY6F8AURijaesT8imEaSWKpQ5x
+wA71Z7qvfh8fQvH5K20h3pGgfOchfOHzT6r5VMPO6fBXnyL3gSpLT9XvIv05UiyAHSMrZwDs1ac
Bms2GyBAyUagYOi0A56HGclu7bvCbhJ24rxU5nQJu6R3WeK6oFTaPB8fsJsLDJU0OgQvu6vsGd8W
W+wCqHiQm7mOt+9bTFE5d2X5Im+9Q1lFp6G7Bc2HPqcoU9kPNQ3Fzac4B2j3Buuj/Hg29YHXQp7y
98qM7GEZdW7N8hRSsbqd2NQ1z2Ymp+npyZDXx7GoxugNQE+iEBXRiEJwTKmXa/akmvWKJCqinFL2
TjywRK77LLjK3aziuXE+1/X41AU5BzQ+fkZvy3juyouwTB5FAr3fi7eg8S+DyJDAIGmNZbPo+j9k
FDRMTXQSsh1ahFjadg+qUjIuHRdTgIu+pOEdgtT/ScSbLeW7gl6Nt8CBfoHz2AmxS7zbr4qfHDia
y9abuG9vCcCFWY9il/oKlXatRsRFoTJDo3Vtcern7YYloWikWOyh3H+112uY7KXwGO49ktTgktci
ajcVGuZ1yujzYlQJIEx0nBc7mpq2PJVipSy8QDXRxZp6v+RFUye5IkbPiNBDYqigUhF1FNmjv3xh
dxr9lLovNGJcfvN9BzYkejEg8h5oopRunNOBxspKZfZRZ/BTontnigNSV8a2LeEN0NcymwIJ5p0y
FEnOCfPbpUEQMUrX8OA2M5v7l77EXZUHo2mV2Ajyz8qwubOYkEZwCbBxmr+8dQWpYQ6/vjSWcplG
DMuKJ73hvPY5+Bt2Gzp2NRRbQIDqv0E6AEGMVIs2w5kHZWU5ZVdbbqnZhfIzip6WO4lUffAjJi53
+5vio36zwfqrc4npdzERqOB6ZXLmyLBJK8QbARgZ8U2q6Ba4th1mXA8soOas4DVrKf/trG6RbKgZ
Txta8UzK85Psjj5dc0CTNMRTST+PDNLX/Z3n5hGe+LFO/1uZUCg+lwJi/YHKgjlInzVYFiQlEYNi
mlYck0R5WDAXuodVMUIFjmiT+grG78Ea4bk3B7ojxd8/a4z+Km+XOqRWBO9Lsi7YDD5oTEMCGYpV
Qc94Y5qWM6zyrFnrLaqNdNma3hiu6s4WDJRK7LWrcyokqR3P92H0xrxiLdYXcAwlrYZ6pXwYrBh/
s4K/FU2oixqfpWZREAWWQZuU/HZ04LSlyV0nhxA/PANmjlWE8cxxGPjRTUuRHb7iXLjb3Vepr7H4
DomCAygpyQyFkH7B2i49yxL+nWlIn4Kzd6xjdvSEkLQZqXZpHe9S2gP5xxCoyr+6SGMM+Fkf1L+N
1hLC5sZ2YG5EH+cwlpurwHE6NDmG4kd8GTLvL/HoGYFkSUX5HD193+hYNFktU1e/fgzqa8o4xTjh
ENjjiCUFsy8QA/4SGhejAV2l5PnQ/GOrn+4WjEuC81/cLtCzQ51p6RH2bP+aCwunwHRGmkBaS7rV
sH3M/R/+JNlJPzeB1IxFM0txwa7B7TBcfj6jTOdoOeVeP9qQtCscf5rMFpcRyXwBjcAkfretWDxI
GWfPNmb4za4tQ9dnJ2wpx/BfaNAfJpkQjUwtoHubIWPc+jLwENrRnn+5OvqAWeTj4e6Xaurc5QNR
e57KmXsAHev9/mDt5d4glwK8gw6Iqfa+7/7EGN5tG/HqePfCCkEfGCDQVT6kak5n/G0yACAxCSNm
OtTj9d8BZoyygk18LSopLe+G0ePEJUJha7h97HfwZ34qQisdwvCXGVR1hLeWFAPwQ27kzbrbDZEr
ExnDTY3aU4VIc8JMpt/AlzTEGucdh8XaEJvWhe0qCMB5i/jiAdv+rwxMt3yAwBNbQtbAUq5natfC
g8TckjvncyxBBIvAVTC8ZMfwPLT35DAQ7cCS0lQfLX7IblSmO7lG46cclLk2jgWYbMlTZtxx+jx8
JxIpH8Ij28pQZiYqRvR0z/SoJPua6JjSeQqqsCKCjdM6wAZVXv8EQhBsMP261bsh+jgfx+gIT97B
6vQn7qJbGxFxHHG7RJ6am/1l6whUShxa6Xk2zd8kyqPwSUslNq+78v3rGraL+aLA8RfiaPYkWkIs
8/qn1/wM+Jtabi2nv6mRCbU/r/QaVgOoj66+CXddygjo4cX9ZNBsbgk5kqU3S6FLiRmEnScNTV6J
zkUT5qCYtGJpSY2yz+r+GyGHE+TEbnnB1LrhDFKabEer//5B2R9NFgv+SXe/IXmN/KSq7GKv5WoX
zxwl1XQsfLenriSLUuuQNP4CPZvj0XQYzjoRevb9Vf6XfMk4pg0zbatnW2kL7ABH/C7pTLrljs4P
bkol0l+zs9qwwpY1P7oQ4w0qAnPZomea9mQR63mpjTceQx581vjl/Rvu+gXMqaMbzSUsWlPtyclJ
Zw0vKFTFm/I7VPazA+vv4jsR0nFVJF+qUaimAgkPsGsteH+D2WFZvX9+Bg6zTXk10wTVxU/XEwpf
UaeA+E4Kl3kxO3g3znRxGk4gjSEXEOMNnGzE7KHSOfPj3sU62w6E6M9rplYdHn5tSJ+XQ+tctgcr
Bo4eUd8zaOw5qMWGjq571viA1lPMnddNPhInpR6swBSh06PI+YVeM4YnQoElWDYvKeJMn+28VMVY
+Gw2SDeIYLL3A1dD5+DXnNMnLCV/LYt6xLlLyXgfSR1uRFB3AR0/iScAhqVU/xTuaOhslom0PHnD
/tC9BHdcNUoIq/r9cfRtbGdLKE79iEcp1Jv9D9U7qF0/tTdoifkppYg6ovaLzcw2zYjdhS8gyubC
vl1tm0w08mrnJKnkfKW8oS3wx2odCX7gYQCvIJX3Fgai26Yn4QbFcPJW3Uc9Xa1NCRKACXVPrXEB
eSDvaoWfyjiG4EsA03Ua8xPsE/FgUpuqSrVGxEResysnOD6N1n9h1VZ2aZnI7N2GyxkNOQZUfzRv
Ug5x9VdLqYQAeq9j93sAnjwwz92WLbEnjqscPbu+cOy+VMUJgDz5HL/42iV00KujPuNV71BMXD62
CP9/Yepw2tvs7uNydKw3Pj1cXC+c5u8XSswc1QTMbWDvidBEFkP0SwSaBkAkRQbZiQSBiGHRagnb
MBXgR01oygQ0zGPrCcLlzf8B42yIHbpOU2rJw6iMTug61zCpdrq6iS0s4hbB6cLvOZH4HNZTc7de
PVgYg08TW3rimbw+fJOgn4e4Oh7JBKnzvyCwyOCWHV8Tcj+UGMxohPOrqhOXl7P9DuNn2Abe3quU
a0fv8kGx9/m97nWrXZbqg6PVtLON6UHWeM/eDGPJ39V/UGDGYvtBfbwF4UjoAtnD6WuQtKeT2499
nAuoGTepHk3v3NxILmkP1RNTngUZFRP413ygx3uDw+sdR4O2oEa3IVCLkaGG9f8KDMOnmhyDVFys
96xQxcKIDBpTW7z0LtQt9QS95HKRJsos+bPO+4o6tbA7qS4UmM2ZpdZyptqNeTLczHus9j/g6MId
X9i321ycrNpzxid9PC6geaRMQ4dTNjGVWuDsfrpKby2meKAx7jJiRsRZDUxh5xLCj6ehr5Gv28Nr
FBsxHfQOAOwjcB6Kq+E/1J60IWt2foCR5hRZH0OD2qmCv1i6RNFljP0oPbV6Chn1OQkslCNGUWCm
OvxjdixpY+LNsIVUPb+6p3x9D4qdc3dzt9NavG3LungYGd+XS7BV1flDoI/k5BHj91zRNVNoXwxE
0C29HngcWPMW4Sovbex9fVCj9+rZLzP1Xs14XpUmFYL0SqfVh+i+9S9HSl0L78M/DDPBPGPlzGuQ
aF/J3r7oisyx+iImmk0rmFRr6CcxcyMam1rHRoh1FU6eWy4eOFBlSxoHe+GD7AlmTiOTZrET0771
TIzTr+9UdK8qoQMYaFoP+zQaGFcst4+6DENP7SfwaN5flxwkkWY11OM67MGCb9a4rXDzU+2R0CE3
Inre4lEmnPyBOb2waUIapMWgaenX5Teh+P/MgYWxjr/IQ/lzIOACujCW2aYFtd7XoXPdNJOJu33F
zKURUuTRsoUJHX/na7KND29wC07C2T0VgLkzBw3MJzhRMTZcb3r3MGNuWLgb0he9EmB4c/RGh8Vc
0NUP9hESq+fC3WrC6ryqKkEeA9LmQZrpLUC/FFSiGcSw0DxXquXwcfOLF2zykV7M1R90M5d3vCLx
f+ykCO917/lckj44HvMIS5SZ3xdA8xvDx+LggrDN6XOJSuObDOlkN8ttSs/r67QcJ9G2htDIfMur
+23mq6Li+VY8w4paRmk4neNpmUJFxoHfPGaPzS77dhXTeZ3klG+p7PHpBoWNheTeNGpp3Dfl5gaO
2txF8ZA1G5OMheqFNGXUi2RLb24kgoWRijwTVeDDqLjN3XaCc/13GkPqkkR787Vb/C8npJwBCibm
YsDHMktUcCKJrnH5Kf9145QFmypQ4ON2Ncpd9g8G62sbg/5ZcPu39BPLw8X7AgQeLYUVQCtRHwZb
TuDfpZ4ra/pH+NjXgmVbaaJA73fzzsIGkxk/TUJX+tewlXnUHLDZfraUoJ+79BcNHWkv3BDOYhDH
7uxCKV9ys/zoJWBx17iQyctSKYAJinkx8X2JGCSJ+Vz6janvlKdqIOOFTaI/io2I5ynzBm5YZ5iK
rft+XcYdt/frOOtm4pcwdR3diubzMvwzVYLRt0nV7Bpdc+s2onhDSCiAwK0bZtHj1kCp5z3KfxCO
YC1iVOVu+O59setgYWFqj7r1UbwkzyjFKqLkzzwHFuL0nybTuOAiyiQIpbhUdbmU8a60qEHcx4dZ
rUMyMw2GpoWTymxuJZNjZsqkI1dvozT6vaJi9LmgeeFsJ60l8lxaHa8ZwRXuqOlpvXrOliNlgGoa
kb6mKaq9CruzGKBaSCn4uymwGrJ7YClsFPwot2emi/TbG/8p/hOPDVKZ+MfVhnKMFeY8nuyngHWz
1OjQOFbDvO2amZMa7YUCKiZeN4+9W1kPhzohvWrxkx8xCcpH45g2VftxI6JBbmbk8pRhGTI5pMKH
vl5zpK7LlM13iZoao3URw+hEQg8eb2eiWUzExBiD3ZgagGuQZsZk5l+XzKXfTOLzcNj/akKPGxWx
JQFLWHIT6kjegtAb7Mltas3UwAlxfV2X6ZCuIMHEXKLySoFP/wLE55oqGGAEkAsMRixGdTBjJQ3a
VZS/R1YsSFYKqBOXXlyqziU2jJWQszJMWjKvgCt4iuUXYN7ehgfJLEW6zCFk4Z9A1XTZHp0VbzUw
oKUlBVlFcBVBnB10zTDuVSVBlGgazkp+sRIxBa5rRVT0BgpkAEC/isyAp+nECa0J6G6ElS5ud06S
gpwP6TSCDPxPqq0HsxGYwJ1tOWlQaMeSFuvKoce9d5sRZGfnZsyrY5IdgN4vg25imKOYNXY5/Z+R
8bSFPbPM8Ol0XRAzJi5Awjbm+fqzIbY9OQDDebfwxlmMh4pHggsYHC+UEAdFZNzoN/qCa8/WyecB
09ZHtFmhpxIJXTadbTwGXUVd82RxK4aZVEAQWdqoP9XlC/Wf2tOj9wnGFLpN/KmdJr0iXsdxTcrl
WONpj+p3SJGhhgxvUsiqEb08Usp1ta9ZtuHr+nskV0aw5PsgDgoAugX+Hx9E7OLxm+5/3mjYgtZa
NfKEwKg9VNyTTb0yzG3sTmCbX+VwIYBk/H7sCUVUTcVA/FlbZS0PFWkzmbGnBkPF2so5eLvBtDiv
GxY9DKpV/jHbnMrNFCyTEFz1zC2K9VCyGU2jNxOMPIqqGXbsdVO+5BHtFKSI2UADMMXPxX7UG72F
qQJDC8I/y3dmzDk2rdPYHPexC8lA96eGiRYw/Aq/0yYT2ZiMZnWo0gVGbot4zqBOOKRBry7q2ExT
0rdMgpjRxjHfKI6QnXAUxzWA7D3+vluwwHflkKw7Psxr2071VvyteQeRXsaAjNrKe22xJDtvnlEi
g+ljqH/NnGEj6tthXhifWXNaT79fbtZvb8GLXgq9cfxjZ/fb9IMoPlMpcONyy5yfkqTstK4GMNkM
3W9ZSJdxa46AHpKVQJeCXT0CkB2DhXuF3Cb26DQD6KJlXzhuNdNTs6Ghfr8p0M7Ok0THwVxgUvtu
qSA6rXMGpPTQmNTzh3PX8+afnK5hqOJI3C+1OGjJlZ28RlZyCJu6T88lGxuVZOwpHddAHQyiCLe7
m8quC3Q0x78f9Ac3L5cLgTQUcsbzdvrmNjJjW6psjJCEy3V6VxqjhEjx0293zOYDdH1CFq3ixSFq
ThdfrDM7JNJv12hgGun/61XCq/dB/H9DKujTZFOqNlpRc5H+b4ZphARpMt6PjZqKFFtlW5D+vchd
YBcFhcNAQeNdHzc3mq/Mb9djjNmCKTA/WjRp0XjWvHHeKyGZF0nIJfRQk6H7GnOvGzoUoP4GEnMo
aWKDhVvFsS8A/XVZHXdHImsYDAYUu653/gY/LwdckL3bdgXo9Rb3I2DsSt0R8Itj7ux2bDi6VaW2
IT022LJREod8j7Y52P3BOV5dACj0/8d5vnyosqghv+VLqQfExPPFe70Okfqgh6gD9qxUOE5Y0R8s
yltWHYlxHLHRxtlJc8BuehSyXykEOVmi1XcCOnCGzR4YSnxkVa2uNgVQHFf7X+dXRgp4wo9h8ueM
LmH6waYk1Cp4AjlNr205za4fXOWiPjt13glqyJo9eLtgl1kjkEVEAUsPHeoNM9Wiq5dp4fUQIkva
v9t8wr3X+avx33v9iFzBciIsXlzSy4rA1p1uToWIhcny/KsUnT90vTbR29Vd9ehNfX8Cv57RtSAO
Ifr6+RkcCrC01bE3yX+LYKuhy18MZQgKs0ex3owyjG1hBXuIU+8OvCDITzV3wXWnie7m2j2ei5Oi
PBZ8o1QqmvsPdEztNUEAjIorw/UWXbh52VDTDqV///hms9L2kGaJ8pL2VLesWh8D8UOnF9I0Lfuj
qhuyphT4sD95zo4cqkpcDriYxitSdRR9ip5skF2WbWFml0wcCp4jg+RaW8/T4oZT2rDXJtdeN12d
m0+/XZI+hIrJpXPXcrNMBFKubWeVbKUndU8Ct4cClvYlD/iqW7viyRnhSpdE+qAgzA3L+sfieA4Y
GZx+YYM1kUqCAPfL81LtWlXRWpF0ZZH1oplo5iRjf65PAAhiSput/6BzOScxqbcyPi0Yam483E9F
pV/S9/rGYaguZZ+9j3nn8tMnT4ykNJu5T5a2oVKZgeE8k+p8HUnGJ+sJq1ZZ3vp8HLLcELlUwu3L
cQbceN9yxcgf0WikwsFOWr99gfGGenm9YW7MuT03mVUXtSQQNXhN6IHpAGaExq/wEhSnJfVuEcFZ
T7IotEFgMwiy5h4Dpnv/51tbj1VvQQ15redubdeaiWjbHE3Ql+JepK2INb13oKwMuJwZ4CDif6xk
C0q+tWg3H/Z6bBhEvzZzA0g11C47ebMZyllaTUBnUTRyZQIeZRHK1vYlOosxeyouafT2V00BLGiO
71dTWNrtqLwWnANcxT7daBUhGtXGro0CNPYn/zz0LYxSl/e5DyUuIGjmlJ+d2VoAhrLmitAvXNcf
zTn1iiR7mJ/1UHWVccJWVkVA1rUsCkpv5xoplbmg3qUg7OHtOASJFDhsBizqjfPDBDekrOMrprHT
0lDR4czdRWtEK990i6F+7AYnBd7Vl7kA+02itW3SKDeYUmQjvO95ow7TfrhKh8Uy57mELEVz6lpZ
PcOdIt5/VnJjX7YUeTY1o0iDgHUzFZjZdqrel/ea+Oo1JdfvBeHrH1htiJwmbSa/5YDwgtCmZAsV
Cu90w2t7wdDtnGkLa7AIk1Ee6FB8d9zdqoLpI0ytp4pKvnqaGCPeveE5cR9VC/t0+FjDRRMUyC7F
o2nJGBFkzTRxqQfUzUV+fCPdlO8+KGK5pW/mM5/3i8SEKX9rS8IGeE87U3FmCLr0FdzmQ3uQwasd
iUTNtcjKHFQxPncd9RWn+KKJ3tESpFnW+0CZt/s5Reo0vwcG84qApkR+AYnK7n2K2kwxC9TSKHIm
hZOUOQSMrOws7KcQ092ukdAPltSeXnrOD/LDb1T3mFVtUL+dfllS/lwVgT44G5NyiLIA0vtjLH3X
pG9Qbxr3as+PwYyzh/AWRBZ4/16YrrNwuMxN/oAv3ElQNOcVspu3haZD2AWtkbnjmR8weqOCOohb
ffJCxfX05lSS3n1bXuY+j00g6UlLaqosIQSFgZKtmFS2r61Mt56wXgZRmSh4nODFt5mueWG6qhQp
J02T+JmqHni3s3B59DbIDDUCQ7+bkZKrXXtT1AY0m65UksuPrBP4sR9dYuASmNz9IeRU6JMvg6FJ
8y2nxEYEkFjfonw34v8ZhhgPCYHqPLnRN7vEFmZGsGqGBAgBBq478uK46BkFPfHN5DBrT92559fc
omJNB5kNab2Og2ALDndsR2MmV9g30PGCWvwp7HthUUUPxHkt20WDp+2nDhPLEGH07PPXGmR+YOQB
ULot+o05l+249oKz/E58d1anktDdLfpnx8v2N5gYVU5Y637+Rpdf/qsEme197rx4Ju1REE9a70Jj
KeV+WIdsDhVrO9Z7+7o57Y+OccIH7KrtpBjiNGk+XPdou88mqpMj6nxEIowdSvXJYqg7z/ZSsSAg
UKPIt2RBLHLRG4yC83OvbkXGObWWQBtzjjNyKyL7ht+CcBZvYptVzdPNa25aHm8uFzx9P1kTXTHy
Hg5bWQ6DRcyv8e6ZRjBxEA7ZbdZQpNFW2tESAOJpQNnkpiOo+sjmXaKZ3ekPNsy89YY2l6c8lFjc
o2ODBEFG071GkJjpb/tgMVbxd7F4gDnJnlZC1FnrFBfE2d4B9vWKZx2FVKXqOvs/JRvzQYxVIo9T
nDcQtL8IqmwjvB0GhqXpWxq5lcIS7r9XrotLh0rO/jDU47ZcGnSX88ryd9BirDrDTgYAuYsabEV9
pesYQN3xPwhqcJyudiIdoN0paUIEoO1PtKaa9b+ul6mFwquqZQaboR0w2XWmmb5mE8DrWPPh5Q/g
cDIobcHuIe4mnPCQ5l87dHmy+qnQOkBQX/Gd5Vn/UyARQvIURZEurpRVsgO3ZDQ1K+EfbAgTTLxP
EjWie85BkAllDx9zqJMyeLima6SdqQ9Lbv5Tc4bqG2ghbZ4UfxjI6DZ0uZNKeSdEzXyNH0sw/B8M
yM0ROJElkHkS0WUQO3Tt9LBPDi0U0dGBy4WAkvn1f4UcWpbpKOGMthvMO7qOnuwsvaYek4uTzbid
VY7qlXJAzNLEvws9WvK/4wReLAroqu6UL/+6hHbI80TGEY4AfXmtLrFb9sEMCGdUUXdeA+0PABNS
e5kOkqKEt8NYCW3L3tvCVcQcD9eTyU5zQCIvcgOZy2qqT57KeZt509BhL2twJfq8ob3iA2q7hT87
9Atp2UZ9H/Gmuu6OTZw1XtEW0i59GrGBijVlnseNnherRAEqZk7tsOzKpWc7xKRxoSb3rQlktvCi
1QlfWwzwST8g6+ZVm67S1YF90a9JsCuK8TIbDQk7GD9mpkgDl6jnLwk2UlqZCrCDaFFldVxLX8oP
3tb5pLSQDzXKdoRCCmuTxuXgP3sN2kEZStqE3rJRcnQUDwnssEtAWDVTN49toXL2FG7HRu72RUzN
u179tGz/FWkBZywceUe+S14kCRh/LkIUBKKGeqkZJaU6hyxn8iw+s07X21YfEpmj31RRUJUfzasG
E1C+dc9fKvRhrhMqf63IlXPA/kQ6UTKAROqXhsE19OmTXXY/I5lMPkc6IfjyUyRlvYZinLJJfzGm
jAxPdrimeoGxvWEOkF7IYxV0IoQ+aUcBmZkbt9T4wEqDs4HlLG/uGO5WN9ItP+M4gnecaSHrk2Yk
lJSg2NxSuBNCPKMq2KbhqzTnfEu4fnzp7jTDhZHX5YOHmHQEUQbZkvFQMO4QJSEWuZzoYDNV2oti
+lqmUMuJpE4FOQm23BLcdQs7mKycOUXdsHFdVmisti/sohE+7ZPZlnfVvXS8qqJ7vIsGN4OuIOLF
6SgLn/UVq1eVryWTKtiqzQvxCxE/MyO1vhTPz5MsfDr/e0YOlxK39GP3+P3jFvi9kUKLuBkzO81f
GujQMJ7JZGsbmmhspCgwKcZp6p0FpktfuykOLv7r+aVhfMeUvYlpmOPHZBqQFmkoY9f63BIs8gN9
uMWO0qtKmwnGxC8RnlE1igMyI9lp40An9aCzlAm5qWXefqSsxp90gkbpm1LF2RUNkhOxRQrGN63q
PBtBJBdjabtzccZ1MjpM6eFslzsLyXG2sW5Yfft4c9HoHtqN7Yu2wr12CwliC7HyVjPuR60UQc6k
bDvGQsMmPR5WM2L03Vwd14LUHFG9IFHEPD3KL+k8j261oK0cYxprlVtfgkW/FRgIULypV/yA9NPR
q0aL+C+w0Z651kqWjjLsTMo6fFgNIE+fP4JZAQd3dDP/Usib7LsOpVlaOXNxCdS7+u3p0fzyl1nh
dXRYcwa5WdCXM26XjYjrnky5MOC40PS+laX+ETamYUD3E/sF0cAeCdkv3ycGpQKx/6Tlyt1tospx
Q/G0fggK2dgoDYlBWT5OWKP/tqAyfo+A+0+sXbp2vyjkNOx9p7vBrgM7sJjBW4dzYHhJ9VYbsTZZ
u+TMXNrr8A1ozdg3jhOjiJ7nT4yIYPBiL1TL1nlf/VGVdNCzlpIebJjZaDY7naxLNCJgCLI6yb/+
abXoA3KFmDCnrZYl0MK3nAUXQEyfOP1P+cceclDJJSmm8XM0yJoh9NojjHFKpkxd1C3tc59m4Guu
Esi3Y/UIOQNt2EqyXMArvF0b5ckffocoMy34Njxawngbn1weqfCYCI2pzn3Emzev58a+CwUu3EJ8
WkDbP+h1naHr4BNENAfE4iynN7+KpCn7pEg5Vsbqx1e9REvBQ7eRtxg9A5cKh/6KLAb9hXRdodhr
kNKds0imfC2eOTrjkSBbYViY92ZZFFV2ASMrfRGdRmzGNVXwHeZV+X++vKjYkCHDGfwQR8QdOOID
vw9vqUV16rbFWTW++Ade7qNnQvfd7NRqUgrK7C5B4gAypDdW+fcOQzzlWIOYOLdeNrsHDFQlnzd+
RGwc4v5FZSmJFes6E2SeAlvPLek0m3Pp+4AbvNrsMULn01pkcT8X4Kzwu9oK3PS8MF2R+/Z1YCkK
4PR72AKZAcNQrOBi5JYYRTcx7eQgm+zaLEDXRMpa3/+rSMr00aquaNefZaW9MAar5bJTfRF5Bjkj
UjZt4s9W73VgqmyIhSZQQvAEgGV3umPFzpTKQQsJ0EAwCM2tYeJiybjk4jgWTE8B56/O/VbZUXY7
ru7DQe0SQS8b3QIfQwXTgiFHFOPN1GJbTzsde+ZOmlMlXC5awSrVm7R1iEDJRaJs0pHph3cymBEv
RDXRCaUrLIi8q3DNADF11bSr1TfHwoXqS7ZkUQNBC3pNfixebGncmolVV8xqUIqscwIvzLqR0HBH
hZp+gdYeMLqDRFmeC56edwFQ4NHKWFGyHLuMs1EZ4MKbWS8/ivQCrnJacStp4mhVeUv2cujayuZb
ESIOgNmO1LG8nbstOfCsK6KMiK6AMZ0Tcjp7yXgNzhEEiSIQ23ZY3W2ESk3NvG5b6uJou79Q++vF
Pm9EmemOtlhgKWcsY0Ih0lBs2Er/7w3nSIionH0+ndPs8+JvWJobk92Ft9X2Rdft4DGN8rihR8X8
CcaYCSKPSaBBwnbFNphDHeSJBr4kLKigNSTN4OlGPZw1dYDIo13l+H7pf3oRt+Fkqna392AD5w0M
pksOBD4notk60wDKnyvtlw2T1DGoihq8KGGcqi2K7HCcIegSl8M+QqxOUP+RIugxdrZoGI1Mmn9l
aK2tugkihQY8M43Np7PzWdetu4wqnKWoR0waIP8J1qw8BAx2XQbSp4gRNfUy1tmNVODt+LoC0d5U
xRYZwVsxU1tLU3+DZFZGgg4+LPd9mFF9FgczYqzhLps5ntWfI3fAH3CsEYGvR6BFOPPI6lMdB2rj
KXHfEiMRKZfuWjNSoN+L8EPJYUeolFHYiMVcr80sibast7j7q/h/6ZQhr/gufHzG4z9fjxng/urH
INbCfdwhmCOIFAEXRSI2vWu+gPwpBmOe8Q+fGITtSOhfQxQc8XBRS2vBFLuBSnZUFTBlSsB1ogFp
lw/xKh+bG0GnVFIFWsn91T6TQlHnM0vnaykYeD8DpQ9OhuqcDnOAjRP8SkXR21bnuaQXK5RgUVBx
zy5S2O+cDDG5EbKvYRR112+BG97gaxBF0P7KRIhf6h0yi9nzgKPQtINgiTeFqEMrIKAcYRrbKByK
9zDD+Q83bVA9JzCYO26PwEipjyeTUtNi0IUHh8GSXyJciOzmiCn5N8fopHgTMLVFgjNmnfnZ15M4
WgE8/C+Iy5xGwuQQykaK5x+oB+AmhQUkyooq1yBcxWuT9zwD+lSx99VvyGrdI24SHym0d3D2M0Ts
16/HLa6YyamAM7esaG4NFncmyliTtfS2p0ww5GF0UEpk8bjqpT+QZm8qYXKqxWoAigyDEa4f80i/
dMOxyaiaRIT9ddPO0cQ2gXYIp3q/+5cUxsom2gFCtM9djsd3Tw0oP/eFTrs5z+60CRrrbhBYIiAB
uVvtBQfua3Gbzwgyb/3K6SBy3tgD0d4Pjf2u1oLtGQwyjBJYn7pfPuwPdghxTyeSBwGOiK5ErFzT
nPHEELomOtbHta8UIsIO/7UnyTQXp0j+TCQAmCEzje9cYJ6frMvDf7SF4J1A6lwyrmyecmwff6wu
+SJSp6uqCkU1mGe9wgcjwOkH5wKiTkkkNOXs/yvsX/vvnVHF5zOm2PNm3UguD1ws2PmP9ieFy8kF
c+Ob3rB0UP514yPze+HRku9LEUQF/ulYhi5vz8ibr6Y34nxES/CzkZHnYeLLG+JhQ34lttJYCahL
k8f1jISb9HCrSh0S1E1qsImxNOkA0/tTv9I/bPXOT1kZ9B1D9QQaUHVnhhtIdrOfFMXTZu6SplDz
nFWTXxjvXUwUImsfR6GJ7MqcJZpNYtbQ4ccymc/csbGXkeA3v9FBRbq2aaBXQCefpoHaohe4ekj1
P0LsT7ZicItzix7TMeuc2vtybfe/JMJnj9o871hRmPpdTPsSIzoZ4ZJTJKPooCoSh0pchQqMUhqJ
8yl45486QYazZPShhNZa+vjtRVVq+KbmI0BmcyhXmM6pKZxIum4/3AVIb94RPrxmN84NUrn0aZJV
aOmR5+KxORkAJUfXEUNc7LmSeijH5xJ5d+smpZwthcHnSMocijXigWe+ZpqpVLeYiG/4QmZwooyI
f/WYZRuIDWJ6vz5sNNFIYIA0TWsiwBQ/x9zZGhZiCQfC1CxtjNu5LdTuNJRMF3ELyVQ7W+XB17fB
orGKgXwpMGtm97pyZUSQClclh4flN5VmTOqufW5XxpQZ2qJugIlCaYbSQyXMx7Y86PPcf+FJno7t
NyZxWYCBsrMu8PRv798amC457fxcO3jtbU0+aqQCdSwbRLrL8ezhGS5BT75ses4vUI4by1deCkJe
0NefDOVT9v+XD51UIZeclCSi0XP39SvfaZ+jqVw9i9cO69ECpx56Y7nhCiF2i2Ak2tMK/ymG1mmi
4fpW2+Qw868DX0On7C2RJcJVB19VmbyJNEnxCiK4FbJCA7WZO8JbkSmrdX7Kn4/W3A2UfKfCz+oG
7o+0Y5+QDUV+MAEC7lbV04arD59ayRwQ0Q+NLxIJdZkjcAZ7s/RKe7Y763Zncnm+97jS0PoPLtpi
+SAY/tVeohu5re0DzLK8PMP5Mie+GQW6Yrw8ocWkS4avJswcfb+igXpIZnXUod1UurF6AgQmpSFB
fdE075aryzRCbVSx6+733kpx22KvJN6JVmTbui4iRmCLAwtd1GUO5Oq1EFLnzscPfoYLjUZVMgmI
7oi82oWwRi/8vsvC48QB3dzhSJpIgfZjtbEbiObLMcFm17wIFp6VSE85d1oj9Jnjc6uPMKGUzkzW
SaLTnsgOT4vG1iEkwZWGWnodlgReubLl4UeDQyn/mJrQVyR+GmMPmj6t+2jhlDvq411U2Int1PD3
dfiqTr+6Mw3FjNP4lRrTkwpu4LR4Bp86WGWGE9hVpHN16Fjuz7lakSDREIDpL6SMrMcDQMbgIQ/U
hI4pIvU554yVOaLIOVVLc8V1H8rL5x5AiWWaKkOdLlXcuy0la8bgen8cR7UTLvQ9u5Iw0kXpFvF/
f+ij1C4CV7+le7pQTLzAbS3RWYQ2jHsBKsdFtem5EWhTiYOSjSgyIOYu7LuJ8A7KSTEDaWhPxZPh
uFJAGqLz0ISDsNW1A5moZAL6ZmWbzQPcu4gloEfsEUyeXAUK4CKPjZQ3iXNACpCq6N3Iohc2uU1M
laubVsknR9lfi2HOX8oZau2OxcDazXZhP/GmJAUt45yUhELbX7ODe2JTJxWRwbpw4bxowBVGzyRR
zPnyEAWOIN3WR7UV3xdq74egRuJab5FRRfzeUP/FxYbzImHfxxvL2pWNtyUHUbsbcckK2yUFfi2D
9rV+ZdXGe1bPWufIg/FiZz1je/0IkIO+R8VPOdNxjWjoTqMDHNJKgfivLFqCACJi+KOPZdwDxCPx
Endg8UgwjNzf7+Nr5cPBM38nnHCenTBhcz4NBON5uB9h9HEYr7fyBIEmf3v8UM0y175XhFFuS3zr
JVe/eLBCDPqo7DpU8kFxI3FFSnbxnBcn6Tj0mDbfJdt4tP4jwIvO0+rmzMAyxX2NqltL1a2TfhUi
Klf5edVzt9VbrYdVdnDwGfeeo+QvDfKJziGN8RzTQto/2CSNdjTrtR6bQbn8c6Q0bcABu2q7qr4t
6lAAmr0szE6fMIiKafmu9lM809QWTtSn88iUKWtw09W3L90Gj72BznnLkp0YME64Wm93rFU4kKMI
0iSBNg0kALAaHT+ld2muK8Byqwyn/3OYVsGc8R919enbvbMKK71BcqogCalIlqik/BKsM9rqyxVh
oQydq50tj05VHmJ+twhjY2PYIqHKy8H6H+ORb9cdYGO5dWRywvsqMynfj9RRuCZ4W81wPTleU28Z
SgI/Yb2fWTt4sNUC56DREHyF93MVDNfAbc2kLW5aQJbktjQQEyvcv7s75BtK+qta82ybfUqmPdeo
ruq44il+luqixdKcO3XXaKz/ELNGNuD/xG3+dbMWdFuYtDp4Mec7qXrXWmb3dJvzX3D1K7LmALNd
FqvBly4Foi2mS/OlrPr2v3+T7i111ULnm/LGWJtTYSlSgmt6UEHrpTvRiTprEW0qdy9Hurg9o3r4
F3ofw8ek+mruGW5zYIq7e2tdtO92cYjyvZEYzaBBBA1hUxJLhUEHNjUdWvTGcbSW6z0qas/V8vR4
GfzmJyRc4u8fISpmW/dztkCXkPfyhBqBlPqC/zpiB+xeZ3/6SqNB9YSKMESFbWOjxC3Dj8WHm4DW
AvcUNFjRtDG9nt5xlSicBR79Ktbvjsto8PwxiL/Vfz+k5DHA5HSFna/8MWPzQHjmyWr90kBsG5Ay
8NxDWl8s6qa8t/lr0xdM8hVSrgz3w9gYv4gX7GHIWkJhIkEVVesiqfMr3EAtC/rre87Nag4f6Bjy
USxRgRZvAFvAaATsjmOi1h/fB3ER0cOpVYr8Ur3NlgLoyi45z0EYw/WyFtJ1BzRWCGBrLKuX23Je
1VErTRJamojwDHKn5Yoki/E8NixD1vCL7lEh77SnPigxKAoAWOYdIzfLqL/TJqNDW+wWUZGTuMuP
JE6k+DlBkyMop7dK9tQ9IC0D5NgcdIixuRG+RjBrVGl2eVe20ajNc/IhKZfc+54J/4Bvd28Fxj/F
SwHeiM/5ea2iCW62b8d2OVKE0d4bBU32nrli5nsvwsZCuCxUyNnj84/6wdlRkRV1HZgbwYppOvx0
jnPKM5xyqNzJxD6CnbM9mdh3Dsawgwcu4aGbFfDEvc1B9jnCgwWf9BeSX/WmYGr5f1R7G6Qr7fc5
f55lYdgRRWTIt7OJUNvjCHighaAZOZeW36uMUzraAtJgFBm8kZnkv2RVqG+SUo+v8OicsSxAiYHk
f4OZkRQXPRZizhT7Q284qAaex4tyZWqprPxSOW9D5gbJnv6dR9iowyw4422ncz8OqCQHV8v9U62c
wHi3eG5+qb1hKJQTCImNaCxW5lcS+g/EAQHJssDHBKRytRfMLkGWrNhyz6iZ1OXGAQRHvflm6yiy
8SstzEfvtIF4BlTZglvrGOw8233vppyHjFs+0+OnEXpWzV1TFFqx8R8xdHdOJtwN84LbmrHubKzQ
hufeRiIYeMlmHN/rvK7TGDmLQpY9gjWoInLHIRdz7BmSuX6oxFP9ykndXtsHSIPAuJ3xIinyFvzI
ZtYE+OHCVQJ3EOal3D/fAsYQ4wjqEAX4wGu/dwFpu00TlIpTJWSjKx8jFc98IZbIeJYSgFCLfB9v
49z73z5JX6aqmiTOilAjJgICLJrYIlwy4u6AV9SzF1pmdHPIA4ZsGaomDjbUa6D0RpoRWoCmDcPm
txMJZkYHLYxNJas9w2TY0oL9FsXbmBmAhjvZLPauhDAAZy7wMSX2tihSmXwXsQAtsC9zQowC6y9Y
n/gBQAw+M1cn3ZeLGZ5uvFLw/jwgT6UIQF5KIM1Ior2VqikodnwNGM9qZtAHD6xaEyxa2f9vve9C
0ZuDVyfRRHfL0ZQurOfU6VbQUpUTYMLDNh4vwh/3rvDv7euiKy18ab+8bT1k//FdvovOP1beHsVg
V/k000B086Y9tmYlKGAfNi816gpoVM0OzYarsSl6MTHw9Y1mVlm+EqvaJ/UgK9r8axanIx0co4c8
sportuHDgwypVBH73tjnKyNpmZ6Ngj8q7bNdpbLCR3eyKUt57FLy7efBvO3AIo3cyNdjhoc9ofeF
uVzKWpYpEOxTO7OwDpjc7WAcDZsymniuIRlOxIpNC3e5vyM/6VkAx/wv1B8WfpK1EK6zwV5kvT+H
Rkbn+o+CrPeYwbQ2k/hYMWmYAZLEs6gI9tJ4AWFGzx61zaaLdMoHaZ8ebKNxTPqJdwQ51sMSrzzx
UOGOHkiYycShE5Uj7lztTtf4dL/jC1lR58bwwhWZ4Hd4UdCoSXRrwIpM4Ku8jf4GtTyOdnKxRD6l
Y6c9jjCmoKiFriTQHjymIOx9YvNGR2Uon1RcVpribwboUTYaw77cANI7HcVCXWown/kYMn9aeKxE
vcl9S8PihD6VmlkGjvBVmnXKEkjVpEcfDA32FTxNtKEgmubXKRv9JI43QOWau+clidaLdcq6d9ud
QBKTQmjRzs98vGTl0LCjLTMABFS9InoKbLfNwHJtQx2gj5tqGqiHj03XsGqHFjtPwKR2Piog/BYt
EZazN9YDjSQaX9ELk/xiLEdEX+i0U9xT0J+6eFi7dD3bALuCS3YAgWZKzfgvffWvBwwW6EqHnhoq
8l0tmYVqHL8gOG6NThVz/hfeG5x/POwwXw9VycxUre9w6VRMyOo3T8vx9cIfaTEjIg9Rm5ygX4Ch
fh+zWXjPF6B18UgPdujyDqNdKr77HSWS6w4CwCyjctBX6kmf31gvvBQSmqqW+i12MbcvNgyi5mzS
BK6ygXTOP4FbHbjO/K494bdFt8KFUBdIgj1D7HRGjKhREYLSgATM/hElqad7tKZqy77p2leXSvTg
FfYvJ+Q/wM87dhRkY/yUQNK7PeV6xLbrDIFTywlz8l6rHjW9Z5awZKqnZ5uJq4V9ruiwaIAPHLQ6
/lO83Nlq8vLvD0YifumMOKkR7PP/80kbSjmTQGoeNsjCF4VTBMxfFOpw5Tvln8h5Glg8rCeUiZNe
Fu2UBkhTXFcsZuvdFyM8pbdxwd66Hhm3RF0rnU+Mb+oqkiKHCFcrctCG8xM+PpS9LG/GhkpxdHfF
WForPcLCaLBbSjX19abR6nAp5Exa9gNkQ0yShRcyork9GjBYM1foANxzHYaTWLuz4bT0tK6QtlIH
NByHlayooPhEl+/qMRgbeUOEzG/iAEjxTYf+GdwUuD9a6JMYJG1S3lWgVek37aDHq5iwFa6WJzcF
TCFTI1DsZCX3vgP/YpwecOq2xm8Q8otSOZS2xGStERV2SnEwGW50xy9aP6dutccdDTD7AOgeb6c0
jtompeMTMgsapv+RObYG1uQ1/RtY9QF3+E1MlyhJy/+ODMUpIqK+Scd1rsgMfdUSoC4NDeokn/EP
F3395JPBVrJTrAmLesQfxP4TrM2Nwlh+W3/QJGOfasWzAOIDl1VBkhzAvRr44keufT7f1htPa/Nw
3sVq5+2R1Ab5h8dw4ZsBz1M46EucFdNfPg60itUV05ZxrxNMald53aEoBcKqvw9rNydOXq01xzQY
uq0YKPevODYGyd3j+cONReeWjX94RevvrsRgAwnsua3cgGvqpLZHCn3qc4Ifb8Z6j/Tcxgj10JFh
jbfnAM9aqGWLdHxj/Q0nd1cfDAPjvO3gVpB7bJpMNLFy+9oiGoan8WVFlLJThwZpfK4Pv7UUlabP
QbA1I6QKIEDqloDwYLGSzYTb7Kia57a86V2KvOcjfLxIm63uONLsfY7KRQ8lYIQU1OFn645wQ7S/
RHYuHsT6DMJwn/d5mWQ0UXuM+ongBH11aEhBAZHdJUu48TgBJ4FNZDHEn3pPB+b5RnFREZs/CHdY
536hxkYll65EUJTphiEeIUuDhJP7847MB7ClHJbMK1cymj5mvtafYtf/yvhn9r0n5u8x3Wxget8f
zvfGN9O4TJy2sMaUA/0vQL5MF4vdYr4K672Wsa50mYk/Hwsm/MbJzfqNVElVZwAAVczgz9ijopJ9
0Nr7gjq8N6+zR8kf4QDWMTZMxBa+sMsn9BjPs+JZpiOobqwc/FGToDQ4/mAHRqpdzibbC7mxTu1p
vpVnbOzIlXIbWoSORIB8geu+5q3HcYSqE1wPHOjJqjS+ga59GFO757PU04zvDjEVi8xGE3JiBA+r
Qx5YOIcuFul3VZxGxDe3eU/hI+z860TTWuNkm0MsraqP+rPoB9PaHWwzXC9y6PQ0IVWNZeJKvwU/
rmq/ILTjXy6BX2w+dpKezjLc7iongXEWQYglVq2nVbuUG5Bca6uzKNpl5eWlBB9IkL7dvaKxrb+6
mu8Ks43VzVOpBocpBv6ovPta4xT4ZXR+59CiBqfJF4HcnWPRuxlkfdR24xJ0jnTsgLpCViaG4lA/
C+JKd72Zmwbwkh3atI9Suf7AJJmvVr/CJgT9YPwZXYog2A6hyuEDiTsgazWLiohER7XU8JPvl8Ne
S5n0xrdk1BX9jWEzvH3tF+vVm/f2vFeJuTrgXB06fq987X2z3NxNHzk1sUMx7KOTe1LLHc7LlHgS
KQvX+g9Qk+SpZ65PX4wN42TqkozsBPaYqUqMvwdqq7xQQnWgFqKlPlBb6HfAB21RYfBZbOjA3w/x
2TDDvJs/mGxL21Z+BRnBt205WD0HtAiPAByYhRGc0LKKtxVP9tHy90HzuUs4HZidRFoD7LL3rIeI
9OyIPqfIbnyw/uhnwOX6uv7BzAvDxgcPvij1VrfbfynOEkeIKaN9FrifmAUS4aKc9RNYQljHWAnC
FbYyPJ/Y22J1dqekbGT6ENRAPno8dslP8puAnvZ3KOEz7yoDvl2AmEXSBKIJyKJMtmnFpF8GWoJV
mV4x83awQ+PwZJO2USJdQ0aZHuWWDvdWPjki2XSQrivzcvQDHMQTbuDR0IvTWUhvt/F6iBeFFuUi
yaJZL8iyQnp3lYZglbF4J5FW9YzaMLqMieuiQNmZHc+UCsbWJfQjnvBcpgQvQOyXK1ZoxgEo+koo
6/0E/E5vbkFJuXDh38JP1yt7x2s8vo8559bNJXGrY5T/C4ESA/Zo/zaNCWYQq40qNNXA8TvFill0
swO1zuAiH/iny+Cfzdk/Ga3LrCR4qzU34Jhb7AeVILypfVOLlKgCxlLVXPV6qQrAi9Qwfsngejq6
e6UBSelAyOfNnJmMEpafb/w4GnSnUl0/rScPiO1Ao2P3pEHIrTe6X1sPG39qRuG6EggOJqUJlUjf
Hfgp+fsvQ748MMfyQ7hCEs2kjKf7VBrVgtmec7WiVfMvQC7Y0KVbxYA3yRKGqgE9dDnZh1yP/OTN
RU0voLJ2SsvzZm4Y/6q2qzwiM3a3vGYFR10qYc24gtOC6oj8xIwPG+RM+mwiWU3PjcMjO80+c0fK
5FnhY0j8p35Ht5XYQmIUaZShpnLaWbtSk1NauTOGDizchSbPhDgIJlS7WZIjY5eR19reWmPquYJy
TF2eyAvNeBXQkMs47hpk46xtdnMe/v/YfFlRWO9hpYyrU21eRhrkuO7BpnhYlw7I36T2GwhiWf3n
DT4mAeDcJi1QQ9VJTOUUYQhBOuNvxhY0ynZuGwf4itClphiXd2xL5c3Xm44jGq6S31t6RdZy5pmb
bUhfGjuUkzEEoDqqeL5JgM7q1t8h1eFnloDGQZnIrj5r51cfIgu0UvnFmghyEqvzuXwKNXiCm91C
EUrBqIQLWYgxUX/rAGNYbaoR0XMc3JCqT+pE85K67Dn3l04QOFH0rzM7s0iEFsiq3dK8nXEZxtyJ
y5NnxK2lVWPIfGdkpHA6a/F2xE4WsvKp/rrCAf8I8uJl76ENWdKzruHSybEkDyJ4rWemKAdW0X3y
NRWJnJK8J1R9D5E1n2xCytaHIoAbgkmZIu1Uq3kEVi3iJSdgIwfX0oraZUqcNgUp7VNEp6fkplir
9hkCv0vDpEK0V4W7DaaZ1n/xlPcBNM3kGksF2cylakU3Vh19+7g/rSOlDVA7cTY7KAHACSj2GpDo
tqGzByWcdbsgdii9zV8k90d3eSTOq8JGvI5r3QFNdpefwxNFf9pMWTTzAucZ973unSoznnUhbsXr
L/h8T/BEGqMMWo4S2pZjirxgriPgEBbSqoDYS+dgREiSiKNNdyEf+cGJ4U2zu/miZtS9ODWWgsYY
GJ8NPuBrOO8J3TTmU/qpa8sWpYqIUi0c0emkIc8xINipDhLdmXquyH1WWhchZKGw6X/HOI4xR39I
CFqOabKt1+AITE/N+QKlrBG8KVQz5suRFh3IJU+qDXpsw8eCIXX+FZiFnwn0Yv2cxKJbPC90lbso
0MmSXwi6mATEMr8x1lrWXg23iSZlJa8zCpuufXs1IwiGOxu5EsUBW0ck+2x8SzAwRgI07F88+1qq
OrIf4FqtGRQqTj9TAx7C33D2dq0WkndYj/OW5NtJkgzZoedLvX1HirPuYwjwmqaR96YdNbU0Gec0
h9tjNg6+yrSChHT44o/n8wXWRUKFemPk+3rzVyMwTDK1LFQByokD5xYGrOiMYdxYhKPoC738x85i
uGzMBx/CUi2yXOsgZ8YZKnKqd4EMfGlpcFzLCX8/VNp7DBwjgtanGqW/1/7B/yLhkz8nSMnO+6QO
BbRobhnF98PEyl/sRwlxa953+K2rz6pUe6Q9Q4dYWRQEHTQICqdoGMET6N8ukydTFzLl3rO0bpC7
qbJgQUK0cJj8wEyxFdl2svic3fpD2LZ0x1U/iEz2ojlreitzqrkScyzk59bAm1JboPWEDxc2DSH7
XPyVTUAa0pBphIhDhrTiF1muplGsi3xkNJvijJ9ExWi/4MfL8yvJM0QfFNYm0StzJ4fUWRdJeVau
kuuN9HjXChqzrC6hG17k6gz6UgpQssIDMKmAda7V1oh6lR3IPrkyJcColqxWf0LtQN34P/3gouE4
d+P9OG5HuNRxufL4S6H5ARRk+EW5xMYAFl7jdj5laMSljWJrbKdP46Aj8aChxtxFqXNOlStIS/Sh
qaLJdRDWT5BVfljBoC5LSfwcWB57Gb+gQnSiH+MzEwHx/BP1tbPOZB2jo4DCidcoY1eDc3dLRwAr
u/JxWGur97o0tphFwEa+2FkCb9W68A7Y/JL1CXXV9K5IXlnzmRf8/Lx5DH43JpTxmf1HnSa211bO
qIj6MYXhWGhjrzXe5PK1sS217KN0S+GUyQORuduJAdKGkgLT17XHi8JFghI4QsA0vbPJhxe2NwSM
z3CF3tJvd3WsHtV7xlcRsd4Jd5EztyZGakaGj01foc5g+IjI/VrGoDpw3YcXrGsCRkYi9xPQvTA2
U/9KleKXt2wuKNxosrMwS4tWDboPMdLEp20eVUFudx9BEKYLN5RX/qop6XGQmf2/WGXtkZHmltfW
90sBt9GhjItlvUpgm3d895wl/xebiJ0xZZ8nQub+VlA9uHRsCEZDJe1AoL0192yN6nnJO9/MFmUt
1ALrAKW4mCOEATYKNU8wA/52UZj17haWslPBgqYiY7yO3a7tBjBbItTUaKXXn47qfodTXTPGAj3i
bWzNm3IVY/noXB3v9s3RVJ7RHrPNyt+eV/z+4PcJ3xH83B5Os/iVeves5pdeJOxIqa1eqxmRwgNU
3/SP185tlRlcTxR9KiK0A1AQdlGflPjmdAIytaVD1EWI0IN95E7rSDNurjc66fiF7WC1GYFp2WQH
txyCEBT+FDGva44Oqe7TjxhgGwj0nyXpMdMBaQK0lmvtfMfwGfNV9BsUhscekfNra5XBijlHNSoy
tcm7lPGmCktLikKahWRp5XEA6pMG9MR/AQws43g/pYCsoXjcqUb2jtpiclg507OlZ7/67eIkz2JO
wSKbFcbMM5GMFejwjm6n4BI15dle06iqn3qU9P1m56121P55KQfVmrjOBOk2vEbcahX69oAY9agh
m+OEaLZH5g2rhavwDWnHT0l+PKeOUPQfsLqWx7PibkWRjouSggVY+Zxiwu+AiGE5KpKbSzGvbDlT
XKMCzhOlmt9TyavI0FdzNnvGUWh/UXM0lBGTyy92Av+mN7oBPdve+v/zyS8LLSheqp97Km4RcSFZ
cl+mbchf8YJRRQQmUxOwKljr+rVY2bYDryruUoMxaeG3uDJwhhn0u8wDO+cckM7rT/zZCQyMpqZJ
giFmdqsFIOFSAf/eKZ0Y2/h4pg25vEQvgAOoO4mRAe186EefkpHbYetMvAf9roa3mw96MZgRVO8Z
l6Kr6/2uEoALa/MWr1o1bRlCruCuE7Rqf+y9jBUKoJBwe/2LfLD4XzGxoLujOUMPpJBGOQ0D86xC
MUIfZHPtrUHg4wn8JPCJsw5Owp0IKfdJPZuSq4nv7/4aFXgS3RJCmJ6iML+BNXUn8EI5eCzkqcpA
/CeF7Sf9t7CKq7AMlMMEinvhh92CwN04RDbUkKv9I2rXpnrtlIghAZzgLOM/5bZk94rRXiF5rS4Q
pfpAoePaYf1vaYYct0rX5bs+FuG3bvqhG6vHZIW4W0p6YxoCRs71m1ZIXGa57uwrSn2hRaZ5tI7R
m9xykR3w8H5pfJ6lrYPzdMqKf9t6E86QqRB8HOHSNEIb0HpSV9qAzq4NsEgDzdavj6w/JjK2xjX4
CHzQc7Nk+FkFqTDwLJXixWlfEdR+an2k2nIwos1pQ0fJfA9DG1OW+Q9K3QRIFOL5SNA4eALwy+zY
GZW2nq4y6dFcPxYkT4qw6G8dwpIAsYDGvHNLaGEfK3kV+nUi4xwK77cZiZQxOsZjjf33MTQQ5DNb
TQeAT2D50i8SXn1gG+q7P0mGPMFVyzO9bXzYkDvxWoJs9z9LlSmiF6oZcx2Mohx5iLbE+umA1Pdy
7uO7abEpx5by6X2gMMOoVIbf7yGW9Gg27Ee2dFzBBAelu2ljqU4qxpfBaMpBQ5EqiIJwo5ZYiarB
lQRLBJ506LHu8ysir5XypjEbAxBFjL5bifJs+jyUVxtwwRu4/UX0Qju9Z34tYwz0uPkbU0hY1PYV
Jmvq1QjaqbpRvasyIJMQIwNAQERe6tX+RsEbSNC9/I3F01GECjUrFyoy5KOzIqSF1aQ4LMwxRLhm
PAfFOvrsYpcj8P7mpiSazWLauiT4auNV/F3k5Z3kbVde+QC5rCf3uRLDGBO52x/cDauVyUkCNlM6
Mw7sOE7SXt2gPuWqcifCdsetQXLFr94TsBGxYljzAZdUtyJec1JK5xFmLNdMAz9AQTvIld/8bDmV
OW8BhxhnCjimzf+CRiOBmx9HOPQhs6tISlTFjSpWQp41o5L1bbykpnshO+j15YYDnERJUNMfNTe6
D2FJY4qw0yfMdYz2/QPfMcN/9e9DLvdC0OIf795lGS/lVDTbyjR96O9CpwCKzM7aZrHhhpvjOJQN
JztuNGildnKOjmPCfw15Hk2zcUFHSDEbhWoUOYd5fj8MepuXTZrL9nxK6s+kyp+wReyjtew9Jgdt
En3Qy6r1H//KC9/Pge87QmjQICd31q88HiBhJXlUoPmootqwKEYSnQRHjfp9HkZtV8GQ01fX1p65
blY/HYrP4qo7waq6Gj1MFhJgQdDzh+R/xVg2B4vcQQpPG9nQvQ3QJR1R2DnUjg265maLRpbGFmZA
paV9FxU2bsGPztoSzqvUS5MFseBSebxcDKToKf3UTl3dRBceRJHz1mw2KrrNSEd/BYVwSST8xmSF
c+f2Gaoe+BRzcQeA2nS10k6fusN+lU0vzvN6aiDH6A53KPvECYbr+QAdQMTW/tBr4sfGdX9+Tr/v
Ifr7CKAd7CIItq4KVsW0yQYpo+qPQyKN8/suyP9S9QWvJ/t2yBbLYomLcPk3hQw4BdMm/pxpVwXc
LWqr0tA4CRQ5S3f76aKljJ4cIRphwHGgcnZF/jh9BDBoAJKD9cgAXFDFD5xqDSmUzuclpYPCkqMv
c+1tVDIlA5B9s9GiSmONBQv3djkj2Wzeby7q9m2puT58whIRLsSysuBeJJZVE6NGCnXKsX85xSK8
t5zkO9N93hh7vIHmAzzW9xW6oWGjdWOXOIiIPbLw+cKxO/OBY40OR0yJoLhpNGNiZdu0eq0Wrt36
rqxVsAZK73V+eBkm3QDvIAe1oMUigmUMbtKcY0Qw8IsSun1dcghnFSPFTuWUkQCm1Jneo6u9Qs0K
ZlSoDTw0qBSehnbAl4yvNpQFmoyHII8HqVDbOtuTsLqc3U5I7fTeUu9zN/fKrvOn3WvkwYVufaX+
BG5O4m8EcA4f4duXHQb8F0k3q7oTtKS2TrjbR863tGxCtN2RphL8IyfjA6X4LPIvOOERANGj7NEd
jYkRm7gzHWMe493fiH2zJsn3hLreB4cxelzR9bRQbyZV2kZ5Is/HlpfwtWBcLyBnPwNPJLdUZkat
HkTdUCx1FD6am4p9hRtRkKZ/QPgUnOxw0sUMtWmKdKO+gTIJnP5E1hF8//P6fpZwo9/+uYBSBQfX
L/UjJaKOzY2Vqm5vlHuJhzE1zZnsVSulTBihAWac9Cj28S7Z1oOCxrkzqkhW7GNaor0aFuHTsbF7
KwZEnYXxgzUa0GBk4hsZY3OXxQahfbAQjy6KqrMEt5VDxNXunTPCV3P5FzhL7cugg8QHHSTK8nVF
3TG3sLpszjAG1g0ywrRb3POFPDmyW1oS1qNe6jG+Z3YbASuYo1s8QbZCc3MT3VxLfo/Oelc6QuN8
7vTGHtf/JsCuIx0NH+vu1j08wgR0BUKZDKHyzmPoFH9PE1PruEW5t04anmdFqgZVlm5pdR2V8ZWx
/pI8KVb4SWoDWd5pAms0xkxjpQDSRWGjRYSq/Vjgm2164DNDmxWok4CNG8clf46IZStsycqkTY/v
CDwev9Sc0xpXHmGUcVzMFmjaJyyiA4q30x2W11IcakOMMWXagiQqh4DCbWDyMGW8aB+wdERMthPh
Qh2vQ9xRIIWPmMzInLFxuWhqHJIz/8Bf7mEGqSLGTQ5peWPS9DBFqfaEqnrh0CFVG0+wuxhi7nMS
EpFaIVckcMsGPjOB5Sh2D9AAdNQmuFKCNgeKEorsfgAA8hbgVjsArBaeJR4rjKNqlIuoUTwUUIV8
NgS8UsMS9CHaO1tee3v4XppIee41ISKv048tySwI0j4kDDk3/rC9BcW6/xGrM1SEQlJ5iMrG1MCD
Wi37ShYmuQ5a5zcA9/rPMXSDyRo1LLGZX783uVTmdYxzVFEKZwH/YtEOymgQ0pe+6valdTvLRUNz
P+ahZ6zAjsoWMOt7mrN1d50Cazm54ULuzsSkjuSjpAFCNBFgWjspuIUqYEc5e1tP7/huc33a2DqA
QmswON9XcWn5h+OyuJSV8iBSa1QxMBqMUrlqBHHGgelyCIkqocoPULNFUo4q5WFzHjjyevgLbEbc
t+9lzinHeZDFyzZNYkxTFFgIzo8kn0cZsepSX3cXurTOIug6IKfYwc2yvSlmhlDKE8tTtjI11We0
lRipnu05CAeKvJmYHAG6SdjcVww421W+blgQwmod7G1ICrAE7Li6/n9R0giHBG7dDNfte6L6/U0v
KcZLCnfffe1gnOxgBwAzUoI7wI2X/UNgs8UDJDYtAo0KU/qKIcnJqFurFGK2o3VQjNW8JNWTqfyd
fC+VMBwjbPqO6rhdE8AdlOlwctEBnx0MzzJ5hCorsiT8r9NFgsfxypbBSygoENVuM/zrImhDsB5E
8wnsN63fPlU7oLvT77t3Mic65G2pd/Xb+Zb7IrEGQcXizTfUi+ua01hh4w24WIHMJ/6Q3VBnY93l
aL/Gv2bMl7STqsdWeKeyjEJ9ilJ5XHaRHUsWms3LChnfswH8ZkG0JQVIqH8r3Pfq/QdrqIhVNCjS
79TfZvMmQyiAp9LW8e3iPUgvHUSc8wVf4PqNR74eh93RDI9+23DMc5LZFnAa4VWYejfPzXXE4cmy
+fR5EfU6TMBHziL8KMDi+4Evowjcn2jHsrvLXMfFwSky/+SbCJudTgRm2/yQL6Q41Lx9zj6QK8Mh
DwHBK4r2gUz8/oJD796ZlX7HMkgykrZvNOT2TVt/Sb7X4fsqJHECPuf3nPHM6OuIg4hy1SSE1W5f
XoNOaoK3944hSdCn9HiGIIepi5IppLkLPdOFNt1AqlXeYjBfdpqSaDqb/EEb/jhro7O3a07YtWED
IGqT/l6Orx5QTKRXaJ7VKSW4uATdDoIkP4MlfvtWc97ivKJgq8e5tSYiwtoEARoaUztpblLpsb++
ipUeV5mV/c0ctppMjTAR7A4HsUkNQbu/cVDxOmeplZ7zXsJAplCDtwf9nNRwGdMDYcBmE66S7ntD
8fhMBCIM0u7RTO98ufRrQYGIOS2qyrmsI21c6O+3qP4KxGSZQ5ctEYNVTxCozdZ+i6Nb68bmA1qI
DcrnN5pUEFZwWHaCAT3Fa4jSPFvzka6eYZJ71C5gSjmMCa+wCBP9qSApMdUMu5r7YPpn6E1v0zLg
umfrivj5NWoj0B6/SGUQfuLwM6CeiWu/XIckRrF/lH+/BH0alM9cj8ewbRNb1MocG7EX2leQEq33
BUZ524EC0a7BBVJgmy83O1+kGZ3VA/2iOoj+ZamJcUn9Ey7N49Ce/EoCrwxmHm/unbe139qcq7u8
o0Z4MAwktXheGx4PRndfc3n9AgZvU+Xd9om+CdLo7ZPZapfengfsU8gTmyn7IH7pk1lrtfMi3+zy
fqcd2G7n5ECTBQxM5ttDmZA7cIdpiQZgquBNprh41ZI0mBA1LLM6NGDRvKTDNYRDK+33dhfQsuC9
uJNEEcBQ9QaSzMj3zkYMvt/DLCL3l99EcUfRRgv6kO/uV34eVWBaPSi+nl0qqhCaWdD7/otWgTLQ
Ie92/jqYWhlrDLKj5np8jC3AWdbId5asshipl9O2MLOwS1vQ77mAvrouoHwW0BaPWuY6jNfTkJIh
dvfakGVnl9IbUsA7CmwKofh1RPcW3SSHrSEJZXUumoImVSCst6oHf2aI2yTnO9ymKPJKrqg2Zep1
XZK8PjgMIDvYhORBviZUDiKLXmuQxQAYPNJx4x6D3GIdg7LB/8UFXnCSYyMgiH95IoWnWQ4EI5lu
mkD7hv/1HvUnHKF0ZMX1n7oc/wKZyKnnTkBuDjQ1ySEljaiBFS+gdcv+sbrQ9wNkFQphAvvlA0ii
L5q1ZTZtlvztZKSgXq/90eFeSDKHr2a93baiHhlCI83BiQvHy55BnCTi/sR2717yC4RIZxs+iLNz
87ipaX8cWk/hymo/iShqWTfSrdH48iAZosATcFlwGZTMtS1lVAMLcW85ozVrxS9sRpzKW1ox+Ss/
H3lpXINdJLFjAEFiOrd15zYr0EHrU5ZDrR91Y9+1deD58PQEqekzyu8PPbupnMWw4yjHpnst/8oK
V+pDf9e7MCH27/lsKlChWMoFPPyVW5JKwllR2eLicPw4RUhlyGzSXTvOGQMACUu0TiqwuUmskzyw
4vtzx+GlzP49Er+aRHGighbdsRHuq+IRiSkKxK8fbWlYhCufnQeGkLA6ealPUL1Et3I/Pghagt3S
Ym6EQwJN/qqDb0+y45SSk/jDSy7cA132x7mCkaUeT7qFqcIPX4R/HPEexi7GnEK2j5OJ2Yk1oFcm
GKSjIhmadSnRrLjABCDlJJsDhKt9Ca2z4oXXUcQtf/kLt6y2zAM/Qye1pLtUnOVjPqwUnSp5ZMa1
9WI4CJwu0xV3QYHo2my1J8II3v012GwT3RC8ipwl7KrWjUeQUbor2fLja+xZyr59Uu4RWt21wTSy
uWqSUBMCGcWy+Fhpcx/dD+17xJXknmWBuaTjbmhyJUNANPLRro2bKN0Gs8NlJZFKdetopt0uUpHs
NJxBoAj1VALgTCHem7qm0zFNzctMuaUdwJnxmN+588sspUlvmIHMFihBp6Y5QvcTj2bJByKyu76I
GzTO/6PLq6ngh86kdg3zX3ytzpC/mgm7Oe2mVkWrG9Dq1akP3l9FMRHyogAmQVi5YjqfcH+JR6O3
pAw6Y8Xd66gM49LYMjqPxJQ7r7XOTjocOs19uXI9GqpWpwc7nf1JXQgab0+6nHDeIjdKJuB5PeXN
0S35UCEDVBGTjqoY22uBoDZit61ivLa8dPimSLhIV8KzOI6H3KD6g1ix3WpRnJTuK/W10zGci/hn
9SQ5PMZpooeaFzJJeCYdoNIXF+ZHna0tuFcxCRtVoNvzf/bOBSmrUwSVofVM0WgbvUbOjMJHwx9B
KoNqkh47LUnHa4rOsSmqf0j2ZPU19wv16QvuzsEZHHNe/ozDi245k9G9HHY/TAW+nHL/3DPctq2O
06UEgZky+oq+ISlHb3cXLRobFZ+W7ow4cLUOH/EkVsH4Hz/CtrBublt0f7pncLHMsKOb2EnlO+bt
W6oZCYIQr1dPQqkBnAvLGh8hHe3Qn0+SNdarrPAAg4hOhpQKU8dIVwNi0KH1k2WvnthArLm7o8ii
hxf7fHUnUyYYDY11MDDO4dnaX/M5H3rX0pUH4eg3Swf0vDUfIFKkUzQQ7vCCnvRekE2LPGZkhXwT
i86nbYGwPQb6aSd4DccuoTxMiJ1PHnkSyTF/ayDpoc6pOwUCZzVvvYUqqUgffezf6YFuHjFMdj+C
1Hcr8fPA3/5rF6zobaebYtfMCgxMZ8iAV6KdujDvXZAQ8GOmXpjzWXZJzL9GpV4yxqAubYrn/nY8
ijKf9rbfMvuAuv31Fe0aTDR0pKLABkX9T+hLhYXz7QysqRvEYmWBESdJtl+N0Qav2/VjnRvfLPeA
B7b931o5prUYZurF2zMACti3M0Thl0el4PZqLDxTTbfVyPaVJM3tg58cIpvT8z6dmdvxXYU88s/t
Nr541XM9WJl9+IBX5v5h20NB8GCtuvTX9Dudsc4UmOHZh8YOJK92RY/GnTQLGqRoiZh6xCXAiHMv
9tvDtE69UjClGjS1m3bMFC6vW93YtvhtNwLjdMBiGKT8sA5D3zd134k/OCMdkhY58vqwoujdjd9f
LGMxSRshRg7AtU/uTSoByvBVQXS6uC1zqjfLbutojjjde/gvjM4TV8b0BT5q5eqN46JLVBF7GifK
TVjxoq+IIfgry6q5S55lFGiN74uUNh8Y17ihJMILzbPN9ymXZDWe0HyzZwNy0ENMe7qZqCJxWjPi
6Eyt1YK5m9Ly5pI3YV9z8kaLPZIezw1sG+4irevyPlJ6nvGnGdIDMVYzP5ewpFsz9XzSl6ED94dm
P6EbjlKOu4wXcVgoGa4hijPmCN8SWxq9WciE4AOBYWEHpDsruUARQc6bxJqcwpoapAVJk4dLt4r4
PEJTqt0Ngellljz6KI1XlDPuQHLsFmzm3gZnMSAqNDDTEpa7qlWEXL1O68ilGNoIysaQHoBWNl3d
W1IUs06Ncf/FQoN9+f85MdXH+P4rmZPZWHOn4/j1J3end1oC/7Te29kwE6MNAzu8l3RJzL3Pn2mD
P8lbw8aO+rPkwpC8+hFbQ/cGY9eptaZyDgJzXx3okFHhJmuPmbFPVzfX/yn5wTPRZGCBZN1fRNGq
wd71Vu/U3HfNKv/lz+5aAhEEoKBO26CuvoIXwuZz5KCCTwxqGDMzwHXU/uRquIJjD6C6l9QsSlv+
jUZgmRwptT3UrLyxtgYOWPkXExyx+EFqjWAcQaRHdKdTW5dMPYwA862MQlbjz/aKXn/ItINVImRM
mO3nlgKG+e4Ip2gYcnRK+oLJPc2a2yTqy0lzJM+tTq38uohLnxnPIY/M/CDYFGv2ja2JBbr3obJ2
74G2uYbkwCjyTbptFVzKaEFLB1gYNAoKw83SvBblq9G03AKPom5+O1MmqGSlCU9QCgrOO0UBkHJJ
HkHKsCSIsdNimh7VnmvAVgTDer7G80pQbtUHHFr0mNsSy0i8NIScqVpHfdzOzYgpZR8F3/yF4AFI
43T46sA9AAlKZVVgQCUozXPbrlgSirV95u8ZzWkyB1hMNve776qi1AhYaqS7qt//mmvZZ6ctgS0e
kX2ZCyjpokXZKYtZYgvEu9k+aj/R41kc+S519Tj0Ihi6AB8Q8uH7BizJxGyen/ckU+xQP2b+pK4N
SUTqozfzjqScEvQsO4Q4HN84Ejnoar4Qg9BQYxZD0+xBHi6nxeChMXthqpAlT0jaWtPOOt3oAFag
FNaYBFctn9CSBWDYNREEoqI20BaqjGXfFDh3buMxp2V4QCf0OO6y/u/z7AaDIa1PCeD7XBJYCtZX
xQwJbWbZkSOt0A8sQxLLdXyeHraJ/b0HjbjXqeVrEsek4UICqfbMMnBZYmmBXlfoDsOl7uyQvMqk
MVpAh++iYFrzQofKpXmbw1u6PHXo0/jVzVRWi/V2jSTjFI9vdp7ERkTfWG0omSzEVEyfBV2YFVjw
iQc0KiUBXQsdNDT8QB7ZLVI38C6x6qKyjlEV++xj5oHUuoHX+2b+1HPLgpsHtKa8QC7KFh5Zm4SR
q10wzP0nrLoxTnlDOwZnPL1esaMcMSoqLosJzmSrytOgpQ8hqkM2JLHC4wqj7Hvv9O9wvM0Jq01s
3W19+KwXk5BV6vkOfrwSCNSN0SQtniDT844DVxNg0dtVo5KZ+ld1tJZlNy2Y5IMJcK3jEz2Piini
k9m2VUhw6KydZMPXTIQp87p9DT+CZSfICvcnMCO0oAE5jyW88hygs7Y2iqi1mX2HQyi6AaCFVIal
Xrspo1BeZpuWwssJLol/uXW1RM5Y9JH2X7YzfJxLlPpBWW2GIsVPNa9BV4086xRUeGk8TTURUB1X
a93+ZS42PyDycfZLlJsw2yli+FBNUabw/yhGAFZg8f3IgL8gpxdreyc5xNqRTdhF66Tek07itKkk
ZsMbPMvH9s/UebGiTNObrYrNAb7YEdD/fa+g9+k6lVZHzHuBXmhkGyX2FmJY6E6ik0Ri1wCFYKH8
utesZkIat2IfWUMiXYEc4qhdG2J5EeLX83Ke11OpIerApoImPoBL/tCrkPiKOAofepw0LODWsoyn
A9zH0if+BOwi61UPvTYYh6ICAfIVE84b3upGmIOIi5AgneHtBSoPQ60VOA7sMA6TwCbLD9ICWNlY
6SA9fSqhFOHbDCYG7ijw936ROBujFMMrmVKD/AYj29hQZIXSKQFji5TjfrhxNla9ZDtlTa8eMVOn
jckBZ68nZRyLNWrN6dFS2URwT47E7yIUp1V4SFjfRv2AuimOc05g4xiOGGyNkRg/Aa+mF+mp4d9X
vmmGx89c8hXd7pFxIHlKEhHePylybV4ft5Wwxun2861GGlSP+XV+JWH4oWuO9bCl6eLs2M37PolT
FFm78FLcqEmakormhgITs6ExcMnwQMPbUn1kAanJT9xnomseidp93GsqbCaQQQ436bA9QRNpVl8X
sxUgahD0JVCQRHeVW/aQ6jHRQi6VbM59Oe4ZUeHNY7fjgVD4cRVIuwDNxf9dAjZReKC+UcIhH6oo
G7UVAwsjFOUzvbEajNtcBtJeeDEpechf3M6Q0zcZmvq4MrD3vKk/l3xcuYdoblIxcqmmKMcEHXQL
8w78+W5hasaPqiYycfzYUakCY8sWbVCLSHeixvMQIDJQUoAf8XeErTSrTd/hlYNgmC6vasgAsQd9
UMA+h6Lds55WINFjsFcq5unw1WjyetgiG0R/kAlfNTf4wOjJfFmY/Jm5G0Op4rs0eTsV+NyZi0V1
to0VLxCFpLoXXvcJ2TT6zD2XFjehnHONo/x2iaLnCCT5d2IB6IkOPdX3tXiSdGoMkROumbiv3gNI
yDWg5kvZnXcVUnTrhvyq3ue91ZzRs865bbUcFjtPS4WpxczsbP6oZY4T6lGBpzWkKr4m5t8pMq38
AHelStDxtQM295Gf05RMMWkziDNbYMSh0fGJ6WcKH+xYIYrshH53xllyOALzF1da0ziPrk2bXZu2
KwPjMJIQ5b6cyZHOZAqx8GsRdN/vJaDjk7PrTxa4K+4Xx5cQUDJqxGyXSRiTuBPt35VwRDrdZHMY
iIcjEae82QdEM1YXiOaj9a0E319UHlgiVtYSOzIGu4eMDUs+xbjOzQoBMyuOaqIzY8DDKOBsAvNy
URHC5y2XBqc0fW7f8ixSKtvOCLZ+MOVqQoNqtpAZm8H1QtR2aL3gVHL4YXBB5wktYzpWD6IXjTCH
OWzXSJrp3xSqdlG/DzUk09szVgvGWjGtYQ86CZBAl5J/ylnGcei0EErk6T4qBOSEMafOzTiK/JEX
h+v/QvbXUAb0lV86AUPjd4iG9FzKa4Zh8FS7yEv/EVNICLDGDFmD/2RFNZ9SKkv6twxbyid2RDCN
DB/aKL7jfuiAT6pM+nCu7heihEwIguvItw9ZatTThkTPVEyA4cSwgu7mrZdBzPHjQw8T6YkZ2l5I
D11MDJiCxJWQdCwAIcCAkodc6G9Apz6n7uRn3mdES1ugwLQECc55dILaFfgF7SPzSmpghTkaWgVf
+qbuiUR211bbm8EB3CKuS9sk6XBEcT3v+3HWU+XGMaaUCvFT2im48C+HJlGYTHIN/ZGwL9hUV+8j
HfXDinXt4UvScVXuz+9WD8f1S6XdsiEQUSEB03+QdhkL/SL13JwzEdgNbU7npbe4wLye9CWmlYwt
NoRgo9tLxhc4vlT8fJAuO8qrslvTg8apaHWj7rHLWIz32sK2weQxcPF7tXmyeJw3tu9ofEy+IdvE
FXwnBFLquMYaO7o4hmTHvmzvJAh0K1NdaJ/NZ+pnm7FOqrJWm4nb2yqBsalGI7kHhBODNJmZrzX4
wh/IaMHGkTKM89zes/MDKkzrIngHM34XnmRq26k/oUwcaEAROLtwqRmKQ8bHPVLMK/zBaLlw8n92
FbdLqMc+cfQvz+lptMugtSwpBTCui+iEDgaW8BzKAvqN/IqqtJ01t9X4+QtEx7lkIaEECl82uS72
ZoxNbaKS9zF8mPt7JsGz3HV0v5rPg3E4U4Ps4HPtlRGgNeT4pUCVm4Q4YiugyGFcfey7BcZtDkT/
qnJFxzV/bUESFUpktNsPYCchH+9vi9AMFpE9PUAqcHA4AJjQD7qZenLHf7+SZ+OR9mh7U08NDa92
WYXWjZbFmzvL1KTnukhbuhHCz1i+HfQw9zVexIQ2kecWZQpqNGsdTAKvsqvProm3QknNSCMfs7QE
wp3OltMMqfZyJoTCP2Y+W6jigS9TqfAKeei2yNzzXUDx8AATUiSHMLGnL8+bTGYRUZXJYMnTC1Oy
sWNnCQ9o738ywmi8rQ1lwP57pViwdaL8/3Xkuo4eOrnsCRfK1WIH6vhudB/ugXCDyrd8HNBpwKZl
BoBZdQCE67XE85PwmLsqYSd5sgduQOVPcl6eqbskB9LeQboT76Fy6LvYvjmATs64dmlrbF0MAN9L
qwiTKsSj76enNkEw3y19/h2694Bc9B66nBz329+J8boAjuHurMOJs9fvXgMa2WPU3k0BWUGk1fXG
JwTGeQNlpeGo6QgD9lIcyY47du1j1JI8YG3Y94+7jexiN0Eku+lkevDnDNqvSa8GbV7nOFTH/Wuq
3I6Zp6Fhcna/aNqbkgqLI2+29+YwmB8bXBaLdM1AcWqEuWQehzkuoVF1TUACe28hUP3rGQfSeaAw
lIvtOH/urz6CLVrNAirxsnHjOkAatXYdBDfMvL8vIgdFgQ8wvNVZtWbtK+gQeiZ4NssGdv1rTFbP
XnISkfpClKn3S8AtJxVnIDp9lhSsKtL20FXZCQ3PJ3iLz888oBFDOcF9aKhC5Sgpu+MPCGTZ8jRq
SAqCq9PRUU60ukVWD/Ms/3/wPTG61NcF8bfMHosxzgGxcS8K05bSG8YwnoAGt8OiVdnOp+5DpMDB
a9VyCmm2yIoKL+MXcWSXGeDXqXZNmQDne2AkuU5uRZk/DOIyyCNFBrvolKP+0UG8SkG4oB9J3ymN
voNjEbMWXPTAiWPJ9qoFwQ7kgdCqOFlYrWSXfdBvAjRic1ExFhJY6IS1tiVMPbh6hw0MIJrvp7Am
cg5Vj6RMp3zCUOWE27qiI12nOQVFG156eqDQ2MuFOYAERH+/FbmJC87pHi2Df1TJyIg8JvjxG12j
MKuEjxQk0pTuxxbkKRIAKez4jt9tqFapl7/sv1mVsWZuRszTRDtRsYd2+jNbMeBtLTq5z6kh9RVd
8YXNtcGwIWunq+XujHHNGhMFnSCQbl0s0x4YrBaZ1aj2Eki/dq9eriVIs0NoTymfJc9AcnAb2BeK
rf2aYsFYx1ZdzLdYkOgrcvSbvEs8AcriOpHuAtHjT8QPqSUgU+1leIX2p4E1IEBA/bBJWO6CuPhh
bZLgDDM5rJV0mjLo11j8ZC0duSjoG6GxHXueByYtWOQDSmBiIAzf5cG+h3QyphKTsVHaR6Qep1LR
aCKUwaUkb2/5X4DiQE29La7dulrcX/9Cxoi0t317cGEF6laQN50AENPrFwxXx6qTtyGoBmYDA5+n
xSyCsDUCNU+X0oERWanVT/Ca8cFY1oZXYemAe7Gm/KLXy2aZPkaNhhyZa30mt2izWySwIJyxQkO7
x8gGfH70c1kM1pqOfZh45DVa3yjMkdn9rAy9QFmhMxfqWEp4aGeyFlPxRQHuzNyem8G+A/244gui
AKbe5BaTomBc1Qgo9KIZFRtElTdMnOdB8d/PhNSIo1AWhIFaXQ6Xg1Px8Lut7+O3anTUslKwpoVS
dUwAg+M+RKJbUeJQ4U+Fb+l//GZd6QBLW3CnqwJqVQJgD3o4vcbcEKxYc9qoW4QeXlu/a19jb62e
KJH4a1rGUqKwM7KWAJSodnUdhkdnXxHZkqIvvwGcJSdaxIzjKEFP8s+5gigNtrW2oemvZRkOlJZd
/yCvwmtNxJ1qvpn/nXKJaBoXr3lqYCbyzn4MJqsapEKITWkoK9tk/vYJcdx4eWGqT9U1CYH8NXiT
omqS/BrrKqanzPA6NeHiGjDkAyIzvnrqvcbfLhYrVEAR1JvymmjdeVoa5LLKoW01EEU4PjKBruoO
EP9V9bENj4/WDU3a0iYufEMMjrBNSSVUEZD7djyRPwQJFRCuDF8DVAq+Utiq1HwlUC92OqnANdob
K8bJhRFkXQuWAmkbb5C5Q8zxr/v1wR6j5uCyRSRgxkWHPCLxbDKNwRsjcgjdG5UzRPbh6UG3/jQG
KMigyXVLK8gjkSRl3d9ZOBpt396Z1ogl5io4OOOdTkqX/+jTRdBRChWTARUIKxcWaIlRT2M+TKtU
K95eXfEEDvznqaW0ihvxLX0YZ3fMLZywVPzf3OegcZ0Ol5xkqScNOkZMKfm8GsA5XQ1S+eDuZHPK
siygek4+TvCThfvGsRW1fEdTUjW66HEhNE1tUdhypzAORBkw4vdYL1I1Qw7avYttCinrTYImwQP+
iRpWUAzrlNBjZ2gPBKr1/OQSPed2wFOaxyTlmn6aitYzr2d6QjcFO3xiRl7uO8862cJujIQVS08A
Tg25tCn4/FqiiELYr1hPPu/oGfQHckHOfMBOC7x8HrSvVhfUn7gxxOCpjMpRO2u35DqGhq40EKBi
+YPLx5sMjCx1h53P7dT7ZrdCpUjPhcmOtQxr80UKb5+HH18j+c7s+89tcd4ELShvPzXOow+Chyna
K9QYw0sbMG2ZwqyC4QO2PW9dmYXyRHXohGt3F0u4jd/aZ1pP03ISu2aLELyds1AsN1oY4I5VVtF5
PPqir1r+naI8THXwiAbigOlZ+A+keZrZrgZaY33ZTjWttxzlttAtgIP77/LaXeowx5PBdMfb/e1W
ClSjQw0zYwdvhBTNlB2xkHkr/LC7TV7WQPn+bRZ7yuH+nioneEwI6ilLKyhH8k1HmGgBvj2ljQYT
gIZW/sLrq80qc7L58LLl2npSqbFC5fbFZ0dyDMrUgO8+FoakNpR0KRm7sMNJYYDQY6etQmGHbfwb
jVaA9DfO5bBitA6w8W+ds1QzenztZsR2sNu7cqJ/SFWrS9eILLT37GVMDWRxpKyLhPxsGRhtzUo7
hjBMPMXCJrb0VfYyritvW2Y3i4IJhQG0EFzQa+5VqEO+vn+BByr6X+H0wzgyLMuYBgDkOGvjksIU
7IdJ5MX13/V2mozY/u7oqLGwRVPnrMxqSoyl/d2ZQiK+N+64RAXVXdFGG6ddGKhXI4DbriKve7+l
VaNRo1RcDQZa4rEb/NN0A3EtUHbBf0bNPkEQ9a0BAwVq4y83kkFc8vG8mk2CWlp5+vogyMzUQ35p
SCz4wYI8h+c5wzR86Ri+5f2uCC8/T+uYeMo4nQBJRm+NKQ9D60SyJfybVL66XncAQYfBKWFH0XSm
CcddmL52F+i1FngAOYbU8cIOJpFhrxtAe8Nag6rgsRoNzvIOaUqRKtF+XijfiT1zn6uwtRZjqUwP
5KZJh1lnR5fTgTm+b47K1cPL2RQRhf5VSsRl1w4LuwNMngeZAhlE5BeMOZMi+auRaR8KGMw96IU0
nUoU/Sg67oDttRRmzKYgjmymqb4kvOQ9veCQIJ/KzLxWVAJaJF7tKa+3jmQhW419yuHZDzlqZRZL
pLkEtn+dCE18hjLCrmWWXyWA2pXD3oEffRDccwJCy7rcyCWcaCGzQkt1Hq5g61oCAKLOqbDiJGo5
QcaUbgSrvXv8PqnzCU00XS4PzEALXAONFaoaLW7TfknUdrFoYHcOoMfyw4SWFwzjViaaw8Abo3Ge
7EeRVEG0PcCOtfbG5GSvw4wb3BAptoXheHBDj3VxZymHawucI2ZFKUl/41mDWSSNbF38e6EYdzK2
1nWZmnZE7NEO/9rTyIEjYdFPOdWUnTq7z83xgHr845BEz+OvPfdxWkQPiAxtCz972T/mtuzIb94O
38mOZ9YJIge1H1rJyCPFrmOBkK4QZ5iBxBFjozw9L/+5lESrnmErpeEIDBV0aWzxbjg9hqqBdlFu
NdHLlUiqpB+9Idw8BylMjLlUnE6CQzmuXOHHj60Zkrkbllu2YDyjXO57pSObPRp3GsQ/ciY0ceyO
/TjA8ynsaMhlVEnnkLTUTFLRjrsg/rNixTxHaDB5QLXh9BTQK7daRV/8k4/Hxbc4TtuTFbxCTNQk
y07ssheR3uglEzHIc9HK6vZ6isBvFzNif+Btmi/qtKcWyc8HGcLJp2G0ofS1X+EIzSvPcvGl8SPb
04JNyPS4Kkb67ICHdq2Q9EirmtVG1hsl3G8jv3ajXZwMhjyT0hu1+JGxNrI4G4KzHIBXT6Yr+d9l
ZPC6Xw2vzTbSFS8n/LTE4ZMEYz4VrQejLnQ+DD2vpQNdgb89Rw/xxqcP54zEPLSjSvPXzj/CIkOh
FVUbu4FPUem20PWKO2u5UOHHhAmj8Cfmu+uyb94dcNRMkFQcg3IGWR58FytqiJzpqZVmO1E2xM+b
ZHSFA2oTRTNmZAqQd1M1Qrd/vagMosXb6kzo4iw66z2J31m9vuxskkTRkc51oFLxeWnJL9yLzkdJ
pcoquY1KbeRI5Qi46YC/5fgE25yH0ENCdxgKOq+g2ES/kqKYBXwf4S/k5stQIRt7PnKKpN80WgyT
YgucxGiIyOtc0fbOauwepnBorqSFmoOPPwC/b4CL5FexMscmX+nOQLkZhIsCa9JMdY/QG39BlfwN
/h3Tk/ALlppTzynoS+7MG4rqitqAfA2PtMk70UrOtM2ihJJaBY1Ajv4gP6wkI4Fxzs5P1ZO2i1AO
JtsRx9hPxg0E/pYQUMCjmuY2rLiQBZ+HQLqtP4MKzDxCmSnqlpSMo+pg79EbJAPPLm4w4UF8GBdV
9j4MgQDMMuw1TtiClTGz31mCu/N0C1EziliPX6DCNcOaxC1J7sa1bCR537q8jo3Gwsn/K66R89v/
s2/jbY1ByRby78htqbzOQ5K+DYkPZSVI7qWjeO/wzOzjpKaimo+lKPJbSUG4OTJWds4E1XV9uNgo
1H2F/aHXCcjgKO0++faqOWFO75LnP3koZbMAbeY+s/jmU/VCOEGpKTbw3Kq8CdGcTTLJ+yQ7G/++
ncKk8xZYMtOArZ0wfp5peLd5lU3QaPRQkSv1697iDcz8tYvfYRsIY1nxDaHbgIg7aC36vL5oNenF
E0D5FITTBnIIq/QX3SkcKTckngOpUaltzDQ2UeKFwlL7vQcjkFN3AzWP5pSixxgJKvucTnzBpK7u
qrfXlMiORvUiG8Bo1nA6DKgSnS0OVi+lYFb0YJmiEvPFAsywyA98/PKnfElQPN9pup2RjVXRE3JA
kxbEsL7qYMLBv6cLuhNinXB+PqApv9spT2EWPZjmhC6a2JDyp5DLcQj8r6rIatp1Ropmg38S3s6M
/u9rpwD/ke6tCxs+IHF+acDJQ43H14Z8plPgfcthqwiVLA9FKBo6v7lb3QUUwmSDuOEx5GeUFMl2
9p0UQnwmrrVUhxR6fGpqMmHNXXIhtp/4JEw8i9PhQpt2Qr604N72epkDc107dqnUv7fLcYEGpOdl
jwUg+F9ftZUMJ/4jtchpwrJ2LMIG6V+VMWf+QwFdS0qjeB1hXbeD2jH6Potfck2SvYgt+RyMEFCw
YWktIoiSJZp+8RXGfxgS6JFF61tc7bp3tutKAeBUkhwXsebeyP5EStgmmTTlaeSda9uyrr58TOdP
t5X1illJxDdQM6Qo/KEt6jq+NQEMxla4bb1uGrEAeJ9buHalutOKSa3ffoYJ1cJMg+WEDRrOC9Ge
o6FGb2QolHbYbYlT3nDqoLl+4NLkw+uxV2q6er9prraT2KZiJa29rhKkmXOQB2mvOT4cpU5n2oTo
jfOkhy9rqY4TLY1pmJYXaVhEZ3G0dPMEKFQiCkHddvMTVh91CyF5KKq1noSU9SX4tIA0IK9rRq5q
qgktbpKqceGzl5kqkPF2RjHrRjZxYro0zkQM4GUexJ8D9HaVjHgHnzmNjEYWeCxZyG/YPk1tWQdJ
UO9qE6QR8EhbBmwXmBfcDAqzp/ytZIl07ESW8TQsnaDMOCqUIBfW9pBMh2QQ26poChoIgu7IgpMt
YjnaKdwyQR1CHgPYg1uBUwt6CglGPFGQlXVaeBnfJAdTuxl28g2sfqX06HCVdR7sglA8NEHaMtO5
y4QFlvcS46CS57Ld1uz2hVrfZEYRUo3E8ok4jYKlDnxDJEm4vaoaS4z5HvmBy7YwCIN+Pv9DRgIr
X3Ivnx6lK5XyzgIUvZsLCQTmSTzdiMz9jzCZsKz40ydGFwCIb212jUSd8HeLFMkPAow3jQcTCTjI
yOkgBRts1K60bsdwSxu3E6r3KXjJaL/WviqylE/0RtLnr4ov2uNA1utVxEqZwlC0D4axWQkPivOE
aDjAkZIeTGLaTFW/wc3zMmuno25m3khUDk4RyYJTDsJpEFNIgn3+JAkj/5i2trT1whD+NQMqw6F0
cN/ptTVtB4B/eZJ3p+0k0JAO6FCoks+Al542CXQZBt9sFGQJGLLAP29nhoHXVw6jY1rgV0bmLuzl
MfzdZHFLm9BBERi63MAmuTxpo6rSHHPKblXAqii0zFlikieCx60SlznSAgWJ0a2i5saZfBJs/BFc
71GKreC0BwCxyMl5cxZ1minapy69x4wnwbalpAZAiaxeoewtlFQWWgQmOccFFPssbnrzM0aqrJz/
E3SABPU2pE7OF2CKXwCmvxbWiD/QngYtPtRMHp55JAqj0nJkxZyG1xW1CG4WvilvJ6sZKOQuyeFw
BTk2VeJCEQtOye/Mr+aPaIdXk9QmNZslSrsPlhA1ejoyUDfrT7hvPuNsRB+HCVi5eGFt7qzRfNQE
iZnJuXOKoNlmp5VsYOyLGg/SZM3ZL3c9Z6GwfJHVodg6U1ewzsA4pp3Rnc9WjCwDwti/NsKXXVL2
ad7gRsp0nVJXgToLINIze7s06O8Bn1LtsOYeDlwdD3i82g3Zuve3moZ8b6qwQMhVz0wySwZ0QJTz
7EZikBY2Wzz6JsFmsxm80GATamXRPVGBBOG0s1L4cJulXANeklPUP/cpyrq1DhcfE7nvVg1KAaxs
I/3htTwDmdG6scu84Jj/4agJI51LEPXZoxbKxtZb8WLmdZ/s6/pvSbW40wpZEtTHYDhlweoEKUgi
zDX0CVGmg3og+D3QMlRDtS9034jvf74aE9/OdBX1XVg9hyeAXJDZF6zL3iZhBPLa1GpZIA/AWNtG
1Ruy3Jc61nbWrmpyQKt8+s894T7J5tPp8jefwIctPHNwJEhHHsRA1lHtMx0FBD661Q+16AayCQmv
WcJdQlqTULp+U8VxqnGJKDa0OCjhEwSoo8gpVTbW0Em3paNJqos6TPbUTEtmatrqkBLIqXWVIt2W
7ryGN7c6pvShlESmxe50pjNIfsVgejFOwAD9JJKDgE7XPOBj4wd+mo75hBnLR3SdWEkAb2JfBvY/
gI5LDysYfblfyZAILsRGC8yHjXBNnTRzzNhiSRdpyPAgjux6K+Yk/uuWn7jBh74Q8qq7S026r7tX
+b5Jg89oarFVeEn+xnCzt5/Cp5DNNWHcV+lQEBzhDDOlOO392H9MnRt1WpQ8L4lkPXnz7QhBfrEf
lM/SRaN9JE591m0zYLPSkbzcWKnhVW8qcCREkijEC0PeSYkUOJ/XT2ueB9SJQVTTYgGucRCzEvjX
7P674nieiIH2jurSaeS5Ipjy2YC0kycwIKqfX8md4nVOfiZmR0Onk3faBQm+U3CLv6epvRfOTz1G
KyRFSC7JnUVuzvkwvyqcrDuurMJSYN8DGkcTniYE71gTbmLKobc61joBYMgiLSDx+xfTWoFsIefq
LJE5nWrxB5zlQxRQlk6CAxK9NzZXsjHmvPCiVPN405xPdak0OGU3WFF1VRfzKOk4USGnEzYlU7i+
kn0A93aVKHk7L7vJ7i4egYGgC9cWYy3oQlFNpZx5TiuF1b44Xv0823+M1oJZS/WdxqY0knirI+VM
AyfOSWQvvwAIklNgGLhDpJWsZaWVeG5a4H+kS+YdwIiDDvbQ8lzYpq1bzUfuzwGYpo4MFnlFFTuc
hohHGMXCC64t/svwf27TD+hq7wHfdylx7R5NNLbfVx5//jbvq6FE+DMd79gW8nEw0wD4hoB1Ur5X
fILtobCPC47zii1SFZUasSpW5xPL01aUxOjxQfJieoOTaeB8qtvDgo1bvXb39/jyHQ01sSL3gBGg
pa0pkqSBgmZUJedaUmGINAoO430AYcg2wpeqbn5Kx49fISfqMCmY2WChJRuBnqQz09sGgGwmeXcN
u6Qhm6mJjh24nkhNf518ltWUKsSQHqrk+N6/YEqYYPeb7rLaxxYfyUAwkqqfcz0bBBO/lW84Xoj3
qfVZuPWo8O+Vg6wedoAbWb/CPpnHhtNSMtSZI2OhCl6pEmfyFIKui5eiXBtyK9FZKfAwh3aVVI3Z
IYxyyICMm9tAwXSunuHIfwh9Lxr+6ZehxuSOh54Qy+gONsNjzoSOqWH3OdnAgW+Hzsj4hbr8IHgd
esSjNMuvfwCSnaIA7c259vvfTtiorpJy0NyI8kGEqlBj815MGQ4DvsaBDCYynt5k6Bdq6plE2bGo
zUGPCee4tG9UTop0ZsGlXUllgmJlnxiI5MBxZjQbV1Us8fidvqvFK1sG3EL7IGD8QiTTGKMIOzfh
N+J0ngIf6gUSF+jqQhENIs+EGh/a5cSj1YMLiWZRjKnWxVgzEKy4BrR2toVcQLQAkIE7zZqw2401
KCt5dzu0UbkW/Oow8tayiZRckN3aM5nPzqnrw+wuoXoauxjxYMT8EuUKmtle3KdcwMYFOs0Ygaf8
hgLZ4eqDnI+fReDbcWA1QY/UfQG5/MszTYjt/tz6HW/HfsCbPgKzgwWUFzvIym4Wl4+j7IhEpI6v
ucINDjXf1WLVvfuQd35mLfnIWI4bt6t5L4U5D/bkoDV3bsEjyDnpZ/IMDfH7P1EFmyTcgllgao3v
ofNzBqpgPMhYu+uv0rmb29hHE8WUYzb+X+o2COxOhtCgF5ylQOwQR41VoC9vcTtuq6G12QaEl//k
0jfoxp6vN45Do/EpN0YEyDTFE96HokoLf7J3nwjEXzMsBs9FjbST79QXyvZpKJoURJYOyEv/83gN
e5OEz/3+rW1SIm3bFQoOHWjDgpw/hHkdTFvEm+9bMH2Ja8y5t1jx6zBzd/qmaqC6FENvuRd6aLEd
BCSvF/zHYJwwluAdhab31X2oL6mI1S1/ev6nL65I6zUwROpJ7emFyjUlH3tbSoWfcqe62WwmciXk
qusryGVsLxYasbBWyTSd06pbwzOeocNKKzHNBPo+x/oqhgZfL+l6Kw36dLVcNUdXJsYP63vnObFy
yMf1Yo/3olwQm3DuQ7Ic3IYR6CTXoyigfilvAemZrf6mxcTpLoe/vN/aAMTwm8QaZjsvCWfyHf9s
ZTr0eS/dMJMVBUHLmfzwWI7/Q0RhXs+PtvecmTAPomSHjuJJ6rzFmtH0AgGddGgQutq/PAj8/1ex
HCBRe5M37abDcOc4rfTmj5VppYUFtxmdKwkIFYBbOHgqb3motvoa7gFKrkNCq869SMHFFywI1F1v
4y6rs4xyMOviGDu/KyvZQhv+w88ttCXnE3eBUSsjq6tcpvOCRDcw3ei8sAQTZoiwJIjuXlKrq6J4
eer1eKL1QlKS+M/DeQG3h3x3IJC1ElF6HOgvDlC1fEeKogRyLl0gwea5tKCKqhLuRTIlMw8j6gPg
pMoKdbj3+GLwlgqLe9BEeCbhNSQjve+bKk3K9n55LmbfJcv2ArosZ4znstEoB9THbGWHH+eJrkL3
34NXLAEoOLxoXlaee6u8eCqlZ+CUr0LZE9TNB7tY6NCn6vTzlHqXtHXs+T3HshKD10N+Td4LOVy0
4A6IOKbB3JYUmKEBFb7OHpHPHzaMpVf4djn3viaCook/ceyt5SXsXdVb+h4L7eQfi2Ue5SfQpodS
i4PtR+2P7MmFTV7/xNg58Ua2/oqg32wRGUgX5IvGMOMGYuq0oIKpV/JX0Ftsyl30xnTSGlB7PKz5
lJ/E/3AbJVQF9gtxQ1CkJtA77X4JXq+Tb7QhL1QFUO7ar9BtNN7TmJoZRfodHggv0P1DskdyfVrm
owoHnKi1sjC7fgQ9FYigt9qX2RAamKJVkwd3eLAeQ66rtxIoZ3OK78Xh8yusPfDAwkzYXgAMDOpv
Ku7eUNQGyv2LHWDmHT7VD+sbzvelW4pLhq+7IUrMVNy2dZZeeg7lvKi1xBerHWH1oEvkFQIZgTtx
GUw/mAYg0doDbUxjB1JMNcfuvAp5e/nxsdyQRBIKBkX5NeYsYgYAsmsnco5s7iArTQPxy39xWGz3
FwWLBGnbiXfSV03QSuFLK+3w8kUu97f5m16Wf7WC76o6HJtLHKrFBBQpAyqjKYHRf2zIOSQK4KLV
cjlriEBZ3wo3LLMvOkD9DZjdU/NXR7H9NdKOKTN9V8N33s2t3liA4gSEmxXqAQLzC+YinbXl60kx
9LmOwyU25Bd31pw1OcSOlSt7Cw/sd87IukcQ5YIZfU0izM5G4BX1m1fzEOyxqVI3zNKvWQOBdC2j
BRhG2T+/1ITPSIkMYEOzk69pF/JMUTJLdrrRxtOSzopPgLiBuutyjprCSF4d5N6C5dz9dmSapL70
P/UbhPuh+SjVSNwzNRGU4UeeapGzugFDv3bTvhbWRcPCOrYjPnXqXwoFfpYSrNhEqwjGYlXqAZvz
itIEV2X7+tqVcLzd4wS86Zss8dzz7NwS1SjwmvfUjo5XDLukF5ZnGx8LSvoI9YYiUJM/RMejqeq3
9b8InhUaKemjS1LBRHb9gDzm1lhlvp7H/ThO6llsI8hKP1Hfmyto9wBDXDH8QALAJ+WZkTr16m4i
+7UNNOCOcRxFkwjRcuUNtwen0TegewczK0HOJUOJPdLzlgsTjmWcAchgu2z4ofsVeWMks+avcXi/
LOZlCbHl2Hmho7weSgvEV9jzrkhQMX15KUQLqt2hA7w4BD5UoqoRI6OujU4yieoH9MZSGneXogi3
Pt3uaDU7PVYOemCz8IFlaO7MrrSC+nLOX/n/jj0w7HuGL0Xb+GLsAIDEHCcvVJ+n/Pez95Qp/SK5
cw5u7H4OFt1gtyCGeua5NbwyBPZxefyQGbuc6ifWGP1fwaS248j9O/WP8Prg7oWh4X5EEEaCn7E1
jVMvAfrmsxzCxv5wp26fqeVhN7q2FvxVDjjbWpqA5Pzc3vaceVBs3ImNBtxfRswyiNjF5zy7/Mh7
+tvUjg8b2OxK0lUOlI2z8ifylkjSNTFOWFwihsyr74wyWo1LskFWKnYfE1ocyphBNT484W5N2zWT
Hv/h+eaB1JZPWRQ21/hLqwRdOwygirQU+16MFpl0HPMm9yavMr2duy1zyCa10ivu3OscueeD+2Ri
LPFFgrPMCASWyf2vJmla7/5Ph2qHzxKNV/zjUuPU0mNte62g6xkcALK7DnrWyjCTaB9t5RQQZUD+
27eLnREcMtqY2L1/caZVQZKtRz7l8Cg7lNmKfDNADZ6/iQ32inbdf8YZyP87gdya9aQKA3uSySaE
ordxDWgUCmvbDWhm3+DwTQYulXT7TqAXyAu6A4Kfs2J4OgxkA5w3cg3rlH8/Kfr3ZuDyixqtgjyl
zVIHg5mZefbccvEjgB+yQf3fDmV8iwivXrueN8vS4mQLk8dp6BliPDGXbkKq/upsoAWGvtA9uOOa
uev6s18CGJF/JEmWiERgznh4J3HQiV5KAhgl0BZ2PgKYih5suQdhxJ4C3toReA51R2W4JZL7Wk+9
m7AHre1rmg+RQ11nuK77926Fb5SkpTdudoSTezoX3U44W36uRMVpLuwvXG1jSNysMJUz/1I/Popl
HVracKaNRNTX2KL2q8CZNOYV0uQgkAAAag0skESdsyEOrVyT0CAivUL4fJSpGz2CH0hdTDON8S7l
nb9LvPq03Tg6oiz1QEZ0dh48Fd3UZQwFST5oeOnEWYkM+Et/XqDok/jrIucStGl2siPCDlDBwvMP
gwphoqttnqbeNLmgimk3MI1SLpf0SpM+X2LMHc50pIsl3QsHy/x7yhB89JEwa8iZ4wyoamlfCZU3
B/lJMY4u9FU1IcSRDXgCGnu6acHfuF8xYEXKNtE6JVV5+IQfAfmrgK5IBsCPw7XKusgimOTtOoy0
hNh2fcurLVa29339mWSfJC3viUsPahNIz/q+Pm3ACn1oIOasG5dQIr1hp3JMeo1hTpk8+ySHOQtN
U1UA6uH37UpjfiBd2Sau1FgY3F2LIpTjZBAoJei0xW6W7hEVv+RbLnHerGJmyuOfL0Q5fCKvIcYQ
XpstNpv7nqpOQDXMeoD7UwswQRrKDmIVhMa+bEsBFgybK07rbm4wcA1yQEzkq/6TK12ugQoA/BlM
0sGlxmRd4tlvkgFA0wJzI49qKXGYsGUfysGVADmX7ejICbiluL4a+yc5l3bE5nVHdT5szetqKBln
LgSYWs1cMeBVwjS5hvNuL9jwAA8izPOPxibOcrcARpePd1SE/7Uzfh4zcpzQgY5lYs9ExxL2o9qF
Xhfa7PeYfitjexmFDLv83WTaVduMLQ+ce1WaA2SzzUnMnv5Jcn8yAWaJgtXC72RbOZUhA+t2zJhM
6myK89Zx9bEx80E1QMnITD3eBA/16jzcM+cCoYYSf0JSU2f79XQi8Ih7EhbKSb64s0ZvXDtIqRRU
7sdPT7GKONMvjIvymK5t5SzcoKXCFT+d71yFwEmnaNBiNDHFuGLHpA2r3/clLIWRlo847hcjew2i
yqbEAo2iaoGRNWiy4ooguhR8jDQFMOCiwGEK/KQco/QNu4G4nNN9A5GZ7mmtiOQNNiBzC6ZIL41l
HtXqxRsQLGwkfGFPPPtCwV+ywMgpZBF9fsTPHVi6y1nCeXwaLRNz0H5CWj8jKb+uBG/ywP1JD4/A
qYTakd5bsbuTHOGo5uv00BiCyCZx+Q32mwSeGSI8SlPOktxgNPafi5+EfnP1whvRWvEGYDZD8Z+L
p33T5A36snxJi6bGYCesACOXJo190mCTst9gKhLflNcCgXrRv/RQ1ckskYTY/m4c6ydiB22DrP/p
3WmvzjHoMLQMDhW4qihC751RFbTQvUE/RE7TnX+L6fpp5wBF86kx9sUGz7pvLnIeH1BrQdTUFIEP
edaTvcPKxqXRJwxwOGbKMsMU+bHKLXXsNqSlw7cNYlnUyXlluQ61lKXoU0pOf3z//ppyGV957329
AjTbKBj9uy3nFiFcqD7KHXqSy4c+9vJMjyoqPMA3bLqiD+h35VJQq2sDALbQ+5EwkoG/cplVz4K0
QqMbvpCUKR6Jajg+7aAj9ZTkUUWDwD4zEM26K9NBYCX9a5Y/rGtW5AG4eejBzGDdrCIn46I3cl5h
A8L0cGkUt9aIprPLjQfUIJHQ8dBM/EXyQy9Bx9rHtIy60wFYIDG3y4FVst2ztAqbebRkf0NXBSem
AkQpXfpGNFizxEpvYTYYtIr9pv3xanMJWcppBi07oXD7oerBoqBfkUsogoCKh9WJR2p1G6yq37ay
ugOZLA/9esjwwFYgUqL0AA3mWcK792M/sGfq8JF3r5CHSD0iN2cyrqV4ia82Sb4xDRTlY2nFeauE
5HmT0IWhcFvFCH8gQUfsF3Gt8yNKUxkeZdPzegoCyKQY7bVl+t7CIr+CwvYS+SUz0LG7TPeQs8Xo
qZyNWgZVfDRnQ7FVG8nN8FcHH8Xdu/k/6C5IjFqYhhrGO7D26R2JhzUBQfyNMjOJ1h3STAOyy7Yt
ApSpoF2nfEBdvHjLDCrSa18aKqZwWCujU6YV2Ve0Y1uTMO3ibTr1WuOCMFJwENRyA2XRgEeKkXOn
OzxoUyCdbVfHKZV5b4W4O28O/8lFAGCbnlC4Zs8cFicb/cHW4cK7T+eAQjx6q8ImhHq5Q8pslOK8
dYFtsvX6o5F3bG8SItOCW3YCPilhAxNTGT//fuM61liwnZmcytkHXHX9mnHXpdKCLtr2tvc8Y4Rb
9fE17F18SvYDmY1P+xyjDY95JkoWq2tyw66LAf7xYIPNcnq6o1kPmZuW1wG/bfgV4POfXgv/gwaB
rWmv7KF19Hu98V1hcZEdOUploy0fPZVx677rq50jBUZsfVO50P7u/FqfpOuRQxWeg/S4DgpIeYgE
kYW7DjWMQn1aonh7MGPUAO0phc3xVTgGm5MgBxeu+Wq+SUuArUkx+HSKH4V7Ue8ed8rKI7Ikj/yb
SSxvOCbgnKdqm29Fg0WHGUFz1kTIYvVT5aB2rEuWsBiw7IEoyKR7XpJ9EWg0zlL03tvtj5X20QNW
jxsPwummA7ASV78FBmPD5Ji2OWcPydaEc7NRuPndnfHI31hrSWyaXc0h1KchEadl60sCz1Q0LclM
TbZoHlAJiFeZpzImypCyBa5pMzVNV8ukVrZ9NyWPBmjVyk1AtryLG4ol8b26UcgInwcYRNrMp9ho
wcky7DuyQ2+ObkQ7k3MZoeO0Lq11dMM8VL0YuGeDhZTsfag3R9BlNysYSxsqawZ4PrSSeQjW8Sls
tbDAz5KsUQj4ExXoIH08FQd9y2Bo+eflhbbtIrjFWIx4UkVKmqu9ztkPTii5YSvmHhs593XQ98VN
zNCcY5+5bSRUhTprISd174TM54eebzd1r8c4kyWZmZDp7/+U5jKGSJ6GY/5VkEZMJYnIayyq+RiN
ZuboAup6I5iD4eXEs5EZfUt1C3k1Sw9yyXCyiA0W8MseRJswQFj6TQPHO4e5PXvdQHB9pFgyhGQk
ygSrovhs+pXjl00xhhsYU17+gwbafehOy7EDw0Pcyxh4RZfAAJn11HQverxcH7rbnlyd0j4B7vHR
dWm/pgnop6QPpuTvTVaHahSKYOHGlceDJJTwoWjiC3yBKLTxoy4xfuaMCx78J5NPXPgz/4EfFkds
ROnBQNKmU7HKsvPUaoRCo8lspDGVyvVvfDR5yDg7bqo9lBO/0iukfPP8csO+jBDjqPNrUp07OyWr
W/H8NsSuB+T1CZZFbkAE84LNaV9xJDj0yEgTS3NZLyLdYRn0ygFeghMmPOR2xh+i7n2NholMJSmO
AgTbgkkVeQawKaeyLJ9WQ59TsvEIj06aQf+qkX1wD3wYn9ntBfnDQtalD9eaYHvjSjXLeugOWilh
DYfN5yl7yMjdOm/vpKZ1MukjByJtb5ZGLiGZF/m0BvQiqKWpQziwJ6psd0sm8HaOENictE46ZN1f
kcr+ycPe83nCCKsZ/em2aTKcxp3YlXXpFJcbeq6q2CpFpnTgqbyQkvAoGst0P6+ES32eY91jIPQb
giJ54gpG0zYYQ0+kajs4xIBcwLXDASOBRFTPHdlDQhVgtyp9o8AuZ2qoovWi/O8NN3d/U/Gazbx3
LbODxTvFksjnawRFcklVvIQoAqEm1KzrQHff6HIs9S8Nk/bn8ximqoG9gJi1rJP0Z9ywwqcF2+Om
eS9TuoCwCiHOT6X11G4iyRkTCU7+Hv4QqrG/NaCDUcAucfKuc4zRlYr0cv5rS7fG7VhzZf80TifQ
AhvZxlAho4mShPi49IrlE0CQyn2uv/DqWigCEyuTRcG9+naOrexB0RV08q81HTiozS2sjr17njEt
8lsuyodcst8czX3PumE4MkwkRQl9bOz5UDpbsHtToVoQI1CFgiLBcm04TolybYv6nEujZOtOc1va
RaHGuSOV/t84nFSEmfhm3nwWtWLOsTdTQpP1F4xdvrV5ThjU+zlzDhcS9S9o2jfwfmBcUkHSu0ng
+Jt/wDTt9cwwxnUrx/UOuuJYtpFdqrGojJM1PM42iiYuCSQnzfrXm486qLBeqB7qcHMYYlQGfCEO
4pzk+q3VAh9CfwcQ8wRyj0N3gA45QOXDd79enf9RfMahkhKNMXeVoJSQvJONh7tThPMYQmkz6i37
jyg+Dej4tF1ltGQinZ8zcNUQf//awE8Lpw+f/Zv0FCqW16r9koxHvQTf5md6T2E7klXEgsu3o+Ke
2UWpaLEDIYkE3k0LiYtKEkEbIbku+LlTg8xdBEzWlmld8HlFl6D90njygoUJJe5Eh04+DdLm13qe
D3BKP+lfiZZO53XerhdZHE0b8XHgqyklkClpVRNXgk8Owxz4jlXoNyh5s34O5yBpd09yi0mrptwr
JUF3xQ1r/Ia59nTxk2vai2pVBXGK+vl5Hlx7KdEUJBtBcwYpFPgIs4JhMqO9zDzGROTRJyi0MSPZ
Bmfyw0EPFxUYH0/01CWxk1DLBK1a3GzefLI2boZUp1wXVrY/p7SNZ7I6Y01TzclNLz2NULdVj1tM
NSCruO6Gm/rPWtzx9LcABPlVbKKJKBttD12iYVcFAa7h5kQBnCE8hDVJDac5nIptzF6DhwX/I2qL
iDaw5GGpZPoFrwDeQ3B6c9mgvoRsTLSZQ0KEFHAry2CyA0KK6yF9s5h/G/czW48Fr5tpeac+yNla
jhFBWKgZF6itQAQgsVX7tc+8kQhtPPGzU/DOQ1BtQbGBpTufFsINsObwzOx9PzxKmhSH/5dUSUJn
USaLjCFsMEBtyzflVW35Nl0kyYoGkCD8aioay/Kw8QS7aYUwcAR7GeEnuBKkgZuY/GHK3gB5xPqR
OK6tgJXMp9y9tRVXS1YW+EZKrSeW2YnWs+1yZfddF5NmpJWJscchpyzIERXslr7i+V3vyFKQMgxK
ODEcH8fgNTexW49ybMlrQx3xZIVAEQv1SSyNJ0m9cc0khmF9aipTbSuwhbiMSo86LiqR71oDHM8+
55kmW1crFwy58WkrFuY9xu83q5WLnI/VjM22p4ymOJZW4XaIKFo8TaogXjCTXPha2aNpF0h7dl5m
lBd1jsTrXpsQm4KVsgoK8FPJuhGdvZ2Zj4J1D701atxFF9BmZor+KDEhuBSUojlMSB4sSdwb6iAK
WbbX50KlqqH/2dzTUC3WXfJ6fkvWsv6SXnN/5PMCdCMqLh6CLO81l47/d4kTSL3Q7Rwg7KRFYumT
p9yorCioiJxhFLeEM8SGUlUyhMmXGc7X0qhqAzCj7QpotTFm7EKliChAbqbAVbMCGi8WLCM7T0o9
izrbQFcm2TbgoDNBYF3NJwbeJ9Md4ObQeNGZnI1wBcHVdsCifEMWtV9AMp3V5TBsIAeLAMVyX79w
9QO6ScmRFL8d15YAu6hI8CtOTUDJY37FgNEcsR8K1U+MhS1+C3Sob4vmJZdo6WByEJ9X1fR3whXD
u7XrDk1YT2je/T9gTMU+H4exzn8X8/gMp/ji/3xbsD7INy12HQAcevgsZg3gH+NPsQdxJCxf7HOT
hRY4QII+eaWb2ZqpWHyiBvGuzjqhujY7cYWSEvFP7DEsYeeRBUw2LaySYh8Nkiff4qLyepyCqTQ6
URWOKbnCewB8EBT0H4goSc1jbcPIbJM0rdrE+QZm+guKdW9M4dVMy0uDlIxjw85MnKSLoIcO5iRF
zHrC61FgiZV7nPfCpqPjabTTT6t4+iJHjrU80dv3l5FKjyk8hmNTdz6S3Tts+JjAQ9HEMyqlQXd5
sAeeAqP9NR48R9Mf4DbH9uGipt44q6nLXwj48wE1cpYIbjh+6t07TPXLCMPerRgg+JdAIaTUo+0Z
SGIWjCZ9ud1Id+ODinEJv5IYHyNFSe3WJJg2nbV/wcGXju2LXn9l3A7lOPEEP9dTS/jOCQxRRqqN
1shv05+oUx8ah1XpjBtR1LIgjxpcolZIe67fL/hZjlYEQnopMO0nIDN3VUwlN4EG/XSUaYrVmfii
j0U+8zW9Q7rV/zv8IJiJZ8AN+Mi+q7wITE7k/6+jV2GoCoAWeB48X/MNx5Byet+WFKHraj2InTUe
gRA5GqOtXgVgq0urAh8v2kv7g7BKAEm8SsDzZdrxT7MPwnRnrYevjs4ca9WjfoMJyY+t7pccXJES
fL1nnQ/FGy2zxnjTU1s17lZbFxmyhCU+a42UVJck+4NpcC1wSsDD7wQY/e5YSgIC9W6z4pRY12wK
SwKFhDmhqgCWC5PDZMGJa+JDhI+rH86VhZcC0PZ7nIZ50iwrMs7iHxWnsztbQFbmk8lLOegL85Ek
kwAVYbV8jJCJJ0uqdiMkeNE0pHhuTi7pd3Jln29gpTT+JLCaYa/q2yATbP5VTtJm4SuNZ7HSiCUh
bhxOhYf21Nrrx4DhvDxZ+5JSsjOw6Z8kgUaZv6iFAOwU8MmPI0tyr7FofZeLBcs8eoUWyMHXAsrA
ybfhVhyOPkC29KjuCIaQJ4yxt8yMOuuxhlF6au+4MgM/7fWOzt0OFOirMxbdwleekAF+o48+z+5n
icgbxL2bdAgR2sUneffaWHD5O7Rpo7Dxl3kJeEvEPAENqyBXFBuvHgYvdCwvAD9eGRFo9vM3yqPP
9/+uXi9VT/MWBc6AEA8MPDlEcdwNs7C8eS4oK+JuRoVUdzkt4D3AV3PltE6S4dV/4o/3L6cjJb1h
mPORjtKubL/LnkPgk7QTmCakzAWUIw3LNjs0EkFsm28+cMAQylB5qE0cQTo8JTr30oyWua+BEj8V
OsEzj/NJECNovmDFak/+J6CTqBcqJsZWdRGWsnCJJq0nKoV2Bn5Gkq8ruDCHVZg0dLmQgG9UmRxk
FRyU068kxZisFLRvor1reV4Z/oL9THmoQ92A1U5C+rZMhIfW0fOVdh1pcfJVwlvLTvKgQh59Cz5t
tbGV+qtWjkMFv02h5FnUbG0nXvVl11j7hvvp03kTG0YNnU9Nu0y2lQSrBJ4Fl+FQpYqYb0hj+RgD
8gyJGp7X5IKym8uN7lhCn6uG/3iZix5sP/M4VZUlqjk6dx6sXDlvpKdWQJNZnvk88SJcnJSk2SQa
ibun2HkFDE+kvEGeO6t6I6E8nksZRUmr6aSnFqJaWhHuyQdPw6M4sfQu5aEIe47NZhOToZq3wvn7
fhEIg3j3JQX+WkH9MuP85rj8Gz2eAE0QrpLgW/zfuOS6OCvPwW0SjMGs0ZhVEBESTX2fnLH3pnEG
4Ktj3IFNDxFXwxLF4j9HPzQrvHbK3IYezEvy1pjZhSI5pLO2VWoVN/0hlY5rH92qNfPM1mLbAb5z
I5f4gJSKLb3dF5Cq+3IU1osmOFMF31KDbOq56JmOhB2PpOyYN+OmDIZHk0YG7Q8t++vv2iyh1VuZ
2/SCTXihEfTBcRwckb67cstR35x9EdQrlMZ/939FTqZavr1wSCli3LqHe/TKZ8U/7a30/6KcQddI
cFtKZu28SBxXQksmLbktszisqynHJ8BzRiuzIcCXeVtWwul5ZweLTfs0sR1LITiiKYb/lpllhGiC
o3jjBJwj7TfQQ/1uTrd05JbfwN+jZVMJtI/KAt5P/ufxM/sVpe0cEYOs3C4MLtmQUYw1TCSQOW0p
czTtB9bAXPg1iuSMLxpbNEpeKjymuPVdSVIbdN00+9ZrUnE8e8A34Lp9xvb7+Iy17/VTkhmnY/Gb
fKnjc/JfvcNguPOc9iq+uJ5Sn8uJC+kb2o8twvqf7A6IIE+shLN8opv2pUft2opNdYYN1O8QZhQy
npaqj3Pf+eElKC8fNsuvx13fN11yUaSryGNBxQtnXhOudWyrdgO5r/VxEMcwYZ+Fr+5mPX4MyTjZ
Kn4/9NBtROWPs2KHOScZdy0NRB8UwB67YykS5dUVFUaqizeBx/H2y7exJtxMKVuwD1SW5xvQcK3R
WPzZqAfmCQd3wu7nTUzSBjGt+awbC0Wb44+YIAvmXv1wfdAlUYjNclUK1tAiWwFZ737GJ/RG97+H
iZukVcycXQaYde0PTi3VucZTM0yQSPhFIMv/9K//2fOb3Lo1AfYWpj4yS635/34AaH0K75Qrn2Uo
rAJfwxI2xJWDbDLdRMdj6n8RJ95UQAvbaPOBVIn3pwmxf4HnadSGbvCiEvCrXwalDck/DxU1m5Ao
+7Al9h/Y2RxuIvPUuRiEUERtrfn4dtkWKHgv3jwoYtbjE7Xolxrh5ZjVVpqE4cQrE3ZxqebqBDKn
YUpxp7xeGB+2H4HlR/OhU7JP5arbEhcKISGuUOz+6LyxBGAJPScMen4ETjNyhj83Hy9SHf1kAFSA
yUYvvkNiNIoZolLwcDQi9DGDcBFsoDUKuMbRgPj9c+P85Gv8h0OQO5XRdi0Lp52KwjkAQBwjNDM6
mrZiWb/QmEYnsJLL+GkWh/qIF4uUvv3dbGSc3T1//auZg8wCr95Wr3az7l0r5K+WdDXa6KT+SSc9
m8dcoH6cjCoyP87xLB9/q1KCgYdFz1MKRun8PvLoS9uGz4kqDRTv9ru2ao6iBZupT1j1DUHIAVsr
wDspTLyTQF0mwtaLhxVibWp5faOv8WUIyGRsBxM+SD3186V1ux+ZpLJx9Ymw0LvqbsLyutqqhY2B
wDUn0nVbuWHy6UzBBnwcDs09hUoOfLNCOmcHUYvl23PvAcxrQjkh2GFsIs6kDYBb3NriUQTrBWiL
hlk8jCHf0LCwSU0XlPaQc3O3Q4UhgBlk9t8rLFFTLZa44y0ntnrstvVhtiVXuarq3dsq+05fe5wh
VHFb9aL5zZmLSRcWTbGUyFgGOa06E2uTVNhVK+tKzg7bG7p+elWX2GJiZKOfI3G+5APFMyFaJiYi
cQ3lrFq89VsbKcdThYs5teJ4NXSaubnn6nNw0J7Bv9SVakS2AJs6gEsfAuxNbSPvY5ECb2wbIIGK
uxaIElf34MPmJ/SiXUCO95wuRj6OKLZByeqT2OIAGJCAuzt77B4IBlbDTd2rOV/b4E//bKJmJUh1
VY5o6STB2OiNJQwf8l4EjO/uDpRsvMxfkchn/XyMj9SJvkqOKwh0O0ayx6OYrYkvQCrbyhJ6ELTz
tXAjt9uRbBh9tS0C1UTiaEqG3HhJITMV7e9gulobLFtvXV96XX9R0xYh+gYQMquSChQN/kmxauYt
JrJFVissdS7aktAyUESLl18+yODL3LkzuylFhnlhonnA0y0gltOysaVFOg6EfKgh++eAufV+p77x
t1L+M6mbshHAMZBew6ExEWzxzx/X0XgK7bjWZhrzfArEfH7H4xN3JjPplmrY3SzE13ZcddJUI8OH
yRNmRhoTWk0nsrrsK0hJnN5cVIyxQswPciXd0R4K9Uw8IJYWBKjYIpiq+F7wFE0afDIz2gzM+C+z
CibQOd47EOOdibhd+hSFCsooN/vlOouZtLIUb4t0X9J3adEINEF7+P3DbBoToL3pQmmj46XvPKG2
4aAakfn9SI8Xh9ynflSczuLIYMjPG2bnOPxzHCvLTqgg/ciBgZdyrSi9n7sonVokMJLY8HTGQQl7
Sp0qT+MG2VpaPqrOedeFpEE7AqaM4eKnLZ24caGjY2AzfhBcVPSIaeLhM1q+dcUuBi0ChVBr0Hkt
axILnlyZtwzw0ZsAHgXEOnea4CVMJ2j9WyrUU+NqRIRsostWHO3unInR20D+1RSScZf1ZwBASfuh
DFIAny9atDfSBXlJQQ5KXDmFS4n60wq5KJC3O0FQCU0Ig/gMreNI+4RmkIiP3khZZNb8Ddc4yb72
LZYfo6jEHoTy9W7eFvcFe3T7qoEoPh/o+TSnASwkMIJKgnBrduOOD5+DxHfUv2j7RQVHo/j181CB
zaLG1haOF2Sbk3r1VnPFj1ROHb6Ii/Q9r81C0tLniqmLehCb9JQyRafy6fkShojQZ1Ib+z2h3haw
iUbtvnU60kxkb8XByR5+bE716VSvHrBLi9tz2EtZTxL2h6eu27oElq0KEBhh0UYpLQojRSaS6qok
nR0iYAfcOnZfOyzcXehyxraAINbdDezoNNh8+19BF8xK7yxjQA/O1F8RMD2pZdlYiFD3uhwaePhk
a99TnO4v7UNWMbc36eMUkCldDKyOUBvOv/EvwFdeRhjZmUXhxI1VDGjYpRwgKcywKANskE7tKKMn
5wlx2Qu5nYFyMti5fV49+5C+bTUFto0BFHUFOxPtj89OYZeTxFYk482uhkAu0/aQ9nKywvzp+bYl
Y3m5m9oulOZhuetzxRUN0gyihMD3lC3nX3rAhDJuBpC9ujZkiuZAoBDI4cwCmoU7sb1oFgFS6uO5
xWfnU/UATLHNIDn0+PYKekLvC12NR2zFcrN0hYxcY8L5d311By5bZvvI4xCi73OkrPPtmM+cC0jV
fYHY9B1XdQyC2wYX8hHRe5rBZ1Ovh80F3ah0ioBh/58dwyVNZXHR0WX89nQ6eyqo3K+ZrMxHQnzy
+W8bhzftgL+HkyMaCaHnCc/vN+L1lX8YeN/7z3F8zfw5lYtIrGVn3FePPNRoi+IL8B6MjIwplwHp
HuXxq6+8E1Wsr+xw7MuihGDlZYRVyoZJhZ9TT4jCP5+S5p/bWIApg32UKxHcQPFNs7JJxGFNOv9c
q4qstKxWnEdJitg9e/BbQcrIBrWIr7/xJG+Ze9YiB2lgSgOv/Jsy0GInU5DtgS9eEpKmrXt8OIHk
3eh6Hg/5sfX3l2DGc8pKYktbAi+OHuakiUeKUkb0LktC3EOT9621Fl2mgSrVlsTw0+KTtjwi7xeu
M/Uhm4eLTUL6BtCfLjSzbn/49JhPoHcvmMQMqqR4mBmX/8TlDfcVfL2XsmzvAs1idcX09XtNujVX
9NHXt/ZANKUIG9TGjPLqMyVSOZ8QIyu7bEazDI1gjj7exm2pLq25raxmFUkPN2HbJA4Z6MoOjNMh
xNy8es1/skMwY3Bn9nfrLXmMR5BMD35PYbYtPBRw/aSCZ2QGQA/mHdJXwh7Rcvd3QYEtLXfAcNyj
N/PMLiM/tm6ZGIdJX+JDvlOj8K2ltzQM34M9MchVI2BQMKhpdmiyQSd7U/sEZTYKXA7i3V/ajaDL
RHABamoxOWyf1O/KRjxXPLUTSxSofk9eShz+wCjrYotiBjg5qz0fi2wSi35O9szXUAeIGN7/oGRS
hV7/mxPh6fgAoZP2hwFdhmW+hPlGmfGcKgCcsjgaWOOkIS3iJskQ7nyfxzHhN0MlpcCjz9OD5Ish
GEPZBQBJBLISGUjzkdw28bCa4fGfOYfLlOcfqLH7p6afVJa+lqTBkO5g/cWQKrHX15I2iJMVacrQ
7v8DZyG2hTQkwaHa91BoMmw+YzAW/TScXFSaBZbbwPrb1LZn/RiRDtWj0Pvy1DiAVTOX3o41NCvT
C1BOkPBg3VzOoqBx9hd0lpxwFx1eUZeGoUJLRtV8fp61Cfwq19AfVuQl2Jr2h5MaDOVk+8Qm1J9+
596mDYKK1l6KqelSuRjQPM/vFQ8odt5aJqXc3gKTn7/c/7BiflXd+m9Y2FPEOro/xkvsEkcsmMZL
9R433iXzlsFgsvDfnMNlSMDslDd+HoKuDA2a2nSVddrWXEcs+kshWl1XHMFDzvWMF7NQjzVVDU5p
IEplrHtczF6dMZd92Nw838WLhTA5ME+dAb+fz+IQlDkuMn1BzWUxEGvY0Yldrl54xmz5FgZ8hp+F
fr9WmmVy4lT5P1cYK8kGImWoENWA+m+I0mqArkLbTbnXXIyvHSB3GNMDZOeHg+4OIfjKToa6aDvr
DVmghTybCd5bNVh12It2BjLtYBA3TtcARLhWOCiabucrRIhGf0828oIi4S2dlD0twV8STwbS6hhU
i6/cLhTJV1xCUcWvHHvmVS41SP1t4ahWsMaQv1xPOWnMe8NCZB9VTSKmY/s/C3mEvoXrf151R7EO
UBWGLkVBg1dawYFlMdbkZm+LiOj3S8Er0FNEcG8RcSiHLXmz19xt3xGTOfsiJzExSdGD/rRlb4/W
897LieTSofCO8VsdFdKQNISwy5TZxxt9cRYLXijdkqRBVrotjVr0tIBwhMUanJpMe7sIHSJyxBcZ
+WgUtXozewIR/NsluoJCBTkUqul55OElrirxoozKRTQF8+nd6UxJENYJICUsRfbTDLWTRy3UxmcP
8+TfkzHPZd7d6n5ubSFSP2VIDwUoLNMnOuSudC0ntJxbx5pQX9lSfvp1ECcb5C7R5HcFZ8lalHVC
EaUj8dr18bxUWHcNK0ofcCpw0k8vax0N5PUKe+P/B0QwTo8AjL1wY1npSx5Dc742Hmvw3RPDJC9E
+PnkMWl1aFaQz8+mkcKgUASC7cbQEwXLlifwSrqDH9z17rtncbdyvflD7womIgRNeynox3Eot2yW
6lMWl5px+pey9I6X8u2OrrggluKG56J7c3Nwgx4mNtRLwFIcciXa8h1aRE8Es9xiHN5Cy2zIk2OH
mMhZLzcAwt4a7MfqV6O3Lcf49/c/dvpouj7OUjeBb5OKApGdSgyubPtngjs87zyYhbnzKAJXlo0B
x9t1shtAaCQVbmrOPuXda7lI/Q1E8qVmIMlLrwQAJhaUlziUjrFBZs2GwlpGEWNhRqcQb1sKv9RF
PO70CTeBznty93/K6FV8ENxyvhiducUJG8fOLcS1h7DtCdT0RAUBF9Z9t7Ibyruebgwm2nuCw4jE
5+AUql8qxBDF+5GPeNYBb3puYKMUGbjLHvlyugFS8P4Dxw+NPzR4DaBe4pOAoDY/539JVqmczpcN
Ih4+0d0c9Drgg9glHjbmRjqZF9WUoRrKJRZf3UtS5Flm6vS77UClAsrJMfn43+FrieCR9g1sYbzR
KQfMpyylsxvsd9UGLBADWSYJlIG/uEie8COEVGEnC8E/TK/ZuEST3CSvcoY4aZLJsPdcByIlcnIA
SaJ76RGfABTP2fA7Fa1m5Ujxp4ETYTKCJGUgdLB0aDiNeS4ttijvGN1yXW/90hsoZslaSYC+yXV9
8SoV4BiE1RfPO0fINF4mXyp0OVaIRrsv+1AAkxY97gPSH+qfZGESptzYMI9Bek9fkHrrYnTsb0ID
EHcAxwGuI+DIFAPf1rJ5ga+5aU7vETvVu+9bBiMisgNlcl53Sde1LnO3u42jSHFVHzskR1kRmyD6
ql+sr9A/e0BUKthdc7f9UIpqjGPBHK17WWhdn0SXp6MCgxe3LMGFKMYUeZpL8tWc/MN1PJm3IRbb
8VlrYTCiNRLeME/Bb/vvMQ2jCUqUkkO3zToriXGmkMWmCj6vNModJvhx0nkIRyOsCjmE42h/hQDP
bZqm+O+cWI6BQXyjl3A35JJd0EiWYhDUPJubVFFT6bu6jcD3NC/WXgc7yv6SU7JGLWBUPacQ9zOW
BJ7SBYTNqqRRYDbjmkkwpmH4mf1BLQUm+Bo+Wzlf4FgE8og/NPCegh655uW/mvp3zLCQJKi9Y+XM
mJSYWdgCtBRi5YdVSAk1PlvHZgClw4AxnHRsfj5gAo0Be8Zd/el4UOroqm2/3aVTPjrnP21IBiNl
BxVWmeyecL0J1rXTMwilv8tcpJ3rycX4LZjMe80hLscjkM/sryXTkjy6A7xfPPg8tQXP1OegmKgL
5YswdITLYM5rwSstb6xLJRouoIPSsr/lfBut7JZe7gXQ8FVC8Cd63SEZNFD/bXD7HernyshQz4n/
uPfxDAp0R3TtrB3IxjgiUywdVlo9K1wB/o+ZMnOMlWUcBzKIe1r3keXrk+CO09QV1aSTf6qmlgkw
L0HjSHI44K2iLcobzAi/e4LoP6FbH3dmV5hxJMxzoVYVxJAwqon1ehtfrMbjoH+67oA/fWtGqZd6
NL3+E/PGWFPxN/bKCgHBF4G1qWOYsDB/FUi3LUcsWyjK1By4g7n1m0hmntSidfv7CYyTU9pgvSN1
fZ6zy4sk83yo2qjdEzZEprqqu+nZQ3jn1AT0DPPRHxPS/S5R8CZtulq+Gr17vClCyrE8bLIChVX6
pWk9OPWzmmsH6TQIdk8i0JXaP1ZcU4SHIdB2PR7c6E9ivnIzKksfml5IQ3LgUhxm7+L+Dye9+gYJ
Cx4P3Rs1WDWu+mSuoaYzGFTwoP6gRaBW7EfvQ+DT9XrFL10f2Du+WHRbZ5XoI+NjSufpVOWbguAa
mze2ve/kg1c0r9ynh+mudfcl0+//kZVgsbLHOzsD3H7JpRXzXMfe+ARngqMvW6gAxsgpgmhQaJG5
jHHftFWORLPgx8BrFUs3bjnnSHUWn84W84BurvE9UEN+gjmfKAzmr+bsx1zrXv0W/qIi8wl1ZCOx
xkczZ0rvhrr2N3FXvIzW4OkP1O57lycN8x9MEVsg/zkKXy3FJfpUQHiP1LkXSWHhqcTKQpdjaF3Z
+Dhu9wrLhPvuv2Bf3HSnF24GqVNtZf8c2HdATiJ3OYv2uJCG1FSKicPuwB8M7kRklWtw0g4y6zMg
tTdawyCyd0ATDgE6Kcj7JXNhC9u2b2EqekR/bE7xQIc5pocj2GIeVjWzJNlH0N53FsnnKfRhmp8M
zQ2HhRMZjL9DC24AVUC3rjFeqCpp2YlTXLHiCsWRgKZhY0Hc4jpprCM1y+o0zJs35Wg3C5lfdNWo
yCN2V22gM0+xxW+UBGUTUJNKr5xQb06mebF21HZ69boQtY7qhx69BYBCqCXLaNwQh6LwwagVLSoR
gc+kKKe1kEnWiLRFN5eUO3Ng4KeOH1C0HRn1Pr97MoNtFBdxShZzJZ2+ADBH7UWOOKEirSe9giqQ
9miI6AqgfGSLwBhAs6X/xmKJHRr5biLKFmbvHGo5CSD0Z0hIMik1Nq0fNfnNwfug9604Tqri6jgG
Ad6zdYpETvzEoXr6w6DL2oGf6hZtWpQqN3K65Mx1KaucRmRvbz/q+6th4t1JGtsu+Y+goB4gcCxc
peTFzaoRBC6q+hY3VhG0+Fx/osre4zrWcMKFtcWOVeNsF5ctcPBogo3IImOov72KtC2azPTFQKM5
Oyl5/VRWXKO+KrD3pC1rK4pQCMsWfvrKyzrjGqMVvSJgF359UWcljZxknn9jsFxVs9mophzOwd4Q
wFsuUH8hMv9dHPN+Zdsyr4UrBwD07VadP/EeFtwpkTq7nanGRQDO+VlSB2r7pwf9SsDbuMIq25JH
EOXGatBnHMhORiSmtU1sDCCMYBlbIoxrGrJ8MWKpG0DTYY1RTHmUCN31F8ZXTXRYn7dbDoR5UPU0
yICtOzGYPFILVfA+H/xeRYTwIoP4fvnc+hle6S+pD0GtkGenK3jvmJLV9H3XClFUIB4YcqmsjN1W
HuAOgx2LyDKNcOoMihHe/wpZ1UEn7/pzKUdoWxo3vrUD55Yaj4EmIKz2YiKFHNfx07/4ObklYSXA
VXcSjickmWVCr2tWlp2CN/B/rspNiA0y1LQfWmGl8CeeUR8p4rgSoJB9++6omZSk8CMjfVfv6dUa
aPD4bBn2PbEHkxSBIQK0WUybqYSGJkmFu384I/k5Q2YvcRr5xOpFJRg5ljm9YD5l9+d962MDA6kP
1sbb2t1bKWqXXyRVzYqobX169h084QAcjxp4eITRayQ2jqgqN50c3hiTcIbt2Bdl8Wd5lARQjpJW
8ndAJ0m6sYoy2e5xLsByIJzy7dD5rzoNR1nlvx23INQSRA3azQQreOS5FEcjV6xoqEswrQM2DNh2
iOz0vjLHGZflN1WJGPE4d+q6N1dX/Pp2WEuMliSJoZnullHgRwNdEDOzeYd4+UKLh8rE+jN7vCPj
J4QgnkD55wQn2gTycqpEb9daUSZiNhhovPG79PctzAUAyMS4lIUeGW8Dtvju/SU8PkwkN6NA3Q5o
8wEt+V9Ssqi3baj2ry1fCS+bNA+xPoKdW7isyhGA1LzYQcVI2Zbi8A4694yeKEmiGFfrrITT8AOW
P1lAFwfn3rs6Ho+1Ljamnv/ULj1i9zKFvMu6vtIYghiUL5I5/WtZy/78DkdiJF8aAs8uyMamevkv
0Z0tX9X7t5O7mNAbvnhJTHh+oOlC+oiAV2h5t9Ebkj44URLFekgvUF23njs7WEgp1Z4ha6+CtgIV
tuGIHKuJa02TXogwjyGUo2nGe+nU+V8QWwOhbaGO3fdtlgCBPNbjk5BiIAiAJEOV2hKI6W5LtisE
S/9nZPwm5CKRkEslqWhLyZxoACcoR/nqulNlKHDFfPUEb+wxSlNR02J6jilH4RPd0qRmSyGqVZ+2
UMe/6N5g1ENpeHUeXpuCjIpa57R7yNKA52mj4568UCWEOS75h13tJiZNgkbeU1L42JTTm/G0FlF1
W3VIuwNj1gWqFSBZByizMunfp5DpdE5hMPn7ICsiP6tYgJG+CKz9+Xf+TRzqTBkOHEdhXNvPBiPJ
R7KefN7/ugFP9pC80T8SUzwSMJJATy/WlPO6exgQtI/k06WSY8GtIswUTdh7MNMZVbfpNGKyxL05
QFjUvVb9yBWuN+Y22n6req8q+guA57udy5Cbfc9egjKBVeje1a5tzr/s/eA5pEl2K3FNkvFMIU/a
Dho3JKP1LzMGGZKrA54SGU4Y7d82EstASZQ1tHOlItiyuTadFpspG3s6hH3EKpgHFQDGRitrT9Np
jH9r10+Fq/1xlyYrz30A0A7vL2wWZwD3ciAc7B1rrL/kp45850Bxo1kdCHD0uvuW8rwqmxVxlBSe
T6QQ/MBfCis1a6E6/mwuXzcln22/cSD/kumEuHJvMlZUVd/zf7yvB0Xu7HyHtz7Jqyuz+jNJEuQE
T7h/Q+IxPrtQmO30lw7YkGSKBHHi/KNc2P94i0oVkhIxGisbpRXnS6aA2NYDMZsqS2OACVGHp4Fk
BqMrSyqSEN44/J3BxmLMMzLxpdLMAzCf+Shzb40NZ9zz74JSBHWBRIq47rAUlMjwzSSuei3e99s4
3IGbziKcsZ/uzzVgoOSNUe6Y9YZL4zImzvgifAxF9Ex/Q0tZRUmrhwvv0vDSXeDhvP5IxJl34utV
tJ6spV6qiHSJ3Bi5yIlioGK248pA5APARm3bEHt9f1/ptih5WnpvyvM/OQdMnyMWmzF0OSpwK7tB
EIy9YHLrrELTNIGFmwGlFdqQE4tE6rq5fK29tFzqsMkPzYkS9c7E3uPNAdh7JhO24h3FwYTcB69T
A6TI3xjip7XuIkWCV+9kRJj3nU//fM730FrZFUh9KIcvKzQpqnqO8GN9ZH9xo7UQT7oB8Kj0U63k
KGng49FWd+2VJrFle6BMpMFmxadKt0QDtk+jbi6J4KjLFI6eUKibyDR00H8QiYQApxU1p3e5wGR8
VVzAob2jrq/edbKQEd71+50iW9TSYyMmCMtxm6z+OHcCvgN0dYEwx+ppSsVgmKAE+mSDmWB2WWav
3x+wuXiDOEz4vitGyhck+bhdlOYRRBip/QHGRC4QNuk3yftuZojSek1z73psnXh0Y0n2iwj5H7b8
QbcISN9RGxHm2cca378XLmarJubX4ny8K+ZxujCG7S5MrFyZa2qmEZMQHoxziJYEcg/F7t659Kvq
0A33jyba4Dw9aJaJL5mpqzY1nZovWSpzLMjKi9ZJJ6y+4ohLzhkae9WS9+iEVeLXY7fGsM4UKe+e
LWoU5/sGMC4vihprAaV/9WA6nSVOn826jsJz1swpRVGxCwQI2uAmjHmxwfJPIfVv+c9vvOg80OGq
jqnu95jJ70S4nKoiug2zklI/4tSaLsuqoL6pMBZkoEsmbTRx4amAD3aP+LW9vK441Q+fFvVwTN4v
IQ5b+NMVXRzcWY0n3yVS73wyfYSiUstmQ22lYY3ygdQSsYNqorCsyZpk3xFrQU4UwmkEJf9IppFm
QDhH3W37KttRvEoXE/KSaqLzUpdvgmWQcnW8wsld3sy3+AO+nY3NUpj5HYMeOTUijEwZYDdRPPSj
o5TZgam7viRckTWcM/6Q5y26zfc0oJlHmLKFHYE4ETtz1eADr07b0pz0ZHTySv62+lSwqaQShc6O
sSOV6QyIq40tEdwjC0I1ip5cVLJo5F3nDzgfp8djEqx8BmDVY5KLAgLOnh095XDRcerOIZGr2r08
ItKw0QufhwTSRgt/eaTmWtfVqMB7jyaZ8WlZ0qsAmLm4AHC93kC03KhylBfjNafzMFr7spTYiR9W
R3F8L4ajwM2tiZE9VNzbGd90VqWgEMIJ40Qr7UO2DTHfL7gORzwBmxytqx6+zN3Wd0AWN8vxQlqu
xhKsNbZEt3thz4l3YeLFWhWoWWvNvfI/RZypHUKjnA8xPPZDxEy9GJAMznOh2GRQG+5G5Ecx1UzB
zpDescqqmrpqNA/BnVVHFfEND/czu5lCYwmVb/xfZWzYO5o8wH7kPL2PHWpQkrbjkp+3vU+xpXJ0
F9krMXBQ2k2nn4SS6+C3cFW9tsAeQ1wMIzKRpmagQiiInzKddk8X1cQl5c6ZF3zQXjko+9LAfnbA
rY7+Tll5yFggDxqZHZR9osij1CgUJbFMM4N+o/iC2j/tdF+FXSug+A5bapfU1uNpZGa5uWNuosEA
ZBa0t/phTUoKAY4VSBaKCEKqAiKO4IS2I4hmW1xHBJaKqY/IsFh1J5/yJoZoZ34MXShd2dMNydk6
H6xuKipeeY6HZJnZqMW8cmnVgLg4eC8pQ69eNvbOda+o1WjoVGaXFZB68qfGxU3RKt/cAgyE13FN
I5ecTsRpW5RadhQAaVtwbfz4ti9frEYbju84En8lfY7GZzyjxd/p+AW9WYoZZXpifd2oFCEWHBFC
R5Nz91qQKXSHIpWEIIE7v6j3yRPJNSszwKRgViF4n+U4Wnf//lR/ZgTSpgnB0xbcsn73s9hYl0rb
VtF1VLZ2yzGL16LFVKoHFvEPef3JnIq57FSPQilL2W7ibrzOFOo+Ov4k4vYCdhuuSmJkYDZ1Sy9e
RVqGa1iOs8SGsZatAIGrlbBdFZ30o94W+iXclZItkEmD6XwCgPzScTEd6UTm7uKYTzm3q/7Kvvpp
FcjdFwTgt5jTAFSee8LjaAN3LZWosztePnqS5iw8JhxWA/OTaPtTCsv+QrwVa919l0dLlmvWIDQr
dfpU7TwFoLSLebVr8l354RlUNukENTBAxZWCVQB2DDg9KRXG5pNONIYm1W8ns/iAst0BMrAHWPDC
qDyjoAHXsfflFTS9qcs5ZHds3MYGWCNMJNsizCWYAFpL2yLuKOPjvNhcrqconeM7JaoX3c1NJZcj
yojYzoupiDhsyc+2s2v/TvzBhiuz6XriXUQLNodjtUTB+SXrK3QJD7zG+choDUoLOkSs/al3cttg
gIzqyS1wHWIGxw6fMW6dSurGQGD+03qLUyEiohXf08AfmRf7HRoY1vDYEOfDPPX8ZZy9A3QLvQiM
uZFkL+0nv0gwZ+S6jZMFqNkjYjVbQXwXpTzLSGL2ziAC+eD0RNr3fEuYfvCim78mRDe3hmMImJ4w
qEjAA3HnaK22RaFB+FcwxpsDE0xYWy8Xg7fU3wvdbDLh+iBe8X9Ur6/a8yyHEO5GTN91RiCU0Pzv
Ua1DMV/83vri/ws6bJC3Lq4XzADWNluewwo6UdSpD1+w0aOeIBSWGB4XVpxetRg6x26uNiTnYE1l
tl4fJuSW0nevLUCKSamXP9U/mknZthJ9YxhWAs4cFVtno2HnwLEDQJIeDevG4qvO4mGrWC2BjHRy
CzA678tlBI8hfZM+LbbhoHYse/pnu+hyhmuULrW2XfozkWLtbldJHrZnohIjFcxsSlZWuiU1y42d
scc8Y6RrCK5s281CIkjwxAyczoTmYbPBpQw1PvINgXY6K8A5LcTxbnYJ23Txa3hrzUvJKBeHkChQ
5jqGI/KBxTo15lI0B7QPlDdD3y3eOz5RxjPBYrO34Yflq34lgqOss6N4mY5svo6otISyPNwqxiEo
e9aoco85kr/mko3veuhJdNnrafH9+kExWyHnulou73Z6ZR1ye9NYZJ8oXJv+U/MRQaCarJIfpXDu
qR2dFh7nIR/JfEa3ri+wBQIsU1Y1h+Sgm1Iavq4iv7pVI+yLsi+ZY9QeUo3FGvUdFO9QSfxqtbdU
iA9SkGDtBQ39QCRZWj0QPbokaPGLx7LP5j0HacDhXqHhRVYAkJ+3x/Cv7eu0266qymPH9fthRXY1
bJOYo4kIxM6Q1BF1jiPRbOwlputAZ09BnVC+ZjfXFjT8PIwYTs2U4UDry9qawUANpdWoFjR/021Q
n4TkHdBx6HPUSPFnX6NWqWs4mDqNT4VVDacmYzekQbvpFCFcv5UVwRzpRB1Ev4EINxfV9V9cMReD
ZtOwDUTHsI8LFBvszpGvgJ9PgnDQy88T1OPPzcYtQphm5y1Y3iqCyT+BiSrddx4hkSmPmk2cgWrg
16SnC/jB9cC8McF/fGmxGmC7t3NRTSY8oGZLeV1VlK7lyIiFSbk44Vvsx7deKNNvu1dN2nSpVIpW
X0YQ2La3OgwcHS9Nv7AdJVKQUyhwcLYOcqKi2OZ2sJJ0cuGW5D6oLEj0xbNx+1PGYVC1QJ33BmNg
Xhl2jz59CRlFUmVaP9syfU6mBZhMrQNCtqNiqgt8qf0UdlfaP1qA/GDmhl3I4fzPcDdlCYpfFLYX
v+n24Pzef/1EqPfRoypZ/AL9ZzWqjpGCN6iapKTWpPeU6QmkLojOv+rWbU/cU+vCMdz11eeYCyCE
6jDwotpgzugzqemZ0LjKDf5IvjH6ELJ3OdpESYVWs/eRu7G7zs32aZOKuYYdaRthBlosBtiSash8
C0mXtrtcpbJ9Dv473dGShY8fgPaBZzbXkqB3OiedJnFUGWSymQ6uO4eEbKX7biAdfRwWNhZAcm0U
rWQouw3uxFPCnUNlc4+mpbF0M5ZJ/kekw1TlKdEg+ENQZOEDHQSAbEmJ5iIhSi/C+lizHACJlwAf
zIH4bFtFdmTagXL+koSxvTM5qOew4oLMwMuOE1xywMaTmvPQgBnqH1AMKy3PA9S8Y0LdLmCLjW4Q
dKTNwlxyUU00S8TlRLbJd6q9jRcqUvD1Cw9Hg+I7oTVHL5K2ro96gXE2EDsG29zOD2DAzGJfIq/b
7hyT1kMhIyzovT0VJIKF4PdlmxM+0N/tHbN92YmFBbv1AX1bI6Sxzvn8gXl7Z0QkgoAwufhBgiFM
8W3G0Zr9FCXl4kqz2HgGTgr6hE2U2gEB19owWR7VCJ6fM9p+jXlmfV9P6rBiYd4FwZVOY9TeO02F
cjqUuJpMzw1b4dmcW8NXlWfdCoTgEqx1anKhaUks2w0TdjPylSusOzKbXFo0tuLGzfcZYn58QA1j
RXMX7t4fOx2CMPrz24mtwEImHL3ognM1++0S0Kx0H3F2N9/cWIyjyiSd5zhK58KUEpyP2Q6VqN2U
KuqGiAdO6QDPVIb28Fo/8KUrvm7ImhgiiUpKnsNP3QGdjc4787jMEyOKc1mU7WQ/11V7UgfLCsS8
C05vBctvKtuVwRsD2glMUPi3RMlEPCTLrATjyBcYd5tNpYPofqIs1XxLE/tRH26MTrKcfZMA5ajw
NPGIQ4TEQuf/6DFbMNwAYX1MwkJDli9snDsvNk4usw6D9PjNSK1gFB02Ort86rcqIri5FMVL2YWq
X1l6A07TAyXjAL3PNfRDxH2fEmVag4P+gj3bdhcRxiYmHhXN2eRpCf/9epjJtAkXlvhnMl7jrwDx
P1QoMQzsg944OZ09JOhF0+Coc1nY3QeoqjilJhhiOq9HsAxa6dqQK+LZXJ+esk+KQHEgjxVKF7uR
ScBiPdauIBmrUhOkffRPuS3M9YDWjt0bFzEU4sDTCngYxmlMxPcd0kbDIeX+qFzefbPtCa997Ra+
UdVhkrjPeKaDXtTRwwFKVLKqj5vO/raUWpJX3GEk9epnArfJL2vdltvYTsW45mTiAy2xSqBF0ndo
svz+WRByBDzEpzF7+VKgAtWVdHa9iOIs5lT477YIrh9wT4UiKT0QlO3rPVDyG3MqKIZSLJ2TMcrg
w7wq3M608Afz0SzAHjlHeRzSWHJtOaJBrQHxDGoh3uiKoQYUkFg6l6YfaE9X0dP496Xd0YL1JRf4
bkAowXGcJT1ZTvfqL7OnXQib9JhZ7NkZKdlbDf3Z8Uc3+c0Z7KUopQvJKe+k5EFLdN2IvAmoMzfc
N34598C0Wkk652Lpn/kxrfxM+zjKjCEH0ipT9ZWJzftHcJj5iz+JCdDUk9u6VxwhGdoyUZf19UYT
not02SI+do7A6lXP7VB5T+JahmVtDS2loxyQyNwrUpfulrxTkImi4r3/gOyqYkdHb67uhYPAGKyP
nlys70Xskxrg5qihNxfdbU6DLUnswv5Cyp2YcIdvnlS0goL0gp902Z8yNyMmk9EGaYCD7Sly99AY
3nS7NIMVYAlN/rxDzS2LaWXOP45RiF8jX4oRhcm6GUYcthCSpHyivdU+8sZp5krB3x/yq2TbvFJt
DlzPs0vQ8HHXZXG5zHKC1sAlJKSdFlANzktAqMxv3ZhSwBwfii7z5icIcEW6WrigmFYEw7vn2/sh
f/s4sx6JdYQkgDsMHR2hyR6e1x0zPDCyqPpaWMuIRRdPn2q6goulrEn2Iq+95V3yHYMvizW/KLZZ
Wu2i/0HVeIJAMOI3/42sPmqdYkkOTwc/Jv8pjSHIsX1daQIwz7XnRtTZrrKyRl+yjFA54tf1dPHI
4Es7K3c0qoLrsCvtToXXr38M6SXRqc7M5YOs19d8OvmMHNG/71ejUNLGXJVsEERBa11NXvx7CpRN
En4e7z0rA0VEASrg9chvO75l/XTzKuJoeHse/DsbRWKF9rjiStJ2rqZFyrkXIa6HjJH3HNhFEAAT
YHRYvLYz+vQp2WnOmgoV5p5QTFjMA3bdaP5lj0Suq9G7bfrL8J9TITc/EyoNgYxVvCnUAtDaoAwo
9X2pMmBAy3nJgEaSO5Ar8BNSPjX46CE9v2EFajV09yGOTbWOr245buwlrUAbzhTXxF35Kp2dJDqt
bS8H81K0gbqa1/vBgB1HqMDfUaDqJkhb4D+11LxFbk4jG1W9SFVSMt+von2Sau1fAseqUnVjZ8WF
fWq4X1SQkQ5DYbRHd9oWN05KQG6NJg08Wsu8FIJTJAWVNwgtSUYMlTq3M/4hI1FVKivDCvSnMhVF
A/zPxPOCzNhHOohzLSI0jl1ch21sO2BtxpUQ8oolfMjHVBkejeqtzjtwxDxlgHJJz2H97Fw0JT46
44wCJ5jtLMG/3NOt+kIYHFw2VBupk3cyYya5Fn2SShFqySZ0Q8n9NLY92UJpUD48+EL31hLfSZ3b
X44FuCvsOnYB9UW5ALnF1gcMLSd7N8hdp2GXXaVvTFo3uFIDfuMLvfabcLWhZ4PmliDxUAEbsU6Z
Gzqz0rpvEmZSvhn82+5IVR13ItZb9bdsojF/GlUQhrD5nqqBLPn/nscZwyWS9to77Dp4CVzetq2Y
O+vOWUWCwebmF2oOVetdBwSKY43FviwvNghTr2Ux2HFmxsuNHyFgQgDUZ152zdbkbpbDeRL5ji0Q
VDyzFE7/DUQyhOtvsMfzSLdAMNVsYzs2hU9PL8fIXw17+P6Prz7jqGlIoM7KjYWE3+w+nBJcc6s9
MIkIpwHzjxseO51iiVcQbUWSY7YN0nJPc7nyFepQ0R3+vzXy7n4bpUe/+D2ruVyLqwIQhpDnsAlb
7j55F3M9jY/JKoxBy+IJxKpJFMX7z4NNJ367lh8ppefQS5oyaJfOxjMXA3HxenJ6D6A8Dxzz77Of
hioXd/K2z89xLLZ+/32jIDb28fr03g2H6onlBA+Hp0toSXsYXyLCDxvIU0YWsyz8ut4BMPEkjgjL
+GoSi6BIxh6dIHCWhmYecYZT05aQhVcfx8la519eJcQLQfD+ZZwccwRd6xrPWf+py4SXcT2V1xBj
gtkJpFOGyzYTYPk1C3VNq7fGyeJtKx6gOX9e2Wzwq3FAvNiGCZQa47JpdmTKU8CnpxR3bBja4tzj
Ds+nqv2b6ivC/4c33/mEGXMo8GM56C+4wz7QA3ibjhZRimR2jO6+b0xrqVZ/GXzmGX9ngnOCkNAQ
ZpUQP71cM3J1+NTTQXwq09+vUraoLYWO2PdVJ1wykVIVvn8NR6C4k+AHt/EAxstSrouuLavf2Qtu
YKKqr3/CXFY3eWHj1xjoZg6ufLHFUKGR1D6MlFVOQgWKRlVFCsim9ghCsncDGNKv6s/+0GMWnS/a
n2qZFgu5HR012QPKW5Yi8furOZRR/0YP/u9YVgVqvwHRW8XCvLvrXDspOMBFRVr+KXJ7SP6bbNZw
B2sr34Q0u9RNu0cw8VYACt9er3DfqfXFa5HcKVd2klHyj7cRKXl1ItiBRWEB8Ylna8nERaHeGBBi
makGNZoBqjawQV+jIVub26gdzkpiCDsCkjY3t+6VAypYxkcSYqYKQn//oZRAGChFZWwB1y33Qxro
//IiyEgCCSZBgTJM5vmztIdF4yndXBGxNTxWEagoZW3mKW7VUgwxFc6OscvjFQ+Ix4TjLhypIG1N
sImw69B0vG1CYGsJzdoACkZAKPXjPbYYbsDOV3BHI9NVb8CdRoUwtaMTLipkFuChKxR59UpFbcEm
5heFYCJVzJEfPtdeMrReWJbducp0Zv1AjVQfMsWHgHd6ELJ6S9R9qEVBUSH7ol3FbwzhJFbgxSed
0kW/nOPPqeO3ZgUz8hMuwSYuBlAmkHHzeodtMEiKzWO+eeLrBlocv8GBZ5LbNPmeWoYfO+qE0P/j
GEWc7o/+NzwKQ44ujU1JESETVZ8He2V6LK4KSD3VJWvAobeIRLMi7AQVEEUyTcWYjH+O6eEj8tFU
z/g8Ut8AGyegGMKgtuf7uKFcqvhCFgqxbSKQGaquNtPmmWdPvxcDbPWN1EFIiZbMKRRmselKSUaa
0LDYq5Rg5ihPqtspjnMNzVASxiRz9dXO2dFwwrzPlMcn1i8irCy/AUHfSO3+lt2rJ5kp88lgGwNv
pdnLw5IFyxPc44RJ9KJDcLEXgH1jTfhlwhoqox5eKcq94l+TAsLCUEj0tKKe0SKR60FLFcx4trr2
6Hke42EqTINclQVkZjEACOnBxXjwY4bnPW/m6IIqCQHJfemnq8TyUTX9x2oxsD3OisOkKTDsH1zN
ofs73OSTf9L3CV4+YHNLW1iQ37Tc51R+3Em5UB+sJfiyHoVUOAU/60qpEw5i0gEGbQ2RnZsJ39v/
tkyk0+QX5IDtElFLH9PfGbd+o+lV8CSOIwxgfZbFMwf1CHsJMMcTPbTUi5bp09NH7o+9dv6IUrmi
hoI8FwTVzReKXYO1PZP8S0FbfcJJb/G611Pq1gHlQghahstVLhMj8OT4qG5K3FhqpF0ivXruPKts
Ik529es3YJFxy/H8fie3Qx1LaFkC4dVce+21ZylfzP988ohn0qaX92zktbeKDQWpqron2JnA6Mvh
GoTfI1lucwAXgYn9ZuLDv5qUxW54WVXewzcsGXQizNqxGP4P3y20EehkvxHA3zjTSNXpp662L+eY
ussiD3Lyx/XzXw34gFRaUrK7X4/KWZjkZILlqle9oqj14YTqY8loRuiT8V2IaS/cOelgAs2YAsfy
R8Ef4u03wo5g17qy8NozDHdgykR+YEMawBeF/Q8NimCqVXnNyILN8XcnoAz8la/3wyUzSUmOAb3+
iqcdvor+swkEkzTUZeGyyaXPJbGh6yAHTl0bXQNrszZM1gb9rm3C47cpUCJNSEiXJDnK+XT1FSzB
SdNnyVjA2QiV4Xkm/0JFe2Y5QaTjsSw/idGmt0MGLgbht3UjY34HlqKZJPMkX/77Lq980o2R/Gxl
AC3fpgPQkhI24G3r7QZh1aIfln3Dh0evvt1kmjKHcIORgsM1zxtHPO3dHE9vLJZZPm5quKduVwE+
lXorD5PtEs+csufNwYy90kMiVeX5ccyU83q3kVA12ojgs/MSI6crLnpotlUpN1arMCc4yDcF7L8N
bh21ARnka8j0uc/hlLKBu6TbsmNDtqiPwyy0hNowyYfuWeI/bSSXwSLh5gG8HdREudvTm23CYolH
znW3Lj/noI/RSadafhMpu8kqxx0/eq1aWwj8tIoKAlozzm3jZ+QTLbQKNS73ggIxEBmy7gGc1gfh
v+ObTNeSmvayNEV9PxAoMHuWc6lhfVb5fGwsjIxoSs8PEQfwRh6pFLZseBnlZvr5D6ToHFtgsqK6
ooieBYvxoCpr+IaYDeRGLl45tgX74fRgb9zk/K/214lBnwxVesIb79GMRomAKJR/OcQHiVY7f4cv
KWHNrfeogbJ1Rif3O9zQsm7F97g6IVPgDqqO+vQvKgRCuNyoqMjp0bNPTta27E75oC52t3J6u0HB
oOOaXmCdBJGL9IB0CzlnUSObw4qHZbVkQisR5Oyq7VGz9G5vQcIjf5XE+xM5QjeW1iSiLPFxgON0
0dVVOVnyTL65nSlIhV7tqYbqoC+BnYFR4Oo0dUFf8xFNiZ9xBGPd3s75HuKRf4vys6gMymO5uGuy
B344VS+lXr2NudTZFtQzuMkwAbL5uFtMhuTGTzYhTZe9w7eolGpek8Nmq9hZcGevMt5QoGY/nZBe
MQY0FNsOXXq76AH5BpWU0E+/krXHslKfUro8i+soc8Ze90Bmr8jMrD4BKa1GudVt46gxRc2Dn1uB
osoKqetyxZQmoAfr2QofCj7r3K38lroew7gX6E40Xpfj/AHLn6P0jNK5yWDmDjj5tnIPZuK0igsH
xHCmh602mQ0osBapFioZTxz/qw4C/R2X+Ig9rP2DOfL1zbrfREgQmd+DM2bsaUHenk9oqtAgFdC5
OXlZIDP3VefYflWIYCfcWLqWVupyP9Y3Lq4hn6LQ1I7r3+WjORwL3AR2iwDH4k/d0x/xr1epyGiL
WPyYoA8jgzFfJPTt7QDJdnyH2dTko8aXTz5viELLgYJUMmu+PvRfA8ueZf8wyUpe9VDdEKcJ+o/I
kG8JeKaU2M3E9TTvObSJac1s/kdOgxtsniXmkdSIaaswbbttmbZ6tscMo+5ZINGv6m2m/gz4b5nB
xTplcQbnn5jSaf+mdbgv/+K7D+hcmW4e8zV/FqQeR/4mSRhhmNAGYc7RFp3xLsTBWMBF76KNfmxO
szntpCOaChOe9Yb6IDlSgh4bsjRWviC3DLUeJwmgAsvcGE2q2GZgkQqq/MHTPx9WOna53nKNkhjW
dmjbI+dubZ3VPR5tv6SPp7Q3eUthoBKzeZRr/DC7sACzZDTKL/VfAYD7P2bYzi1N0+jrds6vffal
F9U1ydie0wxlm4E94RWY2RCr3LSQezmmDZMnIUrwjQPOKcH1NGqAu63CbRQujK3c+dFsbxZWgZDz
sjWOdQ6Y3sJGk0+WOe0C9ecQLI5iMZR3ZhcHfrSqd8yQmeqaAon1gYKP1BsmpbksTfgmjJG+Qxt9
qQ8sJ4NPFGLnMyTzsd4zwnpiPizpcvEbvhUAegR0LaVN5KDJkZevgVJBmFZ+fr3D1GcrEts/5Jiq
8Us9dVjEDSGc26fSGDoFxXNQ+Gw6wH8BPWmLu+JS25P/OaMF/I87J40rK3jYnZlcndC7tw0m3ygc
mkdQyL9LqT8BjjuYPM5j4hGs/z8RYtAuIPvTCvGdOZw3P1l/NLphnnwPh+h0piBVWG6szh+ZTn81
xanhNdkyRoK3fPEtMxSFrgahN7GtDb0A3pOmASwr0Jh7YhoUkBBpzanQTQ72Sp8OWWaAp3cLXROs
0zQFPkMlobwM9cbhIncUmK/SRVwLWWK800csDFBTsL+XS3S32+gtX0Uir9pgG3MIP7hUT/Oyru7Y
lYmlU4HIGDde92dce2OaCRFvCiZjR35zX0lUA9CrirDaHDCHP0e3CbUqZQ+vT7V48mJ9Jp6JDH/E
bbktoeFJutmhZHyF6ycV788hS2YIK67Ki/jjJOrec51b6sLZvBsuBzau9izpNBwJiYiHf6GvEKRR
So0FXIP0ZlwmUH97GYknqzvKA0wADAcpfRHklgEEgAXa3m9UUqhaMME50ziITmeeHsL+rD0Qfyf1
BvllIe0+zKAvwHKgdjHsuWZGHNDz6SfCn1h/1tABPjYwBYZxcqEpHrI3FKtG4bqAbeV1vT0949m0
i2wzL51QS5kt0PD/zX+hN7x58xI=
`pragma protect end_protected
