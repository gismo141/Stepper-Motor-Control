// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
cMcvIE3hCYQoNi1CKTNojeUmP0xSDSRewnvkFr8y+RRiiofbK65d6dxy8ARXUWby
L7FrqD4D7zzrfZv1AFXWvbo5yGiLGaIQIzvAx59ZxUqzWanzkkwKKobByHSCCVJy
vs1+GtNQ9qKULyIkGDRYXqnjbR8HJsTXZvfa816PRIY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11024)
YIlfk+7UmNtq3Bq9rW5n8qysI6IX9/VBnSRWBv2cuCKjRxJ9Fc60Gk7AiAN8qqOc
qDD3BeHTQoVyfdLsw7KB2u7bQ263ISQD57FIdNfo+WIS4Qmx4q1lyEjn+JnHJQmG
cIJ4ho8QHcy1Nob4ePLa9rGj1NXCmC/u5/YTBoQGRgEgk+znTuQhzQMO3yXESFaB
1O81pPa7xPUj3APBwKIXFkIvGHQF1248kTJTrh1L/NgQkwwEVsTJciJqPj2Cx/Z2
1m+u4yCwk50jBW5CbevFhnva5ieHJ+1/mwuxegWJdS6t/nkM/llPAwv+mMo58+B4
WVxaIulPxdhQttD6vOLkDWQu3yX4MyctaF0f/3V3a+JxJLuT0/9qKnxaxuQBTFf+
f743wPtGM061/nPsgjuz4Mft5a7WHlp1gwL+HHLYSDB1AvvMIZlNfl4X4JoHaMNO
Af1bz3FTvPmG9Nbc1+9MEzfDuzmW+3ehXFqpZNMM3NNga5yM2hS6EHEO02Of/4ej
EeUn/G/+9rGIsk6qLAobD4kfoUoBSWeEysamKuWrQIsFe/WXq7ZmNanaH0ahak8U
MjpUeEq7wSayykJAfEw56CaFiJxhR+V01ms0Wz6m6Y3BXAKXCh+5TRGI5ej6HaWI
x2o2qd9Gh7CcZV3VuZIqPYALUj3fHQCqU+SABJ2eASt7J+nBnLiyRuM+PYgEoarh
jnJ1fgYYxpba6IbvV/nK87yFqCBFmoCaYwDz2WY+8HXnpwzZvn/5CE6ei6XRD0TM
ubpr4Pt97WRXir0qaqbHyH2Bc2Ro54owEtLkmPYbIXwcgRxcA/22TaIw6oX1mrrF
HkQeuc8xsDXFAJnkHc8rQhWdVVIB20ig4H/9JoMYn86a25UT/FgIg+0jFgXD9/JF
SAuPlfqC9vbqF6W+jYdgVAw1QlYVlvV8ZpI6Hp6rSss0JIsOrSr2tg3nz3PLxT2r
yc0t7Qa8LpFP+fajR1nE6IhQif0mrkPUJn74MEmok39m7+Ki1JZmdw3mlX/Nup9m
jnd3l5qFFH2L9fMT9K7Y02jXGbqDltnRIR+3ijVpRz8ivp/uJo89Rmn7pGY1ZboN
u2OOBjT0rPyHa46y3YGjRyxejFKXTrubo8m9egf7Xt7uYFqgGgGsKMeM0koESYlA
w+F3QxiHTIRqfN8WAkylYN7EH0hnnxYizXz3XO5JevMzydAVALnxpmA4zvFddQDL
KIpHO1H+juxs4k4v63M7SGRRLfzd66Z6HwfovlsQR63bHE4U02R8voftgakFO3kB
DBPQQTeth39V/LdDmlWtmjixpuFLIZnGj/tNKZ6SYYd/55GE5E5JgASmnG13Qa58
ndPDHibZbWVbOadM+sT+dqbIgTq8rIYVDixXKdILlQWMHp3OlOwQlR1pL2c+cb+n
1Dv8I0xIDwExIQlUW4exOgHL2EKak2lKRcVMJBHqjy0KRAEHjBGHye0khoGd+lWC
mX8tl23macOPgQozHA1Bbz78WyAth/l3QAodEXEea3nKTiKroYvwCBtTiEASvRxQ
9OUm7xfwvAlhb6JXfrNAWA71QA/w5skpodU5eVBLmldE/qe3wJUY458vxEtKdLle
swAm6kfbd//Zva2KW9PAVkwwDjGEIbp7CpBGNfHt1rcx5EUtKbxgeLUAM+3z0NEo
8Hh5VROHwbULJC3fy4j9edEgiJljSO/cqMDQ7/G++g84SFmkHg4bjVPf4pwbR7GV
LkiusL5a67tWVLDAllzEtfI4jM1Yt8UIoX4V1w3/+O1/IamVDKNbrYaJm2y+6jSQ
ZlKejZfwOj0Dq2D/tJFsi++W05dK+63dTNB7IbrjnqzETjuGdirOlFSBM6hrdRwC
i5qd14bljk4ZyEpuKpQ5UymcD//fJ0aPntjvF/0Dev+V4ywHeVN/oaN+LVXXPMb3
PoSuLDIxoUym/Og+jc5B5nk7WWcJ/dtEdncXDtNuT1f1robb7GLrRxcuXVI6bbOw
eIjZBFwJw0FjqVxbJndx06xYfs0oDq/aNv1IKo6HV3Xh0sdN5eJIE/pcwZifR5Cu
VShSDDFcxg6CuNCB9wkAvC0tvIxj+Po8Yi75I5NnBDKlq9XfRLIh1canY6cS8VgH
G5pdPGIVj8I2Aik6syCrc+xNg8xEeq6Duw8wDNda9JXiHcgVh6s2FGvlVRRBLjv5
K0as+MimsYynEaDfj77Q8ZoXMkjxjrZ0/jxz0KlBZdc2YlEjfBK1hDXuTHPa/n9E
MZ/thPQJ+ktwRijROY4GjKu95pj4iNRb8d7pESzvWnmlwyIRmB0CeGEQ/JX4CiRt
fsVCaclYC2r1ynb3yQDPNL1TRbeIEtZE1+3NgnSBjZQ7Fg1UqpaJ9cnbdQDGdWwB
M6Hbym6SS4hVXcswgsGoSwqsKHSfYmH+JW9+R4NPozAwqTE0IXw+kYoVoyY6xQse
VS5o+o4LL4pidjG+Kf2IJm8tKLb72XZBKWRncnUd6+HFntH2dIlvnMIxTSiEyhWv
b9Og9YgE7NVIHXpV52i7H+w2RJ+YME5489LS9FlHUtvg8pGBn+WPYh2yEEs4Vm/E
Id22kRWSOTA/xXQHAXTleB98cZKNCKIQycAHttK80UmZuM3sajUv4vZZcUiIr7Gk
Y8HfDf2DT0Moq6bvwejV9Mk03XrvVNrFKzmkbDVVWltl/zdW98BYT4GL9/HBza0M
Z8D9HxdGaBeb3IgS7tl1LkSrgltl9oOS1q0/GIuWzM7cyIYSooqDG3v0Je8OKkpk
wYFpVA7mHgDOlr8imXz2tTt+r/Jv1EcTvGL74n/bPj07ZpXm90cxqkG2toT9Q7Ww
UBOUL9zdqxSolfDpu7qSa9POHqHgJVrrvf/ShSA7BcsH/MzEzg1iIiYq/lOn1SeQ
PA2KTJ+JgtD38ZvbtBgfJaSRBOMNfJGIh8UQynHlGNPHtiWSD92AfPVBEz0Rw4cX
n2OVzPzWlNsoNWlkyXn+QiBlLzpgOBoAndvHQTfzmQSqod7pmBsFMEfDkHvs4K43
BC6aL64VHIUHMseM7iZTfh3kd4fzqk6ND5R9Npl9bmbAQYuQu84lD4ja5v8lmW64
PnN4SV6aute53lsnjMG1WaymYMTajpMuitA95MgKUPd/3y9egvAGVaHo7ozdZebK
p4JlZJLiWi+hfKPZb/68MzamopyeBjAaiy4BOzcTJ1sMNcyxKsJ0AqODgF56Szwb
2bp+8nZ12DtTv1iYSdVpEef2xtWVTsoSjZR2VSFGjIWGBn5RM3qOcDCiz+rkSV21
a1l4oXzGvK+smuVc6tVv6Tn9/nnOPfxTw89z3VVa/SwVTQS8P0Dk6JBEyE6sutXR
qXbX17ZVoK1JolkPy7JtMkMxCz2tpoe4D8h0X2kjbMCz/Ecez741r34StjYk0ev8
jjoCMp6O7hdNMdqRRRlfHlAfl6ILOVgQjuagBbG8/e0l9q/ADPee6+BktgTbC8d6
VsYeMCDz5AJ82LrbMIVkKMdz8LA8a5LP7M8QM1zWatHOCne8139oKYq9UDk2scfX
LtZ6BpCKExJrT+VbNnYqrKk4utHhnby7kz6wmQuuYM8w0Krdw1vd0sr5lnk5T6TR
5eSsL9Dh14TATziD1N7ejxMwWRsQygBFTmFyOXfNXLOTxv17x561uQ994XwWV+93
VX8HK7fc+Tgejlgbg6NMlusxQdC2gKPlH8fOyA6K8chPjiyrxjg/GfKhr2g5JdFg
AX6yRwWbMorRz6FZ0SN34tEKVpBbWWe9j+3IJw0dszn0bQw+Q/uFXmXYcsmjEbD4
XM1UWUOJ3v+yD8o1bRqJ5Wevj3hlxfyGpg+yac/c6qsMQxt1scT8keRN/ye1eoiG
0aHtTP6RKwF05NqLGqsx3fMLwAuo/hjN/HrY2jIW8KUnPlnv47WcpPo+obimM+4x
d9Eo7T/kCAKSxHuAF/cWdtjjIbPq9H4hPyO8Ro9hXPKDSv5boJNq/egmMGrimK8A
EDV7NDDZlVrwqB0I0p079N3Eteap18EqsrcnHqcq+TCmqVUgXr9feTCkW1Ps/By/
rKextVJDSzC0XWZ6NtOXJlBLjP83WAUqW37CfaVS4VEOhsqggx9564GyT/EwLfEt
5nMGhcxcFAAipP2xIhDxAE55L+oxnO0zQU46b2y1xS4sS0J6KZMRScrRDi8+XTG5
wPga1pimiNEUsrFB2+XDIULyKMX2EyG1NK8aDm5pPxwH/HHT/fdPf9G1grzvZBw7
RuY3sX6B4R2QDVfl3FXKQU5GVF9ZMuynBklcfbNCCis9yDZ7U0BIJeq/axkBq+rb
dyw0cEhDllYvRytrJ7v74/PzV0xjVOpYm46grg90nt+WN/JFhfYS9SsrGHAtwiD6
WeypxJ9+0ngz9+VlMAErLtVP5KKBRRlCMw7UXRb8G5iVqrxw4d+CVZ702vHEJEw+
U//1HrwUzZmceOYxLfy2jckacBUB91BAqr5E/NptIrZ+4vNkhjN3pCDQ3xkZFZjh
n6XOKPR4C+9Q2wrm2DBA10m2g3BLyMl9a0PlgfEtbvWlGsQUWW35/abbi+Ph5lrC
40hdsYOLVPUNw8TjCtLcn55agtJ4vtC7rHGGyWM7+pX2L8dMEqVS5FFjiHvkjews
qObgg1ZQCDNd00RFBQUpNkOrkaKcMkl3av7Zj4B0MMmZuQmqI3a3im8+j5xtVS6e
L14/EZr23BAD3RgtwW5F0TqOetLW23W1mZubS7d5YF8bYzNYMXKElkP1R69ryfsa
YEszgIPo/0+Gc9Lc4QbebKZwfseG4OYiWWwdWf4oLM6UwSW8jAajeTaqN57tkGhu
mVMM682s3ocrID1RGqdfqj/OTlROumYmmvz1MkGZA3HFQQuNrtTEnJexV4in2mjm
fULECirwD+1p1vk5I7Iuz8YcsN0zk4FhNpy8e0ivibbQqgtj8crpnkXTRyQz+zv4
Lk2JfbZmRFisrRQ1AdmKbHJKGEpqIn0HWrEJqHbMCzd8P2LsNp5HP5TbOCOFVrv0
+WiCZ3G2hbvxGUSYoYozj64ZLFa9FrppgyZtD2LVxe+FEmuCEvX01STKhvq0Vknk
NinfuOOOb/lBBZ6GrxF8Z74W7YEtNR6Y85tZvjvmBxvBitJt/x8L6Mnhug8tyuud
32O8ZSHSpE40jayN5Krp/7LxEhyVQYc+N/vmfa8SfXURv5PggbWKW7JiE/QZrYzX
9/Ax0w8kkflVOYVnZWZB4LJPi6ltOfrVbE6S161R9491AOFEIitV172pjW23tdFi
QejaEdlh5XPIkDXfoNNN+IHKIhP+ybGsBAIrifRl34xUQ3W44I51BESUgQg2gDWq
52ycB9L42Lz4/YwzGSixu5L+qv0a/eLlQ/Mjvr9ZwZjgy/qhZdpGTFTANQnKc8/0
VyHMtr0NclQZhQL7ci2DRZa+hD0b5mu+so5tuKFXfhQrldCoAeTFXv5psq4X9Qe8
FXL4jRCMW5U1qgS4Jpa2xwPTM5uJok+HDzPoasCcxUjXcPHaxucRqFIGB+K2jItI
ZkqHK6dzODIo/6kK1lQ/PXd2+olndUBOxZerGvICrBVUpGt+1le+Vm6WdoooMPXu
ojEAFZ6k2RBD7kit5OoM3yFECkmsF+FzyW/pdGyB1b5V+EBhPeZVh6eJVVhFCMpX
QluWP+/SUSGVMnPhXIYFG0lxkq47ddrXQ3PKGgORLlSzd17wS2DL2NvxvLRbfU54
23tfI908Ycm0nNbHDHlzMIsfnMy282Cfz0WEyKS1pM9UtdY4jh2f99okLlYFcJZW
6S/zHQXnGMNEs1aDcdkb6Wm8bDcxLt58peTeiqZRVkkneJHaT61RCLksHkGhgASk
pWzYQWlUNeVyO53f6qzvvVR+3ElBUVB+nTkQVWmAwai8kFAe13Mw8MYjsMTwVgRz
fO7mizp6v6nV9yeYVb50Qd/W4o5z+emYCTxZ9jnwCSEIIE5/WV7lOrDJzYRIUbzR
CxGpUWyLt/ceWUAYBis0MuG8v8hhXvsR8U9oWPpHuEwCB9DCKr4OuYSbEpLNEFzG
Q37NeoQdqkjdJaXDDIgMhqNNyu8oJKbV0wzavgD7O6TxCXgdzZm873v2HmlZu1YY
U7e1clw0clKhDwevxmcGr1m+qJs5Xm1Sds8FZrUwcVgH6dIUkftzQ6rfaJ49LmiD
ALp4eh6RxDwRyklCUARbK7gm6v3r6ETcALLQ7ELjsn7q03VcJ0ZsoQX9/JyeAUro
rV/0SGA8i33wiY1d1Jz8oZ/slM0vLYlTCTRcGxx+gj9QPNUYJyWh4Z29CCYMcJN2
7D2JIPgXmt5P6tCYULdUgU/NbdlpXeJLux++X98K0D73ixckwhovT9e0MR4P0E9j
eX1Ttmy2b8y9/oiM/YQ0MG9MB58den92hvJnjN3DiiTCfvjMmriN4/ETYQpEzkaA
4SIR2kAGqpi96dBqLFuOKo1pDy5qMngqWaeZyPDhgqs4PErW0cvd6aAigDCAS6VD
xmBaGIwQD5QW8Xo1iwiXpRx7J4dMblwy4XvQoWlv4RLJOZ+Id7HIXOgWwMBgmeHq
BhKEAu6Cy8bsR13gmuhagnZV3ifnzoy7quGC+Y6OhpLJOsQbCG6oxtmOdrx+SobC
dsiQT7vBw3XlhQx1uwr64hJdDctdDdVvGrOT7cWBwaFAE0IkoD9xOsZQMTeAtbVh
ZrFIF6VtuFbmGR0EA+HieA2j6bhlztupTx8Wfd7ObRihRPKLxh/WUuWBpB8NAnq1
sPMUadUSjee1ad3Sa+Vb9cOpjjGHGBIsncaGWxfz1R4uLF/SNef676dsY71jIvAF
g5dLsRtYgWzEPPyKr02GoreycVEEd8LIfghZvM9DETZe902jXdXH4A+6vj+cIn9b
ag7mznbo+qXX1m3tSo0CD997KRWKGLe2edI0T5EKkJDPzCh9kuqxrJIcthyNK6Dz
VQDjQJ8ZftX+uXtTofXYd1tqKv8IYotNAhz8X50gTsPuy3x5EAXezCgivvaBLhnt
N36hXAjgSCdktiMX4Ewfu+sLVWW6rkooMgrPdDfoOBm+kk/Z49Dy5K0pC4RWIROz
i2b++0xbakH3L8jMWjjbefwK0LhcsLWDW6icgYayubR8oiZ5lanUT6G1JXEAAmd0
1FbU/HEMGWFlzBqiUWI5ieJpBD1w4vGsR1Xm9ZBV9tf+QzM4MDLM3q2QO8wbtTnd
QOWEDoN9bUXv8n374YgN89Lutmkf6zS1XQkuNNcYzRUGVAPfsNZ7Xe4hcBqRkgbi
asFR27DC/FvfB62tPpvltmknxYl/5MHF7E7MfqH2oqTLgqO9H9xSHWTKBhZXqDow
p5+7uovfZFd5GGrYC691Xm2/jipkUjcqUayHrQQ37Uc73ubN29EN5SwgoXxrLaf8
eDmTNOBrSvQi+CuhxInKec6nz+4O8aGgINcya5HtLceflzSkFDoIBnJ21GSE0LfB
pLXqe5dl/+3h7Q5MPDeaW7ivvFOovF3N6NQtOwmLh+c7A8iuRqZeB3UQS3iqRL8H
V2O6DYI+eEh1mJKkHPkP75odUCjG4k95zWMXPhSRNi2AiQcH6p+XMou6f6Qijzex
wIZnv4WnK25+oCTE+0cp5u1WxBwM9eETAAVN6dQT3JJ7roAOXQDrpdNHdtYcvWbv
PP1Zkyqy9j1t37e/YMVlcS8757WeYYXJnq5jusTcyHChShc6xXuZViaUq2K6fHSZ
U8NNQuy7pPHNgcSeGiakHKmavWH/iEydEyzpNp6B53GHlECzjYLxlr1NGXCWYGVt
KvU1+SG2qhyhRZvBKwyX4KFkPNNq/5vKNs5q+OqI1jxjBD+KBqOtyBD2PHKYqjlf
LcQxDQJaEefUihG6nTuuL+DKhvv+/Es+ChKtPo8agJHMibQpElW2PEEAj6II9qDX
9lPs/411iqpEUuj3SxOPUffrCojA40zMrWTomGCk9J1CwT7XtuDBl96/5raqsJqc
N75qIjvY8xTQuSKsPyebvCcUpx6z7R22r2dH2mQ7wnBuJV6U0DPpsrxWyvxAflcd
N8NspDVt+gpZteIOhyjP6rzQUjTEdsalqJqpNUaugVaQr5qLZFRDWlHFaFPFGSUx
UXX66ObR/KUU6dd0gVX5GRIeHIwqbXkKr5sorB6Nq424OuRpIZExzKkXt2WB0Kxp
RmHQ791QEtgpH5kD7BWGXInNM5BFJHMlLV6wo7LNBCv7PuE/LMd+84Idii5ig9cS
rFPftXBYHBgBLOWo5veCHrljD9Rjqx9/GOVgGeksZo/8fdFWdUy2QdEcZyOiItZm
FqZ0txz6ipZ52V87KOMaTELm2cZOEYebp1yvRWymSew3HDO4IlCg2v42HSeViDvp
nZYwxpykS+xeXLOe9DXMNi5aKYXmUmKcyymJzWVjzpK5PBQvqqr84G+n1Pq1zKE2
uh1AtU15wrcx0JHlSqtWhnijRmzqlc7T9+Fsgyl9LO75hvXIqUTbzAFO4/03JDb3
r6+zE+bipUjbVftj3nfDC74Ic8zHdTLfeDZg5/m0MAGeQyh8k+ALas/KrVAympIG
KuSuDW81Is0Ec2DH8Rq3fZ8df+7kujxj0v1eoSgLPPDO8JMznx4MWVTvDBjZNkOV
1lq8ia317ypI4rt0SJv2YO57pTMzYh/tJK3zThmKep/fp2keehtLz5DR8XpZ6u3E
mehbhvo0mLuRD/KLa9hlXvPUMb0ztt5hMVHWusufoKBaG6jPeHICpbiekaLUFgH3
XmZzCq45Qg4RxpKpOZYsps7A2MSDj5AjJLzuiCYe5TCRq3kYWCHxG8lrZE2N0XXU
PgMrANr8PXAmjVMcSwW/fWVb0+RebFcVhfMTNa1W9Nflhgxap0ePxr2noyRDazwZ
YXE5xjUbYNWHHEqPK4Wh+AVmyfqeRg+OLFMs+TmeB0fWon6KljygoHLWYilgUcXk
up+4yJ/IwKgDWo268k6RQNrss2x+aydAcwq9tYRVIx1BMJU0QXpTbkEh6wA2SeDu
WiioC71aQFg6YMRPtOhS7Z4uZ/UGn5Rx9llaDMQmzVmtMOLQlIkLt0tBAZphSALm
Kcyn0EAI450hlZv8RD22KvpIXYGX+TmPkL7G6JK55EwhYUbXOZ5JH1BL0yQIdzd/
dT1RpR6kcfmLxpgJht/9sq0GhWkNpk4FgV8JVqmQmVELcp2P3KskJMGMKcCS/LGz
vjUKnGw5nSfHAimYpZCfUEvWn+nHGQe9EwUMPFy9dHRoW8u0hBq8YFWJFDRKR+KB
VC+zFTax/ma94ACEiMlNAS7S8XM6jFnMM6NYl211p4y05IfraaGN7DLxxHnreg5a
BJPtOV9UAIqgcbd3JSbmB7CHd1haDu8wFBrB5Xlcg4NdjtszPNWXYa8LxDFFH8rT
mA+AWdLJVli5EPGYqNACUKQFDZ9E/uRxcFFalbwjUICSGlSix4lHqPfOVh0LWqml
2uwgPzlBaYxlRgGsgmZr91ZkYm7xzn6LofoJvnjdB19m+tcdVcsIqfb3W29Mf1gE
QLabqsXlpIZnUaQNIBmjUN4fBNFoP94M3ftX6ayWnvxC0E/7Z39tdVE8H4EApKKV
hXbq52REmwmjcw1kDx6QqP20THsYjcT7qVpZj6gFXr0+FmqQ7C9Zcr66qRjZOT7I
q5l3hdnAKHEWP9aU4+i9Dm5IOUdaxvP5NkRZNarCuTYwE7qUzw/fFYT+7zM8/xuy
6ggxLnWz2gIQPft/9TKeW3f4ujcH1np8R49S5o+jaNaWIAAWe4CiBITeJH52zjoR
fcTgsI6wF8HDmgJAQPFQCXk6MgKjMEbc4ClCsMydoVgdbGMveKcVsNJWmH4Rym8g
TpSbvpAwF1VyswTixbbEYA3xm81sKKjXx62oL6MQQMLPRPekPWFpuR808dKujUEV
6x7eZOL/Hxa9pSm1LYZ+zd7KH3po2Yv9wzx83Ao03vV41yj54mvfwy/LEm/Vok8m
1+Y+yk605Pjg/9HwLlWc8GrZT/vhUbaMB1tqhGtIbGpnrIrB8Rn0Smz7Y1BQskBS
a4BAEzZ8QEC+KbTs3R1wY1zOlu/SR2N01iMaZN9z6N2VPMtUx6xUyjQ3gsYw/bNd
ukvOpJ7U3xYH2Ub9Gx5uTo/y7BqFsDazKyFl1vUgzM0SNzARkeY1GBhzhDPnR1TT
SWcf8xVPhzkJGSSEbcZeo3XGzznJrMDGRoPVrnvfCBfJRKpmPlyi/5+YI6/Sj2et
n2B+lUzMqT/A5bRCLULT7m8uhLsKrpc5aEZWOPYrYoI+UFR7uNkRsR8ZUyX182Ph
PWdMhf0Ypb91dF2TGi7wroED9pfngsbjKejJWM8Tioxx1ckeZ+aeR2+X45Wqq+jr
3pbaAfqej4bMeTB4rSQrjzdy3/XLoKh1PBxjcp+HSRQBmB7H/uXSYI62Ld+1JOS+
FNgUKjcp6cppp3vRhy/1iu6Jc76JrEsDgPzxdfPv5Fo0O0SQYKU6lM3oiW+f7l0z
AmZn35gRb/DGayrAz/mamN/kATeTxJ3RxI87g/7qd9Au4U9vVhtOY6qWhYIq3rxy
vkpanYavNMGl/axfXhR6QUr70DWlDVd7CkXk8AhWk8Y9Ca2ViRgnEU1dmkQjz7bE
MV2r25cv6xlgA82t7ac+LSiKE4ZhSuW7xCXqfJEugoQ1BT5KW5KnS40RDHTajPYZ
ijVUwYu8Nj80r5Amr9jdS3jhVhaWDil+ACO9/Raze4giWcZO2UD0cpw6NqZlT4ae
NgsUPX9+JBpvu7ZKtMsFbefKI26uTQ2uHlsyKIDwJscAfUml5b6ufLn6MopeLFLn
tylNx+VUwRzSQnIKrgGj8+wbVpreQxhx2Ava7IYBO3FI3DnteYGwJfiNGUqc6E4E
/9hj59e6YangJ9miuRJvxvoZAQKQ23B2c1dNxpORFA9nErlMhayQXJVpSLPdaiay
wIYy4rXKKNJBYykpxolbM5A4TMmX7tSq3KoPTEDH3Yt2QFDySkFLGgo3ksjxNOKR
ihVj7vuecgRDj+4CEPxJs4zzVP1E47/iFfnyTPsGv+GshddT+2pDDc9xPuyTs5xP
nOsi9trkLSrmlJ6Bk9S1u3Bgesm4KgXtzu6jblZu6UbfJ2/aUweErdrVp44BTszI
GJ+ayKEHiEdQGPacfmbwQr1o6Fws+Se4BCa5VJng/uGTOrK/7l+rYN+O96+suwEa
LnJiR2Ie51rK7w4Wrs/KI/H8bTr1qIDavW5DT0QmmWLQQN+IFimP/lh6KAPsBTFm
lnXi51SSs4BxQo8A5T27esN12zzw57yS2QeHdjbbizXZgqmhpVnUMcXela2Oat3w
R7J0jYZhGy4r8Jvtgac59g9GDu3ReA4Gyhk0+XP6bXgnZPHgwI55wsEVIcSoF0FF
mwt2Z/MDV1rZ4sr/n1cn/qGcow9zxqUJtNBSQUl+Zp0zSWziuxgxjX6In057cc+c
ZLi5YJEJv8gO77w/L9zkauyvZ9C4/08B2Doo4EGkVp866HKxaZo8pbe11YtrPTIo
U61yaV82xfiKQHNWcw2nvSzd2hwJtTnWB+jzR32NFjvnmzKn9lVnBEpJRL8qONPL
iyUVhAF5J3QLb3smcVxYkDYloKSwCh0EmzmNXd4J0dibDB2oM41MbDO3GsF7fltR
hAgpvFYvdmS6h0BchpHI1i3OO2uy+xDp9fnnkWF9YWhCJWBKDnCyPh6ZNfiVAws7
FxtZQXKdKZKIZqE8/D/hr7I3f6Y/ynxDdCa11x2dlsp+EwQlsoAQCUlHrvRNOrBX
QXU0q1sEdyg9oM46X1OwHCDhYWE2NuJcfxylKuyamzDw4mt032vt1zqvohmp7tgc
6NsLEGwfMI/tLzhWrfA2q3ldVZp5R/FN50GWlh+R4aNELVYS4xaBTwQYVdBt4cDT
Xrru4GK/g9w/LZIYH3WgaejxYbPDTypKmyZzJLDcGo8bL328KpnyKWYZTmf6WHVh
+oW+uHkZURegyVcuQ5lcIuVJJgeZXNWaJhEhkoDT1n5E3kXZs0im21I2rTkZQcoB
0Rdeu3iTeXkjve1SnFWtF0ACJatshnQO5cHadDbxxjS+DGVShM50Riy7TNy+3/gC
gaoM2pnkWfXAvU/4x2ecvjJ0XN62z0rKYh/2NK9sGiVbXhTHYk/8XXNtVsOk+ycr
9Ej65UI5ImqnxHUarLPi1df72oS6e0jxt1QQKBtzWVByLjEePtulA8hjM2TW6c+W
VHb+LpnqbVL0Tza0bnDJN9jdPEAWX5qrsnvCVXYW2qafKdApAxJ4ObcM/yxdvjNL
q3N+B5y0wAoPs3LhFtzGLku5SUhkDZ1fIiqlEz+6tiN1w7zOE/PghsQNByhoIo8Y
RFJ9hXDdBRtZa+qbLSbYwVdH5F7vQ6CU7pKqqH3bpWPEFjz7vLO/x9VrDftTaaz7
3t5klNA+rk/469cO07wBkiFtKQp0k9mug1w3HhvL+pJy9TY+2EbFotdKFFAJVxAQ
RS1Y8W6D0CrUtYbrYqCLUp0LIpTmm7sbwKcCA/80i/5zKqUwLDGh/DaNeoQfl9+x
+vSbqt3W1iiGPdAMAccPczUxcrPsEnRUIW3efe8UZJ4XoJgZ4PQojqUR3unKec15
SzD7mPahTb5bk4K/LU8t8i3IxP4qygrsPzShSjFc+lHgqhllycSchVHkR1Xo53v4
NiGXnhss6+Tf6mmv3JVHLuqeQ9ga0VzM3BeuGLoDyzH/66IHa0MotrUDXqyoYvud
BOmQNaeDJy7wd4p9bwXKCfjJrZkzQws+g4T0fPT4JHUY3HAK0WyATyc2m2qZS3Ve
VhzzSooFfV4uDCy3Lb8Gs6i1S5Pc/uWpTh6F9HzC/p6tixysp/rmj2yrSW622nuq
usaGMW1Ocr8qLTUGw3Dm8Z8VU1wSnh0kuZgOg1Wn5PI+9h4yT+tqSOi99ARKIcJg
fgnNjOEy6J56drx2x6MstjUgZMzB39plcU/N8P9jO+RkhbW4N/CzwgcpP/sOIMY7
TAhuwPFTfhrxr2ZjEAL+AlnmOsmqIJ4RfyuN3q0+LpRE7LAoBQr3H/G5nBgSw8sN
v2xmSHnztXvpCQDdYn3naTgBKl8ibfmMRfXwjygKnp5YlitCf4JptBk6n6N42ExT
CrxmW1hpgEMLiJ9DNEFS6683rgiQ8qWv1M7usVja3+gwdPQO1sOHGLT+E61+sMDJ
KcT5ScYOvKfowldLS+Gpv7JTJVBXRJ5mM00jq51gb7pFzrxmEzqv88hVnmoh+dZX
lCg/o5Y/Tna268tR4UB87bJIdk6k1o6WsnlU/i1u7BEHgUbk9DWQKmAV3OyxN1K5
h5rrRCPjO03TnjkyeEc2iu+DLQnsvytUoFNtfkyhYA5Ir03kDBmuREzOlpByvUMn
Plp8tAkxUzOOnQxBgCCUYpVeyaMLvugO0B91Kj1fuXP7gesLtSAGyl4G+WJulMnZ
oJDvqhuFGqKBireriA+YVg7XnL7TLsjjfJ4XICdK9Fc9XX7TLROoMMKa3RsfSzTR
mbyI0KWhMm1e86seGixNJjy0saNzq01ZkKWs8cNOMIZhJqGHMbttGFog7TOIrUUN
M0hnGH88O3obbnkfI5PTYiSiXQ5hyNMAwAjOoPBsHi01jU2vQjMtutLM4J7IusKI
3muBoApmDEQkqXMxVoL+sR59/FopQx5NVgPHHlAnq//IHj5ja3Au7yZeuF4tUCzg
vgYEJG68yRu1BQuqmhtVahOdPMDZ7xSwr77H5hQwJWheUlf17+jOpodHjH3dHBSe
VqPQTS0mELhU0vo1vw1Sk5vhhANMQXjYF0nZRA+X1NCpdDcfkgFe3+5Ho4a6Pbgu
POA7mpgA0By50inzbj+z5RTNb4ptq6lqKOId/ge6zpp47c0jgjQ7Kw4DCeyH8wvA
PQTtni1UiZ4bH1tnK93+TNyJIshqW8Lw5E//wg1O7uI7+Mft4x3PlHfeaRCCFbmv
EMJ8oqQEsTYtaeswtZqRULApjHbx90C+Los3eaZijMfk12eofcdnSLRba+ryKfuw
+kfB5BKMKzD8O1w+/GuXZ93DqfqzZA08Vk3jnfTLgDUa2SNR4//yWIVCvxdvkDYC
bskAjk/B6AEd7JmFkE+I96npK80vvFIcA7Qmmxgt29G3p+qmVUJJaAuEplXmoNVv
ZDM+h0j/XxOHodE22toR0LFJUVGA4vJZKPF3nTBSvuDxPJtmNN81OLta6Cl3ifcp
66OpTstvpYLwXfhp+dZQLKo153TvidlnSRrvWem/BeXUy0xprAUSEdyq+zk0SdHJ
lDu+65EgkpMPZAk69YKB5iraqqgq3PmqdM3/zXC+VLsepMzFVgKEmaDy3S/UjYDN
CowixbW5f4V+3cSe3wcf7zXtDEEdsBrZeZvrHZbCDGQQ8QY1070wU/7iCAvqetNQ
FVNK9+QVEPb2+YY9UnUX375mqfGcFAkOW5zPqI+/DFbJj3BRBZ0DGayErSvojSUC
tslhrUsUES4F4V9Z1PursxYLjeKKa/Q8e8ktElwRiT39Xe2dQUEDd9U8T15vrirt
oc/bzARKVczjCFfz3egF81XGpWNjiSYLDxWRNUtqsoCJKdIed55kGkp4Bfr27rnP
t8wB9MjDdIfD+g/fRXmDvz+vr+VQv/nMAHTXktS2y8d89tN2flqNRu8XljaxC+E9
qF8gR+TV09BPwTuTQKSo71Tv5odcN7nsrxDoOX7iOZ9W1vyJsiyUw8RKxWWxO1DX
bwTOU0UCdN6q/GlnE9DrPl9Lg4OJARlyRGPgoHPJW8Q=
`pragma protect end_protected
