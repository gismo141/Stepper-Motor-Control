��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�>	��h��H~,
�z�*�M(�b	������LV�laD=tp8F�6�!�~�\@NQzB5�1�kR8�W��7�����e6� �����ْ����5�}܇��M� f�/�_�p���Y۪�^�ow��PS�*'��,e�/�W^j��������ք��ݜQRiZ�-
�}u�d�|"4�����fTD~e{�I��ks�W�oKG��]��6Du������V���r@�Wcle5�t��"��a�ǎ����"b:ٯ��O�A���k���֩y
�^P��}cC5	,R�W)��ɑ"�C��Wh9U�sɕ�B{�T��'���Ч�k/Ƭ��7�kֳ�q��	�c8Y�&s�mCM���lZ�~>�f7@��(�a�JL/��������Ly���C�2g�& ;���ս�\w���Hu���4J4Y���!P*Z_|޼��1xA�/���m�������/&���Cʿ(
��,@�d܈�K����~?8�d���s�s��c�8܂��l���SX��G2�`�<Tt5iP&JP�2�8|�1*�)юa��А�t������p���������7?}�s�{��־���l����M}�)� _
�o��&pPW>���X+R�T��<�V������4�\-N�����U�g H3$#6
�q�֕�,Wz}��E��ۅ��Zdc��(���f�6 "4����a�O̀�R�mrM��?��Cgh��7L�����43K�ե��Ƈ���3ylc���}�Ū�`O��b��R�|t�����.���!�F#�0�}.*:"���|�����Z:E�\�d�I�\Q0����v�֯w�j����Ć,{�+b�Q~�X0�h�(D���p;蜁�!p+~MP�O��X#-t��f}Ɏo��`R>V>�����^��]W�X$�7ˀ����KҚڥ�}��7�����*�דyRQ��#[�H"Q+���A�ÿD{�@�
��LH=֜B_�,g�B@P�S*�[f�y�1�+b������N��l�e(<B��R����(�yu�)��?����O]��EW���(jʄ��t��G���K��EӮf��_�E��vQO�e�ƻ��mՀe��L$�$�=���dr�:�Ru��lJ�]��Ʃ+Q#F�o����X,�'do;���1�~����-|����Z/^�(�͒������B��[�d3�+��EO>�/�'����H�q[�lF*@jA�o�P��y%s������y1�x���֫T ��2B3����9�T ��'�9Y`�s�r�3V�l:|��,cX�(����t��2w�osG�q�U'� ���j�wM,6$K���.zsh�G�1Q��a����H���l����x;��\��b�\���7��[��=��g�茬@X����|��K�cg
�0~;J�쉫E��c�@��dK���NW9iZ&��������rdy�����8��6畄Y/8;L\0�iu�IE�K@:��MD�k��v��o:@�b.-�6�?�Q�`����Q �.��څ~�嵨�k^�@��e`Z7�Q'������Y��L���]���V>�x|�vR�	����N\�B��L�����_�g�:�[<N��v�%��{�s:_���K��v�G��z�c`�	ma���v�u�1�<64��:d���3[<6 ������߳�V�tX���4>lFx�i�d͏$>e�60f#��h�G�lR����s�����4���ZƤ Ќ*�b
�����,g�A*N7����f~ �-��+%*^*ʀ�d��z�#�Fͽ(��4���FYa���5oi�.<� 7}{�̼�P��/3s�4��64�(����!�)g%ф�bwG�/I��ծ�����]FbR$��O+� �T��c�Ég�S %K!t��n��
�zZ'V�!��kU��|��i�n3��;*C�:���ܵå pE�#�*7���CT��+��)G�$Dxĳ�M9xgx��
�B�+n瀧��N����*��HE4"x��/"Vu�������W{�z�S����}�#�A����4�tW��ވDy�"�T�&5�	�M�4��x�o4����(��#N����랉�JCdYB�) ���-"���L�.A��Se�2�UeP}��A�fM��U���̐;n*&�oR���{$Ϳ��,�4,[`��M9���dC�i�؆�$��:4f���D�D��9e��a(��da*<����P��͜Aa~5������r}5��Il�u�Ԙհ��h��o��lR��bs�#(��q��n�Q��[erU�Ob��ʓ�S�i^�%,�E?VWM[Pr�L����{ [�b�9Q�i'l1+�}�#)�푇�D�CK�_?���]P(r�7�UG~�����6�ڐ�d�j��wt!��~N�2�T�g|�OF4�ߪ�O@pz#�)�G�=&w��-�m*�o�n�2�3��?����-3/h8"�����<� �`߶0�pؓI��4Zwc0��'���hR����[����sɒ7�?<b��?HS�5M/'LM���1�,c�m �Oj¿Z(H+��&c��h��9��w�KՊ��R�V1���:�E,}�I���Ӥ���<-K�	ꖪ&x�)���5#�z�T/�{�Li9�T�� ���y���D�ӔQH�ܖg�=�j�&>5�H�wHjIh�\���S����=���0��������{9B�������u��+�J"��	\�%l_ZɎ�ѥn��R�bk���M񺡘N�X������xR�����R��|����,�,r]���0��`P�_]�@ߌH�H�[܅����34�ᕦH�f?�0EԻ��@��V2{���#��3@O��7 -<v$�����E�ˇ)l7�����st%�n�,lr�5�
[���HW��*�q}�r$�@4� ��NR������k���='�t��t� ��C����hI'�q@��r�q5�|�C×ڏk	���I��/׃v:B�N�O�|Dm��b��m?�A��$�A׉<��^`���6{�}d>+		��.�9��W�oq���DX���&�4_�.�;��@�-iwX5�'�<��p�S��Z��|��l6��C.�6��9Q.�b��j˙4b���'�ƚ���z�Q{_�#��hS��\��Ə�\X'��+��G���$�`CNFhC3�D$�ꠁ����.p�x.!�h俩�s�8$*������e̯[�V�s��':�OY�-���6a1�#�_���lhrw��5��+�ouj('�+�ί��+��²�dG��`�fS�{r��Θ����*]}�;��K�v=��;^�C���n1�������)��T������m�X�Y�<'Oe���
"�-bI����YB�haH�/L���:n�k�����7b@{�����+itk�Xʎ�l�@p��$Ԍ�3E����-����]|�=��4L�����xi�R����lqߡ��yƻ�@hw��A�J�TD�s����s����-�l�Fb�Σ-�H�F����
~��Ѐ��f<��x�m�Nr8K����҆2B[�B��9T�T�FP�QZ7�؅�䆻S�'EG-'T���wJ���uf�<��$�а#v/`)m�#����H������I8,�8���^(�u{�n�E�EF���U�B4��;]���~��r�:K��� ����Y��q�u�	X!��^�s�`�N�+2��*�ѱ(V�E_�lG�-4oF��������M\��/�H;z�L�!fGm$��<��Cp���qm�|�+ ��rw<����3��?D�7��..8�>l����k�ѩ�Zc�����(��q����9�0����B����$�`-~1M6���ƾE��EN�{�Ľup��c���4�
��-��S��<��YGa��z~Z��`��.�Q�PfX��҅R�w㧂At�vN��c�e�����ė�� �u���5Mn��Ӽl{���N����&ak�Kx"�xƻ��!Ж�q
ȱUޤL���j��0C,�R}+Kk�O?�(������%�=�v�pP�ښ���:�����F�S}K2�A���$�2os<�x�W\�<�y�&=�ߏ�k�	$�H�d�a��҈��Q>� T_xލ��r(o��H��^_$�w��@]��������ɘ츃�U�=mp�v��L�(�L} �A �)�+��&e�U5[�9�y+PQ��7ʙ�W��O��%�K���w��$��Gm	|�Je��6.��@=��T��X����]!���*f�}�:�{����8h?��BUE�	���'�k��@&��O�(k�iE����^�vW� /��id�ec�8,�2��#�?t.$�݂���J�[� ���%���I0g�QfR��L�ʠE%�'�����XBt"[#���U�2>2Jߡ��#�pE���~�+V@�8~SL�ɥ��/[20�I���l]U�c���ҭ)w��1�mY���;b���������H���T
`ћضp����"Ph�J܄T�Q��sk��7��jp���Z���/u��K����@����P�V�k�2��^֦|�Bq�����K�j����D͡���ݷ�W�yJ�z	����阐2�B>V�Z�d�ԳL�i��Q��z;Uo׬Zw�gŮ�"OiR9�j(���F�7_sh��}�l����	z\[�.]j�
����O�k���q쑶G\�Ϥ������9AH/F��v<�ֲ�����S���!1B��X|�(��~ˎ"��]me��U����Y�IՈ��Q��+$�]�3�Ոk�#_/L�uR���ߛ�ؠ�
������p;�¹4y^;ʊ��@tk�^���Z��6�gDp���ϟ0���S����e+�g����T6QƢ�4b,W��g[�u�W��J �B���]w�z���e�m�I]�8�f����fKԔY�^S`u&J��"�7��ɮ�]E~�����I��^�\�:�7"2���[���E��%�xܜM�ǔ�2�?I5'��Y�����4�@J�d���r0�D���ȔRZ����-E?���ss!5uw��Gm��d���ٌ��6Gx+��(��]��1��~��b1W��SSv��47��.h��� �Ns��/9���>�<8Lc*��.���ԊC��he��b��� �60O��:��>p���R�04��a�Y
t�^{A+�@~�9����x������ꆪ��P+M��%�bІ I��>�?Wb���`P���c]ծ8ڌl���p9 ��鸑���U5���N��=#�����;o�#g��^/�ʑnZ��ߠ�S�~֥�IY�j795�EE�:�vʍ�����J���(�h���`-Y��?Ё�v5O�@է�Tp��FGg4�Wf����qӢN7�=ɝ��y'	~��#8�M4���C�N?��{K�2�v�{�"����e�"���Е��H����#DH����)���G�A�ѳ�:��Kwl����3XiKu�F���0���5s��&i�c��jU��We����l�M��V|�G��r�o�/0�^끑���d&x�u�	�aG�.L��L�f�b�uM䈅[�Li�<��ymxzG�z"�k�~�t��8�\%� �9��\�e����4�bD�����)������1<�R�F�34)m��8ι-j� 0��@�R����7C�r�p
�q����	:�T����r�W}�
:i�f���kF|?;��]��-�;k�:����ͮ<�\���9;�ٮ�"�I�>�� ���-��]��Mv�./s������f���E?
�ʥӃ˥f�d�L�]���23L��pr��_iEj���/b��	,�0g�At5"d��ɗ �猾�~L�Y�ӄ�+�~r߳C�nHfĄ}�h�� �n5�z^�����2o_�WK�Aׂ�'	���qçoq����@�}���+^��e��,� ��Xd�Y(�9�.�Aٿ���v�ڌ��_����0�Nw����2os9K�����,|�e��b����]a kv�tUލ��!i�7&���I#c���%.��.i:�H�D����z�5�lHV����y}��`Y@�N���!�viP��Ǥ1�t��eє�q� �ቘH���e��2�I������w��W��,'3���Q����v��nf+���o2�BȂ��������D�������F�������x��� ��9���\�m�`�� �i��;�L���:��Z�r�mHK���)gj�Y�αp�Q�Tb]�k�>��<���p��uҼ���4��B7?����A��2��a+g�V���*k�s2�'c�:XdS����x�u덺�XOG����w7��������y�8��T�<%�~�
#ܾL�l�l6��Z�j��Ga�al�KWa�@ŢD���?S����X��,!|���B��UA�F�Y��S��M�H@�a�gE�H�3K�؏_���6�X+MY��X�����ģT��5`������i���K��ƞ'Q�N���!����ҳN�I��f��K�ńs_��<�[�B�:�g�̂�vh}�������=:��jj����0��=F.��[�O|�/3��s�o�|��'M�#Ӳ�Z[�cm�y�"Gi�t�^��^��14��Y�?�I+���<��=ϗ&�L�jJC�Yϭ��鍹x�W1}=���Ǹ��2p,C�n��fP�C���m��ky`}y�
sI��F#�g1�UO�X��'��F����cP���tƳ�C\�徥u46-�9&�|�R�T
�oT�������~�������p��
a�o��3ZoJ�����O7(��ə<?�0t5-cc� r'�+$�X.��4�FtęV<��Sf��kCMn���w�XF5�U���ڈ��i�կ����Qt5պ`��l�7��R�q���,�B�������W�Ǿ�%������:LU�X��J���Qz�@�2Z�3j�)r����;P�YeH���cN������Jr%��6���e_T9	O�8��LWA�zF��]��x8k�#�Q<������_�n�*��3q �@(��/:?��:�JM��8ק��y��q�U�:�M�WcY1��
�O�c����:u�\��� wKA
x��.���r�Q�	��5+\ēA��l����-xf� m*������o�WR��L[��;�4}?΃�U��[{�Pb��⩅�����}���G��1D9Z���C'��v*X���ԟ y��m�K,�x����Ѷ�9F=:�/��t/�u�Twɮ:�@������[p��|3Ԓ��� �2��`�;���Y*�E��p<k�VYdR��d���˕1��d�Ec�N�I����6����w�G��ٯ
h�S��,Wqt5Ǹ;qMP�|)�������9��n���]r�����=�v���G.$�g\��Lf#�')j�oH�� ��=U|8f�C��<�ڻ���؊=��!����)���P}���V��-*������٤_�<Jq�[�o�bB6*�Ac� �QD��/�_V
������bD����-X�A�0h8H�¦�鰈�r-���U,Oo����`�ۍH9H	[H��.y�_o�t�ݾX�U ��2�����>�!%�VT)�$@x�k��hَb��&R��>�z�P��z{񤐱!m��ң20m��P�Y!X5���4׉�fv����8_��
%u��f���A���?���<i��}���%��dh��o�/�y�D��v��(�NH��$����%	vۡnt��!���s
�y�f��6����*_�<w����x0J~>��fo�J�f�(�L�<�0�#��v.p ��0Ɔ�P3Tˡc$���|w��,	U��[��D�y�A�N��v=7b�ӶS7�	w�~\B�C=�+�s-��4�ܴ$�|���?D�L�8������SF�u۪A� ����z�>�b-��q��V ȷ�9��F�0|+6�u�M�h{�$pE/[��#���*�#ks�r�i�.����//9z�p�n���y�;���+�[���5�,���<��Tc��T� �?���;�:z��G�bs�<�.�S�jn�w�hD��1�|EGs���ElOu坓�G�2B��S}pw��!�PƱ.��Y:�Bh5%�Eߥ��=M�{$�D�[/�mê(�������Rl� B���2w`Y
����V�l�Ⱥ�MQ���kb��3�R��󗺈T|8�w�����ۈbT���t*�K����bO��<x+q�p�R�=reSϩ��n��?OǕl��9s�n�L�U�	TVP4�kڤ���!?5��]�`�%��+�#Ƒ���G�T�b��ot!�呐��db�欧��z�".+�1m�|.�'fD�n��96�W��N�,�٧�oƳS}�w[���t��_�6��S�2�M���W��7����U��kI��� k���(@�
�tT/��'5)����3l*
���Kf@�w��ܮ�5��zY��䌫�~�Wk�,�����8re�}^  ��I������L��.R�Q�Iǥ�Z}����dV��#��!C��h�3���	&��H>1Y��[:!,���Ȍ$m_n�"�+��'	AeBs�l)�E{��+'�Y^q9?�f1��@ZD���P>o�k����
���WJ�'�|�1�W��i�m<��C7���N��KCvs=	���\��56,��NW��K͆Џ��.�*�x����f~{��]%Í�k�I ^��O���A=+���h�i�vU�����������؆`�V��L1u�o��N��7�Փ�a[���`	��g�p��cM�v�	��p�(Q��q��1�J;씑ܪ�C��G!|a��Aht"�IN���w~Y����Ox��É���>���`�<�\Kgp8�n��ߊ34g���B"=VE���D/�}K[�4�~^>����c�):��^0֛�k�og��;�|8}�-&�D<%[��u3�<�v�L&�F�&�Q*Yj���0�� %3~��[�<�ר�e[%Z)�	�\�{�lUE?k��<ZEKbj�hіّU?�T�^��i�f�JbW���������i$�kE<�h�WB=�_(<��AM�M7u෠e�8�����y�R�W��ID~]v�Ջ��z6��<u�O�3�r�z}�
��5[��UI��Flp�ɅQ)D�ߋ~��S���F>b�l�8�R
��b�%u��`�ݟ��pߊ٧�hg2�W������f+RXQ�ɻ�+y�C�]�bН�O`��-�oͽZ
b��C����=�DB[���|�܆/�)�R��R#ᣃe�Lk�3����`�+:\�6x��P��s�Te?�4KO�Ϲu��!4y���JX��+ ̓��^��[ߵ�1�]��A�ͪ��+�B������Ca?P.�>���`~�_���D������?bk�Z5��py�N� Φ��`��C7<�X1'J7Y�ª���Ï�TB��4`������9��#� ���ER@�7������$
Ɉp�gy��G	���������V�I�=o��.�]-}@�0���Kۯ�â���{�R�LB�"KI"���J�����N����E�&ϋ�'����)�(0�2�w� wR�,��~7��*�S��8�2�lqE޴Qun�DiIx�D�^��N�5P������D#�l���������'(���F#]���QXv�Gr@d�Fg4�:���M��]��41'��QR���Nܪ@��z�*��lQX�^�S?��F�M�AӬ2(/��Y|�1Q����
#�z��d݂�7=n��$�;�|� �|$����ߥ_�ᐼ��!�񬦱H������;������$f�G�k`���G�#B�,48�J���ᨗe� F����(1F2/v�ږ�{Ռ=q0a"si�,�Z����.�sx~�ߡ�v��a��1Ŧ�bPd�2=a#Tg������'G:�D�8��À�?�I?(:��$#���u慾0NW,>h��+�ލn�a�j��a*��FLM�.�*���7�!ĠٺG���楅ԏ�SW��I�?@�z�[�TH9]
�a9��w�+p*�
:��ȕ���&Rjd�6�\o�����G�O��ѻ��W:��%�{��6b���j7����,��!�l[�g���H�ʮ�A7ëski��L�l���|=�#Hz�Y�����+To�AƁ=[����2�x���~�,��h����-���+�����s�V��H��W�Y�%�Y�SD�\s��%�M]��
�X�g����ev;3������JtKJv����J�G��X��Bi���Y���T8�DMp(K^G�6��A87���b��o� %���A����&r��]�_�u�S#YĢE�!�N%�ޮ��n@�h�OV�$fG)(�p��0NMk�k��I`{�C����:����S�w�O��4��%�����G�D-b����6�=	]GA$TC���9�^R2�r�����I�ԑϡ��glh����)!\�z�kjt$%�\*G���e���R9�k'ͷ�E_����0���1fyZ�f� ��X\�Ҏ�o�@_�#:���';K!�i�)m�=ې���H��K:���]�lM�
1-�� �����ww���E�v�o2�l	�z����$�ZL8�2�u�I�7�(�˔OQr�-K�卅�N������q�W���bv�Ǜ4b7����!�l�7
6�ц�u�A�P��N4=z�m�7�mq,'j��ܪ~�LZU1h�o�t�6���@�c��x�3�v9?�U���TM��w$K*g���MYXu���*�IaC�2�d�巢M��������?���j��3ڴ���}����m3q�yq#�GM��nȘ�ЙL�|��]�H��î�Yb5�h*:��-]�:y#���8����5��@S���1� �l����Y����f@!#�J� ���k���h.���f�q�<Wt�c�ݙ�ߊ�σ�����o����3�Zn]$�W�ƻA���)�`�I|�iX�.�W�Cuf[�[7P�=��"�2]�}h�gOTN�B����V���UHV&~�I5�
=���b�F���t�Y�ov|��"��,w�
�A쁌 �P��L�E��*�.��QDvr^^�̸��65�N�P��a6N� �/_�+CS�XS�!9-3�x�?b����p�̅�Sd�:4{~̉Ġc��P��䵡�����C�N��Yy���OՖ��pr��qaU�ef�� �_/����|u�#��e���ڭ`N�Z�r*3��8<a~�H�Q�^?�l���+	�2��zm�I>�b�6K�z�䬷4s������sc���m#w��e�mE�4��k�1���S>�C�t���Q}��֞� �q�Z�ɒ+�7G�	:P)�|��#}|��0��"<OWއ$�[s�<��Ў�����0���]\B�-���1u��WΎ��w<�l�>,�d@+�){]����O&��q󌶟�*Q4bUdq�������6��r��mXa.���)8T5x�F����LrVgf��e�&˽l|�y5|��,~�3⡴�AB,Q�p�:Q!�0�U�Z���&�~����5k��6���[��N��c��i9�O�r�@�*�{���n�.Y�ޑf5.&�=��L�)y�&j15��װ �Ŕ*6+pPG�l#~v�H}�2���:-�ҷe �L70�a��b60���ņ)߅�����R�co�CNփŴ�����a�(d����W_ce��i�����^BԦ���5G������eGL��<A7TrG�d�u���hʒ������Z�tE�9�8)��6��{$��n�Հ�؊n�_9��0�Ψ}_S�25vr}..7>���c�\U^a�]�A{��[}��2�}0�}X\ӝ)�A2�N�E����D�kR�/��9�c/�UL�0"�g�^�m��j���9�鯪��Bl��(�E��`ؒ|�6���_�c����2�c��p�lB�783oችMj�r��� QC{��C�3�C��<��:���{P���%~�)�>��Y�1,��8��02��.�V�/a��qՄ�[�Q��}Z���������zAB�?6�����v�H1�o�����}��}�)$X5�L�R�H�-����� ��ޖ�$K ߭ZZ��"�t���z)"��`��k��3_1�do�ǐ����CVU�<6@W*i�.-*��/佲����^�hgPT�q���1��G����.��;S%�7�+J���w ���H��tH<�����O�L,7�8��k�E��4��M_�yh1��R��k��� LI	�Q}G�����ө�<jEpϧ�#�α�"K����<��t��vb�����\�}�C��$I���1�r�o���~)&.�4afw�4!�ɔ /`����=��>x�A����p�)s�����Z�%�g�E�_
(��[�.�bk�x�t񎨝�ɤ��YV���W�z/oE��	��J��;���w2&���U�m�)��VI�M���F���+��$Q�_L��ޅ$6�%�ۣ��@�Z�RO�8q�����.�`&Tp4J�L�ַE߉�)9�����s�y'͗�l�썎��'�1*�S��JTZ�.�|$�)w箳O��g8�2#�ZRE
��~�]w���
l��)�F~<T��]�;�z[�AI)[-n�c5F��\@���ٯI��9q���]׋�V�_t���e)�>6��&J���*�]���ߚԝ���\ON�9
��o��O����/�]�ah$z,�e�1Y&���X lk�	�A��󓻹�"*mDh��Y�D���!��2vƫ�[�
�x����������ѻ�4mA&��J��X�D`�8�^}�C+(G��G��N����Ht�����w7ʾ����v��E�A����� ��l'��`�8Ss�"'�^I�Q�p�yN��ޠ���Fh��0� �I�w��?���0{Ȇ�Q��BZ���Ȱ�::q��Z����Z@���kH���Y�~X����L��8gŕӒ��ˎ��<Q��ϵ>� �[�3!���%Z� ���o(���qg��Lwh�N�DN�!���'��? �'J��&�\����{�C�	cMw��A�l�r������-PwKSP��;RiU�p2�ґ�,��a��K�Y�˨o��t؍v��CE[�WX�с�C&��p�[��t�k}�lP�!���(�}%��W�?{�KG�M��[,���ն$����n�V${r�c]��4���u�	�D��B;;pJ7a2Ay��[�A����F2	V�h;�fZ�>�I�R(���X-`�B�{���1��|뙹����d�m��n(y�=��=��iڌg�6&�$U��/��ʒ�՗��m�E?EN��*���||u6�|y���\;�v��47AR"+A��RkCwB��[6|���Q�ܸ$X�G������E�{��D�o���E��X��0q�# o�;�ޅc�֖Y��)�6��T�?��0��)I�s2��H��T-�R �٬��=nD"�Ҥ�	г����ֹu�ǉ/��6��ف��Apn��r:$��+Ysٞ��^����x�����1,���GEn˻o��:(�q���U&��+�!_���oi&�\�׸S�DI�/G�z��o�E<a�N5��e�x�;�I��J��-?,˪e1w ����#y�h��p��g��\�����=���~�"�DO�f\�3�Sl+/Z���𵺂@�jI*�1�J���T�n�j^��[��Y~��x �=�蕺�8�S�?��H���ýwI�!�%�����塞f;��!��Q��C�K��V��S�U9��<��g�4l��!ֆ��8�#v�L>�,��V���҂�)�[��ov��݀zq�5:1�7ZO'�tD���?�P���%<��c4d�}��#BXa���vk"$j��8bF�SJ��C�O��j�̸���ee�X��ES� ؠ`6�w|d|ռ�b��W���l��N���d�o�.�6e1���\l[<���e}��6�I%J�@xk���u�S��X���g��JS�Hy�_]p<Y{��\�����0�L���������-yO�9�|��V���@��0��U�}���mv�Z�!ʨ�Xh�*G�eqe����d$�\`��=�)I</�]�k&��S���ݍ��%��eBfQ�nu9OMy;��J����5�2e���Y����2ލ��G^&7w9?� �ւg�3��]A꒚hO�0?�D���{lT���A6�f����ud�8J�1������r�A�qF����|]E��y�|�QR+�ia�+������_��¤~݂��م��<�E�MvdP�8��}�d�;b&7��*q�~���	XI�S=$E'��Y�F��vuE��;��؎'l�>��KS����XqQ���z�ȷ�`E����kS�q!4�#M!��Q=V�2�\����OF�L鴺�d�����2�OYם�p\}pHq�(�%}Bi�&`���>h�Y^Ŭ�c/7x��4�P�s�!V	ey���ߟSN���>���H���'�5�����|�P=�9��Tk���:�;3a_c��d���ΐF
3��6�.D�Z�!���>��C�f.��l4Qs�Έ1$�b^�� Q���q4���y�`�0;=���rUx�7�%
VJC�H��|�O.+��C��D���vh�&�c���i�<E����[wkS��U��.X�ܼ�l�-⶯#����w�{0N��C���ˀ;�gG�7���	��T��M]��),�Ty6�q~���0�����D��[�V�7�Sz�.U����T�����2�v���W+�KZ4!ܶZq�ȼΒ�@���_
�+r{��i�gBJ�(���E��$J�^oea��7�4t���q[{�)�Nx����.H�������L���Ƣ�!�]v\��	1<4*_ �X���{�Dڦ
 ��ي����@
�X��iqW��z�h�gU!�>���b��L�"Wt݇k��-#;��RgT�bW�F@A<)��**]4�6b(�A��VvEeYkY��دe��Z��� ��yX���$�q
��O!,���ж,;*k
)�U���|g�����P�hL=�=�l�ٔ�
�&9f�Y���u�7k^��t~u��5�����|��i�����', �ٚ_j��pP�����Ɏ��On��e�ۑ_6[3I��8��3+�^֩�Թ��_[/4Z��1GqZ0��V�"]��;z�����.��U3��5���1ͽV��^���s:���1b����ȠN��@ qg�|vl��%��{�����J���.�ۜ�Ɠl��ߙ�b�OY���ә�O�;ܻ����vfH�Y��7e��}yz��d�@=$/��\��E��0�GP��"۰@�K��ws���Z��%�2������SM�qJ����A�)9�~�*H�-�����j1$Z&]�R(O���>_%Q�Ű�1c#�"�Ҝ��]v��uϙ�Ə+%Wgx�T�����N�U���/�d\��]gTV���&�ZkT�����7�x�f����jJ�T�"�l1T�4��-Y�ZT�"V��I���
2��ϝ炝
*�h��`\� |U,Q�a��:�-�Sv2�3Wwt������>�fP�C�垺/�#:Zn����0�t�W�Cɢ��Й@;W�?K�N"G4�J�l#	u$�[ʟ�� h�,����]��E��f�O�s)�����b�f��td����x>
��M54��A)��P���m	���R���a=���y�t�����$ T/M��ߜ8�|{�$)穉C!�����,���Լk�B-Ff�.�*9���Z�PK�9����ķt�����HQ�'d�� z�V��Ig�Y	�Q�����pPK�x��La�zP�/m咥(~���xf��"v[�d��G���P e�@?Y���t�Jĕ�H�[��)��|}�v��0��0�7n�'ý.�.3�ha�RUΘ5��_�¯�_�O�w$k�	�}Y(���I�Z�ɣ	���}���zU��L�*�/K�� *�gcg߹���e�pȨ����<��*C�:�u%�rJPLڧW3qG��/�uJC!��{�526�ʄ��Wv2�5y2d�4(*ˣ���}~��!�̪{��ʯ�_G���8n@�{�|���:W�m>DqX�3�]�M�(�w��/,׎��ܱ�iW ��A�)ѯ��%8�<=�CV�L]\�W�d�{������kI
��y?�d�`F%��f�_0�����p�8ÿ�j]E~<9	g���� �J9sy��L@rЊ�b�	١K���<�U��̝�Qcjl����/�s��D��C(�nA���hz�qĆ���6g�~!�oo����`m+'��
ٍ��q�K�%Q��`}���7m;�����6��P]�@@��!۵P{�2I�S,0<��"�����b�
�������k?�T?zwS%��D�Pшh���9H�:��C����D�����C�Y+
�C��r+�:�k�%��f~kz�F�C\Q��z"�h�8{���݌��''ю�PU�K��ǑH��B�vqO@"�n�j�/t|`���8$H��wr[�.�Dw!��r�ߖ�cM�
E�{��,?�[<�|�y��b���I�jZ��K��e����+ޓk�#&w�a�/k"���/���JB���O 0s~ݛo�K�Z�n�(�h�TI��g��S���U��F*�I�}�t��Hk����2تB�����/x�Ε�W���� $���7��~[႕.��m�(8��O��ÃA�,u���sԞ�	g��Z����J ���(���7��:Yd�8=�xz ��g>D�$
��7R7���v�.��H[�&dp��	�xr	���<�;҄��Tp�=��V���:���r��Y!fK�E�G�I���V�h�}�M�Y��H�_�Q|��k�B����bb}�=��Hֹ�}���3����{����B8��59�>f	�o�+�ӲW��D���C"�>�r���N�+�QD���USa0�>��_0r���U7�n�|oe���z�?L��K�'���OɌ%��Τ#�.���+|���e�a(�" ���P�u��_&�̟�A������%��A��L�u�׳�b9��Og�;�0���+�H!�����*iD��QfZ۾35�q^�m)��:��4\q߲jǔzlT��'�B�(ΐ��\���_�]���۱����M��K��sy��9��pa䉾"vt��:�U5��"^��W���,g��-h�p�nJ�z�¤�&�`^������&8�M��Ǜ����I5�:[�^��8�������x������I��C=����}�k愐�>KaAc��&��?mպs��ߎ���tV��1A�75����5�*d<Z)H1Wu�E�R&�N��f[��;f{8̻|�I���?r_A\���k0�T?������*�30�o�X��i�H馨�]��+Ѓ�A�����H�������r�WA�oo�����5��
�9�^0,~_n�9��� �������9�"��ݛ��s�غ0B��kR���lɒ��z*�$52����jr�2����M�	�<	g��6ıCs?�߱���;�&^�9i��Ase��q�����U&{J�&��\�"&�����E�?���c�j��Qf�8���(}Wq�Z{�K��`�/H�3� ��RT�WN �����dsШ����ْ��c�]���(�!
NTN"�Sa�mm�;���v��ȹ@7�lm@�t�Oe.��~�5�b��eT��g0��T������>���h>�������0��_aZ\�<`�[j�I=p� t�=���Ҿ��=
��O�R��/�jo�Ey���n�r띪��xj� 7/O�q�0I��<)%(�C6T��}E�*��)���������*��(�h�U��q�Y4�[u�t���\9f�i�d��^���4bM�?����h7�H�J
��}?-�� ��
���@Rj��7VB%��W�7e"2H��y14��|�@���p
 ��xzqV���f��.�E�y����rP�d����[�~��$ߤ!�6��AA�"rt8V���S"\nU�`��?�1��Ts0^D4kE*��L[@�Ӥ��#��_U�2����� {���8��w+"X	�_���MD�M�a�P���>�l~���$u�{��fo�ouv��c�������&�(@cm2M*����E4�՞\k���ob*���.L�[�A<��J�����H�"����R��N<n���9g.���Wg�dS�g�I\����0إ�}���8�<�]�l�	|�xWh���VeǔB��v@�����ٯ�Y3������y�
o��j��p�$*|q~�1����׀ŸZ�M?(;�k�wu��Y����>[zg xR�k'�h���-��A���׬g��9&�d�՝�@�x��q�\��.��ڸ߷r\|����ʔ+e�J��I�׭:IK�ar��w�PF0.A�KɅ
���ۦ*ceN���ءvUTw�N;C[������9;�A\�늮/ԕ �ά�;m�bn�9��s���6����^�'�Hi�7�ISݲ!�~<w����"�63jY3�)fTui� �>�n3}��#|\����'ux�b�E�ت�j+Կ�6%M�٤|��be4n�
�H#�����*������:MH �:ؚ<�TR���L�_%���`�K^A+.rCfe?����%��7.G�y�2w-ӡ&gn�ɋ���ݖ��XA�Ŕ�e���f�?�p����]���C���MB��UqT�^�ĴT�a0˓D�������Y6�d��2��ߞ:��O�Kߐw�9��Y���{k��7�C"[`�h�L�cM�d���w.h'd�����[��D�8�(8��C'�'��[���(lQ�r ���+����=����,�0��ih᷃����D��sې'�'ES�)Zd�����f닓`7�;����QЦB���)~ѕ��!���$����(5[jt�h��%xe-����Z���b>o�#�l'��Pb�B}����u����S��,�9FAJ�8N��;e)�S!	�t��[!t5�9���5�(?Z2�| b0��р���!q�qs�p H&I��{4ܾ����������X��
�zѯ�s�H��⢺�'"�����|��Dٚ�a��Li04*�q�`l����K�=��Z�j�Q�5��
������q�u���B��	���J/�;�LEI��R�� �_;V�y�EP��X�O).�O�%�A�,2������ƴo�!��	�"�^HVi�"�H��Xi��K$8+�8�M��k~#�mJ�����?��n:��z�_g����S��m�p��H��s�]�8�zk�Pe��䦈 �d4 �h���]<J��}:Im/���\x}�)�6�Cw	�Z�`M�\�g��.C�9�a�(Y�}��&9t�̈́ò@N�4V�X@5�vFuJ�I�*��@0t��cf�5k�h�<:��(]K��o
� k�K��Y�K���d��x/+�K�r$�F�� R�ѫb��f���s�lΊȗ��T�:�k���*�k�;�獗m��:�Y3��,��5p��,���tL3�l�:�t�;�n!N�[Y��D�ej&:��.�6�ɷ�X�I����n��+�Ȅ��M�c���Q��b�#�8��F� ����[y��kf����t�f�w �C�'
�U�[� ��KF���_ ��e����T+��ʧ�g&j�������%	NQ	�
	��xUh���)}J�.1�+����^[��l������?=Z'�.�Vu������/��i8��ǟ��p�n��6�Abam� j-��i�s�c�\��k�BbA[/4A�SР��j���d.`����"�O<?��"u�FZ!�u�����+RkV��UIk�E{��� =�So�%� �ݦj��ϩ��<ز���2F^���`���%h��o: 1f��3��L�qIM��������΍Y�	@TO��pG�;�
�s�ՀlK�?�6f2n��s:���z�)web~�������6�K\oD��z��w*�z_CJ�<���8Ok�V��V��u���h
���~F�Ri\�u��E�ř-�����@�9=�+F�)�ԡK���_�Um��1=���e<����͘�&�І�fSJ
{������Ҫv�*P�rs���I,Ǭ��)��ޫi8��jc��߉���,�Hx/���	<�p���g&��F=���&��0��]X�����ϪQԍ��<�]�	Q4I?F=(ɧ��X�O9=�3"��eG��Kb�;S]�Z<_�#X9�mh;�{���ڍZ��HXw�X@�tG�c'L�����E����5�y��~h��Y2
�45#V�u�P����<m�m�N�U �YH���/\���#|x�LMy3���#�FѬ�l@F�� ����
���
u*of�}�}U��%q⯹�9����@M�#6��B�o�Ӥ�����p.W
-񚹍2WE	~Ǿ�f�z.��h5ɞ�������KJ*F��R���s��7P�*�Āp����c����T��j8b��/%~a����HqJ�\�|1}hF,�Ҫ��w�&�˒����< nLe��ǘ���B�WG�Q��,��=�����g��K������x�.'e�-fP@�iT�/���� ���7B5�����y��wAD�L�!]B�sr�J4���J À ΢r���-@6/�f=��"��7�M����F��]�դ=)������=��ФĂ'{p� ^��?�Q�� S"������,,g�1�Hf���5=���7[2�ђ�S�ڣ�^�al��b��_G�TӰF��
��*$A�S}'8״�������$	a����y���)F�M
��uc)׊Ʈ��g�8'ŧ ��Ȏ٢W1p��[����,�.%��:�Py��vͩ�%�(��љ1���N�J��&޴�*Oб~H�!q���Y]�A�>�\�&_����r#M��m^;b��<,w����٧΋��D���
�������`����,�jn�:�HN>:�ζ!�U���Q�����<z"Q�� 2����w��:�N���`��N*����������1�)�� ��`R4x�"�Mq���G,`miߊ�H����	nQۗ1������&jD��}O�?�p9u}T>o������a�W�_��7;�R�J(x#�L��*�� �IR�j�L�J*@���S��<�W�����)�;�Lω�'�<r~ˏ��MWt�O4��)�;79*�V����ń%�����'(�>����x|���" <�׶�-0B��x��L�Mbn}HzI.��p1�������6~='����DhX�Sѷ"HH���p:wV.!z����2�cǭ���re�!ƑᘚG�O�H��Y/�Û�AKST�ơ�[�19��㿪���zL��M@�p�m�G�jA��Y��	��]���Б����.��SJ�j�=��*R�of�$p��q@�d��"�ӭH:��<�}�k��aX���N~e>6�~����v���4�PT���,-�X�r'�B��$d<�W���h�X2 �s��!�|:۬��`��+̔���iQ�X��e:���R*�Ɔ�����ϫ�! ���&�2s/���JU���t�pFIm0l�m³Ӝf@��
��-ߝ��n�o��c�ժ��n�Ӈ�o{�r~.���ݳE�$�g �,�x� {�G�U�-�ᒷ�R���MGx����������R�B�K������4����#�!�n+H��<IGQcAX�o��6�	�@�Q��l
�!�C)��k�ʒ[���Dc;��o� �MW��@���$ugEy��َ���?� ����&u��#;�y/N��N/���A��ޕh`"�L�b:T�����O��)ԋW��4��9��N���t@�pY��v0�*��@	ks5�%�>����i6�Pc푵Iz��m��R�5@P�[s�ۤLџP��D��������,V?0�_�$@��0;�澆��IO�2�8�f���;�n�b��]%Y�T�i1��^�k�,"h���`컩�w��L�����?|�ӥ��Q�Z�ۘl��)a�� �(�,��K�{��l�\�!ÇA��:����]O>�0��87d�U+__XnT��;C�*#�����>�W���6m�?�l�{JtT=Q�ʅ�[2L�ְS���x�H]���s�-❟)��Tt�b#��P�Sk�/�\n��9�N8��+d�?2�s�"n����Z���¾������E��Y>I�d\��_�v�ő�{)�)�.����P�#�x�/�5��,ij�ɯ-)�����v3w�1�M�i�� ����h����f��"���o���/<g������fb�[�!؀��ʶ��*�i��d�+��`K}��� ԃ��aqf�MY��"�]�Z��\�骭Ҋ]�r���x��B�����(��D��	�.���"үaD�E݈��t��IԖy%��N��o�C����ӡj�1�wf��SCQ�Qly��f���zr�7{cC�*�r��D�Lx�ʗ�Pu�?�[(n|`+&r�2d�����Ĉ-�n�����?k������me�s�X���Բ������,�8�o�ک
#���GoV(��*BFsLN��{>M���v_�E����.��K�@U1�e�C�&.UQ��β)-�~�ɾ��Jn�p�����flXp��4������ӌ� ��m�`�n��)��*���X���U�I��m������Q�i�r{՞�]Pp#9�(�w�*��g{����`�5\v�Z^�)��+@�:3eֈ����G����+OlBg�p����jPb2 ����Ha��2���9��П�J )�����C;"1QFY�����G�~��'���N�_�?i�Yza��1�P��H��']���@��u�%e�ˋn[� �ޖ�1݃�y9�]n��8%�ꈭt�gb6�7^��+
 ќ����V�3^J&���bV]�b�n�����Nz��c9�ji���v�f'����K�>m�]�g7�T�:�/	�"��aG�e��pD�h�!�8�!<~(�x�u!�*�W�=���cm��| ��0��ژ�7lQ�����stZ#�o�"R���y���.�ܡ�� �J*I�3��ᰳyk��R�Db�{dU�K����#D$�Q`�mK4$DG����9&Pc���}��`�P����D�������Ҩ:�X���u-<����R��
C�f�>(���k���?�i��Ø�Xշ�j��2�'m���8��(UH�=�Vm���pfܐ$����E7<������,L��J��t`g�9�|������`lZ�/^���->M`�X��Td��l��B�R��Q�l�#�� �$��^Ӳ�,n���X�岦g�:L{M$>��A����� [���@�<3�W�Z^�~R�|Ό�L�}۔,s�t���H��Q5��z�^���m@y�o��<V�!����d�	�*:jz�_n7>���8�q�L�y+{6"��Z�ϑOI���G�DPV�Hi�j���<�?k#��yov�W����&�Й(F��L��B2$�r­����j��B��i����{�諛�ßǑK��ҡq���V7�&�ι���ɾ�y�?�Ž��d4.b"��`�:E�޾�ed�5�M�0Reۅ�X��u��s�/?����GyV�jrDl�t1��s�:��������<Y�)e�W�Z$�NL�oj�0g#��%�V�4u��6e)6%z�	c�A!Rg�w��qJ11O)�����?ɇ�)�V�or��e��&'�(�=�_vc�W�8v[�7�C��E�����
�[�Su�Х��!I<��"� K�����ɱJ[�z�@R*(�7BYh¶������0a#�o�Oc��,hQT�����Z�ӓq�����9c�k�	���Ψv�/mwߺ���(�چ�q�ս����V��U�&ȁ=�V�:v��Pjl	SG�jD(�����v|7n�t?FN��ǔD~�,3KM�eHZhv�??&<H@�ʨ+��p�����?����H��?�H�I(��
/��J���<�N\>�40�WQ�E�#;+>UV����"�ų��}�Qu�\`�>���
�K�"c<�:�t�q�
-�a�3Av͚����>�oz/�ʹ�Nw2V�l���:����3i1�[�W2$�i ��_�����b)�U�K�J/�VT�)�p��qk��1���'��6����z�P�ȯ>R3E�*k5���e�>.\�!'�:mjD�}G��i@<��s�0�yWҿp���P�<��H�*�	�Ҹ�1n�3�G�|s�-/��[p���k�ӹ��Y\��t����x�{/�܆��Rd]RI?�[�0�R�a�Y�AW*k��8�jK��d,�A��+��3{(��@n���N�_�� =r|Y
 Lc �QB�?��Q� R���Y��*J�����_�L{j�l�J�4���̣@K{#adܑ3Q�Yo�Fm�o���#TD/'±�������#�P��T��*�v���	��鞂,]i����n,�P4�39��|�=���-7Cy�$VB10m-�i��j��v.�L�%�yW�̕iVTUR�(]�R`"ޑN9�L��fU���C�=I�<#�n�t����.(���>���RgQ�;eȈ�lx�7�(L5�����S%�W���Qk�.�a(&��Ԋ�s٩�Z�	u�c�TϺ����{|R�д���i���,����lesg���I�*�.�����i��EH�tg���T��|��jD��k�N���h�n$����@^W
�o�&����'z-�cT�k���p������w���m5�U�df���A8VF�I#�?J�����<,k?�6��������ő?a͛s��d>&���� �A��J'�K���o�іƭJ!e%3 �T���'Ah��3k�6$gL�1��Y9d�~����0�����Cf�kLß�D �t�2H�H)�BA�, �F�*��#K·�ko` Қ�;��^Y)d�_�2��$�s~�cj��
i�e�kE��ۿB�P��E&��Vx�թ9��&�h��s�����uLO��v������#��!�]�H�fy&���Mk9����覄��E+PQ� ��yi ��U���ܬ��SQ�q�QΤ���;|h�#���+_ר�^�z{5��M�]�<"P���R�N��p,��r|)ߪ���6�i��W�35�t�r�Nҭ	F�Q�|�299% ��֧��!§{O2�<;���<�����M�� v�Ɋ6l�eս*���p�����.Ǵ�kL�]�g?�D�����/�j=Ώ�c�O�'z�%�|O�o�i��$�er���7v��:��+D�,7O�����R���NL� <�����R&v�F���Mq&���l-�o9%6��Ŀ�%��
�ѱ`)n�E7��ST{���I��3�Եj7��S���W7J�w{L|�,m��X�w���o �Ԇ��=�.��٠���!�X&?���\gk�R��{�!T�g���f$����0o=1��3˲�ux�\�|�<�w�cC�A\��pk7��������2��N\{����f¡%7�5�7��?�6��
�ENӂā{�������M$koAb�ن�A	�D��B�T�������T�3l5]:Xk*z��E73�E�yck�5���g �����U�ǅ����2r�^�l��,ywve���2�O��� �s^h���5P�t�����K�В6������c�5�5z��K�b�X��2���H8S�с�7�է�8���{�e�&��&I����y��- ԯw�{�-��]�0�N�Y�5_R�!r�]}�1 ݅��Z�R��9E�/�g�^f%���� ��7�s����'�h %�����h����,�/�D�.��>J���X׳
��X�w�a�~040�6g-��}W܀�,h�'�wK&�/X��cAk̻� �	>��z��X��b��F*{	rC��k/R"�"��_9�j��ד_�?���``���x�_�kS�C&�����'e]־��Q?^-���N�E�Vi���8���O�!~��# n��r���6a�5��Z��#.�:����}�k�X*s�LcM�b�l�I����0{�9p*mmz�o��0A�	(QY���4I�9�� �ŵʩ�ij�.�|������Y������7�>qbd�?����&�����P�s�Q[91ܒ�?���r�;�i����ږ�����FKW�^�4����Bů_�N���Z)����V˽b��ٮ-8Q��q>4c ��G�n��h����4�5����1��a�s�i��-��f�>��#A��l�s�5���.ٲ.;Q9����1G�1�N�i��剀�<f���H(�	o�M����O�F�9�4������	�+���@��~�Zw}Y�Xg����;̏���g�h�q+z��H]g�9oZ�G?ì�=��'�FFx�*>�8�3�T�un���;����H�w��m��5����%'f��pɧ��8I�ŧe���/�n��Ԍ�T�I�����ةA�1��Jc�g7.ú�e�>�U��T��S�ab���#J�'�XmL��{�d�M?;4�;}�lQ�u?(-a9
M.��B�����8����6���>(�,�*|�0+��t��V�=��9W�T1+���t	[��h�0C����/go����3���k� ����V��"�k����!�;Uw�*"բ>�{_� n����K�ӛ]�kaZ�u�y�a����A���H��C	HO�Ny��Q���S���ԡ�bP�G�[�dx*d]�+ͥعhC���B��\ �/H �T�3���yꊔ:�&��Ow�#0�f�w[�W����
��5��=EyT#L��WL�`M}N�V�-�4P �9S��5n�;;ď�?�%?�0x�� h>�=��UpЕ�����ގ�S4M�*w�6 �����<a,���S3��&/4��T�I��,B�Z��	�q���3t'R	m��XsO{6��@�~�~%�?l�e����y���}�\�Fw����C�A�}�=������dl��7;WC�M ���O��u+�m��go�+W�}g�&��h��~��oDo��B��2���>����$�u���ִ�>��xݷ�/�)p��8p	!eG�Ĭ��[�&7$�N�Q�u�����Û�=?z��A:dNx$��eY�{�@
�0���p��yڴ<��ڕCw���q��A#p����N�yi��s�oPB��	S�K�:a����Q��j��26�6Ud�7��s��i�1c���Gà �p퀦]��5�{��΀�K�1V��ȣ��U4���#R��fTk0<�Ǔ�Vj�[5�;T��gگ�
����m�QrZ��Jq�3��p�Z�t�\�b���Q:;zx\Ȇbݚ��iD��u6��Sx�������g�e	m:�I6�;c7ʻܸn���s$�By[��7��Y�N��`�#�v¬��-���w?�� �Բ.ć;���lw#C�4��B�:d�}{Cҫ/�'�G��&ݗ��w�j�&��"�.���]��h���%u��w/�W��0�u^":"6�B����ȴ�Բ��)���T�LiAii��=_�-s?w�\a2�þQ����e�)��M_ �Zzs�Z�B�-�W�vc���WJ�p�&�+R+^���+R!�ͳ&!�<�7ۑ�V&�g���:i�A�K��G�����}���V]}�"2l�"Q$X5��[-����ikZҠ�=�w6��Is���P)c�j�l.�񥣰�k@P�w�O>ᾴ�-v+P�u5Ux.�D-�78<�9O���>������u���YV�t�FM�>��;�\�5�9�r���0��4�}�Z�5�Ad���O."�,R�t�� ��)�"8��u��c9�3��&pd6P�q�ߞ����N���o���;o` �F���
�ނ��bCElI:I5���b���5��*Λ���M(㝝;�Z��݀
�W�4O?7`L����M5��᛹�;���v�^��w�4�e����T9���՝�hQc�/�g�C���B��3��1��8�}3H���m!��R�#�p6�K���E_<�.�%�c�ZJ$�ck�({�#���Y�nt�u�Vl9.��&9�s/�k���;͈��1ă�:��Z/a��N�r���A�Bs���l��db��&�P ���%o����$8p��>��#=X�|W��+�=�oj Y�n�E4�!�'1=X�S�阑DO���Gk��w8��T~*l�U�ةp���\��mU)�n�%yQ ��	�����H��6��/"{���Gm�:�5v�L���,�S�W�b�o"��;!���=#>��\�giI&�>�̀��Is-�9$�1r���کC��աi���Y�yvhD���o���|��I�a8sV �K��jD���xM���ڨݧ���X �X�G�mm�i���_�q��6���Mkn�;n�����w\6HE:+3�}� ��x��g�R����╵��o��FM(~5ٽ��O܏o�� P��pڭF��N���
��X�_]���DԼgmjy�'#	�c��{ثA,thsҝ-���:��"�d)��A4vk�o⇹�ԺO8h���*���0_�rJ�� ^ki�z��LnEw�7�1|�o5e��c�ڍ��x�zH�ƑܭcD����d/WR�_�yBs��p(�
����.z���ylx��΀�vC��������'o��x����3��!4Min�_Bs���{x����C�+�hΓ��.���\?u�);�]�Y�� �j�� \�#CVǌ��P�F]bD%F�f�����0$��eKL��1�,�U���|�xH`ܻΌ��|-~�%��?W�(��k��*��>�<�e��W��.f����g�rN�V�Y.� ��m�`וq���ô�x�����cV �P#7�i�-K�7�  ��e����3�$��]�[a��	��r�L3��άf�E�5�=x���̨2�-�5��@��Y���,����r37�r���_�@�{��p��W�Q�J��?%���E(��k�M�d���- �>@!���#?}G��6PS�V��@��׿��@�I}�0p
�r��hJ���,11���֤o�D)�ȹ{8����$�X���Xq����I�}A1!bi����~��OS֬�x_�������RѢy���#j�Y&�e�qʂA�t�&����)����E(@.t�1�5�/��"Z���w��p���
���B�>���"f��)�
NM���U�O����"���nS��1}�8��|Ztb�v^�u �ϋ��r�٥�-�Q�Dn�&�| 2���Ȣ���=G�H��I����O ^��ͣ>���C�oP&���lv�|3� �.ɛˬ%����O��pWF�g}T<��� ��]�`�(��o�l�,�9��mV48�q��
����P	渞BlEw}���!��H߅	�>�BH�*���2zpZ�՟m��8��qC��CmwN�	��m���D�
.�?���5��	ÁE��Wi�$�s(�-Z�È_��s����Dz7)Λ'x�$nUHF�����,�뻇�֢]�����w)�GLg��@�����V���'0�b"ߘ7��P��N�s�E�u�lFʹl7Է漌���P�T��t���]n�5����f �L��<�/ƦD��%�׏3��Z��'�/�q���#�Ĩ�ֻHA��#Ka(�ͱ��g�?-�C�sv,@��11����A����^��9�Q��RF/�Y�ó��f�?N�-k
r��z4HCBNy(I />$��qMҰB7�GY��m&�(�׺�v.��*�yf��d��w����i�`]y��G��U�ZPjv��@ĺ�^��Z5������J�_�ȹot���S���K�,�i�,�r���+��P�k�?��*�@PF	^�S�V�_�<�	51��.`/����84�+l�P@� �JR1�� ���l̓�p8��a��I�*Z��]����o���J/M���X0Zu�������.�[���xB(=2�*,63����Lv�Vȳ\� H�Am��q�����~�5S������3��ȚU��ĿDjkK��F��wTOfx��+lf�/;�_.�OąO�kXg��3 ����_���$����C�\�+���O)��	�9}K%j�����|tK��C�T�%��z�"�n�l<e�@��HT�:���/�+J���Ŕ��k�"��qZ�ۏ6�j�����zW,8֞����t�_2��}���0q���:�	Um��X�@׋�/P	f�<��L��f�)[��ө��$2�����ަ����̂���^ׯ�r<'�F,����"�<��d랒�x�J�򧢳,F%�B2��� ��9]�8��J�2����~��pz�4(� �?���+[��#�W�a�*�2ڞ�i���
EH4���'���I����w�Q��V������.�I�S�b��#�Cl�k������Y7>Uw=�<�t9��??� Ӷ޶|Z��av$-LS�`4�%"aa9T�z�h��h��Oh���b?nL)v�F�"M�L�:%�z��m��<�[ }eV���]ԡѪ��bP�c~��|��֏8ݼb~A�DطPR���Zt���Tk��F�lѤnf\/B��t,=���a��q��q��?�]��ᰇFW�$�8ǔx�}���͈d_ér��>�x�\���٥�4~慾�4Jt���<���;Gsc٫G�?�zյ� ���\�UL5����Iwж��9R6]���>�ȏ���X��W�,��%3�LVB��H2!��Q�&�sUNH�J	gFz�\}�]�1���q��0�i�9�a
�]�R�dWr֕�f��1:_�p������l����m�%�O���Ec��CG! mq�H�3�yA
R�pbq+�c	�2!��I�F�uB�p���U4�u�4��-�QƤ�aZ�O��0��<��植N�qn�� ??B�!�~Q�7��Pw�F��F��5�6/�Mq-�`x�pǺ�ҧ0�U�̤�O�)I�H(Z4~�!�Kw^{�o��0{	�#�1�g�=�)P=?/P�*����	�_�-aʵf�(׷�˦��C.��KBӣ�;Q��p�d�(l-r�q	T�`�XN�%pn�P�2P˰�MQ�d��A7����Mi����]��:��w�k����Is��	ȴ*��}K����� ���#��T�\H85W�dA5�G�Ճڍ*I'<�ν�6��x��i}�Ҡ�����$�a͜2����q�O�J��POF,j����hf�HLL/t���_��R�$C��Aw�gi�������h��SFi&��XWN����(��%z�}��e��7��v�c�)�O�� [��;"'�ZK��+�ǘ0�m�a�����l����0۶w(�!�Q]����o�"���l<p��g�7��qƇ���7�fvZ/�l(�ݕ>��b��{Q6����ؿ�2���9r�X(b:##^D��g�����`y�����V�{���L>B��U�%��	yE�V��G�Xx ��0���T�����΄�tgJ����{N����A&:>��;y���WF��3���T�9�q�a��ė����/˶���&�.�݄�A�Z}p��e׉��"2��A�f�(��[%��W�h~<�qvρ�����z�=�c���~zy��~)�Y��w;���ؕEp0��"A�).�wZ�l�z�s$�6���n��^���Ē����՜"� o`'��M^z�%�Ӏ���AIso\���.Y�4as.�9��X������:Z������ϐ��'����7p4�[rZ�c	�d5'V��̮V`c� <���}�T'H$������s���Y��/�

�J �ㆽZ����U�Q��l�݃UR�+KTz�v��q���Q��:e���}T%��`��_L�"� 7ү6�'�Ȭ7���Plx�ނ4{�����a�w�����fNr��nkz�Ϳ�oJ_�kX�7�@������$�*�����5� 5����J��̻�j�h+��neW	��K���R�9<fK܂�uHK��i���@�mE�Ý�X}&��Y��֝�F~���R�׀�]���� �[-��X%_J��Ƹw鴅�Z�kN�kNҿ
��θ?%[�؍��f���hRsΫq������M(~��<+Ђj(�&����`e>�.��4��y�L��Zf)���$?�C�N	Un��w�;�}�L2(���N�]�N����g+O��>r������� ;&�]^��wݴ���"��3��A��3��!t�� �J�_���9��s-{�Sr
E���qȾ��߳Ĕۂ�3R����=W@i�!�0V{!.��TS�#��/��vԵ�/����@E�dnT��%�!�t)[Peh����H�[���b%w��;i"�Ɋ�����/N��?me��t���2ɝJ�
6���9��wo��eM�̩j=�ȥ�x��'�+Ph���a��,Tr[��}!�q�#r���j���S+s4;̼,�ʻ��.�+�穴̕칤25�~��k�=t@�Ȼ6R/lX7�z2(�1I����_n�bu�3���[zΜ���j�~�<)�ٵ�j���P�W�2��#�!%�E G��F3��W���>��W�?߂�L�x�{9������')��w<�s���|!!��Y Vƶ����G�J��h�pu�la��h�f��JJ7)����t�_�3e�޷���Ϳ���>aȹQ��x ,Jg�^�a�v�ɍ5�����eZ��I+��rR���:[t�L�NN1�
�4��H���s����8�g�&��2۫�ͰP	��g|1%���2�,���>Y+�Y��т��;�́�A�zu?<�-T�){�:��P K�BE�����DP�;��4LYms�f��%.�11KK���}h�3�����*�U�0��0#e�c(�<��t]��åi�\�H��H?�@�㖣L?AI�y�'�x�Fd��64>i͹0���"��K�g&�B�f�Ѯ�*�ȟȯ�Ο`l���k����A�'J
x��R�9�Q�pDr���p������?�Pڄ#m��@�c&F��e�n�׵�c�}�V˵�rX3��\C����Y���c�o���N`؞N�`���&oA+��>�h��g~8�1�ρ����Cj�]�"��4��B��2B.T^_���1��[�S��5�G#�����$�z��]_�'O�N�����h��\��_��-�]{�_R��d`x�����t)_���$D��h�������1 �g/�V��L��n<��8�,��IכZn)=�m����xX�sӐ����yd�5gPk5�r���{2��|f*´���y��g��[z%�����W�,FqD������!�<����W�V��أK9�D�i���fY��"�M�@����B��	�r{L<���mO⿢J�&\څ�^��c��ʉ�Fܦ�3���6��"�C��e�q�0I'��[z8�[c+�ƉE^�=-�*�O0/�Hd��Y� ��˪�}�V�U���'�%|w��+儩���ݢ錛}�x��ߛ�Ӊ�f�"&4���`�`�~����>�	�G�T"���^�2.����YI��~���U5��Kٴ&HIV|�fi��T�Ik�s��� �-�� ����W��ƂX�|�p���ƣ��=�é�qt���6�E���YT" UF�r�$q�H((1�vy��1���VC�L�j�,����ﾔ�\|+R���}�&�t�S6�4H�,�Bn��H�"	(�g ra�����L�ȀҚZTɮ`͛�M�X��~r/VE�`9Y��N�9ɏ �1��@�C�����tcV�v௜���`����Y����Q:��7�;d�H�κ��G�����KhHp�E��������[��|��?���4
1a��0!<	bDJX�8d���!���!*�
	��ne�m<R��*�d��#m$Z�e��7∺`{�v2S��!�2w�ύU��fy��N�J���bݫ���_W��������͞�@H�H��$V|;C+��+!|�EJ���?�ݧC�Ny���0�d.h"=k ���o�Iiɠ���,�����	dS���EVv7~�����#�����ݥ����gte^�+ ͊�����`휗kLw�����EB�ő�:���0��h�'�^�-?���W��?#���Ԕt]�H�lx����՚|ެ�����`-4@�n�9�&�ݐ�a��(5�,˻Q�a6�2��2�Ǝ�3Q�Q�/5�B�(�> ��קp�	���%<o��P��pKm�'qOY�N�Q�H�k�a�q��d0N�ژ-X> q���C���#c�KP��4ԯ�^�8�A6�%A�-�6�Np�ɼ�+��3�Z�}9�5���h��X��`Kʎ��b��Y��b�Plټ�g��7B�S�O<&G�L��Q���lZ�H��b�B��ڢ���GH��d���MVe*bN�AF��V�Y�\?��H������@-�y�5�4Ɖĉ=�)'�0��(�Me�M۟�h��!��  |��1�'�탺�i���s��p��T��~K�&�� zI"��7 :�H�@5A6�
�$6e�y�tx�v��ڬ<�'k���v�����r����V�'�d c�' b9����b��2�#�JK����g⨪؆q��.��q�պ����h9�u#nN:x��~��I�0/aTƼ��7���n>(M9��C��"������}�u��q ƨS@:���x�*PNQ���8z������9����1�wu\M{!� ,58N��cv_���0��!=_4��&�����3m�C�,r�tE�Ө�z%�T؝&�u�m���P�O|�|�ӑwns�������'т�����J��-�K'���{11��C ��e�g�g�:P���L�tZ�k���R�]��d�~85DSm�C��/�M�a�,�}3e:���?��3+���[=��K���(��8�B*3K:?�|� W���bX�G�\4x7	Tx�>I*��o"�vd?2E������Nh�"�{���f�F�n��S�֯���h���d��k�k��������seI�]��*���l�t�7GV��{�D�!{�h g�~	
7w<��9���6s����p��ҏ������]��f�j���wƧ�e����ꭳ3��+2f0�K�Q�t��4�6Q9�g�qO�j�S����,�m\"@�x��^A�&���B�V%�'=�K���b(tɥ�'��`���1z�<�GYg΢�ʑ�����R�q�QZ)4^��l#�2�1 �W��-��9A��q��?�u'��{�� �bH��rԕ�m�����S�bͿ.i����;���$�s)$�Y�urpfK��:���w�^�Mh,֬$,�(�&���h�s��M b��W���
.��aӸ�����b�ebw3`M�h=Q;�~lQ^��l��6�:��5��EIG]N�kRA!]���6�&9�ec̶�T�j.�jQ�my1G���@a��7V�c�&9U\�Ht;۞�=J�;�RȺ@5?z{L'���-�LGMP�+
�f�w����T�!JV���$0�h�HnД�R��`��
<��i������Q��Na�"p._+q�htC<FU�
0��D����DD���M�sV�y&+[��9����@�ț�[�X{�T�tOz�r��}���#�x��M���DS�fl�Y��ѯ��XF��8e�{9Q5h�����
Z�D�B������f�؀8����R�.F�#��� w괙xQ�Ȥ%	ϱ��Zu��%�e�nG������񙙒�$v�H��zM&Tbo�N�Ҏ�Et���� �{0i�0�_�e3��8�������27��$F�i�Js(������;���O&���N{~y��L�&J�#~F�%��ݲ0�*���;Z@�O��
,�C�x��h͂wE2����D��y����xњ�W�-E�b�T�Z�Aqss�F���Ra<4
���6Ürm�l}�ݹ_{��6��P�#���^;^��J�h��LRI�^�0y��>�yT�bz=���U]�'��M�@���\�ۃ�*�퍪��ӣ��x�����3xQ�����H��@��
�������w��@���������f��d�kSY�}7�֕e!D,k��K'�������I$���i����!}���L���Oo(�QAф$�>9�X��&O�����K\�pH�J�]$U��0�5�;N�X4O;Ks�u�Q�4&mι
�?O&���"�CG�����5?7T1�B��c�tEd���h�5�'��"L�Ðaؾ����%�@$`��#�8���
/�������nUA��
�Ԝj��d���o���790{e��w�D8�����n�ٴL���x,--�l �V������,*���09jW��i��+�Z���S�=K��(L���������
��0>���eʚ��O�n��O���
3FƄ��kl�������$e$u�n���_t����8��pKxG���O���
@1Iya��^~���5;�_��Xߘ>0"E(pY�z�A6�M.ub�Z��+ynf�O6��@�O�$���Y2T� �D����4Q���w|�C����u��mW���z{䒮�P4)��w6�^���xT�<hs��s��)@��_"����(#��|dR��G3�v�},IFxQ��@�w�H>P�EM�1�ж:ʔո�WQY�퍟6��F0(� 0�>h���N����P��P�l�@���mJk�lR�C�0@F*t���MR7�d�q�0w��t2?u���K��Ÿ�s!�m[��g��6� Hr��2��fj��W��/�:s#NCm��R8%�q����8�y���KJ�f5��f��1�W�G�C0/�-��DGRȵ��v� Z���Z�e=eC��םwKu����j�pd�*C�q��g�a2��ٱ��pM��&eu
��jf����or$�94V�i��&j�^ �֤�t�0'o�o�`u0���`;���;�R�8��$��2|Q�c{+x�H��h���|���$��Ij��o�CA��$'c�h�At�l eb���j?Q&
I)�B��Gr��yB�jc����s�������dƯg�T�L�}�۰��?Q������iL�׶'�S��W�B1��7~9� E��`�2��u�{�H^/LB/%��syY�|b�B�k�B�*�DϴRf���bn����D/,k1������]�L��|,W�	����#���8޽�	(T�t��䀧�lze��ɰ�3��#��%_�!eg��kO��|��s�����2�Md����.Лl>��j:��CNGo��at��43�k�B���n��)��\C<��I�����4�����vB��(�S��A�$��cX������o-�K�S{j�hb��a��2��yQ������x�S)=�:�	�o����������-^C�u��� ��mPB�~��t�s�/�BD�P'F=K�L����fQ�ǿ���@�/(b��č�խ���hG���`�̬����*���*%'��L�X\�ܫ*�3� �} �pl2`�J?8����(aܔ�-D�L-�1��X��\"�X��(�O%_U�n��U9�t/��
/��V��A F�"���#W�d���4�e��s�d٥��J�o���`^���3��@F߂̿h1�9���o�7Ya�U�^�I�9�����:�)FJ^�.c1-�@2�v�6ޒ���O���C�o�;؛�4��;�&�<� O%uMP��WM�#��*oH���T�Ka%5�����X����`o�!�բ�vt�t���4�ϸ��cd񷶥;k��L���a�&�\���O��Eof�g�I�x�����3XpZ�s��h ����x/g�w��JD��H�F��4�N�Ƴ��
֡ٯ�=$�|��I���T���#����MMa$����9Eki�sE��}�Q=����12���Z�v��zl�$j�S���!�w�
H���%nZSp��X��{�S�f�!CC3ڠ_�ۘ�ܪ�����f���2'�yj��^4VyU�D���h�&\���'���e�. �Ro͑��/7`�,Ë�
��@�4=�x���>k��7������*��9i�&Z%LD���h6�xf�����\���g�D�>�\]HӼ��G��R�(k���m��p�A��-A��`/�����"��5�)�_��>�!�M;.����^��𷬲�E���⣿�o�z�(?��I��|,Ϝ �������Ή\���\@3D�!�;��$i�:�Y%�	�2�I^/[sEj�����V^�j���O��ݱ�n�X��� ��ǂ�����B8�jobK�7 ��J�e�s��m?��
pX^����j3Y�)�g'`!ݰ��_�^e!�b^��#��Gg��X�[��ss|�`��G�5�fk��:����H���>���Rt�7Y):(V_���*�n���m���7�+��DoS�yP]k��ڷh�2�,�0C�1����/&~�;]��%rs�w�a5)=:ys�-tb<J+�oO���=�]���\�g/�굿��\��$���Ktc����ݓ�'V��pU�m/��r6�{��WtbU~���
S�X��%�EUR�ԧ��C�R��AG�o 5�IW�X�M#��/.,0k���%&�*ۅ/"73��t�i�rR����]s�]ج��q1����L-�J��bh�]<���O=�r�S������iZ�\�]$Dm%���$-��y�{�/ډ$0��e�M2 �m�f,��TwMIt�u��bC�~�C��N�g���M��²���v�/\�2��x9vMuu)���	��`��"��%��� � &󞷫o��t�����2X]Z ���״,���l���X=qr��
5T���O�/�X]5�'�d�tY~'9|\�D�p��'�NՓ���`c�X�0w�c���q���ز�t��䩾�R_��U���uH�\��1{���eE|�Z�5�oK�BUP��79!�q�u\��i��/�N�p��^��&�O�(�����
o��U�JO%����@�Θ78%[:��w�;�(�n����C�7�P�����ُU��8�aB^a�����5<��T�0nB����Ȩ2���c����dm8K�o�,���ػ�w�5)0�|ϮNL��v�*��,�������=��cJzP�,���+�<7tE�iY��"�ۉK�q:̹���m��u+�࣫��Fly7϶���c�B�E��_C٫|U�2&��L���T�e+X�*kq��_��s8S��JWGk��ud\���1����b�p���l�XI�������j<�U}���W�id߫s]��Џ�����W��,}[7��F=]	@��u����v�WC˵�'��[�661G���R�W�Տ~�ȷZxx����T��������)4�tQ��B�x�A�C��G[�^���_;�:��Z(n�ɀ����5�p��.Y�m9��VPwrj8o#-�9 �D��VhI.@G�~��`��6c/t�P>���u ����p���Q�o~���j�����쾤�@�p6�3�E�I����	t���cv �H+q{s~��KiAZ!�в���1���Q�W�dn�@��،���L��t]��cVa0��0_b����I����@�a��:o�3`.��Z� W��/��c���y�D3�xqMn���B�[�̧WZ訓���:�0�F1�k�:���c�vF��g�/3Uc98s^�$��':��p Bo���ՅQ�u�e����7[6j]�G��z����Y2��(��u��=���y���']pJ6��' �|�z�tY��ʇ� ��0�g��E�����A��Ho�(��%�U��%}��3nϤ+������ا K=�-�VL�؞�V�u٩�b��z�v\��E�Hu\;�a(��X�ty%�di�􎹰�cE�ug͍�Ҩt ׭ab5e9��6*���(����=;�`����M����>9B��d9_�,�D��%(����T3�.��0��=��E����(��j�#�Wgs ��ʾ��X�a c��~���+�FƚW@c��o%�
�do�պ��� ��f�7i_�:�{��FUeI�;ߌ��:���|Tnl�3�P}��Ї�r $���"9�)L���;&�
Թ>�:��HVx���A���c����
]gǘ��~��d����jC�0�U�MOg���Kk-:�`�eGK5v��~n��_�F]!��Byk��W�X�@��rDv�	��eAw�N?S����y�'B�h����#�-����0��4�BHKYʳ��*�1��aYy#G%������/�D�]U��S;q�#Z��8�&��rﭘ!h`���⃖i�l\n)0���%���(��G��.m1�f,�'���r3b_�"DG�?�
3�����⋑h5��n����En2�������[���9�����Z �ߗ�� ���
��Yәʮf��5@|�J�i��uX�G.�&�|�c]����o��n@oS�Axk�ڙ�r&�D���9o�]/��Ṗꜥ�3���a�AZ�r�d�s�Vh��xU�L�F��Y��5��&`������a�z�m ~�|�Q-��]��`YU���R]0�ͪF#�g �i�m�R�Z�i�|D���5����Apdg�q
p����QtH�X�
�L&�U�\�u��lW�p��1'k;��`�j́ ��A:��]3�L�)	15 �\4�,���?/e7�rː^��n�7U&n�2�	����s�4�V�����'Æl���E��;!�p���c�*ƧS���%-5�V=XO�:134M�������`"c�	Y:q��è�2o�f���w�Ĥ�|sk�1rј���]�i���
V.��r�OnS��l D��4;(�qV��`��U�X��"��Wa�_gi�9K }�@[��\��C^l2mY��m����yd��\��V�"�Bg�V.�������{��mq�-�%�ȶ��b�rn���	g�Z<!F���fz���msd��W��z�.��V�/�5iZ�_z�2�������ex�!ʗz��ڣJ��7���fLB,�?'�����!P(}�B1:�̨x�*}�D8�O �v�H��&�W�� ��D��a4;p7=���i+ĭz#�Gc�;Y
Ƴ��ֻ�m>�̾g_^E��D8�L���	 ���C/u��2G� �=Uc��#�����t�[{�W��ͧ.G�g���ͧ���e�yY���aPwڟ���w�4�d�rH�*�v�#���;FK(0�����l���є+�O>7�Uc��6��BX����6���
�!�E^
Ƈֵ3Gf��w-�q
�<�TɄ�pV٘��ϔ.?��n��g&���פ��U��ZKv�mȸ|˒,C�\0�$�i?�RުvbXB9y�i���n�w>ef'�xc5s�$]���<@;��.�Z��$Ƙ�������#��{��
���(k�x��of0w���6�c�u�c����!��3�4vj����C��%�(l�~��%����jy��A�y�M��d|���5 �KP�
.���b<�8q�P{XO�H�`Z���vOr�#��Rﰬ���S���i=�~������<��a"�螞:S�{�^��]�2�$�QoB��;5��GB�Z��+�_y�� 2}��������hF�
k�q]�>؏�x��"�W�A�<����%RR+i󰲚�<1�!d=�-�y����λ��I��XM�HB�F�V=���O�!��tרx((9��B:�[��O}�x��;���f,�a0zLφɨz�b6�s��v���M>ao#t�8�� ��,/ �6�W�o�.�K*�F�&`|ls� oK�>�S�uFM�N�F:/��X)Fy��»t�rE��e��>����M	e�K�IӴ1M��q4����������kF�Uq��{�|�ȱ?D�lе��p\��1)�=R��L���]`��6ϳT���PFiE<�;�������v��b��ö���$�XT�+�o(��W�6G�+QMFAh�-�F����8���-�	�IWi��x��/Bܞ51һ���K��y�D�g�lm$-�ӕFu=`�����N�w�|��fJᬆ;٥v�#����n����N+D,`�)*|����� P�ΏvxI�\�?� *ٖ����<^fG�B��7\���g���~��a4+8O�CEf��E��u��#|~S"n���禤ļo�u���S��दt�~�����9�7Q��7H�G{#�[��Y9V��
ͼ�qe�s�h����E�Ú�)��j�Ǿ�[tT��a<��#y�p���,��M������48k�t���^V��j�	3.�ة%�EgP�� ד	\�WKߞN�.��#��}�Qj���zk����R(R��%R±C�{c�O�g=`�b�Q*ag�q]9�V����H�my��/�St���rG���ZJ1��r�w܁%���9,J���Nm�V�g��Eq*b���^+���D��Wv�,y?��4X�Aѻ� ���T��	��`���%U�$\���W��HE<���F+o�(ɓ����=f�Z�k`�Y6�Zt�8��~s�˸ކk�\��E7*9�<����4<ѯ������ô���5l'���:ݸ�TQ[�l�R�´K�H�m���:�15J�U+��T���ݍ&Jk��(����b���;�5e�p���N1`�v�М��=u��!�ז�$p�qL���PY����[�Rde������t�r~K�G�C�7���P�����#�5q���'�g"���C�0�U˹��jR���pbh֊��<�rĖ�+ҝ�wJ��;��(�<{�<�eQ��-��&N�0&�б�g0�3��@�8[�q�wmd�>�gKv;������/�k�_��b���/:�W]@��j�����ス�T�d�ڌ��)ބ�x��TR�D���8HxE�!��L�\����,u%���4dh���ȥ/��� ��� �7t5�.S��������nY��ԗE��ö��G'P)�H��:
�,Ak�H����K�m�
+�����s�d��
��*��T�[���ɵ��p�*��٩��S�b���;W���>L`�������HXQ�W�� ^�otzůg�@��ZMq$�T������m]�(�6�R�g�J#���g����avp���sF�(w��ⷍ�Dng����2~4�<�n�.Y�S�4���t�T�G�.	 ����0 mnX�$���;è��o(������U�U[��^S�+���1	�k����Fb�Z[t���K&-��|4��V[�O�V���c�b@�^$��D�5��D�Q ~n~���o�gԍ�{��FD�f�`�#�k��nu�;��hTGpf$�>�:{j�]kGg�T9����:H�u|fh�c�jR���Q������k���3�~<@��p�����nۼE%�1�'���7�ᰋ���^=GH��$�,�2��}��r<��H�v�A05U�Ĩ y�:�$��/�L?2?HO�bA��t2�n�H�s挀�c�b��J/��ח��y[��Q�Ƭ0x�4`;��<��]�cO�Nm��j`�UV�z��N<u�^�&�w$�I�oa�L�ⴱwq?tZm}��}I�����lD�.���
O���g��.�R�M݉���p�y@��@��N��S��v{���n0�j��?�v�tZ���Y�e�C���R���ʗ�촸D!R#�G�(�s�xrXG�ڼ9��:[��$�.��Ͱ,x�:J!p ��MÙ�CU �$j����vW�=#�kѵ�Vԏi���X�����NP��,�A�t�-2l�	�����b%*���xA﫝b@ݷ�n���c�lh=g�1���E҉��� }�8�+�EiV���f�f�ot��fl���%".�H�~w�-O)\����:h`:�ʳCK����O-�3���h�$�.����X)ݰ��b?��~ʞTF��u��g�D윦U %QY�=�= �c���,"&c���".�����K�~��Q஡������+R���mr[-X�k��z7Y�!R��
v)z�m楓dO�{�z�!g�Ŝ�9J�X����@i�iO�;�}�`}!t��4�f�U� :J��(��>�ZX�#�C!��JF�S���^ҟg�uQ/��sfв�*�`������f�% 5ն����~6����\�-s��F�Q8s�J��%����A�vؠ�P��h��%7����gV
e�S1s��r}��!��}؎�VK`��<�=��a&�@�J���Mn4A��)KR�f�߿��)�X�veߏɴixJS��ے�0��gVZ��(lT����!ؖ�I��)�����5�o��>��w�ߢ73�˄������z|X�Ԙ�W��rKbT�u��`
�q���PF�rwS/4/1=gh�^��,0�{���Ym?�b[�f]��AK��Q����Þ�L�7ߌx�r�2����캰�?��g`>7���7��!�J-�P��r��L}�z%WDo���If�ʔ�|ĳ�?)ܫ�3Q�fX�N]?�d�'�~Z�U�+j`^�>��C
���Ӟ�:o�7����!��x_F�C���-
����R�����Õ_'�Iւ$Հky^Etk��$uq��Y:��ό�MW�G<�d�����mT�/��i���-��:oO�l�}��I0U�Az}%'#3s�Af����_���"�e�Z���p��$�3����]�&�Ad���B����~�[�G��X
���Q7��[=�lX�r��E��q���U/�(W�T/�V{?��fW��$��?��Q���i��_g����]��3+r��T��BG��'4AK`����?8�/�+n�0|!�y�I,���R�jI�Kd���Zމ���P�� ��.�O�sW�!�ʗ��R֑dՓO~PcCy���e%I�2�<�~�Q��"�k׿��W��	r���� �v�:��N����C��Z�Upq��)�����:9�iq���?��s<�8H_�-�����J6@,w̓��� T���G�װ���t9@�F�(���7J7�|	�:E����Σb�����_勤�@�f���sQՅ�%mG��۱|`+���T���0[}�7/� HK�H=��鰼�@��%|2b�OWU�wG�,d}p�H�_�ZJ�vuLԽD 54(A�+5V�3x��ݿ�=�:G�z��|����JKY�����|�zFK&WO,��_��{����p݅�Ïi�@;�uyo�u)5�S�.jl!���p\%� �=�U��	6‛A�R�6zv'Z�a�>su(\�G�[��N:�s�D]����"dqHz� �tڵHÓ��'�{4dk7�y��w��l=��}~b0w�B5��@��ߝ��=��ww�!o��Gv�U�x|��ƾ�л��ҽ�%�"��j�_���|��ꅶ- �Ԧf���ը�pTL��\.�HjŤZ:���q�]�&N�c�"`���й�� m��~;�t*AC�ٰ�YD$�P\�<����j��V�����4ן��9��R)(�ُ��⪘a��bi4L�t�1=��s3v^w�.��.���t�J9�b:�YY��O�QXD񗂫J�3r������4G�y�����ݧvL����Ю'z_�t�ps��J?ꁏ)saAC�sg�p�^Δ�A��`4F]�n	|�>�A)�ɸ�,�@�-�m�^�?�fy���!^-��b��]sŋ�����*`*2���GD��h;�\�;S�O-T�v.��_����ɓ�����i!X
�#Ȭ�Nh%����kp��iijJ!_j��o�?��%,xt#i������]pnsJe�f
��'����H�2n(/극gEQ�7�'���h��.�fl(#QP��Z��%UǶ�o��#������B_�Omr�]򺹨�W��j�º�s��׏-��y��N}�{��� ߵ)jWe0�>{�=������	�<�Ŝ|�6H��2�������n -���G�����g��"�9-�$Ǹ0�6�=�!��c�����g�KյCnؓT�Mo#�g�lRT�EgDC4]�3�k�g{��3jZ2��|��g�-9#�:ɕǰ���?�wJ��
�c���j�rYf��&�/��'tF5����Z���$+E���Q��a$bH�U��:C��HM�Q�S�D2�����|�x�h��-�&\�[�n[W�ܷ���x'�S8?�69�+�GmRn��Y64���٠g��;��7T�*|q�-ʵ��]cDN���~2|h8lk�e�׵�4y>#H�� �h����B���1�`Z�NN���hʍ�dv
h��J���Q&R��y���n�B3MDk~�ƠC�ʦ��a>���>$v��gF�b<Y'2�2+��\ng���np�m��}�0�����iu:���d�r)��&�*�#�Y�����R�d�b���\՟U��=E���dj�ˆ���8|�}b��5��4\cQ���ŸL���T�z��6<�5���j����kr�cm!�&6W�5;�����u����Cb{�u����(Y@�/�$�@���b������*c���`B	��sרD��y�T��҈�Y�LGTN���+��"7�s'/y�S�.���b��]ݐA���N�k�2v	S�F��6��G�|�m8�����) }��@�ym�"|3��!Ȏ�i�p|ޭ�]ҾC�Zg3�
5OH��s��n4-`�OIq3��Ij8@K��)X��{TAD���Ri�ِC��)��y����I�_��4^�<�{�u4q��Q{�l���RڒT���@����a�T�/Q�ºs�#l�2�r(�j�]u��|�P�%T@����l2OEqv$jTI��a����b��fr�R�rgbA�	x00I[%�����LV�Pb'4�e�������(�(�'b��6ro�W�*N�I�\��ƴ}a�1�h����������َy�~�諠�v��o��ΌuW�e�A%^���>�(����"K0Zq��O
P��= Yw�"�gǸ+G3��1����0j��w ''-q8��q �����v"�^�`~��Ġ��ӓ��Vv�Ƿ9�?}��*�\B�o����:UK��������NL%a-�!�<�7�j���!�o�.�TY��05���<�?
��X��;�^�٠y�*!~�=L�)�࠻�1� ��G��%@��$luZȭ�P0h+p#S\םK-�k����u�]��O#ϥ�ߕw�Z_� ���>$���Is��2<���q�fE��e�wl6R����t A3,�b<[~�zʵ�M�u��>�v�]�L�0�_FU��53�U?U|�����z�a:��"�T��f�_������}�4�
�� �EE�^� ���~��n䢙yVzjXL��9�n��L���U�[gw/t�n�V{z�e6Az��\b �<�s?%{rqӌ[�w����
��נ��΂/�V�?_�X�RA͔�%��r"��$� ȨL34M[�N}����d���%((��w5��?;V���*�ȼ��s=߆��<�6k7��/O�DRX�s(a�Ǩ��6��0��5^C� `M�w�D1�/Y�$�S�3Nh�ⶔ�Q�����1Gi��Vr�(��9-�<���0�a�����4;�Qʄ�|�O�R�d�Q��v	���ֲakS�M��?Zz���"F0[p9��2�������|+[��_5;	�ny������ ��gPp�{�\��;w�x��C�):Ix���3]�|��^݄D�iR��6��<�g�^�Ry�u��x1��r�ә���7���a�&=a��oB��`,ב�7Q�$y%����`@�.�/���k�+��I4�d���)]�m�����K���	v�	)�VM�c���ຉײ��=!������h��Ow\�<ii�.�MJ7T��Ru��칝e���W�2�;���%���T�CQ)������a�
�\aq2����O0vTG�z_��,.�Յh��2��n"bOM�B�t�R�����t���QM�F��CA_�гjR�s��f^?���7=�nH��WqX@��ܲm|���}��g���Ʈh�9p�럖�8z�h��5��3"<�J�K���D����6���Q��N����<��ڣG��e�kZ8�,�bw�u�[U�L�ֈ�^Gz�FR,�o���K��Ap3�5�*1����S�6�`~	��@xM���+�T~�0�LJ|�CP����d���T���L�>N�����L1ܵ���n���I4ײ�bS5']:7�#�9�	��{`<�a&���Q�yF��6��r$s�2t.�!��H����nb�5�³��jm�Ak�k%�/��:��˽������pX.��f0Kγ��f={t췟p"��i�X�S�A��*{��K,'e�t'��+��S@���Y��{a���<8���ƕ�-07 �G/jU����#&�6(���z��6��W\�]�>��X:YM��y�-MV@�N����w��Îy?�*����-�8ۄjd����I-���� �8/^u�2O �EP�������[�)*����V��ub��z�X <M��;�%g�����b�'�uI&��:`�N��_jc�ŧeI�ϊ��"�EeY��.�"��4>-�	�T��)$�����P�{37kr.�-Zr��-FmR=|�2*��_O륪r��D��Җ�#4��k�&��y�)�Li�����\�_�������^��pg�g�D]�5��6m��N+h�7^��� t�؆�;S(��|���"$p?�������6� ���P�,��Y�*���X��?u��%��X3���湁�=d���L?��U���I�r%���4Su��D�QMЈ/]�b2RX3�Xd�'^��
j���#ZH�U�1��2�I('5HF���M��#��'��JC8o�a8͞�Xq(�ꙮ�ɫ<\9��#�+jf~vp+�fp�2�����<B�����%����w�@g�.� 0�Տ�����6¤Fg���2ZT�>&԰����5�25��s���.�A��pH#�)�}Z��(���ǧ�+ӫsy��|4F���?�j\�c���B����P��{d0�v��\�L�+�~�M�b:���U���u��xd��q}�M>C󍿁�$�]�!�U{E��?3�d�n8b�G�R�È0GS���cj Um��H��,�[�fĎj�>�G��$.���3��2�s��/X]�,ZS�-Ǹs��-Uv�w�"��Ϫr�����E���?�y����.�Q4[=X����t��O0ge�/���#��X�]Pk�Q����Ď�B!�ڝ�N�pYHL�S`��%v63
s}�Y�}�Sم�+�d1'h�7����P�FF
΀rº}hȓ��qՊ����7�o�N�<
Ц�pC[U�/�-�FG�:�9.��R��B^G��O��C�B���]
��	��=i2�ʿE-pF4����k�f.�Y���裺�(Pn�̍�ի6hB֜X/��fF{^�oÌޮ%h؞�>(�Γ8T��Ά�\~��M�JC���:{e������{C�:h��r�
�x)�p]M)H��=�G�nK���G���A�t%�0��6Z[<�n*x�V��Ŭ�����I�� ��M"�*/���̷nXA���Z�rL�Ը�~��� .�\�#��pz���"����>��QT��샇`��6����k~=U�y�3���
X+Q����!�WC�	6?-1��ϭP�7T^���p6l�1�K���t�l�����&x��q��%22ƙ�@�Yb���ڒL�!>"h5��>"i����\14�r�(�����T�U����o�ܢ�rZ����c�3m�`$�߹ގ�z {�6&E	s�p,�#'WՏě��~�O����:1�Dm�[��̩�F���O<�_(�{|�s��J;���-��yw�W]��C�2�ZM�M��$��Q,,��Y�-���0���\�!�]���:��K�sS9�q�q��O���}gz��dDb��^+�Ա�FH���z#i9V\�x��?-�X\�U�'S���tB�~|�t�7~?��L�N2I��aڦnBk��y�Ӻ�D�R��g׶s8�����WP$�����$a�u�Z�1�Oa���b���ek�W����L���7�W���%V���l������_6� ����ʻ��`����˃�ߩ�W9�y�i�eDFw���Ua+�������g����)L�v�*������բ"��w��_�o��� ���"�T�`XM{E��-i�,�� а}^=�����^�_�p�g�BU��hr�2����c�mK��W�6���~=/f�ϱof?c�<�*ųr��W[y�`T\i�����,�Fע=����ߠ9ae[4�N/+�m��p��r��IM�F���yZ����:š������? ���Z?(��^�����t��9�ѝrk�r!2��x�ӏG���ʽgO�a[��}�f�7��ƥ���at(N�����0^y���Tq7�-|Eܫ����v�]�2T�-d:����PZU�i�'��_��H�-LH��H��Y��Nɼ��*��b/�pN���4��M	*�Ť��O%�	\�o[ʀ9��Ǣ~Gg�CT������:q���܈�r9�)��0G$�$���;����Z�y�gdr���.��<���hT�r�No��}�~�R$����.P��w�g��z��w�TX�N�oZ��P�I�`b�N��+8j�Pc$X���=���� )SJ`��f��K(l��jTVݦV�}3bbܤ����w��JP���z<��*x�g����߻�4ÞjڎV��ՙt����E �!0P�Y�7�M\�zi�p�[��~Ez#*hF� W����#2�������I�L���+�Z�$5��`J�~�.�#n�W�]U�R�ۗy}��*������JC�	r���'A�B�kd\�wI5H�
�
�4�KZ��z��l�'��+�ލ�1����V��,!.I	(�Z/ٟ��I�)^�k��_�iZ>�ʚ!��hC�����3L���w���0�'���f�k��e<\wS- (��i������1��D��/S�%�B"5WWĻx�U��Pn��v`�VYUA� %MQ�(C�\�j+f�I�D����H�[z��^��a#���`�2>/+#��4͍��n��->�i�,%}��g��=��H!MY���Z�.�5��̝0[s�����U�E�@u:�敥mD}�Iر�5	�`<�����i�HM�݅e=Ʉ��<�;FyΙj���8��B�UM���l������#��n��ՙ�r������t�)4�y��IH���dҽ0�j��G�����JaH{ch������w��8{�����4�E��#���3Cm�.�=�����s*M���i0p2����Sߤ ϟ��SE�$�*��\���m��>{�S9_.���AS�������uD���^{�
�p:g�����M�3�ǰ�n7��V׺z]�I�ݮq-�5b�3���V(p7�'O�C���Ԅ]���������"i(hm��Z��(�H�紁9gVp��}��P@V���d�ᨐ������~�����ӟ6,�`��+d��8Q2��OX1lw��bv����#�Yk���4�p@�y��}W>Qv�9�/kM�8���_>�΁Ǟ�.`̷�}`R�O<��WR#��!�q Q���<����D����@H�E�|0��Œ[(�	� �mQ1���6�]���(��d2b����Ey���*T�M��PxHќ�z�9m]iű�[�n�K��:����5Kv���A�[6EΪdE��h�v"{�I�FWS=D�Ap�d0^'�/��.T�;��"Ƚ;uZ��F�K�#LQ���q�S'��7�7�V����&F���WӀ���6�xU���Q�@\K��B�T.c0%�ˆ�J�n�c��@����W�:���ŕ�y)�)|���p�b�	�/���Q*�-?R��7�u���/��p����	��O	���,%�r�{@�K`�
j�Qg�^`��mOFQ(Y{y������Y����s�P�V",��u���u���g�媛��.V����=�J�pdp�M����u���]�����8���]����O$�Xǯ0%�􊱊�R���J6�~NE:�N3B	�ª�+W}��8��(�b�,�`.	g�ή`>Xٚ��S׺?���,fj���ӈ��a)���H�ء�ਝ����.��8.G&Ea��)�WRkG��!�jO�Y[�˂0���1�&F�������d>�X!�'z����[�zsN؛\7!�D}/�z��jL�!t�2;�67 �e_��E�_1�%H�_�λ�Mت������<�u�<7���H�@
:����ͧ��6Prv�6{���)�0w�f^���۽?p�{���͋�_���z@�߽Z/���,I2�i
U��t�i�J2YH�ԥ@�����^AMM�+2�(H!9��_����ӻ�+遢�Y��ű��]�تN�L�e�R�|�=+Fo��>��7kD�Ę.�=����k���,�V�����A�Hq �}�4�ۀ�6l�Jf�
_�k#��wI�9C�D���H[G��)O�o��&�Lk�-F���I�@5�჎��4Ӹ�c��ۤ]?F�����34���iOgnϴR;��Jn�ǽ.��;4�6��T#���s(�o5w!N��_q��y)�2:I����!�ʲ ���}/��mh��[�!i�^č�Z�)�]��2��n��pT���}<G�S���UK{���Z֡�]�Lա��Z9���䈯t��� }������>�7���5lB�Ւ��S6���aw>����䍳��hIhʂu�:*Q𼬎x}�;~�M�؆)Z6���ջi�|eپ����Y-3.&jl��k��H�ۈc���u�[k:�f������=C}8^�׀��~�{*��JƏN�L)Z✢�̤C�*� `F��)���;�,���\��S��|=�l��s��:� �$r˞�� א��;�ھ\�p vmI��^O�l?�w3�,��U��$�P�����%3
|S����3����-�Qn�-�}�P� �Z���>2�u�|`��	�3g� �J�v��eP��dQ�E�䢋������i��:���8����A��d�^Gp��@b��1b����u ��e���]�{�����]�����<���6�#Ez���6`��.�[����Ȗ��v���[�j���֠�i�Ϛ��	�
"hkx���LJ���b#{��i��8�<�g���a]�-����k��b?u�b,����/�/.�񙺼ҕ��0�C�â����¡�[d�� m`]̽�ZjK����鶾<YBi�Ǭ"���#ႈ'�)F{�D4*�f�w_B�m������ů���PH:}yّT����1-!�h�,$3�}|�G1�"�瘏�L=Zpwv��=��V)��ʓ�`P�{k9 ��I�"����/�������Yzm+L��jE��$p�Ǽ(л���X�߾�_Fy�����yHr^��-���s�aC��t����C|X�6{��n�˫$���a����E<��+�V���*�^�l[��/,����.�x�g%�f1)��2?nULq���,�7��������*)���D��4f$�K�X}W�H�ܩ�EiѾ��*���z���)n�z��Γ&J��(U¿:��>4��Ai��^��a��DI�<l�K[y%�f:!��a䳎M���M"�F���(���������r
�7��wn�Ӎj��^��cK����3DhO��oT��K��lNSM69j��Qr��4-n�v`l����Ck��m�ir7���Eu,��9�5z�nv��=�Q��r��6C©�� j�հ���{���'E3?b���D_����������"b��t��� 8�H�,V �S]t�M�>(�n��a���ϚOu��JGy���Tq��k}E���g��&Cf��hc�{C����V��F1��R�Kfkʊ�ټ��^�+�����ͫ�ĝ���Td�
���d���|����_���kB8Ld���m1~�}ds�$�k�,H�
Ƥn�"��?�G�L�^����W��g�|��J3�a�t��O:{n0��\\�&C8#�kg�E9���I�ʷ+ynuϗ�j��Ā����Js�� n�֮�B@�B�[�ʃ_s;g�Mzv��ň�s��<jJ��4;�Z`�!��/�$
�|TZ�P�{���#�2�HW-�g��$p�7�a$J�?t�Nt�ك������bȸXw7��S�إ��Z?o��`dw�`uzJz�3�,u�U�x\x [+[k��K˥ŉ����$���}3�<8�ts_@���f>��U�m�d!�"	���P����v2{;�"�`j4�n+3@�H(���oi�-K;�!�@���J�-t"�V�YC����y��vA�B� ���Q�#)Caw<g������J�ޤ�w8z����/�:�=$��OJ69���nT�U��E/�/zDL�%�+��J�	�g>�<>���.�v�+iJ��w��ϔ����<�烱[q�C[�6�k9nϔ���B�NTZ��Bqƺ�w�@��|z<�^9U\{_�$��{�&� �5X��@<��j�]ҭq+*�����]�Y�u��%2��Q'�!·�.7�$�6���8˾D�S�-�;>��=U��q b���"�pa�+���e ������}8��^�L��ݨ�R�q�5�����~�}rK��hUR��[���	�9A,��!#Jڬ�����#Ň>�C�
�E�;���)��c�ni�n/]� ��ǫ�~�v�qӔ��ed�	^C|��6G��"�B����wP.��va{@�۸zD�O���z��Iy|��b۟*��%Mqًe�[���(/�0L�����kZÜ�eq�=�G.H_W��7�k<r���|1N��B��^�>�)�M���I�q�5|��CZF�b)�G@B�������(Vx�r񳮮��A��y2qE�$�Fmc�ystfR��	o|��8���LC覱cl?�d̚��w;H�	�ջ�����<ίgs��=y�Tg
��Ecm<z=��  ����%�h���grJ���Cvs�\�í�&0.!�����E�5���4w�_�qW�bTN;��i܎�Q�Q�E�L�ËqܪV���̕�
�=�|t��4��}𥵟������._j`���/-�t�K�g!��w�b~��v����u�fD7a;�߾P�v���%�c��������LU�w�+S�!MMm�Y}RH��7_��$'�^#	�jF���$�L�s����Zsf,x�T��G��ƈ &�qIj�6�ZZÊ>9E�J�V��Ux�ݟ`c���_���)��:�k��" Ro���X����n��B�Γ�8�Pl�I�/�����VM�&��(��:/%(�>OSVN�Au�n���#%�?�n�q�q���[�ة�b�P.��*`#�w0��N�ʡ'����'Kc�<��z}�Ή���4侕�װk�h
���c2*hQ4���eB�2�ӆ]�aL��$Վ��^��g�DzsX���Բ�]<{s���S��ӕ�N#��F�'}h=oϲ\H�2�g��QK �`�ߧ��駔p��g����}t*E.�텶��]�M��>���u��M�9~d�;���0>%��G�G���z���ŝ	8�/X�<� ��+U�&��WL}Kj�'y���Fyk�r ����M��w��K;��0Xc;�=߀<���+ס��  ��H��~�����,,6����\���=oA��1ԙ,�GY]T�.�� �F2O�n5��"&����Ʒ\�Bg7�y�W��~�y�*,9�?� � �+���,�����<X�Q�څ.t��T��?�������A0z�Z6.�N���]V�+�v(�nD�8�?S���j��j�
3E-�(������q_����Y�y��U�8t�{E�f��.����*t�ޛٝS���u߫��iX4ު���(G���yk�ն��q<.f�h>+rǮ��(_���X�y���19Dd�(��]�� �@Z.mG�]��k	���_�-�7H��*r���#f�t�YoެM�G6yɮ��`����As���2w6�:�I��΋��"�xP=RZ<�.4vW�Z�Ν_D}�=��>�Z��N���7A<�� d��/�(:�Q������E�㕜%|G��X{a���Fc�x@P���R�����K�ߝ1&õ�Ϝ�T�.a��0]	<wn-7�,i����f�Z�U�1B���2X��.�7�3�}��9�)z�?�:׿��BI��@���m���³3���.r���g�+�M����>������gQP���[�����2�;�F��4j���g3k�mI���4:!y�x����S>�6�'6�-l��U;���y��w����jE�A+�Q�s����|EQ�����UuJ昮�P�`Н/_<Ր��Ʋ�&D"�rbh���.M�3$X�����E�~�B�c^�:��2o�Y\#��0�	7
�`H�
��[���ծ�۴�k�k\��n���wYɔ�յ�����|Ѧ�CR�� ρQ��o��ĺہ�2��&O�I0s5���:���g��.B�&���o�El�(�9NK�4@�j^��c�^���n�3���i��f��KkA�D����,��L�f��f���v�m�?4+��3���C��m��E��!!�X桖󢘡��'	��Y�������)B٫���!�A޾p��:9�AG��<�͛Q+zK�o���h�A��Z<EU����wZ���"3��1"��Q�H�\�d�B�sG���0Ȭ����6L#��q��O,�fOd �%C��}�)�Z����ke�ʃr�E��:z���I���&^L��R�Ф�����*��П�%��F:Υ�4�!(�0V�|f�.u�mI�.0q-�Ĝ��̶�Y�:D�W]��ʽ��R!ؽ��_ZD��%�հh�A���Lr���>~�F`
��$V��ˍ���L����T���]\�|��bĬ����z5M��x�7�Z-�;
?+��+��w �yI�a"�$q�]p�������C�拇�38bWU�D��i2��M�M���ϼt��'4��a7����y<�]t�����;m��� ����ex-��bvT�컦s��U/������/r������u/cB�Ï�)z�_�@	�m�.B_B��n"�9��;B)�s@�V�b�F`�UyN�?$C�Ȣ=/�1���)S��Y_�!�ǥA����<�#��>��L�QTK�F���V������j�zQAG�s.��؃(V�(2���)�;8����ȝ�i�QJ&�������-��$n2;�LZ��p� �
��@�B��v6�3�[\�߾�u�%�,6sVj��qP�˃Cal
�8P]|����i��-wCd�c��W��0B]+����a�<��Ο�ߋ�a��&��3X�N"/�,ua=��Y; 8l�~݋�_�srӘ�6�Ҭ���G��v���b���O�2�rF�R���I�O_�
sL*O�i�os����ˌ ÿ� P�P`�I�Z��A��k`�]C���1�&�h4�FJ�;��e��^Ѻ��B�rd��E��@�Y@O�1����a�7��q�ﳢ��n�Y�d;�i�9�M�_�}�2yU�l��~�Sf`ˤ�|����^Aew�=�4���y�bA7 ��FV����iV_���D���� 1��桾�Y�����Q�^�&Pi����e��Ȣy?��q�E���Y�'�>�`dM��74+�9��Iǵ;��A<�}ܳ��g!����{�iIfqڴe�<�Lsͻ�3;��V�IT��)c����1x"�I<9����K>���"��ٔ0F��FD���zB�A�!/�8�ɱ��\��N�+6 �vC����@Sba�.
%υ�TѾosTK�΋R�U'�ɝ��0�����t�J���|Ά��=�}Xf��AH�҄�� h��g_r���m	�TUu26(J;C�@���D/?
��.`M���1G'0P�����kwV��0I$ɽk�d(�(b��@"�W��s�{�����p̕'���l�FLTyN�u�����m� a���]�_(����7��Ԇ���d�x3��$P��G$���)w�6�-YZ�(*t��F�C��Z�}��n(�I"��RL�xVLp#J�AA�;0��G	�*���&xk�@�Q���aO�O�	���d�PMXɖ�^������7h٤\B1W��*�>��8T�*���6��1�7�+���h �efࣛ�5�﷛��$%�O��Ёw�g}`����h��o
������!)�l��܁?��е�{<��uE���0�9��Y��d�K�U(�WtP� ��"DT��»�e��K ���OS�VJ`�<��aҪQ��Gh�2���ǚ����=v��v�|���G��=��R�%B�/���#����^͜!U������b>�����:�"(>������NH��l�`[o������8����}A����cr>5�҆��	�@�X�=��>P����DNx�����j�~`�S��+(^�7M\�h+w�c
�7"���ȓ9�ڛ�5���;.�q��!�U���h����,�Z~���|?���U�C������<h %0�[���ҲŜc�w���шP���A��N��G�9w;e4��p�R�ǻ�ND�K�w�e�lA��(Fg7/�8$b�M��[3k>�,�g�?L[Pի�9��.��Z�"�ֆ��:�v����	0�܏b�d7�R5Qt�Wa���9Z���8��z�/Zh| ���S̞y�uko����{A�ns$�#�7��o��rA�NmW�`��O������8ujnc��'1�bq�F���!h�4|Ya@�UY��ހ<l��ޝ���"̼Gg�اȞևT��Љc�)Q��	�_94�+��6���hu��a���H�8�o��E���XrY�]k�N�U�6"��MƗ�э�F8y��۲�hDƢ�bPA���)2��� ���ٛ���<�C��=zB���5���)Z���u��;��߻���s58�#�
��4Pl!!Ji�w0����:�wa���I�v!N4U,SU�=��~U���>�)�K�5#�1����j����|ze����x�Z��)ͣ�t���#]p��������2K��/2����
����]G���9��ZJw$���E�ۭQ�sn,��o8��A!4�������� d�,o�"��J�hTk�,X��L:n���{��_��M��,(��ؘ��g.��{ �V�2-����:�������i_�Q�����ϡy
~�5<~���?���+@lf)-ք�v1���=[��>yE��	���%Vv[�|�QȌ�M/��������7�Ubk���>�Ã�qo�[���=�D?�~|�� ��o�]s�M3�L�t�o���Fa�?~�b�f8r�����zF�=w:�C�D�lx*'�.��
��
=b=N����Vȑ�.�t�h[X+�9E]��7B��TUI��.6Q��OT���@ŧ����{�T7;�; ���yB��O�v��q?#�6�tc3|� �THHV� ��0�uaJ�׼�C#����x����8& ��v��:�#�O ��,Vni��7�T�������!��z>ҫ,��'�bɨ�w��/���W��K'���"�{�B#��[�Eh�O��%��W��� -�o��"|����x5�������e}�W4��Y���Fz�|�a2߸}Q���! RG��H���z~}�=�����o�;�6*s��Q7ݡ�{�n�5	��`�]�<8�vW=VA�Z�w,�l�L��,3m���!+���v����)��&D[��?	~��ݠ���C��{eM{ ؃�]s5@�3����2|�w��!Ť��I��ۆi�'�3!�S��Ic`���2�~e�
 ��bݮ�ܻ&���c�ʙ�B��36ߨzJ�=7'�0��喓c�3�;���voIK���s��k($]���[C�ז,8l��XyA[�_�<��_�����ιӔ�$p�^J��A�!���[���G{���yz5��a��a���#�(5b#Q���{�O
Q,��c&�y�[+�o�2�T�4��L=��eD�?j�S1�ŭJvgг���}���X��?�䭽�6�mYh㪙��*%v�2[�K̃#��Q"ę��71H�*6<�օ,�"G����qI�QƢIʯ�Խ�+p�mL�~M[�B��'�LJ���fw���\��	8dEM�4�B���ۺ�۷a�����ծ������L�qtt�xG�����*���#��Sk$M`��[r\�g����������'����	�E����q�x��F��_.E2/�NϘ)o�O�:���ٜ'2�� *�~M�)�01����S{�~�MǙ1y2��zj����̧l��e-�60��I����uƿb �yj�UӜT�g�4=�T��'&�z�F-I��dD�҉�Z�H$*��:*��
ڄ_�n k�U}�u�h�;�:rr+TM;o�a`��(�gDgb�������
��H�w��V�W1I�,�Qj�R�%��_iY瘯ʠR��t�޺@B�ۀy��t�ߍڹO��AF
n�.9�zz��J�[M/�c��H�휜KS�_)�9�!\[u��}�Ѵ�ò/�EҨBuưD������LbW㑼�e X6n�@���F �$�*���mX"�o�Y�����ey�W�>E*����7�D=V����T��O]Pၢ���'���҈n��x�!�-L��b��+.!�\>���ǩ؆/Z�����X·���NO�tw���Yiy��C��M��Fj._�
�$)mn�rǱ��S����ѯ��5ffw��u�{ݤ���M�6b�ǱM쇋U�Ag���Vy�\��|tL2�N]��]�_���/�A�@�1 Ն�����F���T�F�zچi(��#W��7��瘢nY#y����od�?1�_�9�ƒ�nha�[�u����3�8L�u�Ěc\(Wix�P�ӷ���@` ����ų�oh꼱�3����,Y(��mx��D�\JӀO�Xjm�`l;#X(U���?V�@Xo���lI
��C�e�xY�+up�a��Q�g���ex��JŠE3{q�6*P��_�YJ�(�\��fQ'�&�����[�hs��8��q�]p�Tg%��xt_PpH�L+�e���{�ӟ� �%��x�!����Xܡ�I����\xf���AQ��'?����iӔ��)-������:�o���l}�ؚQ���a�|Wz�cU��}q=ԍj���4�6p ��a��Ss,0Y��ܭ媂�QS�!n����`��Yأν������`k2o��c�x��Q�K�� 
G$�8
 �A�h�l^`���K�U�U�Fh�k��	��z?A~B����:���	|�o~W��~�&�Z`�9w-�.�Di�wU�R3�]ʶ����2�u��B2��D�y�z�)�]�Ik\�m=Z9u���uZ����pN�,<w�[�e2�?��jV��:�fpI��dN�V���3E����u���=���Ґ�!�r���iSI���7�^�^��ϵ��!c��ͤ"�L4Fer�I>1�@G���aD�!�����-T\dpIw�C~6��0LV����0+�.����2�jǳϸ�>�f�l��`��-����H�8�V��E稂1~~~�˳x���mR<C���
�cp���-O����s��t����vK��am-Zk�=�R��K�+������ܭ0(P_���n1��VڜLo��σ"�;��9J�iLܸ#% 
H�#7��X�m�:l}�X�S-7��#��ja�.�ɡMa������l&���6���>+hG���՝&���Gɱ���>�����ɪp적DŮ'Rz��(w��2�ŗl.�<e_�=H,�YT�ӿ���]���4����;�����+�2���d���õ.��)�Htvl}v���b��'�����e�%����<��m��Hu��ь�/G�X2C���H�()>������� �F�s/x}���,��A�2$�5���o{�٨S����c��(Fa\�2<�J\�J�S�����ɥe�+�p?`��ߦ�[[H������&�� �YR?eo-�v:����#{��¸
5T�����.Ir1��t�|��嬶|f�ĘV�z�2�T���Tve�d�IT{U�A��O�h��2&
JBcp!x�-��˶�]'�b)���u��o�T �]�ID����ԋ��w�����z}#�D&�bMcdu�f�U��*KO�aC� 0iX/o��aJ`h�|�q�@��5�n�Kn��[(�\�4rS�Pە������빥S��7�+�w�˯u@�c1)��+��H����Ҭ��q_g�����D%�Z_7K/�h�x�H�wT��"���]ٮ�s&̬�}�.�V�������SOe�d���uQ�Ê�6���'�i{�5[GQ�ݙ3,���R��f6����ة9
���T�%���ld�l���T�o���w��y�dPX����\��_-��(eV@5֠/��lp��&6�i��Խ2�8FJ��2�:�-r��.M�&�x#PuT�B9ಇ״AFR���F�wiB����?�KM�b�A�KX����W�}�Z�c$[k������m���KG��2Kz��}��ڨ CW��1��X��}�W.����ZZS |`�����S���d��aD8�	g9fB��V�0��o�X!ju�r`��9��p:B�Y�]o�������?�`ym��)A>gNӽ9���n�+��J&��vK���3��%⍰��Q������-I�/'��+B�9�2��Ǥ�ݛJb�෰��e��s�daP"��������ӛ50�����&��ݝ�W)������w$�}hw��5����dg����W!���[��>{�J���q�x�.�����LS@�԰w�1J �%7|c���YQPr2�(�Uw�Z��H�#�¿�T�;de�%��%<���{�"/!V]�_J���]�VPN��Ķ�� �
��uJVf6�"N��ܰ*tI���NN��Ħm/,�~͑�����Ԓ��hm�h�h������w*�	E��DD���?D�=w�����p�񋷴Ǵ!���@���j�B:�$*�:#P��j�vF��F�X���R�� k�FE�����lH���
q<�!��Ci��?0ׅYl:c[k��/��m?��1��c�~M1��u��l q�dg�G6Q�!�˃�?���˹^���.ȃ#��>��/ZT- ����yM��˷�5�r1�;�����`jE�̛7��Vع�Ɠ���o�ގ�n��0��l"�,���w���N
�$"_J_?���
ؕ���zj�lCw�1+�5i5t�w���j��u⽔�}��j�A���	տ�Z߳�5��j��d��}���$NAdEXC�NI9)n(>C�g���j��=�����+����{d�V�T��b��1��U������� �;:�I���%��@�ǰ�}�/����� �aZD�.
�Iy�KMR#��
���Q������>ڡz����Q�}�7F�3�	{�.�cw�
�L���w���|�R�O7��8Pd,@�RrD�����������B�� i��j�ܲ(��q���.�d��GQ��s����Ո>r�܇o��d�͓�4��V3dA`x(�B���A�Uz[��Bb���E���N�4N�ފ�v?W����Ơ���7%�4��7�;����/~�}�,��f�U�@��pH��] C1�K��ڿ	]�ބ�=Ḧ!Y�{�_�2��JfZ��2�Pl/H���<�ET=pşgU�`�ntĜ�+c� �Ԋ�����ul9l�f�!�l"����f�8*�TЅ���|��/���"W�'�a��as�TH_�lnj�s3���B, �<�ph��/uI�lhE��S�c{���1H�3/yb�s-�\���&�F�������uY�񎲭�PB�uˆ�XIiGB����g��nR}�5�u��sˏ�v�)g�ֺ�;����2��pPu�� �1���S����MΩ�	�@'�Z���� ���s(��$k�65�{��O�3-��*av���V�5]�b]�����j|���S��άꑡ��M�6^7}ֲw.�ł��������x*�� �y?�j���{��@�舎�ͫ��#�>���������U����\�����Y&H�Ɖp��)~�*j������/�x�g'�t��J��1,-�c[Եg��NRkx2�f��Ε�����b�6� IC����>�F��[�:GW�P���Ɂ"�Z~LM�41��7�+J�M��ܪ
w�_��=wW�NPfݍ���d�Ns瀲�RLc#���c��-L�Wo���P��S��Z����G^y������F��Z\��1#g/v VKa�t�st�Y�E���~�Ax��T&����rCM>jF~m���5B�<P�P�"M��-����ۦ4�Y�9p�
�!��&��=^�a��.-������L��((q<�E������c�/½�s\R�W��U�z��n�U4�6��v^�j-6I�Z^�
Pl���~�`	�v�/V3�KcG4�ԣl�KjW���CS�R��r��cT�F��s�-�t˞L��2^]-�)�N��qD���V�R���_yt�����|�_{b��͜�ͤh!�W:�:�������&�Sǜ�.�T	�F�$H�*�aW�#=��qT�M&+��z��e:�L�W������LM���i�_	%rģA��P���4�U5��ѯ)�쾢��M�lާOȎh�
^��:e}��
��r�>�ؘ���j:����=	7����=�"D�����1��-N�;�z�,���D��=�&�r-^�aǍ�::�d~�iG2��
w߿�8�˥{\�KD�*����z��E?e6�`�B�3gW�I�^NӽbH�%�`�2��Ewq���]b�(�Sotfބe �l���IUE�ű�%�)���A�
���F���j;/��Ow��k�T�6$��P��8�l�.CP%�n6��%�ʰ�˂4g
������-�f�����V��V���~��Vc伍����?�+���Z� ����kq�@fH-��$�
0$��K'α�^M�"v�sJ�U�Yir�y%����>�E�	�[rr��6���ExH7�A,��q4,0���}ߠ2��8���-�8�f�=�`۷�R7��e�ȏ�~�hzR����R���J6�d�+�&l��ٷ�(�9��@��7�t�u�	Q��$��ʌITb��r	G HbW�|��l�a�\-�1�삳TtG�\�XAakZ(����Z$=|봆�t�hqC� /�L�'M�I��Q�F2��a�^� �H�:ԟJ9�=�Ý���ԭ>ߌ��9hDP^��?�~$3O�P&�CC���/IV�,V^!�b<�N-�������4)Sz�ڬ(KA���,�qf�e��w\	�с�b�>1��\ �\ΜM�6�\�VU�"�Z���XÉ)G�i*�=�I��'���I��zO�+�>�)�p���R�J�|��m��қ�Y�����B>�b��X��:�a`
z���d���R�w�r"C����q�n��2����󇳔�
x yf� ��B9�p�k��銆L�"�y��R{�(M�4k��U:t�):1fw�֧��*��)f����+��\Z�=Wݚ�H]�=Z���~�CX}L���7WS^������g4r�;�-���|��E����@�A��wKL*�]{���/�f%���Q������c��	�Ql �FB1G�	!y�Ǖ�P�yW�+�Hɩw��<�. d�N�˗���"C�mG2�ܫm���c+����X�~�-vQ"�@�:��f�캻�+��l�����-v)T �Og�:s1��;9�|@���N��HY���y^���e��g���{����rc\?0I�����]�	�2�G�`�~ed��Z4-��gD���w�n�̙��r���fn8��<82��rJQ�u�+�*�Cb��k� ��Wq�dF���:��L��ɭ����w��˘���ߎ1���:��#��������Y�C#�к������~LJ����.�"���"�kt��,Tᴽ�LH�������w�Դ��l���3)B7��13�Gԋ]�'<!)�5������ٮ6��9��3	��![A�>��k��e
	�H�P[��H����l���D�]ǈ��K�h�pPr�:*�q)o��C��2]�u�@鼋��S�P.Bf_a�\�y��`x�J�E�n]��Y�j1��A�]����=M�G�Ux���'��8����D>6ǭ[>�?cVF��o��	���CXF��>�~� ��]�2��Z~	� ��K/Ս	k�f�.y5���E~c��0~S�c���O�|�NC����6'z\1Ӷ���zҷ^��C�7	CO�^g�!Q-Jİ�n�h������h�Dh;eS A;���C��Q����|K ��˹(�S>d-:Ru�$�Su��[���
�w=�`������kƀV�@�l˚��t+Q�X��p��兎޲�����:	 *�ƍ��R�_�ժ19�F����_��*��d��u|	�)��}��~t>���"�s�1BrE��8�F�
��������9^c�+���4晀\8�VJMT �a��(X�v�C�h�-�WC�io�F
X��OL�5����,��E�gc|KH�	]�]Z�E�� ʷ|&����沁*�2+�$��ХC}/��qF	{�uZ�|���;���+��[���|#w�����
������K ~%�N�r�#��	�NF�Po:O����!��<����X��@y�(�u�����Ά���>��@���}h8_і��:�R6w@��:2ԣ�l�P��@k��@����i�r� q��B5�_�a�uD����:�fH�tP���x��!��t�衭H�,��!�?%�k"k�,�H4y�l"����HT�}�*
��X�,�N%��p��,L��;#�ɖ%G/r}�����3B���/,J�0h�l+f����wg&#��#|����!/n��>���Dy�1N�=��Ъm�fR���BaP � �8*h���?�o���e��b"�b��U$5uq�@��/X�%�z)����D/`Di�U{ٟ�*��1�4lTvW�VA�d]6���9�� �ƨ��ځ[�_�L�2���I��ٟ ��lꂍ�
o�h�Spۂ��b�&$%x�t�l��c�[�3%����� ��ն�p�x*������щ�R`"�����U���z�;�W�>����E�l���9C�Ȼ�lY��AXkI��n�6�ƍ"���NWV�q2�u�n��l�E{�S�lUU��GI
[�=>��p�^O���<���$j%�e���t��VE��.r��
�S`���'Gy2�NK"
?~���}v���:�]�|�I���yѥ�PCYu���A��
Ź2�{��E6d�7�9���q�e-K�EK۝׶�����\�ky N$ 6������}	����#�D��p��r� �{LY�oTұ2�o3��J�݋��1K����Q}��v��$GD����m<�h�8	M~V�Y9��Bݪ��V����p��ax�.�,x�8΋m��yR50����	���?>R�rZ�"�B�<փ��׽A^�)�ߎ�ğW���<q.p����2PZ�K���� �Wf1>0p��f T��i����V'L�H�SH����OzQ\����Z����j�L���+����#���G�g������q�4rDZM�#J��AH�;���0h��Ã�C���F%��~�����`$����w�АG�]iPd���K^"�y3܆��e�&e�M���n�-���l�w0h�7<�G �Z�|2�뭔��-<�wr�e�Md����⑁�����=%�M�(V����HN��I
�?k.2�d�(R�L�_b��ğV�M�Dq2%Ԯ.��>3U�(G�b5�q�m��
Yq�?]�6O�k�9�"?�v(B=|A~�]�
��B���/Պ��+��)!y�|�e�3����,���箬��`���Q���䟏]賭:�A����a�|l�i��KpR��{uXN����S<:����8�b�Ȫ�\�`�g?�4�s�2��7L]�}&'�AS�*����>��u\�3l��U���� bz��c}u8�4�ܝ�ς@���K�PoZ�=���ը�'�r� ]��x�%����<��GS�J���؛��xJ-��;�j>�M�c�`v�F�U � ��M6��LV��ı�bjy.x�)�'�<��kk�n��N��F�g�]$�t�x�Y�5|\`@�:��e>�ú�mJ����h�ؕp�53�VT�O��zF���t(��nO��th��A�>�9,���񶀅�~ZeV�Á;��̗e3����J�z<c����-�J�Mo������C����&�sh�M���M	��u'�Y@������ԋ*�RQ��>WF������}����?#�p��Ν���c�$te��C���{�5q"�H��"g�Z�:g�>�s��c[�*PѶS�(ASf,��*\
�ˊAL��ϊ�SXUh*�����ݴF��)	�����,�@�P�cʏԧ 	�����R(5��!�$���<I|��8^��'�u#0����v2�-&���]7�.^�Z�0�Ӊ�c�nƐ-<]O� �+g@ u�T��'�$�,���1�ƚ~�S:M��̼������k�Eb ��r���H�����y7����jMk��iw{���� �zi�z/����/6>l�0��$Bg����ׇ���g�I*�j��~i�NDf���M��$3����g��+�"g��1���6X\x4��{nr|��ψ�K#j|��O�ji޼��l�iR� �x�	����'��6��Q�>)U}���eH<��v�zL_C_]��q��6���>ߒ�CR׸E )���(�Z��5�N���8r��.H�
�L����}N/e�r�܉��;��"|�I���RujS~�a�o�NW�n*[�|��'�4c�0�]�HT�`�=@�
����oз�T�1|�ր^ <�prm�J��4��~VG �����n:��%�3�N�?��H}K䋷��Ԝ����H��P|
�;(fm�<آ����7�|!.Q��[8����vN	Mn��PFn��E�uaI̠��w�=�֝-���H��#�B{ˠ��N!�DR��L��oD��eU���*~1��ؠa;�gdt���a���r���U�Y�3�d�[D��`I\l#�V���Q�U.�N��=�e��<�V�ǽ�����0�]�V����起�$�&A�tz=v���z�orMގ3�
��<�?_�丐䋼u[$�ۻo��Ŀ���A� ���ZՐE�^j�! 50�|Q�O��lr<$��1���;�ЫKo�B���d������G *�N�,����޽̂��4�S~P,�$��5WlIdA@R����0jB6�;�B��^CY«��wh���cQ�%h�����5��<^J���I�G����Ǳ�!GeOz3ݺi���q3E��y�I�tT����n����vmee�Ȃ	��4I��R;_�Ֆ�7�XvI�=`ǆJ��Wc��Q��W� �ܙ
��2�<$,���?�X(�e�:���c��ԇ�B�--����k���qJJ��9�S-f�Eb��1��RB@�|9�P紵�G ��ْ�*�U�~�Q�X������ƚ�tCQ����5�T��/7]����s��$e��;�;_+�-�ܷ'���K��~����˵p}�d���������lЍ�P��cSL��p���A�H�G��5��o��+��-�.Hl�n��MR��Q�v�Ж�>��2 �q���Zpos. -���L�ݺ�$�~H�Ȗ��jk����b��|f���\TKp���P"�޸�aS4���I�=�� ��t�WU|��]��� ��$������3�.𻴤���H ��|p�?>͆U]d+��dλ+�ٜ%"6���]�js?�Ό�n��u�|@"�E���бb/o�"�DID$���'ɱ���
-t�����*��?��!Ξ�t���j�z��G���wq����P���l�%����� �0�-�����tv,���c�ǈ��}��8x�l�!�y���W m;��F�����̚����Q��dZ���`��c@��$lM��+���5�z�扃ɂ�̋jp9��)�-�x���>l(,�)�u`9��K����\������	k���m�v��S�Vwp>�'7TJ��P�{��}S����K�7����bJ�ͱ��E�n��bݾ+��:hك�ZȐ��#�����56%X{

�
����1�Q����s���1�1�4'Yo�Q�,��W�.�}4��m���
���#~�@���2�y������n\�NB`�_ͤ�\��&�Ҍ�����]T�w�Ɠ�cU�,ʝ�;�� ���"7�c���мT5l� ��y�������qq5��E��tqzk�����f�-�
��7�A*����]�J�yd��	��Ǡ�,;����qU%Y�5��8�gjb4����6��(��a?H�c���������2��G�ߋJ��
*��}�/|k���"E{��ct:�uv;�H��;A��mc�`f��m��(J�-��ב�h�"�L���n-2�ſ�x�#�	������O�Bx�N�Z�ʃ*�b�朧�
�ެ"���ҷ�`��"��~�b�WjE��q��Ф<�d��>��9�'_�*�Rl���]���ͫ��n��U�Z]Z�f�F�����q$����Q��vve�L���f��0�9�t����Dr��b��R�"�ߟ�[_?���K��1c�m�3�c'�,��hLf���9�n��t췢P��__r��X6�e"��K�ЁqD�Pb���f� ��b<u:7��DSt�oԾW�İ�k�c�����r��X�3�7��8I�b6��̃	ץj�$ĢP�2������G���$�nM�Vk�5�悛^�6�����Er۟3��4��j��E�{GH��m�H��S�E�*�^HP��*�x�C@��N�Ij`z@о��l
����	.2/b�lhS.j�}8{�Q%�-������Gɮ���˼��}u�vFo2x�(9�O@u��[3�M�G���x����)
0��a��l�8mKSs��U�����������N *4��Mz�C2"�F���QeŤ
&NY����g��5��L��uI�e EDǤ��a�����Ȧ�UB8Wt�gڅ���b��F�@��� ����š����8ʛ��1.,�F�JӛL�=�6�_�G�FK�~Ob�U**�;Yr�Ph���H-���ӄ9H?�T���6����8���M�<$��`�ŚӉ��٠�{]�������,p���K�-��	�H��#>K��P�r�4�
ZC��� -@�oe���Yc�J��/���k-�D�����@�������y9Lwn0��.-��uQ��L�eg�e�\�^�KE4f�z1�xOf�):��2�	Ϟo=�q��Ix&�R���5�- ��+�|��q #�^q	��򎏈1]Yq�������|�A��5������ �-�T�H뗩��?�fpW�'��V��13eFM%7����h0#'z�/�ŏV�����[~>,HQ��*�|��to�W����.UWK�N�n˥����L~�[�K����
���C.�M����?f���*�=���������z>�P�q��l%sC]��"N�<��	οb%?��R�j4���dI�!~�Ѷ[g��kZR�[(��-���TT ��T���n���&�W� A�Ȣfhuo���
1?I��G����w'O ������9�p"��}?[�ʴ�wwQ8n� �:�H�ۙB�o�IC�>K0��}N��O�m%���s-(6���"�K�j<��L$�~ua�A���.����U4��xWv�6$<H��7�ms<s����(����=�B�O�����RM[�t�GU���Ĵ#F����X^��3+�*. i� �XZ�vm��P�������`W�V�ɴS	G�]���L�!��u7'Z!�P{��C�J���4��{�(
آm�~C�(�o�o�gD�#9{�_�ݜ�4xeP?X+*�C�KɆ^���֘�#����˖b�K(v��9I�  X�Km��?OQ����&��,P���=���*�_.�g�����f��=Ρ!�����%��u9�K~nҋ�Q�o!q%��~��X���G"D��Rm�c';1��@��a�};)�U��ƥoЮ�I�P��n+4C[�$ ���(z�E���J=L��SY���g�Q���O�f��{�Xi�:���\�w�b�ȗ
�t�^U.�����߻^�rr����y� /T�Y�����:SR�4�T��j���N������y��u\�ߗLY�J����m��3�3Td	bdP�OY���Z	8OvP��2/&�>�-��V%p�,�d�q�-䧉S�%fy�/_Y�w�s�wU�$����<���Geņ;O�c3u SY�(S���jo���X�=��t��5	�&�Ψ�t1��`��3��6%_W��Q�����[��ֆ��C-����..lG���>�r[Q�	T�'�(doe�d�	�)�fiMh�iN�R+p�=I5SN#��y7&��3��^���z?�0�LE�w!���L�z����?�h��e�=����� ��B69�01����
��$IҠ��6K9fNIR9JO#�I�����:K[�V�-gz�c4����!>=�|.β�L�r��<~��k\��Q������?ᔁ��A���ѝ,�`�S�-��V3�?���n\���J "��vIc`���J����a@e�I����^�����,�L�b��X��}�g01��ڞ�N��|�����6��ԶE��.lg�Z�R��],�l��!'����mRW"]�E�yoI�(��I�7#;c�ky�N��
N9a�vr����'�<M쑂8pjd�|�vp�c�MXډ,�(;燜Y@P̗�ghED��N�L��W���
tUv+�e��J\:K8#r>(t��ʑ��d�O1���pEv�XB2'euWI�o���ӑ�]��A7T��g�i@��&� w�����M�%�	x�^��ڷ!����;ݣ �x��)uX�1�S�3�d�@� ׵��ݥ���X�w��,)�% *�ud���o�{;&�pi��nb=3��>/�rX�^��d�T�G�����hd``�'�����	��+��`;�Q渖���I�`;��gǑbRNB۝�AV������8�Z�k_{�p�od)l���r O�	^���U�ed�h��6�O3����2�o��ˆ�;�)m��ؼ��i��xHӨ�����!��}cxfT-�+`����Ĥ��Հ![�Y-E�I*{ERM�c4r����Mԃr��NJ�,nP�M�[�F�ܓ��o�Ny���EMjmsD�+�CJ����q��_���4hd��#g�b�d6�c�w�^��t�&ILm�u����4u5�EB:�)"P��x������a�`�t'��w),	:�c�0U�$1��b�#��AH��R(x����s"EQ(��3��w��",�{����ݜ>��7���'�%��$��.��q2�Z���~Wj�`?�J�1FdA�S)�,�����}�3bTh��祛��T	���#*���z����Uzt+iYU�3xs��A:>
�Q��8&<7�bQEi!��r����"�v�Z�1@h]`.ݍ���e��ɰ��D��nX����`!�'���='#]D50�^�	��r��1�Z�ٛ~L����i�o!�����X���&��w�7`kb��2p3j-��凇���|�W�q$_k2�3S�:dd���]Ѹ|�6���(h��0��T�w�Y ��	�(��O4�BG~�,w-w����mR��;�|gn��x�§��s[m��� t���- L3.�������a�x��P{VR������y�plcpo+M<dtʕd�����&�Y:v�/(#�YL����l�4f=\uL��0p|sX�^�TS4UKZ�E��4��$�~�*1����A
���1���#�5(�;m5����_z,���|����:�Z���z^O����N�b!/��C�u^i�-�ũkV����1�d��'�'5k��*��?�|�J,��o���ͻ ڮ��3�ҽ����a�=|¶Ƭa�n�]�@�T�	{�R֗����W7��suQե�c���V��׶�]���*�ߝpxÔ�O���sb�ѹ%K�[�T}��"���ʌa:`/�o��o��d����W�%Ͷs�v�C-Io!���X^��PL��2%���f�������G ]��E�5��/Aȑ���X&�]uo�_�y��Z�r4(^!���&R��;`%</eJ��*�+FȲ+gp����11��b���.'��CU���~���0ݽ�	B��ZM~2������Ey�E���� ���2��O��FK�H�U�<��sX}V�4X�/7G^��r����o�|6\J��g��~Lڮ=���n�G�߼(4g���(ᄔ���~1P��d/Q)��0d��q&!��:N����%o�?O/����\K��fv7��0�7*�2"vk���:����V���r��Y��"�gKq�W"�,��g���z�s�0EIMP�ԙ�ڷΠ�2�ʕ�!3�0�ߊp6���E�ɵ]�pl�sT|ɮ,��G��F�ϳ��<N�I�`���b,��C"��T0�K���|na�>{IG=}�\gڟ��G��^W1̹5D�[M� �F�z���r�+8���zrZ��߰�������%�r�K&=JR��a��G��e��c\9�k�5���������&�|IF}�:���ԫ�S�K]@�.��j�D��{��GVdEM���`vd��x�8h���##���g��E�7��	:�V��%$-G� ��=���+�4d�����nэu��_���z�
}���*/r!�T����z�6ӧ�E����ctU"��} 7U��&ؤ�A�:�z��L�AZϗ��U� t�vŃ���X��Im��t��#�Ou�AK�I��@���[��[�1�&H[�$�Hh��A��������T
6��lN�Z�nm4��
rؐ��H������������lS4����X?yӥ���3�C�*`9����k�~x��r�7�4Z�@YF3:v
���"��[���tn7J���"|ׁ��n���L��Pxi0ln�������JK�n��[��az��ۦ�@(���Wɛ5k�j@��dG%�����v�$��.Ύ�P1�v'�pfu$;�8Y�aM�ާ�c{�8e*����W�]��vy�79�#zW�L��k$�Ԝ��cV�d�ly���Rt̋%K:'ڀ���tKyI��?���$dU<<���ܚJ�Q��H
x�"�Ǳ~'ZI!���T���KWZ��O��T�<���3�%_�������i��{����5X��C`�-����ef��^�k=;�N��d��C>RoT���Qݢ�����p�Q;vI񰵤����>����;�r�������D�[|O�ը��=F]��|6o_�+u1��!X�g�cM먐���F��\�S~�Nr'�E�| jb�;<�2M��9�9;��bv�~�H��hux����iK��vj�T����d3Ҟ�y�6�sϦp�AaiT2�ݟ{�^��N�Ӈ��ރu.;�;��ca���ݶ|pW�yIR�����W\�h�}���L^^��f��ݿ5�U�����Fܠ�Xc��.�}`<j�n�mx/����BO1�[ͨ��}&}�G��I��Wcs�D���E�H��d���a5�^:a�
�Yh��ѵ�g�P&�dO@��+qnMRҼ�t��K�q�$������s"A`�BH�bw^�ugj�Y�LȬ��5�)V���)UK���p�e|����fH�WG��B��@>Ҭ�NF2\���
����MG)~+X�/��¾�IRKΘ}X����;_J7@�!L�b5)�%��c�âɁB��O��!V�B��'hn�<,���&g�<�d�KL��Π�?F.ٟl4e69��Y�c{�=�� ��l�l���A�����]�c����V�!RD{ώ��>��.��]aj�~�l�����cl����xV�%1h6��P�����
���`PE�k�χ�k+;�i�G��&3L�!%�ݰ�Z~�y.�f�>kRH#����%�@5�`���ҹ��(Vt(|.8��E��3�u��п\�<��'>zh��R.r��D�h�6J�/���-,��! �&�ozJ�E8����j-@БD]�����ѓM�PM&@��e��.����u�y�(_���9= ���9��N��uEᝣ�	�D���b?�I�0��}p��.�����	�2ҳ�ۘݦ��P!J�!R�����_"��	�R����O@fﺐG�x�-HuɫC�yf���� �=�S+��\4�*
��@��v#�0��A�ToT�P.���PODc�3o�x�1W߁-����(�Ϲ�<�n:ۛ
wb�)
��;�v��4����?���J~4a3`m��;��Ҧ\�?'�/D?Kh��;�&c�z�p2��b�5�ge� �(w{4=+�L�o�-O��������ceaT@�̫><K�].��s��5-#n�@�3�"�?(�������9`��϶�����o=eJж����wYP���R�?���&??s���R5��?h�� �ӣw�z/�*�v8�A���O^X6����.�w�xuzIk���{��<8����4�@r>`xWR𕦈���=���"�K[��~�ǆ�A��R�K��;�s���,�KX7���?,N"�,�3K�1���v{��JcѮ�Ū�غm�p(S�I�rJ�=G��m��M���q"���;;����E(1�G�d+G�6�.��v/�DE��Z�Djyk��
T�]z�X������_�z��E	��x5%o|^�!��}ō���tK ��SG�Vn,$.�D[E�(��C$��s/���V�U^��$K=�c;��JC�������5��to�T��se�?�舅(�� ؀�E���a,�|RE[+1@�R'�DZv^��E_�¤D��.QkX������u0��E��m%�ƏZ��ѐC
�YQ�&� �j��*_�i�3A0��:oa�9CZJ�l欥6� k��\q]O�I�+�?˷�)�R�Ƈ�kVmB���-�/��~��n�r��������|Ҵ��\�7�P؟�M��tD>��D[]!��ʔx�w2���@TƳ����W��������.EEo��V�-zB�Y(t����9�w�D�#�����[֢��j�N���&��\S`/6\�C��b͆Db!��%��7��#䬙��g��掬���/�,�H����e�PP ����
����ʣd�)k> �6�|���E����,�3��f�G�ޗ;;Q�3�|�(RU��S�l�eW��#��@)����_���1���S_:sђm>�3���{�8�̂ĹD��e~6:�q��Bq���WE�9�����J�(,����9�$�Kj��>���3Cv��0ij��FŌ�== K�Ή�"rU�@�n����#��$�R:�;�K��r��a$�ő��[AS:`52Ű]ߪ��r:�ox��^*F����>�*�Gg�q^�<"#�Xs�>�JR��-9_�g/�/����E����Dlx�e�Nx��s:��+���1a[���Y;6{����x#	�V�DÕ���Cͨw�G0���>�,t��ZCߤ�Y/�,�W����+ݿ��N�:o��u�]��v��������ŕ����T.����?�B��hNt	>s���@����v���$�|��Q�}��3�i��3�bÝC��r-0�bC���	�J�����S~u=r�!�p�:=���e�dc�M}�W7�Wf�:�>��Z$��S���
����n���[���A�;�@�E=b��E��Ir�%z����-��λ�(��ƉDqWh�+ʆ:�!2���A�U1UZ�H�Nx"��ws8�i�כ�����*?bz�͚$�]��Ibs�ol~�"��Fv�T�����:q�/����%��*�Z�^"nYQ���.?MyS{� �n�]�c���I�+ύ�����`?�@������LV����B�%6�qhӣ=x��f:u�p�����dX��� ��p3a�
7���3�g�(
T]�IK�D���l�n��]�qbJZ���7_�v�)=Y�A�thE9lz�܍��p�Χ�5(�A��8.�V�S��_W{��4����0O��x58�"��UR1�=EڇGA�	h*R/�7�Z|mݞ>}|������e�fJ��0w��V�zp��(jB��Q��h
C�a��j���� �hL�ci^L��lQ&N�G��΀�TT>;��D�8}�1'm}�0��q϶��k��J�'n��j%ډ�����*􃧅�[Kj��"<&��{�sH���f�n�Kq�a�/�P������)5�4C/:*h��<?s�U���<8xY�m�e�	/�8^ Y&���h5Okp�[�i�k�%l(�m��o��dl���n�/�Y�2P%qFJ�Dz`�1YZ1 G�t�m�5�.�[٥Pyd��J �~��K�G@-y��F�*lnXg�I���8e�o#
 F`>��@0�e��7x��e���/��6���������͋�9�	�dZ&Lb���q��:������������w���t�Zf�?2��ʥ���x�T@뤌&x町��m�F}r"D?4jB{_k���-
8��ܶw�١﬿�T�z�F�qK��$$#k0�I׮E�	�%����z�b��M+��vrpTLc�-幽��y���af��%c���@L]��3r �a�{'.tO̓C�>��:�.Ω���	X���IT�mV�WA\�t4��c��w	�� �[Ա�}	z(��t���D��b�A��<5���z%�_e�s�������u�0���5�o��Op��6g0�s�Mn���%�;҅{����6p��F��-S�=�dW�֡�cMگ�r�#4g�[��j/��V5�.8v�!�sM[�Ʒ����?�Z�P�2�ܱ�<j�\�:��pd��r�|�ρ����s	�\�W���e%8\�J���-�6�'����C�5��ǄV��c����:WWh۟�����ǳ��ʗ1_iq�!�۷�Z�l��cz�DUOǪ��˘M�>����.^��O��2���19�b��"�˷=��A$Xq��>����rK�W����7�R�^�������rw ��E>�<��'ł`��fVk|��^m������G��I_i��ӲUkʛ/� <!c�[�Z���u��<<3y�V�J��i�7(��|��zĕ��8>���=�~����>����w&R�~�n��^��)gp:��aAW0�~%�?M���c1�)��	�����k ���w%'�En�%�p� �b�N�[Ze���$� ,��]v����Y�p��Ӝ�s�%�z�f�9U`6#R�|?�����O��Dv.r}�澓��s�j��1��Ԉ�`�>����e�f��x�]m7~�gn1.�т�9������p����$�>t<���p�M�l�׷}��̌����3�𜠭$3�A���g��-���P�\Ǵw�*\Qӕ�Y�\I���h"?�۵2�	u�%���饈�f�	��0��߫#��n�؞� ����%��Ͻ�
ҞF�!d��֚���T�q�[��ʶ"[��q�r1����o�l���t�@>mhC�g3(6���Xn(�>X�=%;(��}u�B����<����d�kkHШ���`~���e@m���"}���9S�qܨ�Ӿ�0�_{���"�4�]U��q4��o�:���Ǐ��H�*����Jm^�{�mT��Y��e:@�ڏ?�&~�  ҷ�-}��kp$����wL��u��R���xV�a��$a�w�ɵۢ�dy���pi� �밍���n9
�����s��P��G����f&~�3RD��џ���c':�R:�`��
IAhܸq�	�ܢ����#{����߾�苳��W�RX�ح�>�����*2�&5���L Yi�;z#UL&o���� �M������(�n��*��wǰ����wR����	�X.�C}�iNik�/�Hj�x|���zq���+[4���@�����P.�kx�%�%���<�.�����}d:��c@�Ӑ.�}F���-��].��)m�<�g�^�ʕ:_���N1h�2���f�����z\���+\�ŌI�_TNqj�,���������u�BHr�IK��<a�Ɠ�u�v��;U~��T�y�v����%���hC��tX�U���b���ܨb$'�lKLH$�r��wF�#��'���j�t�gE��v�k��E�������!�9�ć_*�V��C�����a��BW�W��w�TZq���]�O�sJ�z���~RJ��n��K�ۤ-���z${ǅ5|�J��O�ϟV3��UV>#"�cV���T�P���Ӄ�-:xN�H�o!卵�縉���'/��O�hgnO�����x��ڵ��
P�.)a�(�#3kz;ǟ���R�ܗGHM���0�H�e�%J�fj�w`X�N���>��1i?1z촨p��O�nf.>;([�i�)�cl��ȇ������z�w�;4=j��������*�5��O��
�v$�%"��AY60����σ�����X.Q.k�6�e�2�|<�y0�N��Hg�~��)�����AHi�_ض�F��i�v��%�^��42�/�<�w��t�Um�j~�.�$�F�4⏛�	똌�k:̴T��娤������7A2���K�m�m�Uf�ŀS�����y�bt�+�l�͟��KE���	D��D���������SF8@����p��F�3�ţv@2���Mw��ٕgϛ���=��	�CNc5�;[�?��o?-����8ٱ���P�tT���vU��H:Gͅ��&�*���]i-�<�~N%�i��4vu"f����OJ?��N�n�.#Uaz+9H�ë&�c&)-��Y]��M����ˀ��3`^�Y��v:�h�)H�?Q�=,@C�� #��TD�vtP1SxoG}Iw��2�R��$�m����<���0C�A��ڲO lx�������*�q`J2�t�A���|5l��c��|��ͷ�/	��]U��'I�����}M�W8�������DD�0A�8)�h���,q�zA���R8���w��L����*7m�١G�����gӘ�k�Li�h0�{GԀ>}��'���u�[z��g�P���gl"�TA'�����\��A+�����ߣ�j���L�aI���b��t��W�jF�,����ɱ*���cQC�9V2͆A�G��{�6 � 3�zQ�2OL���F~7I7����,�j7��D�R
]z���6�숚"�4&�7��}�1�ε{��#SX�����m�1!���9#=ݪ��\�s��wg�)��*��F�WE?I���@���]�%[,�4Z g���7.�N0���e7r}9M��Q-
��M���;��9l��2ڹ'j:C*}��0$*TfnH��lF����/��̈̄ ����/S�8>�xf��w�ms�����k��&��b+ߥW�����-���WSG�X�c�*�B��m���Ǻ��%�$��-�����ynB���9�����7y)/�������Z>��G�T�D�i����T��m�Dn���8,��X%��Pw�wO�󗢆F��p�θ����BDM=r�u�����3,���w�������e�+�c��r�/|٠�yp�Q]Z�K�#g��D����/Jh��	RO��ݨ����g��F�,`͊�z7�]���&^x��#��nX�T!nI���kװ_�js �=,�&t�K��E�z�w~��!1��=j�'赉EP�#&�Ͼ�n����g`)F0��~�]C�'Y#$��R1���*4�(�+��R2R0i�_o|�3���c)x��Tl}-5�^�b87�(�3r�����]Q}QS�뗆s�G۱���΍���0����U�s%���k�8��P�@rO�S̴F<^)���*�f[	wJ$��#��8�@f�uH��KnIL�:����/r��ӷ�M�d����2��~c,{�?��V����X��X�X�v
�Jd)i��m�Il�n��b��}G
���3�q��_��X��ű|w���*�����:;M3��sUa��z�d����,�-R� �� C���.4�Ij�e@�-�Ɲ�:���)�e���dnjݕZ����F�hO8,?O4s!Ψ��������#�,e�O��1r���j�,U"y��8�k|�Wx,�*1�q�xA���L�3��)*��nQ�$�[�����$�0+�2�A���؋)P�v��˛�5$?�"�#�ƀ�����5�"���x�$_�r8@5��Q�yր?��)?�3TÝxD؞�>�a�K���u�P8���WG��H��
t(�Y�fz����C��p���L)d�2M���K�>fz3�^?xVB:�%�qy�[ښ��M06H��	#v�υ�����A3���Mw`�Df�@�.]�9�Hf��,�lG!G�gC�V�W4���^�K��^$]biߙ�P7���S�guhA���v�)�	�̮���͢�fm_���%@�j��w�;'Y��/�4��ђҘ	q�<��,n^�B;�����m8:������\t`ց*��e���?ȳ�W��,L�QS��q�PQ8���0�ׂ��`*z��������(��_�`�X����G�́��$WH��!�i(�-��64B�nfa���2�V���Ri�H@٭��*P�M�e�<|^
S�2���U[�07��i��':�ٸY/�UԜ�>#1gy���x6�T�*�_k�[������!��âԯ ��%�~XW.{k��"���=���ق9W�ۙ32�ٞ �BE�*�L�8Ͼ,�5���~LN.ZD���uk�;��I/p�l���x]q�J�]j=���S�_r-���x��� �1��J�G�3�y	7U
�꼬(p>,8@s�1�+�����CV�������؝4a��@l��Gkg���)E0а��w� �ku�-��H��@�f����B�	W�o�UFXR����7:���5>h�be�Yv�}�c�Í餸Fkc2�o!�UGo
�l���tD6�_�X����le�z{d��wC�j0�[��dE$�l���zΚH4��Ζ������g����d��Z��[�Q �G�p�Cw��ᅑ��Dp� 7~U���@�����]����7�SV������ZQ͕������Y���Tw_b�o�<�C���n���J���#�#4����(v�n-#����Z����]ʯxF��+�KR�!��bUn��v>�E��+�����IK��r�t���$�ܠwZ�$傔=P��Z�X�=�da�v��t�]��@�u`�K�)5"	XX (�پ�S-���Mk�5��Ao�N�^uQ��~��rt{�E�_��Iz-�
�����拷ix8v *�;S���v�keNp5L�y��7�:�Cޕ�qOVb*��6yp�KVӮ;�i�F�k�io4T|~�	%C_i0D�]5n��].�O+Ds��w �t��E��M&�@XuK�V�!���k�`l���T�2�GLv��4�e�MZ��B���q�=m��3\y�j��T�@�x��C:G5���80u�1ԍw
�mjn�C�>p΢B�!���s�:R?�{�0����x��m"�)�|�h!p�iN�^���i�(���pe�I��[� �P�7������5c����11�M�}j�>��ā ��n�#˰*(�Q����qW�*&�M�=�ڗ-xR'k��`2���U+�f >��`�I޴[l�*[�����»�+Q[UVtmhH��6n�7D�_Y���?�?w8И����p�{�D�O�<�TH�}��)�3�K��C� �. ��]h�á#��ץ�mԬ��22/v�ɏ�P�g�*>�_���g��4_w?��I�f����v�<�Y6Q[Y}&�o6z7���&���ekS�O�m��qI���Q�D7e������xUK\ q��F?���ʗ^�iFP:��pc	c8s���t6)e��r�X`��Na!���延�$igJp���*F/���? �)�O�����=g���{���ެ��ɺ��O��A�W��;b(��]_=���Lt}4�/���$����R�x\@��(b.6���D#���}��'M.�n���k�Fjgg����Tj:�~C]$I��<�(˅�DP�~?�(��"���ޡ��q8=�o����t������ع��w�����l>�~�� �Y�;��3�8��?q��[��{� �4@U�^+2Hy��S�3FM�2����2C���ɶ�o�S�v���dH�H�1='�k�
V	Ֆ��d7'6d��xn�v�L��(���q��� ��N����⩋����س��:���I��m�j��f���
�<t�P������70�—�FH�b=Ԉ��ʍ<���'[[��Ӫ�-B_ϳ�� ���3[oM��g5��0?��+~;mpr�`�c�c�s�Fs�G&'%�?�-އ0��m�O=M�T-V�&ߊ�I���R䦆�;#�\����F��ω1?���=��=���Ζ�Ӳ�Fɦ=Vn��S�*�x��tA��U�+�k��_����c��vJ|��rֆ,��<�)y�=�'�oj)�Ydr:|��M��q�� 5H����Z��s ��`#����wY�%�ؙ�Q��hKa�R�ۂ?d�������W���f�p+i�2�p�EE�����-ٍjB:�Q�0�!��^9�:��p�W���C�D��#m�w-Ǚ$�Tq���=����#+4�O�c�B��?�A����?���Y�,�6��a
5lG8��5��)"���x#��:>�&���\��R����pr��������4�V��c�3�&�W�۔}�	6Pgf='������ <�?���9�2�h�­�L�^��TQQ� 0��i���\?�S�j��-w�:�LV�O�R9�d��p��jo������:�e�y��h
>��typ�u+"7-����b�Gj�,����-�ʩ]�iäԒG&N7�����1����XAY�Nb�*]�����1���Ze��+����#������1t��E-�/P��8��E2��O������c�!�a5�mE���O^*.�9_YJp�MT���I0YmQ�/��怒����uą7oZW��ۆ�~�-g=5��1;17[o�fgtɴ�n�X���Ŧ:�=SVN���D����h�A�*W-x����m�E�#y-��k781-\ҋ��� L�|J�L�}�n���|I.�ba:QB�Qf��$���L�]�d�fx�û��e�{ْ:.9����L��v6�ϵ��,F2���[�+؄��
P�xG��a���[y
!<'d(��$��B/��p��Z�z��!���`��n�K�B%�I��|��sDD0��,�F�S��L/֒��o��ט=ͥeo~���#F�zؾ��p6��Z	f�>��N�E���7Yϩ7;2��Ac8^Ss9���kh �}��^G�j~L��|��-�z��4�ӎ�sABԕ�W�8��H�Z�3�{$v�X�o�����G�[�ѽڠ�r%�Ȼd�J��}Ԭ���$��A��N�?F�ՑA.5G�3�H��0>�������J�k��D�G���N�(�x�6 ���x�B��a` \c03e�����_�L��c,����I =�����g��|���ه���N�u��Z4ӝ�+*��}Y>�[$�=d�^ M8�ނ�kL�>�/ׄ���eÀw�c���ת�,�ӑ=ً����n��������T;��yF��٫e��ܥZ�z�`�����?.0��P�b��{�?�k��KK��b�oB��\��&���7�9�'/%u��s��1���|^�!���`�]ʯX�SEc��������I�n�C�?�Z�L�`�u�S=��:σ�*�6ݙ������ௗ�y����{$��!.�x��$�%A��3D^L��N�6*r�-���Ps����
�%�h�qU=p�<+�Z��X��2�6r�G�fl8ɹ�nCX���68\�w'��O�D����EZ���A=;~_	挕�����"���ó�7��e�eI�^_̂�?���}M���G��nLy��GM�ДFT��ǿ�)Y[Cw5���	�/����d<L�o(�� H��ݯ
ftZcj���}lZo&��)�c��zW���)Ҟ	:���+S%�W�Z������2A�s��{s˟ɑ�A'[�.�S,"dN�7͞�j��唐��P��H�Q��S�m�2�w�PC��_��D=���%m/�l�?���^/a,�'I����+ecќ�#<M���"��'w�$��%yqZ�rZp�$3��M���O���́O9��*�"�l�7,aV�,��=�u��m�}���58�^�(���Y	%1\`���?dH��i�߬9>�9�9��_fW�I�#(S�I]%��� ր�(��(�H��ڇSB=��e�y�s��y��V
woڪ��"��HQ�c�V�f'��H��I]z���پ�����6������;��"Y5�����"e��:ɡ��8d�w���7koρ�8#z��y.���?c��X�)B�5Ozv��*��{N�'���܊9�T�W��c�����J������� ][Tt�cHE�t-A��-��N� ;�au|��w���g��v%#Qn/r'1���ޒ���\�����;�{ L���X������F��?̉�Mkc��_����|��м_2M�ý�:
ńF�n+�b5�%�^a������(x�VJBTG��%�%\#�0�~��J��
r�*����P��O]�ӛJ��>��.<�e��f�`H���Tu�5G��t1�J��/�%^�Pބ�+C��o
��̕�;����R9B\�_c2�9�R���[��ku��VT$%��Y�~$�L��}�{�SOi�Q� Qc�A��E/A�\1u��4��{+`	��O5����IHtM�#@�LH���)���jw����CU�Ĺ�����x�h���`�����p�r�@��L�n��/�`����vnc�b��N<���E�8�"wG��^�T)Fh��I���!��Kr�Ng?e��oL���J���d��6 �p����>gU��6z ��$/���~8DtQ^gZ`X'�^�dm�G�اc�
o� �"6��I�̼ј��(�=Up����qz�"�03c�����.�+|8�ͫ���@8	>a��>�����i�s�U���J;߬�~��Ɗc�����|'@4��6S��/�g�cݗ��x`��I������C���Z�i?*tRf�	�X��>p�{�g�}Xy��CX����9ȟ/5��ߏ�
Q�Y�v���,]�~6�[����@�[8�t԰�l�a~�"{���7g�.�>��2`�N"��v������2�+Ȇ����̋6�!�Y1u��f�%Y�]�4����ǚф���׾���B�P�+l������$�,`Sqs�;�)j	d��,&�D�`
�Dh�p78��K�b�a�����lIn6$�GD�py�'I�b6:�����g�@���k�7��{(�Yq�m(j �������`�U���(=���a��_���<��q�ԷQF��}��]Ƃ��|`�s|&F��'0��ucL }��'�����$�R�������ߪҽU�����!$	����ˮ!�A����;�{i;PK8z�pK��I���FvYI�L$a����܃���"˫��3+�~b`�(qo����x�A�^�"w%��5��c��+᣸��  4l��~=6*ݶ���|G0YS ��wS}��M�(X`�7s�1�M6agRW�r�td��C�y[�Y�:@y$��,;��}����ߋ�S����z�	�ʌ�oZ؍%;X���ŉX�]:��I+:��?�xNU6_��t�7�ʵ���#w���g"�,47��r�B�ј"w�\m��D�����'gh����^�ЊV{�O�\y����py����/����}/j�ͷ���	���m׉>�ō#�vlG�i0bvJ2������(9���(!�����C����w=�����x-�4�e>0?���o�#!�Pl/i~�m'u@'����^���'j��ߺ��tT�@�Wk��|�cax�ɑ������}��2	Ȥ�AmҒ�t'�v�*�ط�/4@g4�l��g.�#e�L�R?���ߎ��z�0ͼ�ع^:�d��"H��r�l� �u��I����f���m�=˭$�o�����b��8�޾c+����W8[�P���ĥA�~��!�Ca�+K#u9�!}��̾Դ�����i�����N�Nމ�:��$;l�eq���<�Ąv_eV��*ZU�`{CO�le�3�Q̈́���}K�`���V��W���(:��\!��#۔�B�<���Ӣ6=t�2��_���i/��k�~<���2;{J�~���.�%X'=qR����B�F�W� h2�o����>O�-�j�Ŋ߶����E�[���F�~Q��s9���屸�^����Y�6�>�����؁H0F�^r��A����� �����h�و<�p|�E�yz���+c�*�����c���w+",�u�Qs�IKx�`�'1]���B5�qBxcV+�B$�������̅����/������� W�8A�Y��"��NZ�s��G�Am�i�v���(�0P���E�΋�lq��=H))���Z6Âμ�������$h.���q�\�%�׊X �
����Xǟ��T�j���)�c����'��n[(Sj�,Xe�2�C��
]�8
sH�KBx�NX��.sʭ�1wFT�s�����U�?��+!&������l�اт������͊��ʚ�/ #;��Y~a��ðGĸ�/j~b���$�?���w#�+Tן�>l�&�T������ �J�WOl���	D�ٶ:U���~K�_�EM"X7c��Y)��D���(�T�^�c_��)�FU�f����4�Y�ktHA��3C>��������bI��]NR�z����F2iW�%�^�%例�`K�ÿ9g������-_�9;��jd�� 1i��2���v�*q��PP�R[kw6��j��r	��K�<�2�"�~���Ԩ������[��kg% }�t��p�P���o���Ř>qK~k�V�v7���aJ�v�G��������ZI�V�Ⱦ�Q/�{y��ET�TJ�6��ܡ� ���ef�E�1/������r�|��=f�΂��d+�!��n���G�?.B^1�:Z}2 ���v8��a�Z��yX�
;b�88��>��TͲ��$�`7�[?=�������	�3�|�V�����uU�jP�W�T� �CRPX�ll�@���������Y]	XZW*��׻��)Pf�� ������
��KP���Մ��C}�Q�p��%#���R�"l��ԧ�f���Z���h�j��ș A3!X)|O:�;ȷ��;15B'�H�$GOC��������2���['%�An�����>J��&�-����$�+g�mbe�Qd/�B=���EK����	�I�&���6iJ[e1 �=�k�q�jZy:��� �ŕj5k��ݚ�xV�-8jQd"� +�f��4�m7iח�LB���\Pz�C��V(��kO^��6'2���b �)�=H��ҕ���0P��Y��##�~Z@��d=ifL}w��j�����VY�v2�����&9$�_d̅7��Wjj"��SAd�( .W��$����d�m�J
g�a��>��ں'���(|k���G&?�v��VO&�؆گFVă�O�	���:6�o�G�5��Je�ǨO]��CH��'���@��v/�c��V"�p��b���s�6����7���I？y}�(f!q��Rx��#n�Z�s�尪���A�畄��F��6��.���}_�*�2�Z�K�����4�
*�K����<+��l�r"�i΍�"ͪՀ��ۀ#���#���1�k
P]i�ͅB���ٷm��F"���/0�Tg�̼�oOxR8yR������ǙF�����sc�t���4K_���ɩ�V~cW)�N�e�@����&�j��E�~��O���C�c[�ZJ9���	�p�m�4�� �l7r\O�����W�8��Yf�M0J&���̾�=��G)��W A��/YMs��=Xk�4���U8,(/��?��͡�9Ǎ$�ф�SM��Kν:�mAp�|��v�[r�����yx�!A��		��66
Σ�N��-�	��9�տ�C��<~qeH*����B�
��3��wȆ�7ot�}�����F	�0����e���/���C�@^�uD����i��V�s�a*X2�L.���"�D�Tlb��C�o�r����V��\>#!bk3hU�+��s��3X�$�z�b%ŭ�3["8d��m��ER�j�d�ϲ~��(�/�ˬ��3w�v��R���[(��<-w�1z�QoT̡��}J�e�m���gLb��f�i7r-�8���t�`4��R�\���MV��
�gW�>�Uz��4��a�+�#�œ�� л2�7 ~�f�K�����Hi/z
�}N�o�JI"z�}�\��\�|@+O��c]�|gR�U�h� �,]т]J��dy�s��l�u96P��vi�yU�yS_b�]��ٸ"k�4A���Hn�rP��]�C��؄�I�ٓ�̓~S�v/Vu@iD��7d4 �ie3�I��� ��Ew��1�	c�d~�B�4P��q� ��0B�T�A��^�O�\k���:��aG����RĆ�RN��h�QD����L ��]	���-��M�7��aS�4�`yw}��ɓf�-&��O�����q�z�'y�g���G��ӈ42���D��Öf��O�S-��%~�j'�
�/�SJ�`ME� ��g9��ȦRa�0��r}	�8��qK�Q4�����J�&B��\��p[&q(\B�E+�5j�g��s��S��b\C��rW�������y�9G�u�&������>����(͕`�̇핾b�������p甼�A_iI���M!�2����d	���a����/ʯ�¹�����	�-�@4��FL�[�\��}�= �p3����Ȣ�&��­Q���r��[�S��S&p�O�%q�1�8rlLI�9m �CD�,1��$�����'u�E^O���w��HJ��Պ/�*��������X��,��N4�C*���F�<��;�oC�j��3,�� �-p����uU>H�
�KS0u>�}]�`��oR��z��};ܙ�8q�є�vd��+�݊���eU�T���	S����w��C�&Y��$'�O]X���x��@�!�*�9�}b��i�;�,
n�i�HH�����yS�Y�r��VEbچPZ�/�4^lۡæg=��\�~)�}Hcx���U�m��:�P-Ձ���k���:=c �"������E@c�a������}?nG�7��K��J�ҫT�d(}��;���ʊ�Z��x I����[����c,��R�$Pڬ#p4F�XL[;Zm 3=Cm�H�q��_���W(�	q���*�n�� Z#��R9�'*:��U��r>�6�{o��������k�1$���i����-�}�d��82"c���Dp�Zo䵫�P��<��RLӦ9{��1��Kl6�v$df��I¢�S�p��i7�=;P@)_�����oReK�.ؽ
Q��
��w��q듧���v@�O�|���2�Iޜ3!�7`����C1�>M8�L�nګg�Q���bԴ�@���v���f!s9Hs� �."�������H$��P��mR
..�|��=PX�*7Tcr/=��Q��	\��	��rX�,��������
��fr��Xaޛ������l8ΖO�k$V����.���1�!)@6�馅?Dq��\ET�-�@t����B��_���?r��0|�1mS���b�<&Z���?%�4��98WY�,��u�z��}�Z�CXX�--���wztT�{���jܺ��2Gj�z8�&����y���oC�t-\݆��|�6���bX$�7 $�Df���5��Lc��H��ԍ�~⻬{EG�os��4����la�'uX�F\kr��.x�q+�M��ޟ�zb�O(�8�}@�1�@o�l��ȤH�3���1��Y&���Q���(B�f/�Gko�͡��J�yzV������z����̨r���T��Ͱ!8+�6I����5⁷A��:�0M�Ǟe��,`%��w��~�	��Ĩ7邓�:*�c�&��-�\[����71Tcby��Wܕ�r���������'�4jNa��)e{:�	��/��ډ��s5lX�ܴ�XW�t�+(�TR �*�}<�GTZ��Kh�@�!g���I8�4�&ss�Ry���D�X�����n8��7��l�ˍ���:��`KyMmƂ!�Z"Jo�K���?�q��\�u��z�2�d���h�]��5$��[X�N�]�8���C~�D0l{��µ���i@	j^]k���8�݀���\P��	}��C$)Mr�|�#{�b�Y޲�g4����A��������-1�����3�$�>@7	%����L�/���`��ʊ��V�vIo�VmlAu��$�q�8h�+���]��9�z���yD�`��]�XB�W�����p�����^�ҵ}ĵXY��O"9SV�,K�Sao��
�K�K	~ʴ��s-ͭ[n��51�2�*P���;*
�zw^'�?J��PE,.m�ȗ�˾��V���O�5"d����j��9�>lEU�o��l�#a`*enx�X�������/�����;���T�E����O�q�xʠu�	���fljs�����1Cg�ZҶ�"Gc2�$p��
+�0��$��7D�����X�}ϝ�6g�)uc�H^��z�0�9X'lb��%H1�,Ee�b�?�T�U���=�B\㎜ǝ�%]%4�k��a��v �괫��'y)j.�K���	�&���5IǾ3����V��L
���Q��!ܮ`�NE�7�� 3!rY{/�}��J�B-���,�N�J.?�N~��~�%����bK�􌂊W@Z�бe��T_ǡ�G'�M��!���W	|�XR�f-�Q���EcKh(ּvT��n�G�B�s�U�g@��Y� Do�r���
�d���E�q���j+(Ǘ���r�q�6�J�7~*8|VG��q>��ïz�8��pR�?��Z@�$�7�Y`G�`�1@G�6U������z���<��C�$5���U����fT���~̯W6r\p�0��vp�G��6	(gO�Z$ږT
�&(�.h	�ـ4�dq5�nHӑT �zJ�#���%����oƧ�aw��*�Vt�2�^�*qi�/�ٶZ(����&��\�ԩ�|�:���@L���(y8m��$�N� %6n0�C{y��B?�O=�*Q˪��tV���G��^�	����D�c@*��zPr�~�yh�p���_�M{�2���Zl8�YU��i):�Q���v��'V�<5O�:a����@�Xz��34��t#�3�Z���P��Lˎ�\Ţ�Unu�<�����������	d�W�ryV��Hx��-�4��5+�T8�m��E�;��� "X�l�F���.�(d�xhKo�MC'zge�QÉ�"�-}R�>nY��$��#i�o��x������L�Hc��^�M2u��,�u��tX�#���xjg��U/!B�I3�~�=G
ǚ	H+��,�����qlkx-	���۪mg̻���=�Dz��T5r|=X�΃�dBF����h�΀�E( ^��3PA���e���}U&�9�w�jsUA<(.�rF�P޾L�o]H�ssCJ�l���؞��p�PE(O��ϋ�]?&c�+^�$�y�=N���+���Q�
�g&m�������@\�O)B�"�,R�M��@'f��S���s?�c�uh>E�B�$J�r�Fx�S�]�00L��+��%��J1cR�]?�{���_U��e�L%F�Q�;ǼX�F��{��_��4�mAB��#jM�w�ŕc�*L&?���t��^�>�Y<oW�}ð�͚�5�i�	�������Ù�yB?��!�J��cl�v�t��7��r��a�R��)��1�˔�M��b "��S��8~��-O�&�C=��l�ڇ.!�	��L���o�kV��
*$�]+>��/�!�>ؐ�a��lYD��FF��6�-!&�kb2֓�^��)�x�	`=4���1[;i~㺗1'Q�׎#�WN��wRʂ���w�J��LctB�4��|��e��C|a{x���'�}���))V�OƎթ�!�;��&����/�):�m�Az�Tf]�b{N귻N,�� O�">Ϣk�{{[7͂���"/p�>r�+O�*U1^w���Y�ع��c��SY���4ӄ9A��&^��%EʺB(�v�
��B��.��A���Z~�LA�Ϩ���YK��Sً���C>�nx����SN���՝�j�Jp��L��P��_�H0V�8;�\)�U�m��ß��Ћ7j��
��$eWv!oҎ�'7����+?Y{����^��ۿ�=A�Y�H�ӗr��ݑ���j^���9��� 1���\5Ȇ���JT*�Lc���,g �w��l��}{E�ҽ_�H��K>�p��f8R�ƞ
��#���C���r`�n�9��l�N���dSMo޼�e�]�i�)#���Y*���nN�5����}�)E*֟w�8)�V�L���� ]p$;)B��H��h�J�f�8~�#h̅��x3k�(�a��v4�i�u+�����|t�$=(�ҙ_=۽J��vW��*��T�2V���tJ�ʩS'Z^��v�Y��uH���1��D�X�GF���DX);>�ޘ~��:�ɨ��ey�a�R4C�
e�o�|�?��(+����>�߼ܪ�s,��Z���t���N��,���>)[;6_�ݮ���B'��*�:��?���|u@p�h=Sn~z\-q�q�{�egV)��;�]0H�ͷvI�-�|Г9�x�{\��^"��A?��X�0�=㋇����8 �Jd�����M�����Y���s)����L�;�ݱ��{�"�I��
8®�j�1B�y�	��*T����I��!���X�� �Z^���+���M�������<\�v:N��/� u����a�?���XTáD�L�>��}�r�Q��G����A:"{u��L�/��������$��*�Q4�����A��h U�^|XCc� H1�'C��T�e������^̀�l4�}��3��e�ְ@�}	����b���͊�\ -k�0i��=hM���a�R��*��v`��
���W|���VgYg�[��,���q�/�,���C�B�[�Yܰ;�1T�ƠP_�'EQRL�^�t�̖8�@[ +/'�J�Ȳ����9��@ �z(>-j���}_�$��I#}�B�L�8?ո��SG��6ۉn����y�0�Yq������zy��T�ȍ����Ic�N'J��T0���:���^�v��4p��𒗺l $#9s�a�vt��������y΅���Ÿ������v�>��J~ܧ��#4�����~1�Z�6EFZa�UH��LSTA���C�b��ӿ�N�-�qƩ�{���C������-�������j�l�M�T0���
'�r�&�n�	�B��i��Z���@�>MEI�^��p��_G"��w>7�*�7�qm,?��qEy=c���#�mS��t&�fޓ窮�y9J��5vލD�=���[��!�� 7u��"_�[��L��~�q�aU2P�Mm�����:&�:�eg�;��*0
�N��\+�۴L��[�8?)7�ެ�V�=��dh��4��6"���u�u�4��o �]ac�=�B9���6ѥ���؏\�<ֈ����u2)����T)�)��a�JS&�	c�vw�3��	U�1b���U����&C6�h� ���>AɎ��	��P�̺4��V���K�ߋ�ח�_��ڮ ���*c��Bᴀ�I���&l�{@�\�:O�RpN�}� ����.k)X2���$���8�s�)��r]QC8���\��g��]�ݵA[ ����%�J�xD�����(����^աkX���=A��\>`�p�H���P�ˆ-��n�3T^N��Dι���V�H�O��;S�y��4�#���Fo���.� ƴ�2�S�U��7p��ݺ��Ҧ(�" c��̀]����\*?K*�z���l6��޸���Y�+����@�n�)2R��XϞ�D��h��RiQ��)��Vm� ���jJ�:��o:�؜�)Pf@�A�@`�l%��;���\T�	�]�rAs?��J�U3�g�槏U��X���p�U�
Nt�BӬ?�dAe�S�_��𤊝�
͇�I !����))�*��O��
_%Z]8��3���Ew�+��	���8%X���8�	ht'���5^����Ѻ�ۋ�=eZ���~��MVI ���Z��y�%O��5�l��~<6�E&=q�����1=��fH��Ȝ������
������Ղ��@���7ނ�͋�D�n&@LL&�u�وBt9.�mm~!��1lU�l#3�ו���_x��Ha����U�7�ĦN��UI�X�W��=�,�ʯ�ʣB*�N�`,�
}8���m�0�ր���T�y����o���6�F�]�i2�I��]��U��O�ڶ �z쨳2���'�̠���C�b\,o:eP��<���@'�l��/���2���ǵ�^�gk�tdD;�T���+�Kv\���_��5x��v�	��G�+�J�/)�۫�seG�(�b����r���뱝�J9����0h�ɶH��j�G}�~T�t�cyM()��ϕa�� .
�d}�.�7f���z�=��c��F�N+ɺ0��<����fмD\[\d����~�[k���X��%1���dЖA���DZ=�x����7�iG,k@����K ���X���1��4�dX� g���^�+܊�K�'u�8u�Y]kL�V�t��CF�R��\��u�^zND6��\Ed$ H�2�E���29'���@�����)�&��k��ؤ#ӗ�n김��z�Q�-�e�w|9����'1v���[������ah=�^�w�oM��eP�(1�.C���"��;�hs8TU��d�F6K��ϋop�$R��ţqR�ǡ�]<~��p�w�ZVY��6�`Ŏ���/��۶�r�v��@�d��&;A۹��13�(}`�����xo������"��,
�!%Ї B�#�G��n�j����`��XΌ�)׿���嵳@�.K����?����;�p��AsF���d	�$��_����^��J�$�&/�D�z�g���A匠���5	�\���4�/����wwB�L�B�Ól���B��w��o4�EL� �ڱm�C����|��j��6�
s�k\�7w�4H� Rs'1�D�V��~�D =�������3�*0����"��<��NLF6�@�Y��s���1S�Z���U�v��	����>���$M5b�9�MǤ&6
�����O���C���3]���NFB~�cz��p��ƚ���H������������N�X��2-�Of~}��gLw��Cn�?y
�t�ݦ�׻��mc��j���\C�'oz	��o��1]]s�D�
�Y.h��[0<�x��s�
�ΊҼ�Ro���:�>��d���ȜꈃR���� W?N��*\֡���/�P�T�=��J��F.y��5���j?&�'U�Z��P:y�_�0���b�{�� <rŒ�O��[��`&�����t���5f/��in(�'�+��_ͦ'�v���mr�6�ю��C׫	��i(�Z?�Y9J���$��dRLhȒ�����y�
	W�SF�j���T����0��yd���)'E.�D��9�rN��V	|��F@��t��f5 Y�&ߓ��)<��H����lj�7�;u*h�"^3�T�p�����*s*�j7x�9��h��;�N�a���&�������5GWSdtF':��C�gŽ�C-�ku��h��[(�$Y���.-�+��c�j��'�+F,�h�2�&5�#�j�s����	���*�ZO,�g��"�8�����p���\	J���BB��+<D����Ed���dy^�!�$�-R��ʁ%�R���C@l�d�ts�˃p�^���,K�a'�2���;z� [ԙ�u7]�HU�J���� rl{8⎹W�:z���pD'�N���V]��6�^����4��Ͷw	���c]�8��Fy���4"�Ͻ�3�9NL���5�j�꨹ԕ����2�_�$�\��Sh�*�#@JM�Ȍ6
H��=+#��Q
{�	����&NL-I`��B��e��)*mf�5~:b�$���g?���N�/��VN���v͸C�YN�F�����3��G\�o�uv\$YQgé�G��k�И*a�cp��%�v
x*���T��t��CM�+��_�c]y�]�|4�xz���K�uz�61��$�{��Ō��=�Hd�j�c`�Nk�`���Nv����}䗭��%��VqzY��v��f�~�gL'���D�v	�~�&�>uZ�5nѯVw���. H �Q���4`L�4�ղ���A=�|�����j�w/�=��J�8�+	�H1_����	�o#qc4�X3�qŗ�V6��QSH<,����{m0#@z�&�p7�0@B����~F��q#T_j��9�Q��E���
��������S�8�_��4��L� |h/`7Kvd(>jQ���.lfl�̥_�+_�I�F��e�* ��YO�, �*�FJ�C�t��[jX�/	Yð9{|�:++6Y�f�n�C`����J�;L�,�J�%�Z���PI
kP&f�ܾ�l��5
kk@,s{V��H�a&��+銑F�h���.8�=��������xqP��z���%�[�7\ە�j���э<�2!v����-�)5҆�|��������?�:��© ��J4Rde�R�n��ۜ��f̯�����V%s�J*3R0�v��>�+7h�n��Ϫ4��0��XN~���ֲ�?踭�<S��L,�x��4��V4��;��Z(���M����ο ��+�9rt���gF��\�M��x����)�10P�Vvw���/�"]ި0�d�:6:�r��BZJﰕ��ƀ^ʳO�ސ�b:����C�
%�.,���4�d�z�j�\������џ�3j�E�)'H�g���;�"$��Q��AX��L����6�<���b�}P4��Џc���@q6K��� �ǡ@���yI���-?���9�t������ixP9�b ���O�!��1w���DP�Zv1�����؁G���E(=�<8�@-��J��?�Ը[��RU���/��6flK�K�9wN��;`����;�LVeep�'���&��:C�����6�����]�}����Q��8��u�9u�膸��X	,mq��û��\���?�|��S0��m�#r�E׭x��Y�t��x6�D�"��ՈYQ��S8dw����O��aA���ߙ�a��Z��4��n��
xe�)2�0Qpf3^u(?�&�{��C��o����|=1鷒&+�Ǧ�U�/x���}�2O���z��'���n �z/������eN0>�	p"t�ޕqh�����ƴ.sw_%�6�Չ{���l9bH��~ݩ�z��/��!Cj�e�D �i{�ޫ���#	��v���U�q���i�s�V����Z�	��mf5O]S�5��]�8��o!��X���+��$��0a���`Q_����դ�,w����&���S��ޕU�����o�I�M
Y��&EP��w��]$)h|H��Zƙ�΍�8��+�p��#5��Z;�i�|Zig8T3��wulmt�NK㎣8>�FFl[�-�og��ޫ�âV�&���t���a�k�8��e� �)%��M�p�P9��$c]�T��x���!(�~�q �6�X?�[v��^	�g���\(����tq!���f�J�L�g��_�?��N���rO^Q8*������ּ��*1�i�������#�<r�	.8
O>%dm乧��~�։��n	�F)�7�-�z�i�MܣF'�4>�����`V*X�U��Ϋ�s?1"I�N�W����Z? ��n��/1��Pm�nriº�:l����3]��|ᨘMd�-��*�ײ݂��x�>
2�dݒ�4���
�il��JB{�)-@W��)+z5�'�[<��%�?�L�#��j���Fm�,�m<B�k�����ˀ�y�Q�$w�8��X���e8�����s�|��>� ���l����Ѵ�J��	e������j��~��\��l�g��/��Ⱄ�[T����Z[J�6(�E��%�{���]�w���q�`�g7��s�$&D�V�h+r�����Ww[����K�k�� Q�c��s�f��x[_4Fr���ӳZ�}�41��ֱ�Φo�N�k��e_�;|�7Yo�Q'�%������I\�ȋ(l�=�Q��o���x��|��MPYh�&�V��g��Y}7&��5�h��3۳	��J�_�*t�ZC��:K��\
�&/���ϗ2$�##J�1��d#�E���]�c1��mi�T� �v��Q���S�}/���pj3pQ��Ȱ��i�Bq�:��P�]>M��7{�y�8.}+�Eb#�'�MY�ha�p���y��v�_��s�j!E�j�U�.?��>�XRr�_�[v&9ي�9jݧyh7cB��l�-z�1#����S�+M�9$�2�ɠ\4�qZ��4�*��6o9s�_l7wx�q���aĳp�Ƣ�G���9 ΍H�(c�_oD:��h&P��:wJ�,����Ol;�8�o�pal-�;6Y���A���f��4:c��`�g���+v�)�Y<��Hn�j/oB���\���E�s��RBި+��KT�~ө[��Z�.H�����2��ҭ�L��)�gt����]_Igp�\��Gt]�Q$�N����9�$��:/��'��tQ�u���@�*g)1s;'����=���ʀɜW������
�^"�L�{����]��b�k���4�+\���p=b�h��v����G��T?��.�|�/�?���Qr�R���؄ P@�O�o�K�@B�����u����i��G�n�
&j��d��:zկ�%/*w�@�Y�0���ަ�H��JC��(;�JO���5��?3���S W�J~�Q����:���3GZ 5��cg͝foA+��:mH�I�a���M��P��o�TqUɨ�����H+ސ�{�)�0��HH�>��\�@�_V����|��q�Ur�������g#�}M�����ni?�%;
�ݣAY����Bd�K����hXۦ���-��h6�V��;L܌=s��P�tZ�W�5���~Y�2��i3mA�V��˚P��0���*�a����e��B43���T��8��ѠoG"e˟��y1���AȔ�sFgv�?z,���N#�TgM��:��IH�:V�KBT>m�w���V"���;VӋ?���U��k��|��K�l�dԈ.0+Y�͊�D���F��1��b����vO��N��mh@E�
����x����!C�����v{zY��{�@An^H�fI���ƣ�g����AG����߿'��@���	� v�m���3�X4h7X�u���T����%k3����ib�tF����1�8'lu��H���!H �l��w��ń��J��
���!bkn�g��	3R�Rxh�.���?�^�VF0�X�J�d�Fqًր�R��Č,r��[XX�c��i6��,O=2����1�E�~�5A��6,��52���SY,� ��+�솅�پ����K�!��vȞpn��o����b9��qk���Aa�icAq�кJ��&�V�N��≘kAz����>�r �����tjj ��#1z�%�-&}C�%�ݣ�Yd��BD�/�	�^iX��L㒵tk�u���"�)��)�t���r��M,��o�ȉ ��sf�Z��,b~M�-�u~Nz�fH�\#Ӏ��_=�L�5g�PI�L����#e��Q��,���#�ag1��ܞ��W�Q�i��]E9�_��F��� "ԓ����zӁ��O�ϼtw��U���>�]�0�!)�q����c�*ƒ������@��~չ��.��V�lϱ`B��,P% 4M
���o Ry_wK��lң����.y�� �B��:�ظ�`�l}�r�E8[|����O)�,�p��ҡwO����ց�kX��)���M�)��i�u��Wز��T�0ǒ �)�u��]��{Y��AYz�Y��a��Xo�)��D����"V�i��p�K�����q�ˡp��@�TG��t�� �ys��h�H�Y�M����m�4v�b*��Пpv�N�&Ua������Y:B�J���{��kCU����Ui��F:
@-�q�1��b�gn��o���_o����w�d��S�B��GrU�e����&�M�[:B��x�wh�&��,,V9���cx�SC.H�=�a��7� 
�q�p��rw���dK�l+�Ǹ�O�U\����cE@^u9��,UD�������Z5��s��P�y >��3\��Ek���`�s3�X�����s�k/^�*C���04��fa����_��^a��B�`�d�� J���jR�eB1o�����j+���2�P��ɮ@x�������d�Ҏ�s�{8�˙ ��4�M]��ů���;N�3+�m��Ax%RG�:�/��3�e�#{�OT�w���g���]ݘDi���E�|F#���v�ZR�@>n��y����ŉPo�M�8Z�!K����BL��S�Hr����Q.�q�H�vQ��#�il����ᓢr����U�7Ex��)���0�dA@J��1$����Xv��������իJn�Q�u'�O�yI�<���R��S��5��Bya�0=T+Uk��'1Hyh�����8דG�
�Ow��'�! 6[��C�xQ�t��M(�|���:oO�f�d�e��*�TP��8<��^�����ǲ�MZɧ+�����1���g8VBn�������3�W�Xx�2ƨ��N� t$�ELo9V�` oKF�H�k���#��I}b��B��1��f�db�P��A��o)��6��X��_X���0�XGXp6�N�]��4��ˍ�}�����<��)i,���m�鉎|	*Y;*��;�{������qI"ޒ�/*����y��\9���kI�1�16�pe(�ۄwY�1���`&P�n�/i�%]z0mr,� \h���� \e����8s�b�/ ��,�F�<�_��J�/8����"���3N\.�@L�܄'G��o��1��y���\��X�����{N�3�I�X~��&�ӿR2)�gw��������?�S��5�;�.�z�����k���ȭ����[��l "�I4q�7V�r�?9�f�9fm,�[���_�<����X�����QXWG�H�;!#І�I`;\"Lʶ��Tƒ�.ÂҙX��q��Y��a�'|�ݙI�0685�d󴭉���@��S&e
S���mgS���0E��R>E��wNr^�E;R��J e)ë����48�b}S:듓�V�J�@\h�y�?xnE����l)�9�e�8�9?�@x�)���y��qĩ��(�<_&����nVn^��t�׾T��hW�p�`�Z�CF�3�?i��x�����p�GI�B�x��[ws���$��t���=��Y�s��\H2�o6����]�����D��7W�3�m���KWC��
��$j ���E(��d�KK2����r��O�:�� �j5��r��	��ϣ�hBr9p�*�����D��������Σh�Gf���"ӄR@G�� tv:���W7n$�	Ꜽٯ������*��6a��x���/K�p���>�0]�QY���9����5�R�xC"�7��^+9Д����Ȏ��vrO*b4B��h�!��:r�/ʫo.N�ȭTKҐ�:��[�8�Q����M�>�Q�h���{!�ބ,]��G�T+i�Bˡ�8��~jn}�{4�X׍�T�Nk�Dz�o�T=,�19d.ܷ��J�6��!�d�jpsU��8"/��T�z���hȔ'�<�Jw�iS�������;s��Ҵ ���f_�y�vUX�5	��Ao#2����Jnm���)b��h�����PԄ���	���r1�ێ#�O����,�������t�jt&����l��zt�N�5m4j�v;�vBR�����9����)���Y�,��*-a�;͞��F`z1�|�u\f{M�pv��T�q�s1E���F��?����I�pxe3�a�?��"}7�c�����Q_jrW=p��bW���s��7. ��-��EN.�_���9A�%j�Ӕ뱓��S��s����#n�%oӳxJ\!�I��x�&jN>����܆)�8��2���P����c��4U>`��U[�:��~\��i�\�d����Ɨ*��(�#��y��(��b!�YEFj�	@"�3w��`�+"��xw�9{��	H�SjGoP�E���4B�ml�Z�:cغ�l���)#b }r�ҨU:Jt��Fn�s4C�P��|��-�:��Ut��a�>�1��#�[S1�����g1�L��(�7�~N �u���F"C\Ƙ�
�[��#��2>�hR����Z�W)^=��HOIF���S!e�#�TUST�+�YS�A��4�7��2�ڕ����:�*$s��l"x��˕*�IE�VI��S�@ϓ� �>��QO\I��iҫ�Hm�>HrC`��OR��rJT���j(&i�ɾ7c�t]�)��>��.W�u4=�G :��V�`�J��[T���z:b"͗8����+��X���7p�=y�C��>L��5�*U��{�.�U�q�I1E�����u�k0�abBY�:4p��-�k����v��z�2�~ ����� �Kl�{�T�U�`W�����xJYB�a�̟J]���\�p� ���Q�J��j,�o���8*C5�<qKy��W������p���Vo�}�2$���2��V)�2���r:�Pr ����]��RRq7���/�P2�a������ns3��٪���-�u\��ڗ�U��d�[Җ��Wp�F��/�{uEփt�t��X���c��<L���$ן���.���h/SD�MH�%r��ej	TSwg�c������#�S{�n�E�^c�&�b�T<F���9�Xg�~{�l�5XU��U��ͤ�����;��sb�5[�`����5��*rY0��G)���=ؓ)��I�[�A�Kk���ZkT��A�?�;a�8~Xz��k>�o	������ucް�o��t��u�GU}{E �S�/�l�k�N}0����f��OW��ƭ��h"�_
�c�ЈZB��`�˸k��9��8��Kt�<�Z\1v}��_��h�&����d��e,P9��ɤ��ųMU����	j�� >�<W�8(�S=S��9G��~�M�C�s��	��5IPLoGj���G@��~�g&�-$8p�P�A�`Ν�Ǣ�س������F��B_���E��������B֤~���A����ˉ�cI���L�q�ƪυ�"��1BAAx4�Ԕ>컽�?Z��"�����\�s�DԬ�
��l/�����}*�"��.S��_r��R�-UB��8j�Ӓ� .�ѣ&~��?�Mz������e�[O��n\(5V���Sk�P�S�S�X��3�6To�dzh;7�HD��6y��L0A>�8�ѼI�B�����m�a�&��uV�fw�3f�[��y��C�ǿƅp�F)��鵂��Hy�,B�@_F7~����Kݜmn�m�H����2���P���Y���)���b+]��з�Z5�=�[�h_��ыU�p�阮&��׬/߱�^�\0ԛx����O6=��������|h�.����w�QS���%��N�M��q<5K���������v��\�k[���$;2"-�.D�MY���B����<�Ni&�c��@���I���_jV����q� �٘�Q�x��L��G8y�0�F�n�e�aN��~�j_Q�t�`�A�7�U=����8��۰\H�H.���`��"�q�\�?v�Y��k�x"��8����:ŪW��7�aښ%T�ح@���F�'޻&�3u����
Q�_Y�P�^8G��@���	榖�a,"������I��@�(�-t1���3�p���Bg��L�*g"_	u��<�?=^o��A%[�R$L��:�BK�o'7`���Iy�0W:��nh�(���h�t���5�J��I,��\�Ɲp`�W�/3���P�9��ػ�l�,~KI[��40s��f�3��O�ls�K�
Z��W`�5E�q�"n���S9�Mi!���&��WA���n���/=�B��n#)Ѵ+�<�@w0f���PV���B��3.RYH@yLI�Ha#Ç&P���+SsI8H�i2��ݖ���r��أ�d���\�	Īp���!hYO��yЋ��́,x1l4F���s��N�����X�f��6������i� ���k���v�vAv�0P3}i˚ݑQ�C<�#�Z��PC��õ��5��V�~�7�/X�(gD�����8�ާvœ��=�!�|C;q��%C�Re�h���6;5�d9V��7] B�A:������m���B{j~��4x[O M,�{�B�)3˓4IlK�禯~�����g�v��������b,ǃ������QD�Y��W�:h��?��`����* �%c��|�lV���
ۜb�{�[��Dj�������G�B��>�YN�:��ˈ�3e�A���7�~�'wZ>Ä���k��5��t1���D��]������}wI\�l�%T�4VcDtS�qj�ύ�����\��D�"R�_�}e2'�
'��p_a�����k�C�/�8	��Q�	��P��ས�mI������<��Q�P�h���sv��TX���O���=X���N®e��	��A$���+����uo�ީ���<��ґ�X�Bad�4vq�ۤ����8H �(��*�!��p�ē���w%8��E�-7Hi�)��u�tN7��&u+,�u��p��k�N(�8��g�so�#A9��]�B��N�ui�{�1�@V>h�їY���qg@��u���]{�V?|��C˂Ud���5[�l�*W�$W� �/�`_y���lKo�I�Vw,zE�y��}zir�:�� ��p�tuF���e� �̿�<�.{�.oh�EC�!l!�c��f�;��8U�5;>�%������?R�@i�5�IsV1
�ń��P�o�kv�+�I+X�!�>��¶��~ u �tӖ5��;+T���J�a��"sn������&��#��V�zٗg���O)�5�����z�L�ȇ[Tьk�y�ﻢ�f��x�ƚ�μׯC��A.Rx��"�o���@�F���OS(3?�1#��%2�u���t�rѪs�@���:έ�n�-v�`��WX��&������n�)��v?�n�@L��Z|e�W���$��V������Xp-�5��@턉�|תs1Q�C"ޙ$��W1M��%*�s̶O3�n#l�9�6�ߎ��2�e))?xК�_��� a�����G̗�.�r���:�I��}Kz$�����awJ�(L��?W��R."vO+�`���L��cÎ�Q��?jP�7ӱ��eϬ�FyBR�Q��X;/�>wsEI��x�-�g�IL�&_��o~ W�౦J����\�E�W~1�t` �H��ȥ��v�ϖ	� 8�\D�Ħ�b��FvRрp� I����q��3*�4�9����,R� T��_Ҍ�2���4(��_^�s�b=C��>�l�1��0�$��,�K@���%�د���Lt"�SDJ���zt��Yom��#$MCo�-�K��3}��� ��;�Y��C�Fn���wZ���TG�����f}�艻�, �2��H�����ڋ�˜!ws��#y#V���D�=������ὶ('u<�F�l��o��T��K#�,�6���dX*w�W��ݙF>�;gm��e�Ʋ%o���Σ�-�lz���y�<w�d�D��Hl�^|�~B����g����~�9�C	�s0�Q&�"|d�v''�g��U�r��BV?y�|сM���Y~93M�j��-=*��`��JG���8Q�5�Gv��� �� �ԭ (𧻓��^h:���X5���
�����f<Sj!j�"�E���]$ݦ9FcU�(T+쩭��i�D���O����S��+���a�z.�6m8�b���/'0��+i8��i9��Ƿ7z�Ш�2B8���J��.~�M�	y(���ކ�i���]?@"�l/��6ؙ�ѻ�_՗|�*=Y�>n4��	��!�ҳ]��k���ґy��P��{�̴��o�g��Y���ge��*>GI*�;� ݁?��)�s��ӑ�J&��T��o��o��o�nx�.#�qZ���
�㶯r�!zƅO�����"(��(c?+������F�PM)6Ӭ]�	2k���ktRjfށ�P5+o�I";	 �= 8�8�]��-&
H���ED����F�Tg�-i�3ceRD��7�4+�گ��w0�\w���]a��z�[X�x
��ɂs�F�*g��u�MH�Z��ժ��0Ֆ�2䈬H��. ���Fu�Y�tz��ey�R�m^�ͪ[���ƍ $�>�>ҝ8�6D׍8�ҫ�x��f[�K�֚�u{�J�#	��u�P�ݯ��0P��c����¾M%��W#�ǘ��3Q��A��H3�B��C�/Νro��9�"�k���L $�7��gp�$�Nc�җ�G��?��X�P����_ď�UyX?���r�A�3ȉ�諗bh����E�V�"�����/g�3�����¸�In�«Iw��Vײ�n����9~�C�V|�E���,w�*bql�&u4�,-df�B�Y��BEmV��7�D)�@0VWI�Ho���ak:��(Yc����^9*��D�>8s����a��>10�`m��,�ƙ�IɁ��|V�*�����#s.�\��l��]��abG�CF�0�,�{����Fݙ�����g�Ѽ��,jέ�|yk�f�l��)0�|�9�<�&~�]��K���,-�^��0Z��qЙ�q���v�FA��p�(���$B��$��E'����Jm���/�t��sV�
%��N��b>�(L7i��J����O���BGwe��7΅�����	�|bA��JL���ꚈI����6u�^i�q_�YB�������6��H���}�7�ò�_�������id&ewJ�b��f�V^��)�㎵�U�&�%ݬ�⅒6�xg�ђkU妹�!+k����%i�o|�/���Tӱ1�e\ķ���_�`udZF�sd/���}[�E.�2����t��q�mN���^Q�,����ʴ��k��OL#�!���!
���y#�3h�ɴQ�^-T^��j��`ȅ��q�Qr��52t��C�N�de����'�a�/�w�fvn��kܣ�p�	�K�9��_Q��������Ȼ����H��+�x�C��/�)4�&aj���>9����5U�tO�
>�m�O?I3D��� ё�CΙF�P�zT�z���������K��9\l���� 5k�B�6m+ۇؐ���%>���Dg�e����O��؋fo01`��u�/E�?bozXd�ȯ@���g~	�y�/f	J��=���l7^�0w3W�O�������_Nq�M=���7Rt�9�ۥ�i�E*�$̿
)	�FL �x�V3�.�_���셺 �f���31�Jv� >��k~.00�xR���5IT�s#�x�n���:4#�Uŧ<�Q�i*��n��=�l��P(ן&���c�l.�Se��Є ���7����c�$S΁.�����wd�c�ڴ�����B��p}����6Z�A�	EP��r�c+�"7K�CP!P�ɍ����r��B�Hb�*y�f�5�������K�V��0@��n�b]�-�j%����w�Ȟqˣ0zx20g��d��4u��,�?���3�U��ͷk��H�d����@��"2�u���j(}� aG3� ����a��ټ��<�a��	�w��Q��42#�I7�@>ZSтF���+]�ԣ���C�\G��{���7���̷i�4��ر?2�9Ui��[�	F�3p( �Wn�� ����X|Wq��_a�2�xJ�	E����z!?�ω�. g�)�t�����G�9�>qDj���S��zM�|�~}/R�O�v�2zq=	牢����z_�?V�:�y ia�*�������!�&s��),�)e�}�����B�۳��m%�)t���*HI�p�9�)�ao��}�HCG���bd������=;�x�Ha�f�q����l���`�f���-�ƧJ� nZ��� �ie�jl��E[����؉�����@{��V��h�y��;�/�js���v��o�
�~2��� �?�^x*rk�zC�L}�A>H��Y�W))A��P�\~�W9iGw�jB)|�(�Z�+Ue>�\n��`3��՗��2~��̶�&���<��D��&�9�z|~�2xڏQ�Y~�]O� w�ɔ�Q:�B��͞2o��l��k�~_���nBO,���W:s��w�>��Ua.	�%W_�1���|���9�#� ���ۋr1��Ld�1��h�7NS4gq��l/�]!
�gz��a����B�]���ӻ����ۿ�~|�cK;�@5g����t؅�~����`�h���ܘ��ݶ�I&u�5�5]�c�?��r2�98o��B��,���}����� ������k�/f�9�(�BNfIm�X��Y�3̇r{���pG"��2�6h�oе���2���aSE�~C���#,�U3���Q]�s��>�m��q�;�n�D�7JIܛ�����F���U�J�@IK����3�͢��̠;�;���ϵ�S�����]Q���a�<_?k�YS^lh���3=�s��/��Y���iC{�h�2w�E"pR��;��w����������}�W*؂a{F�Cz�mL�.n�
���&�XE�|�(�Ȭ-���4��q���ޯ�=0{E)��fZ�ue�����̔@߹4������n��)ʲ:!Nl�RF킇�h.�H��9�8��]F�˛!Ϭ�f��,b�DD�8�̜α�ݖ��?�+P8?��"�e�iu7"�xJ�3j^W��[�����'����[��RGa>�2jH_aD&u���d�\�+Fd�s�x�b��&q���k6K0��p�z;��?�h����Oa������uXL32��m�VX
}"�d'�O�
R�����M����y"��[VLDdw.��HR+�s�ǒf?��G"0#ш�z��G@�7"�X˳�ǐ核�B���}� ,�+OK�f>��� �����	�J�µ�r�v�4;��.��	�{�J�"^f�^`pV}qu��|r�P�A1���A���\M��'s�l��ߒ�/�TM�����6-�f�I�*��򚝚�	&�S�en	Z��UB��$���֤�L#89Л@)i,͗6�@t%=&�H�Uy��:��K���K��]��U��I�A<
J�v�qGL�k�\]s��-p�R�>�(��,��)��W���DS�-!z��lP3�����Ag�����N�؝r�y��Mn���3�����/ā�O�LS�R�?��.�r kx��W%L��ƭn-�t�I�Ag�޹�0ߣ`M�G��yT3�9�ː�@��'|*tB}p$M�]�=@dq��-e�����M�^�O���������I�#��-r�- I�j�L�rL�'�&�w!Fb��	���L����&`mu��JSX�OhJ:oC}�h]�Ė[�$9�[D1�.�?"ǜ��c�\Ą��,�N�ڜ�h2Hy���!=�@����QU[�s���@,%��l��۲g��K���
��؝��	!��������)�5�[ݧ1�?Z�Fd�E�є*#B<��|�A��D1I�Ak��t�L���"V�;ĕ�����[�d0�e��&Y�$���b_�T3�s�<�N;ƃ�'V
9Y��N����*�$q��V����Xg꣦f������W�Bw^N(WG���o��EA<e0��e�d'(Y�WEJR����nW7�q� �?<��1��O"�"�G{�e �� �;2_��!=�u�+�`x7L��6T����xv�W�7&�νuQ���T�.�={/�{�IAU�)��Z�b!��aL;gJ�!�l�xֺt{���Dlo�[9w��2�bk��"���b#M���.�O��BO����T��E̫N��3"+0���uҨ!�ʿj�j1��-�Q�F��r)Io]���Z�)���9���G�bK���#R��(S1�N���px��ѱ1\���0����E�%r��T��� a�&�ԓ��aF6\�*��G���D�|_,yׅ���Ց��tI�������u��(����Q�5ݑp�b�q�~���Y��h�ۮ( �J ^�����s~��WwJ�Y��G�D1���K�a�7�}��X_O
�Rӹi[�5%ϸ!�.~279��E�����j�L��B�ކe�y	'�x������:@!\�j@�se}��1)������
"G��q��%S���P�B�)��^�c�G3����52*0��3�}��>?�mO:�?�,�l����܏_;�V����PcF���� �ܡ´&o�(�G��!��y%/t� [h�'�'����6pu�<�n�X.�|�j.1M����+W��mP��m��R��	}[����N��b(uߋ����>S�|�����7`��L�ʽ~y����	N�>��>]dk�*�Eh;�V<�^�h��k�]ff{1�����@ӻ� FcMz��
�v��6{(��dnQ�gV�������p�r!9�c�4�9�&�;^[6��~�z ����Ob�F*]&�-�y>�_��
�q�b��/s�
��ɱši��vT����D0��6�X����r��lN��e��[q��P�{u/-1\�=��;_$3�w��n�:�]��]��knl��*1"!�Ȕ[�������>KGO���
oxLa�!>X�V|��X��������6��1��P�Ħ�q���`�#���`	p��G�j՜�ėf&]?�H�;c� 'txSl
�����a��׶1���m
g=�m:��������R	�ޱ �0�������Ǽ_t����FD������+��-J�U�}�oD��}߅ܿ��cl=W�%ķ�q���R˙�����f2�7��f��0�8898����V��BYyf�z0����fF�F2����\�	5M�a�88�ZJ ?;.q���CV���՝�q��=��[/?	�9>�����rz������r��N4Z�n�mPꮭ	���W��-ט'rT`$�0+n䕖���di��,9��bN�H<�Z�Ѯ��6���9�D����C�=OS�zc��CM��DzQ�'U&o�6�!��\�,I�"?��1�ҷ�n!�����
�R'�liX��uk�׋a�2|)�8�<�~�W)�v�޶�|5�&g��^�)�g{#_t���k��p��� �ty#$%�APQ#�%t'�4�c���
Dr�oFo�k��%z��p����q֓���%��4�������	6�{�8�.��ZV��/�H�[�Ӎe��z�'nr��9�B�Jr�L_ �Oo%oc⌁��I��HBg�`s��ќ�auhoSF��U\sm��^�����&c&[lwt㎎�{��� �����iPM���Sc��j��S�K�Z�G�L�����Z�����d��e��+���6~�\�[�ѾDȝ����s���_I��r&�eB�J%X'��iť�3m�R݁��{,��xY�Y?M�ոp���.V6��n�GFb�J�`!��Q�B�x�"?���r�~4԰�/�Ź�3l[@@C�r�x|����bwp@��f<#�hR�Wܛ��+��o}�$Zǖ(X?�� ���w��GGv�bU�t6ɞ������a"��s�ɻ�M�g�n"n�wZTI�!�Xf���$��i�Jp��NT���~Y�E)���1��;#��)�������u���z��,���#ة��r�X�m��]c=��P��|��`�Dˡ-h��~� ޴���� �Z�n��n6�Xj(�5:��6�4A�		J;��`��<�e\9Ѹ�S ~i��{!�)��³�"�=�[y+�*.G�7���ޯE|�"~$x���Ar?���<~��%Ǝ�~zK�4�O��}�
~C�^�3 ,��K�M�g/𸰂C~��h���~���3'�p��̾���G���{����߀�����D���!�-�����?�� #���v7i;R	��A�XC���%��UT��ĝ�=��b�z��`�nג�޳�l��NI|� �l��I'^�Ilu#�5�R� �Lj��ϐ�;?E�{�')b����^��J�`l��� *B����`�h��;>�СR�.@���������Dw�}h+Z�6�OK6��U,�\�6��P|�iK���=�]�8�f�U8��h��-�?�%G03@k�̚􍔊�z'�U,R��y��>� -[��2:��b���.�}@=�^�4��B~!9J�9_Q�f��	�.�[T��v�(��x���a3�:��d�A�#�ژ��b�z#c���G��ė����tw�E���P��p@Qw��\HjHn��k]}�[W��$85(�� w)����7Y���i\�^��"AaHt�vy$UP|M�|O�@�У*q���hlB��M�g�FY�%sߒ��=��F���r�$9w�{�jZ��h���x_M�lI��C�B� )�t�
�ü���j���\�{֕����IU4:M�n������G҈�ٻN��p.�U[���l_�7���
�	9w�fv]D':��
daU�fW�[Sɓ��|��/�<����j����9����4����$NR� e����`(J��X����V����Ͼ�☺bv�C�8�K��IA��OM�6B�����sGD񺄙�}4��eib�Nc�u(/��F~������6Q!H�
_4I_�X��pC�p����2�{����c�R�<�x|���?���*���dΒ��՚É;�gGn�u�<�I+��Bd48��5"ɰ�ӓ�$�(IYZt�l<�qMp������ͬ�8���ؕ����*D{�7=K909S�@��U�G6���J���Z���+�.[v����1x=||�ś3���M�܋.[�^KS������B�S�~��$�O���U���W�-g����/�==�M� ��а��?�|�x�R��[�z�ҳW˴���*���֓^3 ����zxC����6�B��\yY��J�ʰ/q�2 �U6�Muy��G� ��C���K'4�2�5�f�E 	��H줰�#z�-|���If�=_SҲ���W�fGe(�m��4�6>P�4�R�s�ֻx냞�+�)�� {���/�T腲ł��lcM�W�I'.,�w %HB�K'|�
0i����H8/%�i`�X�K�'�#���DS�G���"�%r#��b�b���k/��S�}�%��.�k(�*�����n�G��Ǳ[
�a�p�*�@2|2�5$w�eF���,=}I���4���ئ7;��L���]�L�j��<��-$Z����	g����	��-Gl�k�ă�i��DfsPn0�u�x`+��	�?����%�S�ƙ�]�L̀E�Ͽ�-�8�0&2]u��H�i��Lk_^M�κ�f�GW����ɠ5�F���VM����{p>I$eX�gٱ��R�����lmc~�QN^�h��yP���(rG���1��`�mdB� i.���17�~��FtSMpG���m�˵s���7}���;��:��>FC�o�3�x�=u�_�e]铟�YF�_�ce�EK�_\�R���5���>d�9�hl2�
>���P�W���h��	��sɊ�翸L%\�6�["J�����{���`���Aiy2�,�X��޶X��k������.�!���lo��\��Ɵh~��-R⃹�eJ�q�b��
�e��ۢ�s]���Hlۮ��sk\!�v�e�a4]O��25f�m��=�>8�_�$녡�V�V�<��������ȩ'�G��� ?��"���������l�G���gh! Ψ�!�I���'{A�����frjOEźc<�P�@��v6�SĠi��Q'
Q.F��K U����ڨB����hl��k\� �4o��gpѡ9x��W�hCR�����n	^Y��;��Zj���]������N�;q�g<L�m��FPY&&|�T�12lx�v_�ϕ*}Qݢ;�l3y��jL�����¨��K؂����1!M#'4���F@aM%pp��n����S�x.�h=�Һ@el��7y����<Є1�?�V��1�n�!����1�B�(�is�����1��;fzN�O8#D��z��	��O�5��w��{��&���.���4�jݶ�i8[Y������>3\��e��s��7��Ч6g��^��v��5P��L껥�˔�I�&{�l��\��@d�ՈXr4���Y�٫�.0��;�B����bM�U�ZHJ�Z�Ohwlz#�o��G��c�� ���� @lco���_�ԏ��M�!���ې��f.�V�\���Q�0����~�f؏b���F����^ߡ��F^�D< ��<����7w!�HkmAY(�L1�GѨz" �d��8��r#�mY�K� ����g�.�o({��+����)R���� Z��]�ȓ�zfl�p��ԕ���ZA6�KS�sn�����*��7�ό0�5"�墉\�b-�{"#��cPR��|y�U4#�Nф8��!��Ryw���զt����0�p^l�.�sųz�۝c<qb�TY<<���(Rؠ�w-�D���6-���ԇF:x��"�!��`e.2*��:��7��d�d^�����S,e��A|�Y�N�u�C����F)Ң��b
u�9>�Ls��dm-��Vai�@����)�X-�/:�r`ov.���6�@��V*`tbhve���R��̏%s�!��fT�Ѩ<� ͩ�U���t�$��+�87|�'�.�Y骦����{7E�'+���������9*�K��S�+�[�zp�.����uY��q�D���������� �u_�t�"��HE���^㈘��t~=7��H�J�x�k�!i���L��f�`:qN�����U�S�t5��g��'qO����0O:��H�p/KtRk�x��F�X�M�uGbo���Ȱf����Fi�c�qOԜ/~$/���˔{�<��k�6�k���`D��ֻ�6.[
B��Sˏ|+mo!��5؇E����=�Ve�e:�W��;2��nP>l�������E�z��_���\q¼������n������ ]�D�Yl#!����xt���pZ�I_ŋ~īJ��['CD|D&�(���ᛶTǾ�^��Kwy�[����q�[%��1���dk񁈧K}�||%���2i��=���d���.i�y)��$��)�%�/��I���H��u��4���vl���-�4��ҹ�6�9uf#�9��#8��(��<��-
@1��PC�Ւ)�����ZI1��C��#��6.c��;_��2=�!��"n�'{܆ �64܊� �C���#ūe�&��~�H.EY4���ڪ�9v�mM�^Z�4ڄR�=S� �������O�E�� ����CgT`;ʇA�Vs��$7��0�����єy"?� d4p?�����-;��{�x�_��MO�@�A=�nM�AVl 漒�=����3���zM��@Hs�Ͷ<Q	!�������	j,ssX�O�!�]�(� �6�<kM:n��4�#�>K�^�ls��-����6��wUiX'n����Mp�(��~hDTTf+j/}ړ0� 9�� z���eň3/�㐳?z�Ap�g�{M����1��f+sܣ)�4K/���)�*��Ck��7��&���lX���ͱ�y��;��O;��n�~�Ͱ�`��ra� \W��9A2ڊּ�g��r�`�����[	R���$c�+^sS[C�^�=��[�m�tf�CF�fڙ쁤�m�Hc�O����1	�����35H�4��@�v� A�q�)BW�ŋd�������q���xx&�����j^Jס���J��go����x�qր�&�c�$�<,���RRkw�?W?�Z��ㄞr�[[�D����D��4����Х��,0�/eZ{Ў����P��	a��G�T[��Ӂu�KhcL��Z;��?j gIj ����`��Z��=�� ���%G�O9�.N�,J)\�����u���y٬ͯ��#I�A��-2U�@�8?Ӓ���0�q�w�&
�;#ÆA��(�W��ڧ� �t_
�K�,UW��H�<v��*��}pz$�)/�L�l�׽��o����Kz������)�xF�k��x�C����S��7J�L�Y����^D�wnY[���4��֊�҄F~�K�)lC_p`:9�,7���XcYK9?���ؔ_�<`u�u��{�N������xo�8���tDn=֟��q�t����d���˦��z��o1Ӊi��K��BQ�b��K�BYE5�eD���Kp:d"��~��[ ��'ah��r�� <m8I�_��j���Db���`~d�/5
��0�@�B�*!�]Yz���%Oֆ^M�Om��T�wE�i>g,s��;9̐����X��Ϥ�Ο�*�{��+K�1�\�5��ڍB�6�(ś��-D���G�c&>�%�g�a}�q�-�S�@���^S��=��|>��9�3|F�5jQ���@�w��6�Ȕ�V� �d��л�M��5�L?�H��Lp�"��*8ȗ�C\��&����H	�;<��
◼�l��W�s�®�b�gr)�R�S6b)����K\�3{����Z<o�jبeQ�+Q+[h�芕YV�oD�kկzIL_���|�i�LyMKw����=��3S����[z�4Fi-q��c���� m�.�v�D���׊��i�{�����Զ�&�*8��rH1�g�is����U�ZemW��(4����{AO���h8����-�A5���g��;����|	ȼ �}��m�G�"(-hq��c��D_�oի�)�6���?�$t�I������7�|r
�*�>�W�ܘn�ջP�+I����4��d͔�cA3w����e���w;�4P~d-������J��+ vѩ�+]�I./�R�pֿ�2�+Yw� �t��k?�C9�_+OaV�Y ���i_�7� �F���5��Z��?Sƴ2�(`ɦ٪�O����_����2�t���T|
&ns���4g��L's��3���f8���Р�}�gh2ۯ��Sca!�L����vɸգ�vy��#��aO�vmy�O��&82"U���d�NT��l��w����P���Ԑ#� rmo�woJ���C H�z���t�`�Z���2�(9������|��1�y9aK������� ��ywBfV7����7�����
�|1��S�I�7q.�`�3��z)ʫ̒�3u�V�{�l�܅��V7�O8�6�����y𩏤F��V����.���Z~��FD�������ؿ~����|�BfRA�&b[���?t�C�������^�q ������f]��z8�߳��*�3�9%:V[�[V��T�Lp{"6���2��;��\?�f{O�w����x!��J�IQ`�Dh7C6�ߋ�Г�Y�c�;��._��:bX�_����iF��͋
n�+�/���Ai�l�<���!KU�m_�Ӂ�9ɑP�j���OI�2=� �"*���t���>�:��o'� 'FLe���t�n��*���+���	I�2O���� ���Q���9���S��|wa�V����gQP��V�� �>�>��7��1����Fn�~��P�m�b/v�.����t|�1N�Q"�S�pֻR�:�I�{��?HI�;���5���>�m�f���hR�vn�;�#U�A���]�H�,��W�#O���VR [0�L�LȚ!����&����|�SV���s�O�Us�Դ
�k����`��T�(*�!B�~C��B�+u#�� J��XNq��R�����
0��߉���D-�ù�EO���k�Z<dD����P���EGح�ኹQd�q��&M�A��:(Y,hg�?�+E\s=����6�`���6�0��p���Y��nB9��ԥ��ڏ�pi��X�vG	#L{���p��=��Rm}��h���/�hҌQ�=�
1�Zx��E��.c���NX�)�$8"�e3X��q�p����%�&Wa��B��l�oJ"�i��8�Vhy��L�-R���q� b���y�k���@�s�j��L	X��ŢŜH#�K��M�!t�����	���lK�P�������_�tY�X�b"p��g�j�uz"�E.���G|�IXg�S!JZ�Ĝq�?I~���G6����{��N:t�^�U�77Kp������p[9�@%�0���U�N-�	z������"Ro@��:i��V���a��y�6ˬB� E�b�4��̅r�<~������+__n��y@&����-!Yh�+iV"��U�Bo�2���<�+��-� +3��y>�(S��֝��oI�L:�c��	����
e�@��������r/w��׮�\���Q�K�"ԜF؎��|J�2� ��{gY��s�۟�a$=M��S���F\�d7ɇ6B��Uڧ�����Zj���!Q*�Q�@�˥�O �UA���@s9�G�R!��K3+��* 2@��Q�v��`�U]�t��E��}��J�;�}�D��u17��WV ��w���$��Z�!0�R��
	[�|��"QσimO�=ưl*ц�q���n=f��t0)�&m�xǖ�A�7*�@�g���8�M�8�X��~����GM�� 6�TZ���8S�p�\yV2�\��ʈ����g�?+��y`�� \&e�eɉFR��RL7yU��s�Y��4�{�7���_O�H�-Hf�T5�C��Wm`��:C㥳z�QM�V��˅ ��ŭH(�T�6��Eq�+�x�/�M�iuĐ���
z4n�7T�3Gۯ��>:<�(��(1Q����7�� �YT���$��;�`</K��9~ �-_+�VTݪ���L�,{Y�X��Ѓ`��+b��C��������&od�&����� �C�,�<@��1e}a��v�:W�X덽�5�g���r�ۀ������[A�@*ٴ��9�����ߖȉ������e�s��������cO���AG���ޣ9)ܞ�/����cyB�[�=�H�)3Y}�[bɔ���8�>f�� !�"k��Se��{�/;0� ^J ����Qd~�G�@x^;�2K6���VS�N��?�(�&n��}ף��k��6�Q˺���&�����-o�1���z_�}�P5�ݺ=��=��O���u��n����g|I���l���������PmA��Δ�}�~�Gcd��	�,Yj�L�&'n�;�||9�1+�Y5��JO�t��B���R��C�b�iI]��f�Aj��< >�@��t抨�^����(�]xw�_��}���x��<p�W�r��tqՑN;���h-��CΘ���z
n�8�!/ �U�Cq�T�xG^�Z�7������������L����<���|��ȫ��F3��K+)�s�08q�"	
q�
P'���D!N���vp�Y֎��%	-4��EZ��6=�X������O0SH�.�����3��$'��R��/�X���p$��3$�k����Ca�!۞��A��ߠF�����U��V���I�ײ��X��S�zg�d.�ūǴ�-�-��6�A�S�f�� (L�/��̬+<W}W�]��<2�|8�
�J�6��Ծ�����7��[c�M��^4&>��aݐ*���b��vI �u2b)�I�ɌC%wT�o��I�;��,ڄSaT�t��ku�n��w����AHqK���1H��lE�J��h�gr+��J����80QX�V�����zy̷���SǼ����[�����iS���z��u.� |ៜTL�_��u����!淝d���9�U�+o��?��^�0Z���u/�20;�r:r�Y:k�!�K�*CW�m���m����ҷYn���:�#�iR�ʪm�F�k��&��_�\-H�J���}vh�����c�1x�/Qkv���%T�u��Mr�i<�5_b�^�}?#���<��.��ock������CZ��M[ս�]ϕL�;��ܘ�>,c ���b��#�惺���Z
��� R�T���|ߗ�s�dE�<@�:���J�FUU���KN�8I��<��Fv�p|/�q�`�'�^�+��;�T�"�_Ѭq}C
~\�l���Or#3����뜮�W��'�}���v�i�ڷ�{N��5G_6��by�K��C�-;R�8
��û�9�8�U��/Gk��QVۈ��f�	�g��~sr��ĩ�m� ~sՉ�W�opx��B(��Vi[h���eto��ذ��%�px~�dh~���_�b���|�^�{}�J�CW�b�w/�W�1ь����}c��Ot\kAA�)��.J�����W�'�(�����j��AG�x���ֽ,�˅���V���T��wj0@�g��9�Yh���P��!F��_�,�8�wNʅ,'��U�>�;�+���JK6�V��z��	�~��44ܟ���I&b���&;5Ǝ�d��^u=eß?9O#,�w�s�pWn����I���疝�1��O�H��G�kk�Zv.}{WiW&�ܗg�9�p�V2�}������[Ჩ�݌2[RG��	�È�؃$	U�4D7^٦��"�+V.x�5�jD�ݣ�P z#��S߿��K��伣�B �=-_i��, )��ݝ4R3^�����$wy��с�4�{,���˿�l��o�.�[��G�$��N��[�R�@:��}/.D!�ɟ�k����178�{c�0�U�MET[cN$��9�˹ŲѸ^kT��#`Q��#��+ntu��'�Nn�K��Z]�`���u?H�UC�͌�6������Y��)'��v<��X{>��{u���10w�b[B��iGZ�(��eq}Ο/;ɣ�م���c#&��.���E�8�PgM�J3m�IQ�Y�V����x��Oe�lY��y2-�X�ya�T�]ڠ�&C�w�6 �c<I�Q�D���J����B�lhՠ�6���V$�[~e�*dUL�����G9E�z0�/{�ea7X�iI�q� �O�z;2j�{Ŭ���r�y�p��=�u����7�&/����ϿO?��W�B��1]�Z��x��/���v]U��ߺGK!'ˣ;�7�Z�d�u�s�c�o
�m�������)0(�L*3��nBi>�T�	�eܡ=�7����k8t���f�d��ρDb�o��S�f�K���j�S��Q���+��U����,R�X`��_�(�%u�6�,�z��1e�h�
��~�ƙ�a��:�ɘ�
q��6��<��.���XM��s�4?�å�Џ�܆5��,��!�b?���"4�����d׮빽��`��d)i/U2����p�"�Z�y5q�p��q� ��^��_�!?��ŽL�7�T	"�YW���؈䔶S�k��"���o��Fǁ�%��[��fX�Ž\����ܿ��j���RyL�U��,��KY0��4˯�� ��/{��￱{z�},'܌lQ63섹�KW�	V}�I�!
=���*x#��2>�frc�Gͥ2uL�ET�U\j��ןK<����2��%`�nE�?��,�H�DF�݃_"�0 �*-	�
������q��ޞ�G�X�q҉-�Q*��}�8�����A.hdy�/�����<�+e��u�͓�4��CW�{��&ur�0k���s_�<�;��a�i���:�r�PLr5R/�k�O���cm�ˇǹɈ����_x
?Ib#�	@��{�L�)����؋�K��&-�]z�� ����9ÿpfq�
)~7wM�l;�]N��o<gx�o<�ذ�`�È���?1�:3}	�щeF�*�Q�<��?�
���}K���x}Dfp�l:���ϝhj8�f!;��j蒃b�ǝhw�(g-]�|���u���a
C�:٢���J2'nֻx�O<7^�=s�&C��І�6�E/-�߄0��Z��-��1��2s�y�h�f4m_�⦌<����V�+�,h#�w�H�ᜆ��d͸c�!a���R�k�5	C��	BP����� 4Iu:Fa�j�M&?��?�0�)�eʧ��9e�I�JF[����z��%�>V��Gz�ީ�UL{y8PE�1��-��/"b���!�6����>�?��GG[��GS	��:?4v����X�lJMfnʮ�bs�,�^���|���*��/*��Z}[�{B��A��2��Ϯ�{�O��jJ�|3i���J3M�%!�/�E�������b����JB����,���"���v=DK��h�X�KB���զ�J�2��%$�["�t�/_O3LC{�}�����z2��{� �� v=�@v8u]zLl�P�^�0�6Q�8L��ڲ�A�s�pY���YgBw�߬�b�u����.w���)��M��M�y�B{.�х@]A��BR��_�}��T���H��E�R� ���WO/d�i���"��^���	��}�bD�>�+`A�	�7�~ni��Kp���d� n���h�?�HG}���� ��n&׈��s�Cμt9�����sVs�n�B�	�j�G�hJ~��-~��9��l�s	�(����mM�L������T@́��j���,2��jJ��Ʒr>g�T�֍���2`�#Ln���v
ĚP��7��r$���mU��UI�H�1ixc6Ո��0 h��j0�&K��a`E��#୪��B�-q�B��f@#iƝXE��pu��5)����{� =R�I����|ۈS6���۞�Q������u�ދ��J��RhM�Z��د�����H���uP��I!C�ت܄WT~J�ٯ.���!p���K{���b���9`q�V�,/�Ή8i�2>S���m��2N_�f��M��lWAkT7��Onz�)�r�,ٺ]�z�+��t#C�A ��B�
A�F��v�t�5~�3����d>��no�\�ƹyo�`�sgR��qV�_�,Z����h�D;�LQ���K*�ғ`�M����a���5��p8��:�qQ�/J���d��-Ս �ˍ��YK��Ygn9�LJ!伥����&�l`�v*ۖ�����*3/h3���1r|ſ�K�箈^� zw�vf�"��])�m�M]�6��Ԟ��r�s��d���8�<W�`�v�4���2y���}�*��6F@������<ypuN6��}WM�6u��}/�y���7ʫm?� ��r3�ТHc�Ew'�_	�0530l�C;G�S#9��(����Ȍ1����b:��u��Y��Al7�׊�n�P6��sR��y��uQ��;�LfKQ�z��vv~��-� \u��yl�"tԻ�8�@�·��r�ʠ;�U���d���(�.��tu�k򭳛ܛ�[�R��[^L���K���c���0��W�Q���1���gCE{V#�E-�GK��p�ѓͺ�C}.��O��C��N^��6��t~���g����n�r��hI�;'�� Ze����/�,r�z­�3ٔ��a��c[�����@3*unȇ(��>���ǭ3�C��w�Y$��~;t�
Y9�T:��8��i^� �7��1�W���i�H��د�5qWZ��&UY.����������SS���P�
��Pt�ˆ
_�m�Xl���@���/2�~�[�#l�9��yTx�6E�[Ӿ�轟O>h%v��ee�j��r����"5�ɒ�� �`u�Gq}��R���u&��B-���:TK�� k�]�y��-}�
FS�Z�Q��V��I&�س��']�g�L7����'������{�{�+�?2�҆��Lv�2\�J�1�ө�y)%�?b ��؆p�J��=๐R��"O�L�:p���G�]nȐu���z���"ڦ�(��[����,O�M��5?�� �G5������	A�y����7��J������K��2/���%[b;Pk��L[��c�����ɃL&��kj�('��mUbۙ���$6�i����OF�	n�<c7���-��_��ڥ)K4�d�S%"1��ox��t����J��ى�x�4�A�����UF���ɞ�O�E�'�|,SCc>3=ې�;�y#_���5�� �R��+�'V9B�+�xoroSeբ�95j���B�n��R��Lz��|�������sa�Cc��[�6O��P�A�03'`��n>�S)���(��
����H�F���N?Y<F��Z/@(4,@�����|�6��D����j��ZN駻��ݴ/��a�!�15ygէ���iD��j�)�A~I��<" �����2.?���2��Te��_�kL!8{ ���,�`�ß��O|�v�s���\@O!���W<z���С<�3�0�8Х�d2��^zX\]�+���g/+:T�d�<��8q�aa~����~�eT|���Y�&�sn�^}>7��t�v6�~�L{`f�!"��θ102MjUٛB2�A�ǃ6MW�p��:e7ʍ7���in���?I��>�Q��5� _���`M5�<
<�?�Y��D.��T�H!�B'F�[/A�t�.�hɌ�s�.��]=���R��4]�DtA���y*���t0�\4�$s�����a�
ze����{�\g�6�G�Eg��u�[8���ͧZa۲* oE��|j�j�dޯQ/Pu�������D��~�3Mo�?�z�aѝd2�%5� (�Sݎ067~�#�>'+�(m�Y(���jp��/)q��>��D)M+ͤ#���V�,#��"֬N�}e���ȤX����|tv+���Oz}Yݦ7њ#U�=��߁qHJ^�>�=n1>E�����[�k����Y�T�\�	����,|�$�c��n	�qE���4�)c�Ȋ1�c�/L�6���XC=�[n�x�=��R����������=A�$�6�QR�$�=�]
��~u��j3�^[NX�����8Ea�
�1�����w��hl���F���EV4��6>��ǣdO�T�h��\,;8������m1�os�nUw�1�/�m\.��ؠ�t���;9��-t�4ء������mEo؝n���ڂ�&�^{�-�����+܈���F��(9��^�>偎���8���l�|��~k�1`g˰���e���́x��LDYz#����"=�z��戌ٶ�ǚ��	<�XG�^ ���� �K�F��P5빚���Bl�7W�tl���^��<���k.Ҟ4]F<��I�yD:���0��y�)H�)�:]��|ͷ�}䋙��-�^Ԑ`�:��Eϛ.Dp�2�m���JTx�c_�D_dYڮ0�=Q0ƼǠ8� �B�T�	0��y��{�I��9_aK����I���R(�[�ـl��%O�-B�;.Py��!��X�&բ���`�ˎz�]V������^�u���+�&��N��j��u�;I�P^���Fof^�
]D̈���,��O� ��3
�`�sb[�ˡU9w�ȑ*�|�Dtx��O�*,j_Uq�F�F���{�"��A-�7�i�\�T�ךe��tk�u��$�(5gb27ϓ���f�W����v<|:u��� P���J;蹉ϫ�0�2�,�Cǎ)�U�(L��2Y�J �<��u�y�%~H� ��^�0q�t|L%E+� t�ԹԻ}��d͗wy0�������D�`S�j���K��EyP]d�}]��E��0���2���NC�c�H��̕�nɟ�oI;/�݋�Kw�9Cu@f>�R�(S�B���}��ގ�P���t�'���#�_�2�xR�����5�����Y�ծ:7�Ev����˄L����w�U���W>�� w���.�A+&@UWgG�P�؊lY�.t����̶������t�!� ��:W}1�h�>��}���˕&P�/��$.we|Z}V�920�B�P��XB����7_��j0X�o��0��EpV(c���o�0��������f�v�"7О�Q��$Vl�����!�X��o�i�`p���|��+a���?�ˆ�.����ԱG�P= �K&h��lY�=�
��F}�V�Ҫ$�skޡ LjKĹG�9YcGRaG�Ϥ��{�3�8i4�,ria�
�Z쁟�ӭ/�x�j�A�Ø9ϡ�7�B�����+6�q����/;���RF�G�<��<u���m�r�U Կ�����ѕ��7��1�͒�ǦAr�>��ÙM�4��/�v�`�ߒB8�$��Uˉ�Zq�q�x/��ǀE-�fP"�O�����ϼA�Uh1�"���xT�"${v^p^����H�M\-b��������X}�~�A{AEkm�nƧ8�ֽ�-����?���D�|��%�n����58⨎dԻ��9��].)�l��FՂ�*GA�"�T]E"UA�Q�� �Vp~f�4��<!�M�¸��X�wt��P�|�t�x�_�P��M�8Nm@�B/T�Ѽ�`�"]MP���Se*��m���јC��d�a|�����]ƘuЀF�5�M��Ğ�Q#�a���TC�@�+l�ǎ�����I饩6E2��Ό��h%�Y�>����9X��@��	�"$�G��~^t+�$^Bs1��>�w~ڤE��J(b���l�=yQ����_1���^��7�a�͖v*�ߓ^Jft��L���2O\׫�
�f��jk��D�a�rLzH;�;3�w0&K��J�?؈�
�0�qq���;�W��џ�A�N�����L ���D(M��l,ެ�G��9!4+�N����m@ m N���!��׿]Z��R֘��S��B�.��a+me�Pb-�;�S!m&N(�f�+��k���hN����ґA%�aSi)�c�*:�dV5�hɅ�n�w���TI#x�{;L�§����	����[O��3�݋<��,�;.�F��*$��WW��d(�Ԫ���H��lfV�H��x��w�>��!�~�GpL��]��nɌ�]fe@ͤ��H
si�l�nl2�W_+G���\�XOBe~oQ	���D&
��]a_]:�c�d%�����6xS���ζw�;4��.hF�aù]����xe�(K�5C)vl%�A�,9�*�r��V���灉�VF��}��9q9��<�ǵ��s9 �bE�KDo��Y�s��X֗��8�A1��$WX$5�Y�ʯ�]��Ya�H�ڻ�:���
A-[��YI���(� u������HQ{�\��|q��|w�˃�S���1�vn/���'m�p��a��\5�|*�r|Sm�C���#�
Ʀ�|H�5���6m5�CB����؟3l�.PD���Y��eB���)�S�f���ǖ�LT�����vt���o2#�Gtw��+���/7x4t6���zZq78��1��'�8W�:���iV
Fb�C]�P-L�r�z���Qr��9�-�z*o��kܡe��7�=�	��6B���.��DI�v�H��dUx^_�ъ�^2�iA��3�]�� EyX�
dG#��J��r0W�3���b���.�� p�z��Ͽ�p��v���xb���WI���$��L	C��f��w��\J�x�8L���d�B�O 	��~��Ƀ\��8��7'�?�܂�	���"���&b�K��zv�H@g!ڵ��f�#�u���RN�D����Y}�ܮF��{���=���h��vB������P�T�"^���6c�(_��L(�������tm�x��<W��/�/�,iMO�(65(۹Z�q#�7�W�(��_��|]��3��fcp0��|�MX��
\����F��R�9��#삁��x�%�Wa�ʟ���`66^�6��G�v�O�єsp ���Q&���ӿIO�6ϸ���Y^��}ؒ�4�x���I��^EÕ0�гAz��c����ᨽx�0��=E̤�WW.G74>���[��˲�{7�S�)��A��ְyP��xJ6N.�8<7�M;�����B�HU6�������vAM��x�'f�j�jmƚW��R:�&Z��7�]�F�h+K+�Z����B�u�g�A���O��z_u�キx����]C�bG}��K#������r�͙0����$��V����F���f�Wm��0c���и���C`���yIE��)�m��J�^�4��^�����(A�NK�2��+���n�f l,9{��hoD�;7�sZ��q�ܙ�Hє������_~H�4^+��
ZO�M��'mg�9�[ќ���*�5l�������dR5h���Ġ,�
?*z؜V�6E/�n�ln�ݚ�A��
�l�c��xێ%��K��7���<,
���%�	B�C_� �r���L��_6�8�T<(Xjx�ݤ4��c/���/�����LxP��3Y��S��:B��VR�ac0�{�k��hQ�b��y�SGu�ɱ�m���B���@j��SkR0�P�b�/��������>� #z��<TO��R7��quW��jc��tI�J~��*=�&.���Y�[�!��|z94�����s;ߵ�{��{��\,���]��u�C%��m�m=�1�����K���r&G�Q�8�	����C�������eß#|���㧰�.м �nU8W|D��2)�D��e��6��a���9D���n�����D�Ab��C{0�J������D�O��0�U���n��n�K�
������`/#��6���^��j�FT
Wt��& �o��n�7�Vk(%�����˺����P	�O�KJg�5~�t��#�{��4B%���p�^�����R|���u� �c9^b*�r	u��c�C*ޗ7�����G�yh�����R,G�}���7u�b:���Ҩ� {��*9(#�s���l�]e����
����$D"u_�Ʊ ;҉'�.ڢ�xK�����d9�n/�KF��ۢ�}���W�V%�S���Q%��"� P���
-Q�Uw��V@�WJv+ʢ�a��eU����nf=�7�!t���v/��7�}�4��(�=^�[iS�FS�>יd;#K��&we��p)ܠ�r�s	��Em��]1j��+�c_�9PP.�+�&�=�6�(��$�T�H����P�G����׍2�=x%ɕΖ� �T4��Ԭ��+�Φ�5R"E��]F�����Ng��/����3	�`q2~� �S�ncRV��٪��q���JEZ��XhB�s}Gog;o��$��N�t�T�sď6�_wm����H�K`��OZ��	��68�-�iH߾ʧ�W���eC���7x<��R{vM�����G�zؔ\����E�@��9-2?��#%�:��7������4��
� e�U�k�·	��F#�ݛ��h<n�Է7��Mk*��o�hf���F�?u��{���i���D�	�ݎ#� b[=]�hq�X�'2����.ܓ��*���}�#%�z�n��8]磼�g{
5.�����;z�JP�|﷕x�狠@{���Ͼ'��o���(U�n�I��i>���bn�pmJ^��8j�梖���}?3���V}�We����X�&o#칕ב,�rM�����k,7�y�0)#��p�����0@�U��'��d�g8�Q�҂	E76+�nn+������b�����Hs}��(; t8�������j�8û�i�5��蓿�GB��o�ZΧM�C��*�׳[S	�S��.� �r�;1տN_|l�*m�Ԛ���1�#�a�H�ݰ�6�"�Z�]Z
r��ٟ�e��/v���s�?_�����@N]'_�'(�e&����mu -��\���U�tթ�����V�\��}�i8[�d�'�- s�i�_]�M���RA]�:=~�9�ʞ�3P��iͶ����(cE�M)z��#u��V��˷"աfk�rT��C����T�c�0��
��u�	��A�e+|�ڛ����4TE_��V�n���Evu��`G���S�������NFY����=HíG!mg�k�7�.��g�s��ږ1�w}D_�����w��j����`�	D�_���9�w#��� ȸHHIwk�7�0u�P��IB��'��#�z���S`�hA?<o`I�l�!rh=���b�:^���b���@���(,O!��.��r$G�����RoNG�)];Q@�7O
��[DvF0�ֵ�]�?��!�د�Z����������5_ F]��x���̏l��U����JQ��T�M��2�]Mn$�M�1"�q���s
B�5:j�(���x���v��In;�H��o�c`ֻ��G"4�a�?�� �N����^S����K�i�e�D�`�8ȠĎ�Y�&3G��a�KЫ����u0��p7h�����ITݿ<��U�a�(��T�K�?a+ �E5o�A�-<pђ�[,�'��j8�$#W-kM2�zɈkX�s)n�B�V����UWA�����K^d���W�C��׿�� a����� �Ok?������N�L������ ?��zPQ�܆�h�2�	�`�`]i���}��E7Q�������py��� 2�3J�	�R`��g����N�皙��W�2���|��	�LjQ��P��{�ڪ�ҟx_凮���6^~�W�k�4)��A�1l�<@�KIŞY�e��|�%�� �jS�QOjS
׊�Y�V��7x���G�9O,j)�auBR=�q�8�E�c��c�Ꭹ��t\-��>�
��ܫתoC�B#��Ž��{�,�l�����T�>U�7��~;
��+j�C��d�	fQɭ�l#���i�\�V�J��@�m� �e�;W:1'����-��g׎�V��m!�{�{��3�[�9I���$l�[_I�,ۇQ:���:[l�c��q�Z�=TE����w=�n%wt��-�k�&5�}��U�L5š�m����ZQ��݌i�;��;�������s�t?���&*R��ꚍ��u��Y��/�7K���?o�i�ZoN�(P% S���=�k�����i�k�&Im��g ]�_�\��D�(�1D۝�.l\)F�������3t�r���M��,j����s$-r���#���D-n����,�����\pnT�p����ډC@V�{?Sk�������v4��p̆�w e��5����s<�lc>jߙQ�fǧk�b������Xo�lq�P�RfX롍��5#f���	k�)�"+K�ʻAlŏ���_�P�0�B^�X}sp���f��Z�B�!���C@�Kz��ӯ�9�
�)Nļ�y�/_@���&�/����3B~hqO۸ID`�˷Uri�nC<��]�8D�_��81;����n1B[����L��ԇ	��6�ú�{ǹ�N (*�� Y�|�Z|�	X&�j����g�,Ν������F1��yl[p��������9�i��� ���w/m1`76;����4.!��FQ,'�vT@ކ��6�6��J�'p	E|-���]ɑ�exfQ����@��]�8iJ�<@��	 ��T�2/C�Fq�8ΕISBT��&:�$��m8�Ċr��{��y�7��M�s��ո���U4"v����E���x=�tk���9��ś��VC��RO��Xg,f&��'5��b�`����]0���V3�P
���žAem}�>ڧ�f(E�W Μ��S>�*�G;�O�9�V��S0[��ߒ^=����.&�`2�z(����h��T#��o=����k)Iς1�zc��a��Z�d������(W��i2��4������!�~L'��l˸�PJ�� ��JW�~\���������:7a���3:l��������8�t���*���:>��K"�w9���ň�sg𨵿��<^�)I�t`����� ��^��p(�`�+��߻;�UA�7A,�X�(�,�55_�Ͽ<�PsB�Tw�3{"�f^Y����
#��|��&�:V{��±�S�����.~R��;�.�e2�:�O>q%"Ro��X˩Rx����Wdo�:�C�v���U�[ DذD�?S��L8y���:�\�tMua�;-������v�`P#������پ,*,߹�Z�m�D��f��i�����ϊ�-K�텤X��S�n~�y�OQs��?M0�r�ig�(�Ă�j��,ٗzQ�6�H_���P{H8L�$���u�)�%�'�R�O=�¸��h���j���ad�U���X8N�4��ֶ$�S��$�-۹��5@�̻��(�换rc�ꂖ��W�R�#��z��
�/U1��������o��B��&uO�u61�`v�	�f)���2�&��ӂ����8��Q�p��c��ԩw�(X�2lQ-ЙP�Uag��e�v��#լ|.r�g@���X�|ְ+� �iC��-�+�O��4�e�#�������9�2���tv%g%~�uޏ��zޞ��ieF-Ii�4?$J�NU׀%����W��2�}�.��.~x�l�(o$3�+Y�o��%E3�?V�q��n����"��~��j%?���Ð�ś�3^&�o*�?Q�/tU�
:�Y	N�50-9ϴp�/�̜��/��`'���H��S�An�-��
�Y/��DEl3��w]Օ��+�<����SU��>�oƌY��yZ��ٕn���� �ڪn�:Sa	��s�^�MN�"ۛ_��ݺݥc�Ih�����9?�FE<-p5 &x���[Aw��*D�0Γj.c���k"P��i�x�6�$�aA�������;nA�3��r���<j8�;nՍ����h0{H�L)4NEAl��E��bE(\��'���,�1B$L�@�hS�&X��K=W�,�_��nm/j�8/@ٿ���FRA�������W�	�#��4F2��/^���<.U��UHmD�+,�sR��T���&:A\��a�#�p��P�����GgWG.�TP��*=�� �bդPbK�9)�z�2r�o�o$��ٟ�%׾��!�d"K��,�~К�ּv}ga����	���A���$�_��rd�������|N�^(%L�Z�\� �%����T.P��O�w�U�0�HfV�i�����ǎ����ƹ���:G�!+'"i�ꥥn+����Rg�:su8�Au:7�=l�Ԉ��x��_��6���J�b(�^��qqK�%�:h9�D��vt���(�yrȿ�!BԿ6Tr��q��%���@���~�l�X���
���WY�m�0GI�4�����h�˒ � �����D�@����r^H��9��v��r���X�5�Ħ����?Q��}��_�����q���jAH<㠧���'�4sj���䐫0�M�S����v�w�y�J��H!=��cxy&A�m)P�[0�x�/�.U�qdr�6�m���n�Qn�v����<v��0�Q�t
��Ty�����}��N`^��r�E�@C��s����G�{��H� p�o�9�D֧*�}	�e��$a�Pe�Bd~R6<ȸ�h:'����6X�Y�la�ȟN�(��@c}Fyyp�i� a�R]���T�?݆��
�gѺ\?�S�����~M�Z�������ɁYg��yhI���նP��[]�Q�i~ڷ�y5�u��{�~�9���F�_�sC���Ps�)�
�߉uf�Fh���V�-\K��6�8<��/�Lѣ�dvf�D�)nsx�T��^��H;$�f�{�
�#�,�(U��C�Cg��@��.ZOO:mqH��[�$�lQ
"O��n�TF���uw����	G9~#k���Y�!Ќ!��+e�͝2/��A�tZ�1��
Eܱ��$"����D`v�iDR�a>I�`X���ti�J?Ry���	�/�)��M�KS�<0��&���)�F�<�ק�L2%S�-'����'��Oj���Ѷ_�S��E��q_B�",��w�mN�^�S%V>�:t�#mMx��Rpʶ�x�L�8��2d��A�)���i�2LM�/tRct�FWc`H��+���!B|I��?"���gU{[�'T͒��n�.��Ƚ6�	J��4��������Y.d�Z��o;�.�g�R�+���,IU�H�B4}�m����+�Μ򧔎fI+�IX'0�V8�[�ti*���vj���d��H��\�'W=96y��]�Ks��}Q�G�`��������W�,�����m�Ғd.�����(�@�6����5����Of*�~�`�D��)ۊ�����a�u:�zD��p���U���anܖy�y\�>�(��!��-
/ܙ����7����2�1��ĭ��W���QU�X��!�J���k-������/Ny����nv�gQ9���2����u�����h�%�"��y>�h3ز����$Z�Q�g���h�m.����WH/i�/	��s�|$	�(൑Q����E�x~;?'6��ZARE>��q7t޽uƟ<%�<��O�1�IK,�����a�<+;;Y���k�y@���]ʊim��D� dGH�|��'���c� w��,,���8K�>��.��M�y^`�^��MV�B�>
%�C�ɬ��Ʋ�kؾ��0 �g��Ix�=x��!��`ms0JA�T���I^Dӷr��O���6�`�H��{CwP	"*sg���*C�"?x�91 @��p�t�\��F����vk{�U�2����zr2���zܐ��9�>ŝ��Q��!��֙�P�M	p��~�'X{��i�������YZ�*�_k�A,ʌ�޸"�
�#C����$<�jp
w��upM.�ɑ���v���\�d8KW4&~�'�_УH�P �Z���"m#8T�(AE�VV�A-s�ҫzT��)h�>�_3�+b;��є�96��9v� 憽���3\�y^��IU=.Vy�ʯ���8	�y�
�'�h�`S����<>�V/��c[IN�҆�ǿC{L���bےj�)l���#0��.��$n�y4� ]��-��gi��� ��	p��?,��$�+���~����q�Ƌ�h�!�ٮ��J ��v4��\	c�.^�8�X��Ry��P!_����Jv����(�!2P��?䞒7�%��^��x��5�1,�
�'0B���*�
KfF�	�T�A��^�&��,�w7u��Ę��"��l�W�>E�I�{�C}CaRQ|��2_�����\eOU����,�.���Q+���n@������~j	ֻ%{�Z��A�XH|T�:E�te7Ś�G���wo���u�]�R�Q�m5ϻ�r�y���	��kqJ1��m/h5m�d,!�9N��0����K:��z5�Ӷ;���'=-�İZ��LUwY*i=�$�1��H���ڟ:�n'�f��mEα��q����%�e2)���?}x�����~�lXeζ�|<���[�W�R[!��\��r�_Fð�ʕ��-<�r�F�)�Fv2�{o����H��ݒ��x���"=�~e��8�
0c����Q����4��'8H�������C�dT/2ô�,e&FJ����B���7$G��`�u{ P�d��P\�^����AЂBMgvLw�s
ve��	(�7����p�\27�z�p[����dF���Ts���'f�a�����{A:H̖�єK=��O�K�y�Z����i@������P�I�q���)�ST�2q��eh��Ʈ����۵�@�DyN��]װ���]n�|�dc9S�� Z�|� %�j�,y׏�4s�,߃^h�l�G���N|�+����z�ݠjO\w����.Su�z�|*k[�&?���
8=���z�`P�EO���R-R�S"VCȚ1$�g*��W�-�=hMYs��e.�"�L&#��)p§�!%���X��3�OW��
w�d��U�P��bH��߭�kvى4dxp��+��ڸ�1]d��7��8[���VЉ��+�;�?Vz'��G�3��9Z�e��)��O���rd4�O!�MFC��ә���T�|��+j)i�V1���j��t&�=\�It��,�%4�Tf�J�"��H�أ0UT�r��_Ц����;����)���ޛֿ�p�<�Q6��<5u�c�mv��Ԏ:Z0��^O��n>���ӷöh%�u�#1�����q���>��t�#F�C-wڅ�e�0��)�+f�nw�l���xE�۠U4=�J�?��{&��Q��U܄-���l�&���Qb}�?U�/��"���h�{�k�N�h�!N6�����ua���}��?I岰�w�����#	��c��s$��|?rZ�9�
%�7]��+)�^T�l]�������$��c�n��_]͕qbS��r�V|(l`�͆8L�)�}t��Y~CU�wd����E��7��a,>��>��t�&�!2� S��͹��k���0� ;]'"�Q���"%���=��+M�b_�]�d�;�W�O�v�K/a���Ԋ��H??�n�l]e���eb��M���5�)1�=`��m��+NE*���s��ë�D4�����1�"{��u_�|PlI�v�dL�S}]<����9�>S1ץ���t�І)S����P�	EW<D�)���>�!���d�`]�(���'��^J��n����ѧ�DpuI���ǧd{hV3�dDŤ�`s�{����x�
x������7]�tD[p��Ζ6á@�x�*�3b-��������n�J�f��nr�MC���$�>`�N�=�j�t%N�E����,![5��-�ј��#����ϱ-�[]=���������m����r�q$��v��u��������YeH@�fw�Y��Г��y��&O�����hрKq!�zbAyOV_u$/�JS���oU�D�zo-bd��WL�7*Ic��f8��w�rY�E�c�~���#�s�k���Q;L��C T�)X��}'�0�{m���Q�\�@/���HQ��GnXP���4k�;J�'��y��(kb䨚V����L}��vwWY�%�0�@��,��+��e�B�h�@21g8��u��w�>N��&X�r�z�D�Ы	�-��_�TM�<<+�+�����x@U�%3Cdv�I_��_�z_���(ɠG!����]�����`	��,�e����fvv'L�o�H���4��n����Р]����Q�B��ց�&�<�8�-�T�"櫚<����������U�cv/�a�蔫���2���d����q[�b3~��\
�-�mRB:8D��?��?<B��S��+��{7]���)|M`�n��my2d�+(Y��Y�c��4�<p�C(����.n+x�"e��C��	�� 7v�z�W׏Qx|���4�E���C�Ɓ r�E���1���D��/$G�5��ȓ��y^g�2NR�Z�Dh=�h��r�]Q�˸:�ޕD�!%{C��aM����u�r�;����Wiz4���G}��/6�M�>i�Ǿ3��`��Ԙ�w�x�	��F��Ñ3�.`y!MU7wu2L�9߹Py����8��xQO�'l�:ʫ��:K�Mt,�H׆�"���qt�ox�g%s�ǲh�\�����.~��:�0���h]
����
����i�����gS_p)��=�:�C	F�	�p1�mG?H�r���4(F1'j�	[K�z}*��w�q���v�1.�����bW���3m��Ks���g�%Ò5*/$TI�=#(�ӌs>h/MG�\������i@aĦȂ��I���W���� �"���}�-9@��"_D=�n奸b"�Өv��7Vv6���)79�*�Vq�[��Q��K�Ta4m}��>����CX��"�D�(}@n�d�~��R��Ol�Ĩ�B�g�h��k������}��\jP��:s�V~��;�a	��,���w�7ݢ}:�o��xL[ӣ׬��67u3`������ 2��I	Gi��q>�+��Yk+�a&���L�LL���~V�k�V�2>��][=�9�r߶USuEv
��b�(�JZ�P�97v����ԁ,���r��Z�:����OPݒ���%��:��̏�v��D8������~YO[]j��W'�$S%SW�S�L��!�,N1��ﶱv��͕g��W��"|L5�ܓ��x�����n�����6����,�ľj��Y�����XG�Gw���J��z9k�������v�o��<�1V:��\�=����9k��-
��_,J��k]�}G(
������J�x�M�QT��jo�]9'�8���q]:II^S��{U��{X��y�̅՟����.�����@�Ē��d�]�%{�cE���c멂 �7�$�� �d	�Y�~ǌE��:�]\w�8��d԰� ��+��,�e�A��y�..�H����~��Aj��G��5!!�춋�CIq���
���C��nXަ�=�	�<�{M$�bk�P��$:�C�<5|�!�Ч����×�����h���^^�N�Vcc�5G
P5p��3���,��$8�-���ڦ��J�,[|lK��M�-kZ���"�ڨ��~{۶%Zه��"$�����pM}�0(���?a���#.~�����Î���q
l�����u��@���Y�ͭ����vH]�z�gfA:�K5?�b�����I�J�	A�4�	`O��-L��54r#�Ɋ��aŴ�^˟$������aR�0����Ɩ��Q��+����]�F����������Y�V��t[��M#�'G=��jH�����P;{oD���f��QX����[9j� �b�=É�2�bйh������b�X�U���]��гb�,��/O��3)8{�}����וs\�vpz�{���)'5�/>��x-ʰo��˅&س+d�meŠ&�#��|7�������p���0�m|a�\Fi2H�]�u�����os�;��K���7NH��e$��1��_ղ~�\u���T{���r�v/
}�4șSb��:�N�G�lk_ y�ݬ��G��4�f�Gv�J�����!*�eb=�ie�S#���g����O�a8ԇ��������Uw��_@��9[���.�FdpHq���.��5|����+����p�.C$Q���s��@S�'2��{}5�+j.>�,h�81*�}�R�Er��ϒ�����y�!C9��j9S�G��dg:�����f����Y`Jkp׺����L����)�t2R�y�����Ϊ��
��ֻ1���Fځ���z��0gTjp�e�*@�h�n�����@��}��k����D��^9O�f.0Ԙ�������B+����('��/�����]�!����_n��`�8�9�y~Lsٲ���a0ݒ����E0@3iP�#��86�et�6A�,�F��6� m'8�%����U��T@Sf��d�E�c.������zIi�a�z͌)���6���#����Nc)��WxFp5�5A|'Y�i$o2���#�]bC-n@T� J�I<���&��g��˷��uR����'k|�9�A���]�ߩ���FS�΁'�*�؋+p��PTu\��%|
�s2�	��嘹FQ��i�E��P�Q�)6��H���r7�.���Q�`�������,gie�u�������׆[,�"6���Ⱦ� �P�j�P��J��TN�bъd��,3�#˰��s&����Rb��ˀMS5OA�5���.��q����v���S�G��ETt��碲�����(��NM��|�ٙ`R���;�����\������H<�����`��Q��m0�Rz��c;�5!���:�N���q�l��q=�vѐo68�;�������("�;s���I���"]򐰶�+����Qt�A)u[���~�%���Ѭ��\Q��LKG�[#�M/��Hz.�!�9~5�C�\t{�.�X�Z��x"���gPa��h�1c�w�Ͳj4b�����6a���ȕq�9ࠊ4�73�*뺗�N���t��`������D<>���ь
��ԣ�)��Lvڮ�i.���FD&��NT8�k6z���fqx�K�U����B�j����غ���0�2e �i�,�bms����x��i�t�H3����P@'N��2�FB�����V��)�;d�J�,�d�B������������C"ֆ��*�GP6�H/w�=��i�Z%s��J(/ȁ6��0w<�D�:�ަ;ݱ�ߠc��`;8^@0�F/��6�uRߝd
��I�]�������L������do��Z�Ը'�@�X�4�?��~	��szl���,=��Щ��ę]
#��iY̆Vd,�L�"Gz��K�?r܎Q'�an�N!p6�?��l���V�
��� � +�f<!s�`���ȚÿC
��0!��r;�_���uVXpa�L�:�
���V�Ŷ.$���͋x�Z/gϗ��BԤA��c�@5qZ��v�#���0`1	�>�&�:��߃�1�!Y�{�p��'��EM�2.�)�~M|��&��,�^����LjQO�w��~�*g����e�������Y��h�؅���+)S�V���Nu��Db�F��M��Ջ�z%�?��ALezTХ/��ӷ��f� &(��S:IH�!�~���㚈`UB���M=�UD���n$=˛�H���8g�j^��e�0gCJ9-�
DK�ƒ���_	�2
�#�k�.\L�u����X
K�F&�xCr�Uɍa�4�h�#��q���I��H��d<�I.��<d|xem��J�x&*�n���/k:�m�͡�X�ݢ�� U�ݸd葳�F�|�]��pN�{��+5m�����5UUu�)�~��^'Å�6�]NoqaW`4��H��c��*�DWJ���_����� �G�J
�� ,ʺ�dY�`���5�X���s#�Po�Ί�I�l��yx�wT�w�t0ܢ����	�s��Tɫׯ�OǄ�P%�H���D@W�]���WSt5-D@�����*yPP�J��5(
���:8���Ҏ(��c#5{����C�<g���6A�n�q��ڄ���P�
!��BA'��!�H��Ry��t���Z՛��6w�?\㟣��}!�.	�2��M���c>q�d!ַ��{��[xR)R�B �����#�����$M�x�v9�,��T2~NMx?ħ	�:�W=�8ؠ�d&��Μ�rH$7[�� ���-Ԙ,y2fP�`�I��� q�aÊ'70�%"q�Y�`�<�<�����}V7�rS�"gߒo@���qQoD0�� ����D�e~Y��˨F���1�
l䎾�ٰ�;����;�!�o���#��ˑ�qBK���5�d�/~����or��l�D�B�5�j^�y� �H%��GΖ
b����]-S�?b�Qp;����L�D�iqc�ߖ"^<H��I�}�6�+�Ե�c��|�C� NC��.~úk����^:�*��@��y��9!RI�W'�oheTm��l�q��ko���zɰ�cO�QRib�M��1�z1�{���l���b��*_qMk2'�@��~�[�&�C��y��Q�!=y�rwjE�a���YkزǬ� ��T���[�!�O�'R<���%��*�˫�z�wm=��J�����jK�y��$0�=�ʫ�ĭ��U���2��H}�w�� �.�ĸ�!x����՞_�?J�NA4��ғ��癔�cW
i�w�/�~_�D��K!�R���ǟY�wD�ܥ�e힥���>d.^����&UC�4CA\Sbײ��8��;Q�)x�Z�d�h��(o�.	Be�ۮ��χ+u-��+bRZ��!�F �.}  i$����c��侽>d�
����i}�o��g��وώ~�p�O�,��A��]eV�c<�t:D�ph�*l�2+~J#�C��D��k�gO���}���S��XRc�AAu(o�&(��Q6��l ��'�,�+�o�dw�+���D�B?{$?��\Wp/��.cp�OPZ��NQt;� ��y�*ߚ����?���9�2)��G<�ۯ���Y�Ӓ��b����y�\�X䷴��3T�}�(�#ra���c'�@6�0����qlۍ7KoM��{#���e��q�G?3ޣc�L�AyB>![)��݆[�{ {>�߻yt	��
�(��l�;Ӈ_�i���0i�p�"��� ������Z�b�=��`F���_�,@Hh"�A o���l�,̾'*Z�fy���Ȱv���I�鈿x�M��B�PU������EKX��y��^�X�1�~��A�����sJ�x$�kR�63e$����g�*�ܣ�W� �&�f�s�qd���PTEW��2,bhC�V�=��c����fKǨof����vat�7Q�B���~7+ܲ�7מ��oi퐁��^wHUn�(eZ)|�/�r�>��Ri�X��v��']�N�?חp�9�pܵմOT�}���V�我k�U���&�F�|��%���F��"�f8�G���<ff�����)�3y����"�VJm���/����E?*=���P[yD�0�:�U~�$��O yl��[m�W�Á�B��8��ih*���ʌ��g�̨4��SI��`߃�5Hp�����YSM��#�ՠ�������7[l��u�_� �B�����6�W}N��d�[~}_c}��@��) ������4l�[��:QT�o�2�����8_�D4@�~�ca�)�J�jؕw$R*{Ϳ�V��
�����9F�X+i�^�6kW��+��E�7>U�����1����E7|���v����R��*�3�A3+�嬺��7?o�
���2�'�X%�����X�/��FP6)p�m�)"�H�c����ը����8ok?T���F`C��{IS#����P�(<�r{�UU-c�	gI'T�E��d��9�����Dp����|�BD)8���D4{#Y�A����dIY�e�s�:8�2��S~	?	�L���7��m�B�m8(`�h���9ȸ��O�mW����"� >�=Fť�Jpث��]y��Jm��@ �ډ�y�3�]�<T�9����y��PԜ�a�t��sea�� q^��j����`7�L:��yf�*�'�]�M�m)D����P,$o�o��eSE��h����D�{(���M�g �����nAB�y<M{�V�	z��ُ�iM�����Fl�TL�>�\�K��Di�4d:�;�rN���4�5e������ȧ���)��jRf��@(���t�
�e���5�0vA����;�y�v���[�X�}�z�	*[��p�nTP��/�ۧi��G�|䯒���8����ߩP8�y�:�4v���0�$��zۧʌQ9�b3E�&Q����6%��'�zY;���x�0o6.�@j�m���Qn�+ll��̲��`<�d]F b��:�-[Ḏ�|~䲡���7Soz����S7A�S��/Bgք�B�sH�*,b�5���5���$6��;쫖���YH���'`D�cչ�L,J��M�� ?^�L2�qP�aF�w��"&���ͅ"�%�`���V�kx ���ك�t�7(%3��%I�-4J�s��c�zYoے�t�F��0�p�|�+��]�7w�֊��\�I�O�E�"d�^`۵�ɐ��J��Zs�����Q��3��_�5� ⇢{~2e�w�����P��B�R"�'2�J��k�RP���#���4UPP��7�˅�5���R��̆<U��Ήf���xE�oe��*�jV@ �2��򀎖փ���3]�k�ȍ�%9�U+����f�7f"k�Y�WVB�vͦ=���%Z �`H}:F)��B.�i�0%U�����*� ��dp���9��\�0F��wm?�4F9&��`��g��q�O��1&�4�R�._;�A���(�Ń�s�oW*��떰}��C  S��P&�(z����)�̅$�%X	�za0h�cz�+��)I6??]-�AW����Q>4'�с; Ǧ�	�`YS��H��+,��
>����L���F�\\<?��1*�L���P�c'a!�F@�і[l��+|!�c?��N�-����i!f�G�<~�L� �U���DZ	��F�8s	8R�Q�J�'�\�)	��?�[�&��̮�:�[�BQ�ЫPFV���=d��[)<��>I�mǺ�]Y~�lW?��Lm�A.ڏt�N:D.����'ц�AY���	%>�N	�'Ј	�.��k�+�3�=�X� �%)ݎVf�u�PB}Q	Y2�/M��<yU`����Q��}��Iw6�P��+�L� ���.�g��}�������жl� �9e/���V��a���ǿ?PԮ3��ԕ �l�)]��ϭ	=*K5�2Q��>���������YAt.+���\du.^�� /h��,�^�t}�[��$+�9ϚZ�֖����>$��
���4�Yn�����
~C��vj��2����E6���AU��6��]�V�l�Pt��ͺ��_`��b k��~�$�d��	`1�<�0�}G܃����-5���^�yў�n.�b:�^�O�VQ��Y���<kH� >V�ޚ��6h���f�L����U���
����p��a���Qc:+�{:�1c ���ײɫCdI�G��ԣ�����ɖO<̃��G�a�.Hퟅ}�3ϝ�_KeN�,����s���=/��޴0�����Z7�j5h�	�HF1
P���(3�Vy��wr��i��A�/I�h!�.f���B�4��;������'%�'��������� ��A=���Q��7?Z_HjB!8������^ŬT���L�+����2��o"#ɔu~�
5�#��훒�`��3�>��K�H��r$]I�e�W*�޲�otx~�P�X��kcs�wǩ�p��ˣ	)�W7K-^su����]_���Ж}uW��-:<#V��av41:�5e&8��@��G^���� �Vo��;����޸���LP/��?J�P��+��nm���^q�E���䨜GBI�vY2��i>���M7VA�#�A�h�&�d�*EO�V�_`:-�ָ��v�&���Y��I,�%�m�4���ȑ�,�� ��D5i�n��#4�/с��T(�F�DQ=!mM-�
=ot6*9$���<��.i��7M�;��"�l�V����I鶡5�s�
�J����D߉5P�p��S�|P/���' (��ͦ��Lxlbп�5�(w�
�8S�pR�8�+4S��]��I	S||cS�V�ba��?�A�sA��
�\o�vsR��J!u��_"r�n��n�Y�{1qh�Z�`��|Q`#m�2T}(~�����nH�<�
�=O�4g�ڌo�k�d'��䉻�H����*����8�9���B=��K�6��{�\��;.6p:�N�[����j`�J��	Jo�'�;2_� �l%�'�>�r������%��Xx.N��ȫ�է
D�ނ�%� �)�T"�1�C$�*�����Oa�3�F���Tޞ4�S���;B�p�|gOϢ*�)�m�x.�+���FIцFr�9B_..{����T�f�1�	�= �q�#�-�qz�c>P7�M!��Qu����}�Ä�����izD�ܛ���a�����;�^b� �P?[�R(��֢
.O�1���娽�h��x&,�Ã	���_���A3���C���E�׉q�<��a���1U ����ٻz��,��@�j6�[�G�[�Xs��$.�_qks����4h6�+��'8[d���Q�G��lB���P��6�7|Ga�2�A������V|�c����Z��D%^�6W���b���~s㌺�#�DyB/�4� S�,�m�*�Zd]����\¾U�!~)|��E9&QE͌n��
)��y�p��sh�<H�ǔ���������0,~s��Oº������W'�b���2��j�Xa���|�?wn}����;~fS��pR�R�AbH���2�'�H�f�����}��*V5�y"�b�ʠ�ę�
&b��T#7���[����]�a&����_�0&�1�w�65�CV�ls	^ԄPc�DG��,f�mɃ�n�|�<��:�k~��DNF���4:��M���W]�{�[�^�a��2��Vgy~�*h7|==��.�!Urb$<���R�u���w�����к�7슧����d-��ф��K�ξ�8#K�zv����1{Q	5����v/����{�$ȫ��O�JFRQ� $����_���V��r1�%�z�Ɩ�틕D���H�D��Zn�֯ ��A�oJ3z���J�����}�Ru.��#:Xo_��@ �_�#��̺"���� �yw��t��]L����Ӧ!��|RF3T�"�8�*6��#0��P�2�=��K��!t���s�"�_�g�]��9b���Gˏ�X��/���q���h���P��E��.����i?���
�xH�^y@�-���K�kc_�@��Ǽ�Qݸ��w ��c{�b� I�r8��>�j�f��O'mK"̱7�n|֗�!E����z�'2�#��%@?6��$�1�p�0�żq��7ŀH%�_�g���uB��]3�W2x�ŉȦT���̭'�ǯ�S& Uz '�Qk��# ��w�]�����&��\�ͦ��9[؏���Y#�ʠV�pz���j��N�^���H�K`�+6:�,D�"�k2���*�%+��{���F�^�����~��C%�R�zk0��b7?v�ğ�
�� $w�۹*u�k(�k��"�q�{=R8e�u}1���v'F�W~��7���%9�R7���_�E���?y�H+��v/�s�`P"Vk�M�E���bM�AElp�����<.��%�sl�j)!wZZ���߃�)߲g�D�jF���������¬`��.��S��\o,�%r9qlJ�d~H9�x�W���#�����02jj��3O��sq:S�XtwF�AЪ ����|�k���)�H�F�<.[�0Uf����	U� ~y�.UƼ8��PU�Y�=����v�V�}!&��C�6pjч��zVY�W�ü����Y�[�g�C�@��7cbY�����;��_!$#�+��H���o�W����8�7�s�@�����ޞ{1)��F�]M���	��b��̝���L�-
��5ޏq jiۍ �����@B-�^�îLu�1�"JvG��촍�G�ȋ�tY&l�'�D�#�O[�ǰ��;"'�rfd䑓�
����{k7GK`��x�^�Cn���Z�h�?,��@
Hd��:�4ë�چ�2%v=�X̎�e��Q��5g�/<���!�*JQ옣'�5���2�ȃ��Mm��Aڌ���]T�X/&*
�kWզq��;A! w7ڙ�=��ښ�}���N�Z��fO �����qY�8/DH���i]�� Fꗁl���ᤝ���YetE���{�
��T���:P�۩���D\C�˴���L ����zlz��\oy�DSӫ��u:�G+.��
I��7>_�	w��AO�ϕJ��Eܸ���TF��G}IU���ވ����������J�{��?/�o��.�$�s2�xw�`\?��Π�GX�|��L���h����B�;�ߏr��#�,����ŵ�M_X��+��(�g��O1��\&��I�58�^���s�R	E�٩�mW��ٯ��	�@k4ۓm��έҏ�ng��/,��'n�;��=q�m�����1�na�~���TO!t��=G�1gD�J�}>0��y�A�{��������!_����L͑~����EM<]���FBl�r�t��w�=�1��&�,~x�3
�S�>�f�i�(��P����y���\���~k͆z9�%k>���2.�w��F�Ͽ�]l����VЊ�"�����cG呡2���ס�˦�R8h�<�ԡ�3-�!�)A���R���̻j/���k�J�����c�c.�ϛ�:s�mɈpX	G^=>��{�B�AL��oQ.��0g��@�|���<��+����=�%�cl��u\��E2�6{F����E`o�^c�A���DoW���~n���n�6�Al�Q�r�����ga�����Z����m�P	-$�}�)��8�v0�C�,)v�G����T��w8�0xe�|��[L����*�����J�k�֊�Ǉ���𰟪GX��l]���Q�R��M�_�vs3ө�$�-��v���nǺ-�+;<�Pwr��!`O�wXɋ"�N�|�p;f��ԟrIJ�z�Z�W���,�V�.��̺�]�h����̗dfD��B(��|4%�5NP�H2�\�K� �y��~U�x�[HP��wyH���)�D���(��jѰkA{�]v��\�Hq}�\` wh�]���2��Sl���L�׹!��v$���Jx.�+�� 3tR+э0��b����j�WZ}�!i�c�f>+�в�nQ�[1JA[�z�[�]-�S��{d�.�4����eKܐZ�qi��U�"��!y<�g�2�A=�G���\ʚZ��w������)�:�7l������G���i�[�s�F�A$Ա!�0���>+��q��{��u(I	�`O��|W�C~8������#.mb^4�s�/�X$&T�+��zhN*5:��	ۉ��a��$�T_����A��
����*8�$��5�U:�𥇡+�3�Y|�Ű����'?2B��O���|F��z
"aU�:�����>k:�0�
o;r�L���҂���H�cE���s9�}L����k��S�(SN�>�&�8�P~��^��G�fd$�vTRJ8\Ϸ3�H��<d7i�t02����s�̛&h���PV(dKb�a���jdy�}��sm�XEM�w�J4E^������k��q��_���f�H���������Վ'�y��[��CɅg�#"��?C�)k
�֠�1�C�m��_�HaS� ��.`��T�����ϑ.�f���/$�~�0I��3��BiU��<)�1�BE�r�o��Z�~#�+8�,]\��!�� ����6
|P�=_�O��n4�U͠Q��Ƈ�K/ƍ�E��c��|��w�����׹�ċ�� 'Mu����*c�嘘EY�Om0�|�{2�����h������u�F{�����o�P�H��@���k'PL��E�1R~�^]��b����9��[o'����j!ͳ��ds};1�|�	��{�z�V�����^Cw	R5��]*��(<*��k
Y�*(�H4���k��Z+��I���	��Д��I<�ц��Z��/\T�w��)A�f.a�����c���Bz�<�}zR9�r��z�x��w�A�yX���]EAJ���W�7ea#�o'�7c��+L�fT��Y�z�FxO�$m�[�#=u����<�(ʓxFE��X�.��dza��'�s�9G<KEd����'*���U�މ�t������7�3r
�i�[��}V�=J�
�sz^��Ģ����߱j��H|%%��w�����9��r=�X��/�<�>C��j6�7�i\�P�!�Ù.;ٚǄ[3�FR���8<���!���_d��i.8ؕ�w���ˤ�~��:��s���bT�+��>��Om�2	
�b�9h�7N$�F�e]k�{ʡ-H�Y�� !����{�\�@�O�'�:���Җ��!T�Us,�S&�.�=�(�Q����§��8ӗM,�r�l>�|�� 
��&���:	6��W�����8����DBI3�cպ?uF��[�j�L*N6>Dq ���׼�ơ�Z��`i�\������R���'��#r��^�� xA�ˌ[eݒ���'F�.Ȥ���EF{�P��[P;D��l�|6pq>-�8�Ei��-���dU��+�k�C�����2A���J���E���ӂǞ^t�$��:�[��᥄�o _�;��޵@Վ~P?_&�0>nY�>R�9�>�7��LG�� �������%�D'�qQ�v�Ԇ6�L���	�[_٫�y���8\jR�t R(�)����:���e;�˵�|# ��檲�x��lc�_�ձ�I��5-/�2�~�_o�A�x� h��g�����>�8�Ӣ���z+�1�*���4�;w��_��O�
����~yxX��:�d_"��Nc�(;Y�FF���L[p&=�qR�����F����9�ao���E^!+�}�I';c��,@�C^��ae���K�5�V.I7�*�dP0��tvߒX�~s��O���J a�|.DV��L���,Lߤ��w`AFF��&M� EQ�ɋ!<��W-k3����1�bFa�T�?&j��$��:��$���S� A���%X1:a�b����3�Β�0�����u/���⬆3"��HUJ��72�%��1��=;
m��Dx��OY��p��&eM�z�K٫�u��E�$��)��]��+��b��J<�@�?4p���K�g�II�q�P�x������7a��u0]K�3��J�8�\4�;ͻ�kؚ�$$ƙ�֦c\�Nd�Ŕ����KO�ph�G��`n"�OW�U�sb0qػ0���'*BU�/KT����4�W`.� �u\)e�$�C�?r��+���}���(B
�B�i�Tz��:1N�P�j*��!��-!$���s��z�z�����ò��73�4 �$��!�W���]��W3qc�g����LX�nv��380�;C�6�]��Y���O(t{��ڄu&o����;<�k�t~@Ĉ�-���n�Җ�Є�4�-2��wfm�9^:p���V5������52-�^7z:����J�'_LN��Ǝ��k�S��]���Y�%���4O�ߤ.�>��o+1����z��g[t�iL[j�aH��[R%C�x��w��� �,�u�Dlv���R`��W���d�e-��5?�8λI_ �ɠ�V 7�#4����DP�� �/��%�`�m��]��=��(UY�=��-ha�م9�h��A �/wNy�
جPAJ�H�$ _��51sH���;����?�����[O�m/��0���յ���W^2�/R�7/�#9�o��
�i����.*�aA��1��x5���U 9�+�aS�S�'iw���Yw'u�?���[@��{1����pm0��>�ɌR{2ƞ�������}�F!�D�J\�	���n�F�疊��L�gk�D����Q����^�� �4ض��07����׺ٟ�>�d�#��$�8�
�<�Io6Y�N�i6l�6��w�GF���z*�������X�U�}���Q������G��>v{r��>����+@��Du�R�q���oύ�#x�b�~v ��"�t��eƓ!�n�?��S���H���jA�Niu�VD>���W�`Q$���2M��m�ON�2�����*rd;����گ/xH�N��2z+J*f���[��u��UŐG�K̤T)
U��"�8�F�j
�+am.&0�8�n���ĵ����ٮ5w1�*u���){'�,�2�?���l$R�?�s���pf�~XH����X�Bwn �|jꇒ��1K�"j�-��ޒ��܀gdPK'�o75%�&��c�ǃf�u	����9�O�H����#zY��3�����a�ӼbW������E7/hW9G�"�D!$�J��J�-������$n*��Y=�ْ��|��@[/�'��w����)R�e��k�FRؾ�}d�Hr9{��ܠ�ϻ��¯���IED��@vo��"6���E:wM�/i��Җ;�;�;��L�S�Z̄��Co	���-�������kc]�� ��y�cj�Ş�xZㄷ��b�� �m=e+ғ��#+�����̃`�<�~�J2���D���B��u��RJ7=����E)�}�i����j�ìF��s����;�ש��D5�ʕY� ��ڽt@PX�Zl5I݊���Ԛ��� ��Xo�������u��٧C�p����Q�EN���Z4h14�A����%c�̻��*�����D:m���iL���9��_��\a�=��qMw�OS�`6�hb�;Q��U,�˯�efAɶs��Xx\����Ys~!��43��Pf��G�a"%n�e�	>O-"^���q@��vZ��ƹ�a~l|I���/%6��Dʗ�Iܙ=��{B�N^q��j���� ����J:�6�|=�Χf�}�R�2u@��z+�e�읠XiDQb�z�ٯEK�%���El �L�nY�P����Ʂ���������0v����=�Dv`W��R0��Iǔ�\d�C�ǒ++fX���W]��\n�ClcTk�.�gƦ�%�>M�#�	��r����n��LX
��.(N�+���K��|hC�NC�wev��n��䆕dp����w��ݡ�����3QH|^<V��=�5�Z�J�-�V�@Ȋ�T�$���е�ӕ;t8֦ۖɂ8��@i��c1��
���b�*�����N}�r;�����g�Z�_�rM�RM^��7)�I�H�Dc�����~9�
�j�$���ȭU �����K�uu��SP>+��`�����}�:��-�A2r@��� V��B�p��� ��=�)M�a{��;�?�N$� ��Br���Dp�c��+���Q�fǊ��|��R$�U������و�q�-v������yW>�+@՜%+�HM�C��Y���O����<�=�O����B0�p��🬰2ø�&=��mk_
�ät�>,?g�4)_-�3N���!=�L�t�D��i98�{�D�ۼ��.ˁ�!�:7�+m~��s�~d�٢-�H��i��?�	ZA{��������2o���_���0���k��$�ܭ�V�lD>i2��2Rz-4�9���]�W�D�J>�R�>I�y':�K�3�o5]	�����t������^&�d���1:��9p�C��`�x�`-{�4�%.fH��^���S4����Lz��*.����MW�&:K%��5p�&������MP���x�V�J�P����C`�IM�v ?os�v0.���C+A��X���N �^ޕ'a�#��Wх{���t;�и�Y[�(�����1����!l�ee�;���I��9�q��t]��g�k��|+�;��fuBf%�W6e���	��Pj���4�ESO��X�Q�q����P�����X��探��U��XL�V-�%��3e��\-W����ytxb&����c�H�_�
,����!�#���#:�z�~����ӂ��D㪃c�wh�����;�v�Q���{`��k��u���ʖ(^W*�2��x�(�U����뽯/c����;�ru��|��D�9S,�J�k� ������Re�VX��������v�n� �j_0e�5H�j������z�ӿ�&���Zc����2�j)-�"3� g�*����b�%�����w)+>$�t-R9��V��>8�E���SJH/5�����B��S!�Tq����x��6������.���� �3��V�x��h��M̶i^V&�ï~�N����$%�_N��Y@n+�FC�՗U�\�RlC_���T�F�>G�,�
P�Ђ��h�������S���\�>��>,�%�j�H�x�Q�@�x��߃��9L�'e`MS��O������,_@C�K���*ˍ�J�ˤW�n��*{x(�Oذ�vp�g:^{�CT�ly\��暙Ra����"�O�C����-�#���ׂ y�*� �vGf�-��N�����l^A[����t�K�u�$)���mmS�lR4@��0�sU�vf�7�G\�u<0�ϞL~L��9?^��E�f�?ׂ;���*z���)q^M�����@J���7N�k������5�`f���qܫb�+�T�Ҥ��
�`TCG郏Z^d��2:�-�/�%��+�ߙQ�nX�#��@�Eh��GS�7``Y�(�r�0����U�J?~CVc�ϋ�2.�0t���!M�Ҡ:"玼>���-���M�~���r�?XM�c�8W�w	�I+�^S��Z0��`���e���NO��	[Ȅr4=,�j��^�$��.vkSEe���/&f��N��(�S�;�y�t��?���a$�΃��#{��F�'M~�,Ey��x�0"�����meO�\ߒ���ٜ�b@��)'���t,�9�(�ux.֢X��Hv[P�V9�w�*Q����x�Be��X�b_���/3԰�s�՝����l�,
.݅�KTy���aQ5�<�C�)�*j�	}�v��(|.��	�$˿GK9��ٓ?�"��5�&�%�,x� F�4�Y�m����p� ^Ӱi�m��BO��-Om𤇚c�Sb#���
N��9$���O�c��@�5t�¼��OOX26�XA����9
�F�"�څܧ�[8���� �Ϻ�T�*;˄�*,�pq߿��v��q�(�0NS��a����Gq�
^�-LbUzx�ߪ�^�1�4'3$M��b���ZC��Df5H��.��Pp��}�6;�Ay�<��,������u��so2<�k�@�1h�a�����V��8���B���8]d����7q9l$Y���?�L���,�:#	*�:z�'di��	#	45 ���4�x|��~%g/Z��J��Jv1CזB9Cа␧�]�oJƵ�����t�Do%(�Mb+��X���P:�'��`h���d}��H��O��g	�M�]X�(�}�t���w�#/3��}ۃ	Pn�U�er�!�^c0x�W�������g���A�k9���D�A��^��:Ķ+0�wl*��d���y�ؚ�;���((�_jN�v���n�k�x�)����)WWi�3����C5y$���b�*A�A��R;^2鱷�*
3�m�Z��>�b���;�n���O�<ɸv�M���m ׄ8�P��u)W�����px�>>V�R�u�76N����Q\&Q�횦�U0����IZ�m73W�ǡ}$:Al����nY��*��)�Z��`#~s���Z
��4EF���6R���0����#�n� "��M�}���N��
�+����V�T�xZh[����(����q��	�\(��7�ρ]M���*�2 Ǳ(�FT���ю���r�����!c+I�A�����hX4�౅���
Q�������|��>c
huV�A���~��@i����bpy�Q����+t�´�!��W���000����b���yu�u	�N�=�m8v��g��_)���tsy�'!27��Wy��ta�6XG0�8a��ݓ{���ӄd��O=h���,��Gδð�Jy�H��;]�����u���џE�=�wi��y�ɱj$Sj����L�C��J��S��5�Bt �7�� 0�����n92/����Z����E���(a��<��N��v�>�&���45$<�?FһY7���a��ଐ�Bd�8>Y�Z�WJ�����Ygj���5P���s:÷�B����x7G3J�"D�e�@��1�Ul��O q%��ZP҅��|r�$���#����dK�?TE��#!���N����+�S�)5<��t{�� ��CZ-uHHd���j/'~!���|z����7I<�=[J�!�B�g��6�_jDp�������ܬ8�zQw�ч�Tq����*q��!*S�A�(�!f;w!'p�>��mae/�&�S��mgG���z���ܧ�o�h�Vh{���F��Cbv�*�_@��@�ς�	$h��؊����u�w�F��~&Mp�����e�fP�g�a��}|���dl�.I�H~�'��l����x9m<�n\�/�qb�N*�_��Ѭ/�OQRw���JWxR�GtE��A��W�3�o��Y-��CӉr6����7O�-��^Gb��)TAf��uJBk�V�dUO��al551���~�M�w>���Y����
6$���ޟ�<��t{��3�>�S�P��>����P3:|�����
@'�Eg'�EN/������[r�v��E���"Ld�6`Y�6� ��~y�D��@2)��JԞ1�xp�jpt�d��VMcz�1EY :���h�t�(q\���]�����RNdc `Q���l�]�'��/�|W0=�)�t�
�ՔF�]:��	�_�U,H�s`HO1����M95jf��alo�����%��7�oL�bڕ[�e��nfm���SpZ=I;Lw>5n�Zm6�u�6�שB��K:�����7�Sŕ���EEP�c�ų.н���%�F�s���0�Z�}�x#���2b�v��5��zo����h�r�U�]XJ�� �}���5cY��B��'�o��˓�h�%c��Q���b>��f��c��Ha��O����G�G�s��?O(�V�+y>�GIo�M�l�:�k����/�_���[�I�M�z��0Щ^"`�d�y^e}�����S��z�eZoF�+rH f�4�x^/��Z�*��gx�W � �ź#}=�wyp�r���k����|�������eo�&�B��R��:�������gV���+��;��������Ұ��W��~qY/�N@�9(�5��I�,H.:��P#�J��@�6�����-/�#U�`c��4 �I-U2���g�T�R��v����L���}�6)�Et��� ݪO|73��#ɣ������,�U�2b�@x��Wt	�rE�;q����3�b�z�9�>�`O��$��xvd\g���C�<��s�e(�<��y��q��CU�:��&�k�s���t䒄+�;� ����HI`O��`�E�cmK��8ɢ��ђ�O��F))O� u�a#{�{y�/\bi%?u��|N{�S�F_�	X�����OLu�q$ڹ[�1i�q�.��3%]x@I�x�M� ���3뜥
���U����zz�!Ď�h�}��	����N9��ew�ԫ�>��C�	N��N�/M��Xi?j�Rڤթ�G�Oų"1=�g&pv�}:In�<-�䳚���9��p!s�I��<2��Ar5XXU�0�^�`	=}��]:�V{�T�]*�od���Љb�g뢫�%S�@W�	�d�(�����L�m��İ��tE�b ɂ!$yQ�������EB�`[�sU��]�9���q�(��bnet�Ѫ�����<AS���v���y6�����l/L�)A�rJ���
�$��ό�šFM�B�m�>��n�����>��$I�ϕ�����9u{��`��?��]��hE
����\%���n�ޫ�H�)���ꣁ��xN�T/�9B���	ac3V�}Z>���8��>�~]���OZ-���e�*ߑ��M�-���a�NfE4�K�&�\�gq�����Q5b�-e[���?gE �I��/��J?�,0�⪼O�=��''z�8N3ӂI���o"�R�n�t��\�k�e��)�E���Ec�˪��l������y�v�L�ܑ�[b{��?Z��-Ҕ0���[gh�Z���,��8��P^��3$h ������s�s+�}���۞�$2�|t%���_2����n���U�/h��I��w�O;���"H���%�ّ�/�+YE����Ҹ��R� ����5Z�G�y�ռ)t �4:�%��(���M4��Mh6}�{�|5��	d_$��a�GDH �s�8���T���Jh���%r+~�>�Z�bL��m�nU��V�#QŬDP�]�D���ʨs��OҔI��)�U�;ul��W�Y�`��۳!����UOi� ]�,�;M��PLʣ)��G)�$87��?�J*<�� �77r(W;iR�r��7uk�(�x~�Uuf��D�cK�@b��n��'�E�7?-�d�g�h�kEt)A,ll=u��D����꣰���֗~�2�(4�H*δ՞n�������-�
3P�3!���?�'7���%!�pU>� ��˻��aw��XW�[`w]B�P��r���IkFF��{ݤ���4dL�o�y���8Ǘ��_�	���g���E�	��ӳ�4���m�=�V��#f�����,p��1�\��ʂ�ne�[Y�+]�p�5i����0�^��z����_}P���mI e���������YH��DQ,�8
##�^F=MW���^`H�/�$ b}�����?���7><��H� �J3h|t��՛:9�8��[����T�qk��0�G�~sd��	��.�����?�Ǐ�I���,�M��^YPnqѮ(��&g3��?[�sT�~�A (�^VKb�s��x�(���"����:���h5����x%�Tڃ��75J���㧊|�	��S���s��bg��vY^�0�߭���a&y�j�X
3ٝ����:<S�^����$�B�\�mހ���j�o�CP��:��(o}D5Li���M��+[���B��JN �I����[c���i(��;4!�笫�0�����3��q⨙�q��4�7z�e�]�� �K.d��G4s�5<�-���Et�j�u�Är���0��ι1��l�g=b9��w��a�7G)�}�o�t^��[zt��B��1�5��2��0��f5?A^��{���:A����NOo���&^W(aA��=���8o��e���:�y3��<1��돲.ӖŌ�b��	3RcL�`�Z�ѯ���A�T[��*�MI��ă/����K��&1��Waj�?e��6���qY߂�hK���_e0�vN�O��;x?'N�.*b:���7|�y�o������De�O�<0��(��1�LmX>�"�@V��Jb,H!c"�c2$�6�[�Aq^.�|�7>U´��֘���ƃDN�rtw\K��SU��U# }�� y�\	zcIU�d��LbMH���^#߉:��5��]�0E�D9E����&9��t��:�a�$P��<a�=��~�7��o̸xS;g+���p��5]�t/.$;��.%<9O����^�,�`��2k�¤ E��S<=p0c�˵�<p:ȉ�p��y����g�]�9��F��ǩzߋV��6���vh	�vq��_��ÁZ[�����T+�k�,�Y~ġ�_�G�]�t	$�n����d-��PW�u�^X[^ﴈM��YAQ��
4YY �w��(���������N���oi�xm��ag5�d�ʱJ��4%���
�,e��S� |2��	�����L�5�������p.㨓溤��<�H�0˃�p��],ۂx^*Mn'b������=��UޝRt��̃��/��@ϕs�g���9,���&�x�.�T�z\�U@��	J'�	!%��Χ.*�4K���Ƙ�[�-1�h�l�P+��NT(��`,ZԜf�n��������a�?Ħ-j��&��A��Yta�&).���ev�oTԣ���ҫ�ja�����a���|�:���'k�X�]vJr)%-�|?^)L���E��PŶ8{:���7J�Z��R�q`/��AABI:�2o#����[�"�P�ӊ�gI��e��w�Ġ����� �4ϳ�7��?l�r�n)�	��k���C�����.W&Kp�̒��a�J"��l�+
��(Q6�B�%���9|C`b:L�c��P�#M�{���TI��x�w�f.�&5
A��Ts�VH�w��B�"��w��Mm͑3�u)-���������O�����۪� �"�ۄ*p؉\��#vI6#X#d�$g�����p��`�){�E�!��K
>�͂�	2��I�]I�
��q���!� ���i�hkP�gen ŏ�d�Z��{'��G�VP�����tB${�Pp������賡L�5`�/h��3���Ը	�7a�`�	�M�0�}��ƚ�@Hq�R���crrIY��l�B	��D7�|-��0���Vs�� n�|�G 5d�g�N���G����M���M p{�r�� ����9���"�v�����6��(Q��ҿiĚ�����ٚ���w���Y"��!T4��ڵ�5�G�b�rWjG`�| b��TZn�fgyܖ���W��и���z���<,���ڽ�4B
��ggԷh� z���󽒘۹�Ǉ"�ys}4����n7�:D'�&�r�JY�ͅڽ	Y�:�҃��Y��u�)�s��^�ט5��P.mm�}Q�Em�|�[���f������^W<�q���4�[}g�1V�s#ᢹ��aA�qeh��P�B�tQ�2���׿Ih�ǅ1����6���.�rC����+����)�QI�>o����)D/��T��<R���0�I�MӎHS��L0��r7P;���^�~��h@�"�	��(��~30���&�-���F$��}�#0��O �Nv�~�&(�'�F��_=Ϣ��{�[&�}���v����g$v�-g5�Oy��/�}�|�� G��y�?~����GX.^����&�y�1N�\�}���vI�s&�.i��e���pq�ᦍ��%t/Y������B_D{��1��	!��P�E�(�%Y�W�}��+hDQoN�w[�;�#�tM�s���B��ԍ��i�=�'��T$��˰�ݎ�(N5`?���>��"=��܂���l*������;�o��o|i����輩�^*) ���:�T��k�X��#���5JCP5��P HG��R�������lR��4�����u�9�Y�-�(f5����7Ё �� � a�AW�M6�dn#2�Xnڽ��D��-�PL4���bG��.�K�x\��+���\Q#�@I�"U�޺Ω�b�'�z�cP-�'�tן��w4LQ�#2�xj!ǽ5���W(~���e��L卹�����o*\F(��$G�^m��K�`;,Vl��f�H�W���DTM�Wp͈ȟ�ê�^Z�[����5F�:��eM~�u�e*8 �nW���L���_Ӝx1�96�U����Юt��V�T�$����`����*G���H��Ǣ0��o#2�-���9���0 q�j���QGCf/6���<3	\�˱��y��$�g��H.>���M��)X�
��u�T���"Pq81G�Ҡ~B{x�.�)���2�}��<C�&���&�"��ݚ���[ E���n��+*���'I���s��P���/�9����k*a
��՘[-7��~6�Pv]��I~/�у�����:��b��k�|��,�p�c���x��S�r�tV���
�� �˵��u6<B�?D���]$C���A��Ę�3ǖ��7JÓ�����':�2ɬ�>�vO��&^S�D{�����O\�Z�|]]gS��X/ou�X�A��f`L�`����{�G�I���7nu�A�+�zH�s_*P�"?�^�呴�F%#C�c:Ź�t(�E���zR���S91��{m��N��8F?/s�0Ծ%Yt%�Q ����+_���f'H����9K@y�g	UUU�n��F�m���������A���WB8��⮲���K*:<h�P��b��ov��O�0PgW�G����w����� ޷�.@[@��u$����ЪHl�"�&Fb������K�Iؗ�9�" u6ג��s#�#P��Д$�bۮ`���k�bwa$z !�X`�Ufd`�H|#֝O�5��[k3����
b���)P���s��'�QJ��a�ˉV��Rr�rp�	R5D�g+٘�űˍG
YܪiH?���@ F����j�*��c�$�hHmQ��s�NB��e>}��!�}�(������"�s=�5g<��W�h�d�O,#Й����?��m���ӆ&B�$�]�8F�Y�.9\�"Ol�g��9o��;�RJo�"j�K�,�U�� 6�R�#�kN���NA%�^���0�aLL_�D��qX��7A'S�2�Ea�]�.��[�wy<�%vo
g�����&�htT�Ƒֵ��>�ڙ���c���0��Jl��M���k����5nW��Ǌ��eʭeL�N-gL��>�0����O�>�������.e��z��(�J���n���:Z=�gV�����Q�ʎ?�?�~���A��|r<�n˜W�6�����)��i���އ�i]�io��a���[�Lu�J'^���R��"�&	�g��Oޯ̹L�U�L徣��w��K=i�4K=N�a����w��ub��D?�86U�y����/��[|LG��Ӌ��Ը��e+��')���K���h�xG;�'�\��EC�"`Q@��L��BBAF,�8q��W�S�l�\t�'K��G7���J��PZ��[�v�hW�?I��)��P��Z%�a�"	gC�� �f}��?#'� Ç kH~I� �G��KTl8z�@�l��I��Q�[�9!r4Q�V7����k	���&�V�;�P�	(/q
W�ߩ �n��߽�'ֹTL2�<H�^����ř,��Zǎ#?m�S|�t�%�|���=���@�IP��7�8ILg8�TQ+Q
�ލ�N��1�8�r�v]��e�+Q��v���.���6�<����ы��HY��;d����)���W��?��	�ʻ����ǐ��/����]���x�]$��è�*Èo�v�~_C���ms�&��)_�H�?��	�L���G�
�ܷ]5D��]\}���fp�KG���W�:a�W���
;@����^� t�YtFX�����E�.ߴu5���j��mx����Z���P �^�
��mx�q@��,�Hf��-�����ɳ�Y�lO�@KB�g���;��9����H�Ş6�	�6N���a/\x|�>��sQ۬F;� U��$�~�<�!��P���I����"�(��+|��x�8L!˺'���Fj�Tn��|����eH�|V8Q��ށ㼛U��\'ơ�5��Z�/|X�}�����e���>7�@�(uG���O���~>���Ӓ"���(�I�d�ó^�F�.GW��X.�J�9��<�����vd��Y�"��Q]J�&�����a�g|�ң���7�{.�E�e]j�	5�#א��l�A�2rX������h�H>w	/Ad!Ձ��u��^$kY⃖f�Y+�l��>�%��%��4C�X9a:���
7VąUe��b�3D�(Ч�"����y�}�F�<gۋ�@�+�;��j�,�	�!|ۚX��N�OӞ���U��L1���x �����:�����0���m'<�S;�o���_RmF�����́�9��Y�ʌv3���������+�Nņ:i��9f�z%��'�ʩ���x�ġ�zas���H���V�}y	0ßN�!��Z�t����v�fOg,^xm��z���2�abk�f�)�[����;�ĭ+�޳&�#�������Q�S��s���|�n��髻�8�y	QЋɨV�f}|�mZY6��(���m�m:����2@���t{E���=}�������%~z{�SR�
���߭Xy���4� �[�?p��Q'"��?	Ph�]��>O��Uo_� ����]�j!W�07�$�e*����� ��)���>E�,|g
`<�ۏBY;���89T.�����V�C��Kt�"m/
�P�:�X6��L�}#eÐHW1�e�"�;N�8}��\�R(f��󓫱tR�y2�Kݫp�+7��
��u�����s�;�a\H��q� ��x�O`���fkq⿬T��,D���KE
yW1�U����g=`��5h�l�g�i�O�k���[�tA���z$�x��%#��~��Mx�S聤3���Դ/���'��9������bRc�|�0A���r}H��R�O�u�����x|��)� t'cK>�@�5��J�>�Sio	_��~�i`��T�z��a�3$�3Ob��8x��6�kI~�|	�q�7֩�A�g[��T�Ӏ��AgXa�٥����Q��eo�<���n������Q})٬��r�@��V�����O�أ$�m��7���rJ;羏������ܗ��?==��_M�.R�eEh�Q'u����Ɨ��� ��~����I>�֛�V`p]��Z�o��Ǹ��r��һ�#_Ȓl{�]'D��Kͅs�0C�!i��<<{	;��w�M
f��%9�/
$͠�U0��Sk��Ƌ���� ��������m�N��{�*f6[�t�-�ϯ[!�k9S����j������~A��U	���Չkٰ�2>#--:^M®E<�֞Q�����R�b՗�\�����m�bgtր#筌�m*G�`�>�ٛUv��4�<5LiB�|F;���V����m]�Ɏt�O��O!,Ř"�کW�2o�e3��zu����6��=Lo4w:� %��	�]-�͎OȨ׷�����^��ɓ����tk``$���PB��b��+��T����OG�`3d��`Px����y$����B`;��k���T�Đa����r�򘚁�?&kF=���bo\$n�)�7	g������7�Te��H�O���P݁������L��ӑ�Y1MPjj�z>���V��e�.�-Zʽ
%��吪ʝ��|8Yיl �u�GPu�����=Ak��e�/�#�x*�Vʆ!B÷�3MK�իw��h(]� �K,�tk��!f2��k:́y:��2��a
̋���D�f;�U#{psDu/g����q	�����Q��"���A�
�.�>�x(�����������;cYm@��&����Z�P�b���o.7(��S ԕ2����o�C#y¸cKCcRZ�3���2Gr�B#�� ��#�*^�õ8�{D�AͰ�+	�W�`�#@��~�Nz�Z�P\2{8	�h~��D�[�BNV�)g����Ϥ��w�x��Cϙ������K�r��It��1T����1���H ���S���]p����.�	@�75y���Urޒ��'6G��}��l���g�ϒZB��q��$�e���{|?z�@"�z.�G��r9���~�2i��8����{��'e�������?Q_v?��K�MXvʡ[7zԲ��PZY=�=�A�A?�K�!�q�9}Ɗ%N?�z(��Mр.9
r |����T�t^U�f��މdݒ����{�=}�fBF�y�\� ��7D�7���5�-�@~_�_�\�c��V�J��9�{�US��|�(R�6"J�&�ŵM5r�*���DW�Z �$f��i�E�5�D�o���sM㕮�u+rK8S�'3��g��θ�/�E�1Xp����
�>f!�$˗G:�|��{�*���e�����i�ܺ�G榨�z���ژ��=�#4Ϳ=�q�~ݕ����b��NC���-�$CȾyo��J��/wh�I�y����M�푰V0b)G0��?�$~E �B�{�@i���m'H�0����G�@*�Q+�q�*��q�x�Ck�K�[ARZ1�4a>+���Ⱥ�� �����|'�{�'�ms��i��瘥c@�a�"r���R�y�r��
%��LǭB�y��Gfj��2�S��d �Z�ް!���
��7a��E�.J���g�ZD�<���^�Q�.w��ZS�#��bF��I�5��~��
|ՃQ��l�s���v�g4d���dT`�3�t�g�ߍo��)#~Q�ܮ��hw73�e+�..��g���b�+Q)��:o�����:u�I/B�H�cx1t���5F����]0#�����7�k�}�������e����ѐ����[�Um�T��/$ᾗ�a��7�f1#<��.ؒq͎�	�B���s�/W�Wn���T�Ug��}�v�HDHT�%�c0�� Uv?��.z2��ָ�4Pu�d��5�L�}sh�����q��臓�o���`[�;��=_|f^�]��mӅg��*�κ�pQ��;��n�o�q�e��N�ƀ�}���r|f%���|4�Ֆ�O��z���>U�4J�/��#� �U���)l�M�Q*s"���XFJ��;���pd<f��ރZWYD��]X�'��-��J>%�iE�Y�og)�}��T��f����Y���T-*���K���a�0E�=]�6�#��͏���ﷲ�3�	�Y��~��m�w?9�hok�X��֞i��bk.�.u����Pa�qH��Ǯ��?
�f��6\ʎoD\��s����5����OVX�����weM��ؿ���C/M{���g�4כu�$@��Z���-�E@���3�nŭ2��g剴����'D����g�t�s�z�R���S�~�1��&Ҽ�jp�T�LGc5�<����y�wy��7�_*G�Āl��;��A�*X��$т_��~�PL�eee��=l�mK�]D`�*Z���.Z`Y��SA���ˊ��e��1�c�� ��1��z�H���:�-WS�l
L����N�|��;��|��1��v���%�l�f&��?X�;?b�A�߇�f���M�P���>�@���Y�Mf$C�HX��W|�X��'�Y��z~J��R"C���"�%>���ۜ�1�;��,�e��.)] �|�J�7�۱T�.�=��<j�b�.J�E b��[����������eM��vw�Zu���Pf�R��
�����2�y��]�0��MǬD;�DY����:p�1�4窥&+�$C*r�`����Q��kntzGd���s�h����e(3�Oo-�[?�i}Ҕ�����l�+���
Qe*�|V}�o�i�eNM̼a1������Յ|�S�;�Ed�s�U������&�P�ʹ΀�r���E`"�/�Z\��nLݺ.�|15�c���k?���Ș4�xabn$����8%���n*���:��X���t:@��Sn�����鯃�x���S�/���xU�>G�	4�A]�*�|�6�a ������ش�l���'�`�����#�|ɻ�[�o.��+a�j5�5�`�7.B`�ӂ�Q茩�.}�Q*EǮ�Q�p�J�:��`�Qm��uב+�D��+y��1O�^e�Ђ�5
�����˵��.����+�qXe���9�;m�OK|� 4���w���o�W.>9遤��%v�E�gzBòt���u��l�w��%�@�J�H��I�PO���-7���*�	���0�`&�෾����Y��V4�l����1^C�����-�1A;٬��4
��ż�E�E�(��=�= �{��\�G^3I���*�}X�&��Z`���`�!
�Dr�ѭ��]����)Tiwd۩�%�aԙ�#<�	ȫƮ��xg�\ڞь�S��D,F��6��O��.��<��w[�͔-M������/&� �AP5F&bxnӀ���T<�fEO��5���'Ld.��-��!��P�d+�'f >��X�R�>+�o���fFKN����	Q����](?#r�	�8H�t]gC�R��r���Q��$�0�>[Y��X�eN�0���4�����17Ng|�p5�r��N'N�ѳ {{�큍&l`�)?"�8�;=��lNV��'�$�$*�k��Pr�U�3�?H1��'��ؑ-�I���y�z6ו��I��c�����M�!��2�x��kA�/�2I��S�\<�����8�/�n��_��̅V��M�{�����B`=F�NhagM��n�'O�*m��,;$�u@�)����7XN��lg&�w��X]��7�PF�����B&�PO�g=�F�l�z(Nw�P~c߼��;�j{p,c�B�6ҢlSa���	5iS����#1�#kU�|:#XV��������n�N�@+�����Th�\�e|���H
�P�X?G�Y3JTv}�.\Rs�#R^+�\fԱZ�����%�{�G0{- �P���C���H��u%��E�*��䧡2k�$�5���$�#���~�y�p``����4N���A5W�d�y���K�� d�Ņ��!���G9;�c�1[����?�	�� �*�U\���T�o�#�D��"�2����6:�z{��]xXV7�lu獃5pF����)Z�Ox����Y��_�ư��������E�����q��C��\1\���6��Oa��!N�]�Օ
O�`�R bF�Y����/��v�[�+1�^ݼ�E���h_?X'�
̝��:��ѝ0� U⑷@xwpw�}{ϛ������U�'��`��ӫ�}��)���������ut���!��O5`��)��[�O��Ǖ'�����n��ʪ���?(4�R*�/|��+�N�~qu-�2h�A���=9;:�W:]޲~/��	��#�(|��U9I�~�fw�N,G�������f$�ҩ��t��.ʳ�y*y@J�K��_\~�c'�!8+�}=/�c�k8�9%Z��$M�]�bI��yk1_F�%�� �w����6�r�]��{���7�o��o[O�*/RB��G�C��8�\�v�	�?Q�A�I�K�oƁ~���2��K,�����0ɘ%V�^��]�BNt	p�U��+�z �C����}�e�����t(0�똛�*��3?Vm�b�X@�o�4�5�7ݽŊ��Ot�UA& I+�S�P ��gO6+�Nx�4�w��O��oX��W�sI���x�� F�v}�T�(�`r%5gq�ߐ�3�
#-w
-��	��J.ә���85��}E�꒓c���^�O�]�>t�_�JVj�Ϭ�{��5���3q�|�	x��=��������U�P��
0U�vV��o�h�p�'�M3鸐S�1Uz��7i����"����0]�t�q	K��bZUo&d�S���Dl���ɀsLܵ� e������֨Qz)s�v�ۤ��U��3����R?q^���#�낫)��x
2�r^q�&y��]1xp���p���C�b9�^!�X*ˬ��wC���+�����MR˯�a�����<��*���ս����$��wM���?#[&0�S
��ɳZ׭��u菖�(��0��;�:+�m�|�����(����^����0_������zp�cu�D׬Aw��n����:S`ru�^��5�;�[>C�����
_aBt|Q0��ڠ�3���\㛸���������k��l����([#��g���SK���(p0�x���u��9;-`�=�ϩ!Vc���0�\�e�T�����j��܉ó���A�崺�����H�<9�L嶧�}��FK�7�]+���3� ��Ҕ|ث	����-�p���5��/:]�*�dҏ�q�A�\��}���{�A���_4z+���p�ī��(&��9H�n�y��im+d��ÞJu�'T��9GH+4�9*$7�¶K�����nBh�tJ(��a'�g��3��7����ی��d�+v?�a�����-�ɢ�Fh��4zq�ނ3�j���<$�YE���5_�&ʔ3!Y���b17|U�h��p�V;_&�N$�n&OD�����}�@��a�	,�"��S�NP�pQ��٦�Uvj�X5b�EV�o-�u�e�:"��L�pI4�5����^T�j�l� t��~����EɛԜ�w�y��zv蘇Z����;\���념�
c�_��Tu�P�¢�}.��A��䎤��M!��j��h걵R�?��5}aS��8��<(��[
�g���"N�O���Jz�O� ��k,��zC�裹�Yi���Cm�K�(r�z��\ܺ#u~w�?�$�Qagi��޺"lc�}�|g���.�61,siܭ���ӟ�I���^LYg�������������R�x�	EC��$*�����Kd�ui7䄊l�GMϣ)Cu��d��_�}Hf�f^��4���N�Y�n9�%tZ���t��\�ݕp����;Z�Ӂ��'�a[Z����$���a�_i
?��pm0��?�ο��1a���S��'�\T��O����)�zI���>*��d�C2_2F|4y��R��1��<Փ�����sBF�1���Q���F�vȬ�d�_2_@tV��8�q��<�d޶�4��}/ݳ�ð^�tM/�*;�Ɍ�l���gn���I|��Umk���_��C�r�1'�x�jb�q�K�c��4�Y��܁�n4=�������V��|G� ����Ͽ��Mq�'�)(�դ��d�D�͚}ob[�]L�l��� �8ih���i�L�,J�fH�GW�ܧ�9�r+)��R�?�63)Rґ)�D�x��CnQ�R���N��`e��\1�"�,e;�?{� ����i�j����������9v ��=T��:��c��c�HK%#�S[E��3��=����ys�T�w���gL��#�L5��lF�7���NÚ7&S�Ĭ�F��G�x����Є&�]��H�.�^�iQ��xH�#�$+p��	��k�� ����ܔ�#��1����կ`�]�y�K8��Al�1E6-� �ݢM(¤����!��D�ƘJӗƵ��j�S�FFTpt�7f��5Cdm`G#��&�ͩ�ƃ�W�kJ����k�����̯�,r�X�'"W����zk7���s�o1�Ɗ�@�(�9�-a�����y�e�#RCrdY�
����`��jѺQ]<y��c��|��w�8�DU9l~/iO<.S�)��
���܊���` �F�)Q,�9"�er�9���1�;*7�Z|:+�B����w��,$*����q�M��D&ͱQ"�#��`��r����<9]���}���ak�A'/0�a2�������F|g
$�����*��(���vP�dpH�"�a�UT����If:W�!��v�IT���!��u��v ��L�F��N����}L�n�wӐ�u����٫ta(�+���
�������W
��1G:��4s?_Nǎtf���S=0:���TQ���֮�o�U��X�E��|��w�'�?��
���0/��ŭ�	�oh�����`3b���~�Ѥ?=hL�O�U���n�zY,u�5� ��Ź�SN9m�|H���H�L��|,b��Q��6�G�����]���7Y�`<���$��>�9ag��'<����i�����̭��,AA2>a�<��S�<4��w��ߟ�"��IB<cP��1�'N)}n{��ʧ�� ��W��N�Gو���E�c#d���S
l�Qf�R�z?��(�s�<sM����r��AR���*�㩀ɸH�G�C4�NM�1v88s�����u�O���Q�6An��0�aa�[�ôI��um+Vԫ��n9H�M4��O�}0[����d��FW.7����m�g&�y5��8.<����e�T�8_1Ǆ�{�\,�
�6f@Dw#؞6=㿱�G������(my��Zk���v�|V�S�SމA��s/
��/��N���!���m�WoOz��|<���ѲB�q[BՋr����Es�Q'�)4���h�$w��yv��C
W��yjHEwe�5��"���XT5�W��M�W�m�;�j\�X==��?�?n9n�{��,j����5�./x67K�s�X������W�0`�����L�2'H:�y�.�����UA>��ԟN���{m�S �B-�h��g���5՞������B�24�YDi�zx��6��(py礮�U�IG\��m8P��]H�B������a�Yj�ǔ$D�vR		�'��i�vs,��T�9�z.C$'�ډK��Θ�=��n�}�#�[��d���_}�[/Y���b���ZGs��B�@���(q1K+ �^bjH|���i_k�]53o�e)��Pxv�|��Qa��,��<ZY�3�pS����p�ko5;k�f���ZP?6�ѽfI��g������U*���^�3����<��=p����=�� �]Jl�tE˝���0N��<\��n��j���K�x� xp��(w�Ʒ�������QԐ����ޟ��U����/��f��[rɳ
��:�s��O�U+������g^q�;���p��:ek���ʀX'�"C��z��7h���_�@�'؃�l=�6�w�+D[���LF�"�ҋ��$M�-Qh|���rv=wϒ��A�g̅��Ɇ�>y�b�\7��[}�D�c�`s� xOQ��9��
*���������"�q}ϑ/>�hmg�c�6�)����az;��F񝓂jC�A�M�_Y����Uk�U�|�G�#��	��ӿTN"ܷ2�O���'��
,�7}�, ���Y��{�ZQ���Du-6��(U�5� �T����.i>�`��ߴ �Fc\��v��65��'3���=��:��ߢ�>-+�����H1�3ۧ���2�3ƕDT]b�#@H`�����c'�����>I��l��~���?���<�=�iR0�7�D~*�_R�	���eײ�Ȫ��9�0Kg���4㽴H�<z���/57�V� g�(��_t߃!f@�����uQ"�2>�T���[+�R�{�+ݘ��n�T��b�)��4\g�9�ُ��p�D$��5�w�����ӡ;���U���4�H<�� :dӆVxO�V�kU�P���b��O%ٙ��� ;���\Sz�F^w�ܤ�3�>�4W��O#����:h�<�-�#vר�QF�sr'�y�0���'�P�C%����K���ؒ{�\۶5KSkh�ۉ�;P�Ą����Ԥ�MoTBD�����?��=#p�t^,ZW�9�}rN��q��.����H�ؓZqa��W���^�'s�[±��5[|��sh�bH*E�	Y����ت<I����X-$�z���].�e(vLǪ(& ݪ'��'2��4U2�_�'��d#ғ�ld�Q;&Nu�aHj��x>u�G��-�P�:����f�"���gnf�""�A�ƶ��n���/ӈ�&$��&_R/���f��`�r�����S
����r�\!X��8���T5y�[fT����A�I�:��2�J���$t��J�I���yˆ�D�S��Z������<T
�/Jb(���|���/�����M ����&G��2���qJ���q��5+�$��vUNã$��!�)�N�f}��Y���j������}>,K�
TS	\j2�b'�LO��Inn�"4�����Eu�_��[Ų���`� �@T�ߓHʨlv3�O�=�X7dȊX���n�n��j ����u�z.���w�)�����X�|N.� �湯��`�tl�g�!�6�ƻR�,����fP"��m)b�w���h��c�?�'<O��@Qo�\���r*W:P�^Kȫ s���2D�qzĝV�܆���k��d�q��|�������Q�+-�3�f�	MA���=O�	�4�c�&8�h�oA*��Ȝ0�ٟ$�iF����)A�t���J3v���<�ɬ���K�5`z�	.�����c��3f��±�	�+`����amN���Y�-���9߂�(!�&��5�����眄�������>�	r��	���}qͩغ_�.|Ю�Q�~=R�褸}���Bi�(|M�Ct�$�o��4��V�;i���	�Θb$:P�pGӫI\d�'
�N��To��6z%��o���1�5�6�E��� ��Ү��]3B�N/|R_��A�8e��(c-�
�u��&���"�H�L8�^�N:�Xʪ!�j�r��a -����q��<�\�eU��7y�5�|��M��(�r?��d����u9�l�_���ЃVX����$��%��)�}�8�vB�d	.^ؓlX�x�ֆ?��M��0�W�l��� ��8k���R���j��	���7�%��%۴�å�F�+7E�5Xo4�ڻH�0���o�ޤ5d(�΂*���_�@N
R_�yU��t�֒�9W��sB��`d�`o[��Tx�^��Ch���[��1�k�n�|.(�8��H.T �I����:�#b�e@������a瘀�*�G��V VF�NE���-rbS��A�O5{��8	��2�Ÿ&B@ ��-��W&)�uE�j۔2��CV���ɗ/����r�,{�H�1տ�`��bw�Odr�4�q�*���}������f�ΰ���W$ufr��'�;��d������������0W �L� mB�CG
 �ٺ���bI��[�A�L�R��[3�3AO��b9�V3���zA��ׁ3���݃��a	���P,tS����.���+���O'�^N)"؜�h���g;��Ffߝa��a�!]dM����ƈJ��n{��oxM��H�?1��2�I�{6iXC�-=3�[")��QY�J{س`����pa�"6�PphӁ@�~��Ѐ�I͠v"�G��S���������tl��Σ[�G:);*3���1h�ە�T��pʬ� ��ڄjV F�~U�����T�
ToB\��j�*ѷ[�2�,u�)~Y�:)��Ja�@Z��P�A��j�把�x������{��1m���j�fY$��W��k�譕����y���S����Ј��[�n�Mm��>Dԕ�<��ՂyWzO�ֱ���[�k��1_�ƙX����L��å��v5�[�;�}f� ���/w��N�8q����h�+����d+��~�Z�������?��>���aO&��g��vh��V��G��w������YiI��@ ��8�xyt��g�T&P��P���ҁ^�C�*�1@YB�V����r�j�+6Sސ�I���];�(NT�ץL{|y��'LB��5}��"76�E���3��|�!p���jI>o�Ȟ����ש�I,?e�P[ k}�S��M�PA��2%��?��j|�Ƈ�� F�:�34+��
د$+ZL5C�M���,���e��oA�]^#;����~�)
��h��ކ�=.g��)���|�:Z��B��:#&����3J�-ُ�zWV��>vҎ�	��j��!��ԬqTI���fu\JS/��n�6���R��3H��`���+��T8e��7�e�&�hs�y<L.��=�a�k��b��a�����d�`������h�V�s��N3T �d!@h�G�HhJA�X�����I������.9#�ѕOl��"�Ok�A���^I�LLvc�Uo�cWIXbQ� ^VȉL/����5����Y�D����t��'c�=�#X=�z�ׅW����<F��D�/D����G*l�U^����<��X~n{��+���Kҧ���\O1���"����q�k���tی�_\�]��xV�Qm�E�/Z:�>`�Sow���H�n����!�ԙ��?OԷ���ķ�ں�g���ȍ���q��1���P�@�̇�irbMH(��~Y����A����m9�;��,P��B��e���2��+�!)�� �u��q�
���`���q�v���}��g��m֕��y6BT��X�Pfɞ�n�/�ߑ�L��D4�p��#%�1Uh�<�I��6���V�do�gxMfӾ�]{-����¢s�ܖ.o���4^��md���P\������@�D�0V%��P�ήy��7!+�񂳢�5A�B5�����P�ЉPb7��I��Uv���Ӈ��Տ1׎����֍k�G��lM�JY���m�����[�t^pwl]A]y��7㈷�W��FPSP6��t��x��q]0�~�"�h�0J�����UIW`ҡ�W�b`N?�p��\�I3[���j@e��!��I�=���X�&Z,��/m�Y��&+���F l�m+i�&ޟ ؀i���NWZo{$Dui1fe6���ӷ�{������w�����%�аP�ti9r����X3��R������t��O
��T$���?���/X�ZRZ#4P�q��"ol�c@ʣBkIv?�^�]�y�b�5e��w��<����lF��{V��N�r�N���kucZyԮ�[
��9y�Eq�RM�h[[��y!Ϥ/�'X��TJhI�v%�s'�@i��pg����X���?���p(�����i0�{�Z�A�C���ؠ\!��n�v`ʁ������ι-sƪ�^���,���u3G$Y��y�p��4�7���!�Q�M�KǇ����B����gF��ֻb2�R���6=��� �Ԗ^���_�L��O��z1��"l ��7� �*ʷdJ���G�65�J�#G��^v�:h�s�ǖ�oY�"��M���*�kW����bٜ:����>޻cB�Cd素j�����l�E�G�Ape
�M�3��?���{Bh�<�v�'����E�=�aFS��ߘX�����j �XY�pl3�^��9X��������w#����nH�7���p�2S��#+x���܂�����ᖵς�=ØFd.�:�q/E��8�9�d�z�:�+��Ϙ}�1��I�Y��v�q�ϰb���>�4��2���>.�h��܇�쁅nz����Xh޽�LlPv���Mb3ֺ	/H�΄��̤��nԨx��;>�}��:����!x�$�
J�����5P�g2�K�6�����v ���֥��~�Մ�t��yV��q^���e���.��/�ms��&Z�)V��̂JKA1C�!H�fte�ٖ�j����ԇ��B��7t�73񩫣R�T-�Q����V��=��pP��J��F���7�D�X�4�����2���2�lx3Ě�eD����w�P��}PG2bi2˅4��W~W�k��^��]eٜ�,��}��֝�QjdL[sC��R����	DU����K���]w��4��Vg͐��㘶*�T@�6��Cd��f}����Xi"Oݰ��Vݍ�ʦ 2����k���/gd,��X�<}�"�Q�9�̘
Š�����K1k�=��H�]�Vc��h���X	s���qVqL~T�|qm���qD[�Q)4���HQ���(�ҵR���n����~ΰ}f�����QD!�:��7�߀����}�_���^t�f���T��oX�{��J���#�uس���� e�e0�L��lY
�~�Q'���w�y��J�.����g�r�h@�|swI%������n�n���p�߸�@�� ��w������~��&T��Q������Q�J���8:/����z�i��h�%��mZ:O\���Y6�|�X�W ;I�-{��>�I�z$�R�*SK�{ßrY�pl���&����֝Z-d{t"�SZ"�-��3
z&�JziK��[9W珆�'(�q��OU��ɓt��RY����p�q2�!I�Y��u�F�����ڪs>ĥ�t��V�ܺ�טُ���N����	�Am\��2u�	#��3g���	�we��F;�����UAG3���`0|y�G:�޵n�H�M���GG��B�=�pm(�A�:C��·=�m>��6~?�q���h��ф'��I�[�M��e r� �(t0g��o��<��od��[CcSM�|�O�=���jǌ-��k3N���SZ��Z@MJ����1e���n�o#�|	����5� ���H�o�J�+�kԻ[G
TN�B3����W��T���Yrg�մ�f�Ob�=����r�}e�}��'Q�"����^{UN?-�tB����+������w�("�_���E�_� %dL��p�cέ�hϒزh��ﺱ�'y}Vh�	�PS�i.��=�dI�1!�ȅ�_<���̕�O���^��Zc��Ff@��%|!I���qO��r0<����h|_е���+���<P��]���X�<�UU�@����V�N�� �MBx�0�q"�6v����.�lDr<;:~���6y�ݝ�I����`{���A���O�R����`�v�d������<�h.��y���໼)G�Ssv�կ�4�q&�X�ڼB6�jT~��?X&�2ƿG�^,h���jp:}�\L�ɒhL�Š0ǲ�%7A @=C͛�iU)�zu8�
����(b$��w׷�� �����'�-�M����ң�Hj�Clu��&�f`��_TFJ��@�� ���BE%�ΒFƀ��n�7�Fv�\��l�Gs1�A°�8��<s�V~u8TR{?�ٻ���e��Z��l�ͯ��Ӊ,�ܭ,�Dd��+(���f�����F��Y��4f_|\�����`����� '���Vш�T��9Th��%�Nt�Y��(� �+��:Z뢼���ϢW�~�?#���ޥr-����JrM`���*ox��Z�c+����M�����כ�������o-�e˛0���7P@�WX�=�@�i(Y;�=;`���g8��1��S�{���;֚�F�h��1���Ƕ�����g&~&I�/Vk�&�����j��1�B�ƱW�3B ��	^h��j��q@�P��Y*	��)�y������ݠ[w�����G�~p�������؎�����,P� c�[�n�36��%�>�����!�BhԠR&׃j&�?Voި�_s��v� >D� �Zuy�@�6EĈ��X�h��xV�O��ri��։��T0�-�����~����b�m+(ò�m�Hs{�q�4�g��M ���ٱޝ
�nA�RI��J�ĈT�qO�4�^}`RC��sЗ��؞;�'�`���q�q�7�Xw�Yࠟf^�I�'�I:�e)�e'���0���*���hӐ	�i�)f*ķ.�t'����n�d���#�D��Z�ձ#3��jKޅ?�����h8�{�D��X@���ga9zs��9�Gp(��?W=��>��l�1g�CNUl��y�!�L�Z劕�u� S?����eA�pQ�P��$Z�:�/�4B����������+X�G<���[�~6qm�Ce�𿀴�x���6�P$΂�=˘�6�H��Z~'��K�W@��YX�	���8(G�ꆔ��}� �D��"��A(h>Ҳ7�<Ώt�]��Z�ګ�Dm�fO�a�:;37�
_}� c�Y-a���#����w����������U��\��N
���ƍ[�#�c/$0�E�4$0���w(�pnl���Na:��"�������eX��(�2�bC��~�x�К�����E�Za]�/ȍ%�kđj��bb	�T�q�w.�R�蠧̸���x�9�ܣ�sf~!T��.����Ｃ���]�R����WH��AQ��l����^��h������L�KY2�>A��l+��Z��]�N-�"_ d��*����!��`�2�iR!�1 ��֛-hC1R�$�ڽf`�tI5��VU^=���
��F��_��}C�$[䳫k�}v�zSehThcG&�ȃ�d������^l�J��ժY�+Bp���|�J
���#6���c�,�����L�ȟ���KJ�C�-�a,�"@1Q�M���st�L/
�:Xޫ�0�L�|���@��
wQ�=zh����&��zc���S<�܁k��4���L���["x�bs�g=�k��](�鍕%i	P�� s�!�jp�F��������:�%g<�!�N�q���wV���}�ާY2f�<U<��,��8�C`��x��<y9��ԬެL����2E �^��_��R�b��Į"%q��4ԙ�sF�����?Q]o<	��:8ᘰMo.��g�i�eq��ԹZ�3/ ����+D,/Ek�R@4>i<��8�[�҇��@̻�4)o?�)�o
ڦ��[���X��֒_n�oY��b�dB�&غ]��?�/��Shۜ�1��Wl}��b��q�-;��&TLn�&���P�[A�@���� o��I��Q(�M��������#kL�`�"+ ���v۷���-\��~6�a:����Xl�������eh�_�e���	�7s����I����-��M�2>�x��'<�+C�?2���W	�gC9��z��eCS�34o�no��L|��v��đ���V���N#Xf�m�ڶ��E�a�Ww������RQq�LoB�,�����b(sC�
�f�s�h|<�����C	[�;#��Q��Q�fg�֨Z����K^��&���vi�ro�y�gK�ς�[�L�u3
&9�QϤ��QEK��{su�3I�J�e��Q�4(e(3���4�2Ԃ�H�/�1�� ���T�ƵZM�I+-�^��& ��,�h���32fɄ�ؙ��#�I�0�2$�=�}��wKF������0���HnA6o�<})��a�D�཭ +���B8q�hFb5s ��8U�Z)ů���yۓ�/D�R�~�GX���^km����;�+�� Ž������kC�4��Z�T�~V⽞nD��=��Cx����	�@���˛Ͱ���7�-�8i�0����rX�!:n�X��Pi�=b�ڗ�Ut���@�LVIX$�2S����k���}�dJ�xE�����i��tb�|��o�@�UDbV��Ǘ�Y�}l���t�1�6n�����k?�*�T�?O���_�W-��3X�Aߕ�O:_5�	9���t[�y̑)��K���b���=����C5ɭ1 �q ��k[[9cVWt&�i>�KE!�SO|W6{�fb~)�w<	k"�.�5Gv�j�^*��X#�6DYu+]a��bJZ�/h��� ��"� ���x�m�W9��P�W��>�󽻿č�����j�T�_�6;6�������0o>3��� �_�ZG�έ0�m���%�@E�R�#2�2�Ҕ�b,݊�!噜�[Eb�x��}K<�<3�PZO�y����vn=w��&�,���D�[�wF�rC祿$H����B��z��kz1+j����H)�t�4Ό�|�!��"*���j'�eN�(�g�����g��.�gˆ��;[�i��^�!�k�Y�y����U��g�'Z}"�$�4!TQU��A���'��FJ�l�7��9HE��OLm��M���Uӫ��&��֘��^H��%�J�:m`1L� |�N��FJk0_Me�&����_�.sy�-�JR�gZ$�"�Ol��^�SG&�\���d�SX����������sr��G�T&rҹ{M�dj ��z������1A@��篘 ���xQ�i@ڪ��g�0��]Q��-�Qi�DCj�D�z���V����GA�.rft�Q���7Ǖ�a�,�~��=�����SWϝ���e�
 y��ʰ�v�4�z����uˎ���͢��u/���G�l!/��@A�/�,�_�������v�ڹG�VR,!\`��E�ߜ$�b͕I;,��'��2�d{J�0Jޛ��Cx}�-%�t�7��s�e��.�Y���"��J�.Z����U?�)N�-�9�"V�^2�9P�~J1���V�몪�\���9+�CgC����.2۟�����U��Y/R]�=��HB��}�bhr��c�^�A�3���]�l�C��"ì��5�����*2m:�:(N�%-���Gv�5���0<��!*>������?
H��߸�	q����e�Ay�'1 ���ӷ����*j��B|t�_�J�^,X��cn�)�?����@����i�;aL�#v��߀Ʈp�0s��K�A����Ƀ��sʃ���&�U~h�H�#�.�~�a�P����������j.��e�	��2\�r%FTQNH���_���������}�4��p#ޞ������E��2`ki�<��h+/8B����V`H׼�ۇ�;'�-UY�р�`�B��m��RΪ{Za�l�{��?��[)�d=�7I�6	)H�\��7XU���������\����á]g��Ō:�MLi8��L(JPU��SXSN�(���Bԑ�ڢ\��Y0-kx�3�+R���競K�%!�V�c>$�f}�_]��*�
�\d���^��wē,�wh5��,3Ηa��J���\��Et4��)3AI#�fA(��q[駃ԅ�_e��e�H@2����I]"��?�\���,��'���u�B�����*!�jt�ۨ*�z�cJ㧡3���d¼X�ʘ`��l��i@Y��gZM�3��<H9�WZ�Y:nn��a��5��A��M5ײ��[Ou����vΰ) ���M4Ӱ�
̄�!n���]	��d�'��Ӏ[���-!3m�z�|"����	CO6�+Pe�����b��Y_��ʮBE��4H���.З�Y�A��kv�RK���V�����ӵ��r� ���B�E�Ph�x��>���d��ޖG��tJOU�N�.����Ŵ���-����`�8�	/�Mks��0��D�2���O)��U�j5�ϑ>�=��X�9Eoc��k:�|�A�:u��H�2�׻xB�B�@�4�
����i�Ф`~�9¢=�r~O�9h���/U�|�كW�U��^�[��?��g�k��4z�]��������~��OQ!�ua�R�9N*�yB0��^F���eS>���0�W~�2�x-=�E��$B�%��1��CW�d�m0���ѡRa�+.5�� �}@P11���*M�����e�L�lxk�@
���s�u$M��+�yC;�Z�0�K�%Vv����pu��"i������	q&�N*��|ɔ-�)n�r���F9|`�a5�»~/�(�BG�p^n��<�L���(�Z+�d.��? FBܖ����X���(�Q�.�!�S�v�B�F�r�7�BW͍a�K��h�����"$C��H�I(��#��A��z]U����msH�
��̜��T�X�P(t\�O-���G~."���v��dAb��{Q��^�Y�u��"@�� �Ɂ�<.g
2���$w��,���q,櫠ȏw+"���':{o���R��
�F��i_/!w�o���r�ϛd��ˤ����?-�@�����'�E�@5�R�d��n��=�7�*�+�1���7���^���$���9:�3�؏1*L��uN��2���a��T��N�܏ph�2V�)p�Y�K7�� f�<�s�n�H����.� �A=�MI,��/�����L����c�߅����2B�Q���[�e�.qRK�L>����r���܌�x��Xw��D||vg�0�|�6y�F�ٚ�k;A_�4��]� ��Œk����=�}��M_خ�L�`��t��ݴ��
��N/�&$�7;jI��U��-* !��,Ұ_a�X�(C�I���e�(?�*�Ғ\=�f|s���X�ĀG:|�!��P~)��kX�q�mg֩#Eb�x�TA�1Bh"�Z���]?8��+�OֵQ%A;��Ap�XR�B�k)"k!	l��瑂���e�)����q�}���b�J��(�-���@d��0�K[�����}���9�5uD��'�hݢ���K�;���>$>��.��V���^E�����1�2�m_�O-��Y��}Ԙ�k��,���l=�R����Xx���HsQ�)V��n�<�v�ׄ7~Z���Ʒ�)b�>�uD�<آ��ߤ�H��3�zR�l����P38aE��w�3p\{͐<u3��GFp^������d�������
 0\���G���b��f3�@���:���d0������o���&B��i�����˧=7�:5���P����'��pB�mM���,�r�J+APy��Z�/��JU	B�٪�:��"��&�����������AbJ�D����;s\��prT�sI���׏2������a��U���f��ưG�i����t޿PA��V�+������O��+�>��ٻf�vnb:"�Bp�^�1�A�-�"p2M�n�~lBB/Ů��'Ӓ��o�r�Ȗ z���P�j���#GAi*�FVPM(�&��b�5������Y����������\wa�U�q����������#,�e�}~�܉_)��#b�82é��
����;��6Uh���/�q��뛴�=�hG�]x���W
��rU��;�e�4,zC�eq�\��]�y����U��P�BY�������xC)�yz#nx��K�������mJ3���\��1�[���@�:��l���n�I��ۃ÷���F�ni ٟ�i��7��֋�l�h ��w2���������,�K@���pHhUu�ڃrF:Bn�X	L'\cR��$.�(�z� b�u6s�-�L�ƨ�����jiݎ����7�~sM���������)'���Q)4���v�B%�e��_���'?���VJ~�ܭ�'59?�cK/Ȕՠ��_��a!�����N姊�������^�:���i�؅HS�#��}�3�$}/5�fK���h��N$I��pK���)�칓&����d����x8㣭<�)��㘱tʖa�e��A��F��ԭ�Bi�{'A��&�=�=�'��n�Z�l��� j"oEuR�+�kwo¥Y��*Ұ��|L'����<�����Ҽ.����Mw�V"]�om�3�������X}�r
��g�~105����=��}�*pA2�`��^�}������������.CR0�H�C�M�qL`�,��i�k'K9�^��n����6��5�_-3�2v�W#�[�bB�1u
�����o`�jI �&��1|~Fn�Q����tKU��?&r� ���Bč�X��6�Ar��}Y�&��;���э�^>��i�?���cɥ�y��+ѿ�KQg���Y*��\�7�d`�����F����fS���?��[���9�4���2��4i����-�k��p=E;��p?���4� �2�.���;SE�4�c7A�&&I��2��L�����U9*j���X�1A�{�^Y8������L�-�U�\����� p�B-���X�d�"9vjS�eX�R�l (�!��e����dg��g�j�W�5g]ހl�W|̋�b�����S8:�5����$�s��&�R&L``�-K�t$���TCZ���,�/��-ܶc��X+��_�"꫇�6'��*�������N�����\w�H:e���:�(�P%��z}}�H"�A�Wpz�"1t��[�lV]{�q�J��t��A�m�f�!�f�''M�]��>�L�.�SSd��Yᔊ=��դ�o�z�?�����?��)b�5�KU�d�lS�Wt�|�������}��ϡ�C��u��h@���ήA�	A2Y��U�QG��i�����+�YV��t]Pw7��VftoS�a�1d�.�j��Cß��ܤ�P��,�m���N�w:;V�+�Z��k�͖W�׈��k�\���Z|�8�dV��R�T��ˈ�f='��PA-T�l�9H�D��kH,�x�g������O L��:�.��+j͑����&�jJ�6���J�3��s� ]�aѶ���	B��L��r�1�ܸ�Gf�ju�����/�Q���TE��������$Q�Ҧ��5c҄s��mU��e�.NJ}c�D�~p&���P%7\½ɜ��!/�/��T���T�p)^���F<�ڰ�do��q��Ol6fĸ]�{t�-�E�_����G�t��;I�y���|̉.��06�~U�%��0��)V�6��w�t���������P�pD����{��j�p��TR#,���tou��̛�L}e[�X<�9+�:[<GnC�U��F�J~�ַdC b:ݵ3��4�l��u�{fK�e����wt"���	���^:����T��DFaȼ�=���d�6����J��W�W�/� ���$�½j?�#t�q,��e}=!Au8��i@��ӳ<��Fq�����a5�����!#��-�!^��#�bCt�,^�3�P6N��|:$�<�s���U����pb2a�`:엢��4A<���5���
�&+R&l�n���:��>�� �ը�"��2P`��uj�h:�Y=��P�4�#��s�F��60�.W9��!(Z�חŶy���;�eq)jl?���A 0_F{B
����d�L��������:�wlk*�Jao�����?F� ��IZ������Z����I��f.�
YIe��@K��I�'t�!��9,���S{��[�vQt��t��$�����N�c��Y/���s,�X_�(�d��jq�l�����6b��%cp���P�t3�N�v�5�o�E�T�m�{	pR=�U*�<���f�i*��p�nZ�����X�?ke���UCϊ�JP��>e9�[c�+�mv.j�����pD�<��Q��O�Z�C�z��3�]�9,�e�3�ц{�+�*���w�`~�@tA���_����V!fbY��\��k��(�<�_�ߵ��<��P�(~��e4*M"�k`�x�_��!�@��e���+s��R$1�������M���r/Ie�������W�U{O���꠱^iؤ��%��1|��f4B���Ć.ء��Y���"NE`��Ƅ|XЅjV��P.��b j�^g�� �2�s녮����'t云�9�W���nh��/��cv��_���k	�Y(����:�j��8��l�nH!�O��2*��In���9K�*�	� ���F>dk����2�N^P�,v4���7�GN������
�Z_p@6��>36loy����:��+��kh>J>U���q�U<1<��G��k˨K���:�s'�����9��}�����W�|2]Ψ��m�϶���!����J�^�M��ҹ�/�aZ$D��X��Q~���A��#7�[�)�[v6*
�Ym�� ��D�ԓ(�k��h��mP~��hՓ��ۼ�`�$��]Z��8sz�ByA�ء$l��%�!������}A���7s�o����#�}��Kw��������4��MP먯)-3`/�K��C#l��4 ?�yr�9��x|`F?��"G���$�zZ�ǭ`R#� vz�Y�˨ѷ��(���?��i�o�	�@Z�Wɨ�0\���q���z)g�;�adn�)��族N�y�L��PtpÓ�|�Ȯ��%TJF��|�w��Ox9������E5�r�9z�~N���f9�Ba�~���ң�H�g�e5�8
��y���8�X'�Ə�@E�����B�q8�L�?�MB/��H�9�rg��jl\�w�F9mFx�%��!L�^�2�P�Ѣ�TYV��ZR�^+ɝ�g�N�\�,�UL�"��ӻfi�$T�'m*��>Fe��Y���"����E�k��w�@�C
������=v�s��X���~�I@�V�`��C2o�u�EǇ=u@�Ɍ�y����v�Y��P�S0v�����c���)���/=Y��(��F����Z|��j4!�����ZAIw]"p�+R��Ȩ�:���cP=���Ɍ�!\��L���&t�k�xq1�5�h�������h����T����~�e���:�e�:X2�ƏD��ozI�ז�u��|
��ڌC�Zd��6���-^�3(=�%�
��JSt@O��&�C&%���!8������\�)n)�3�����_�ಾ)ℇ޻����0ֲ�bSP��I�����%fi�bs`��%{�Y�K��]U�M`�4�2�P�p�y�����_��?�[�*u�*�,���3K�߈ڸː�����R?B	� ��&c�\�8��#>���� ,�V�k4Y�^E4D�,�i)�cPq�,dxe�/"�h��6t)�����������%���RjN���a���T�'���,e-ك���<��"��ཇ�K+ 36�Ѯ�.P�t��������	a�q��i�T}{'?�<I�<*Q�O���ފ�&�� �^Y J3���$�u���-`wǥ�S����Z���J����@XI��PF���U�{ոP@��� &��2���P�%I��#29!l��LK�H8��Q:I��/�3b,\�?�^�*>���*{����2t-A��x�d2v���{b��Oޭ߈?�\�]8i�L�:i�ݺP?j���+��7ЯH}�#þ#�,t0�{�@rqU��mƅ����NjJm@�i�M���*F"����g����}`�U���e9�b4�m�*]�ڽ`�f�H���k[X�#�,�QI)��`J�u5���B��p�Ti�XY�s�oW<s�,?�ŌY���*��('�L��4��(X��.�:S#}�p���cCZ����d�D0v���P�f�"$��=مaH�q.�j�;n�����밡A�`�$�@ Q�k��-��0v�N�l��/Iͳ@�&Ƣ�0�͡�.�u��#�M��h�V����x/������8�CZK��GQ��!�Z�q9��ǭ(wD��9�"0�,90�ł�`G�n���*o�����w���/ǿ�6&��}�M�˞�+%H�j �Ýn�W�w27���y(��S봤�w�8��N�?�iKpY�`V�5iz�bAݐ_5�$�^��}����x���xwi�,u��i^��|��\ ��G1A�����(�qt���9�1�溡��h��La���Za<m��PѬP�p����\$�.���#������`1`YGu6�g�t�H�y
�� ���^���&!����%#2�R��=�(b_�M��k�wH7�B�[`� R����Qe��+%y�:�ô�Uc0��}CT�=^51FU�i}�l�\�j�Y����ws׸0`Bf���^�t�_e����H���ճ"�e��J��k��$�?��{w�L�ޟV\�|9l��ћ~N�����{p��"���Ԓ4^� U��݀n�Z2X$V�����q]uvD����N��7��z5]����������	�f�Ab��0��)v�;��t:�+>F�p���	/����b '�xGb����	s꼯|���lЄ��R��G� Fu"l��%{��;�%�F�s��7ج���VE���S�o��І:��B��w�P�O�0}P\��`�c��Ns�g(��?�J+����<���F�0�j�۴MGѮ@_mNGkA-龭OB��B���JR5U�X <�d��4O�<TX���x�fT�:�k�\��g�>�ǒz��jR�,g(*`��˱~Nd�5aEջo-EXȑ��p��,lH����bi����➼2�9��$c��:��5o��`�Hq8�W5H՞�&@h�f��U����P�L���@�"� D���Ie��::��� ���ć�����E���
�t� -���a�H�(my�	�>�!�(�����d���b�ؗ>02'zl�|<�������q�F���]��]��sS��$�+J����Txt�t���w����}�JA�/��e��v�2��$�N鱬i����B�8�16�j�3�
4��Cd���H5_���T�|֍I(��"� �K�N�ԧ�Y=��<y�u�hsг�|`M�B�|�r�c����9w�U"�&!�3����Q22�Aw� �r1��cgBG������P��с�֯�dR0��y�E����Q�(o�䋳��6��n�P��<(씬�D��KE"�qD�����=q��Ҡ�R���A!���n�����D�'����J|�L	 |�~�DƖ�V�N��9S]f?q��Qbo��/_���$�K��z�����o3��	�w�5܇{�g+��Z�_Y9ı�^ٷ|&�Z���`U�)�Q%�Pv	͌b`���F�R��Z�J�@�U�޻u�_�J����������4��
���ϑ�=WHũ>�^b�Y!�����N?X���M�B��-/���>H63y���c{A�q��h�B�#O}�i����ںo&<���[�r%TⲜ�Q��jF�u��.���6^ʪ=˙9��Bl�m�!^Z��tg�B�ݠ�Eb�H4����2!謖em'�SHmV��~O>Ŏ�H��b�2��bl�v�Ec1k��zE�1���Tr�@<�����PPPC�dI%�{NӰU�j,f��T�m�w�۸`���p�L	�e`��rg��=�{��)턏�P�Ғ"���dw���1��qW�9�X�#�����N=��@K�m^On�A�*�fB'}Z���:��l��������Qr�Z���>�R�û�*f�#L߼�7�r?y�VI(�=|U��PJG��qF"��ĵ��P(�$<h	.ŗ����>��i�*׿��������9=�U�8�s�&��,�ZʓRҐ�E�ݚ�r˟� 1+M�灘�P��䤢�F ��p��p�\,d\� }���l�ha�O�E��)O�\����J(sރ�X�|�|��d��.�Ϻ�Ɉ����72����oR����E�d+R���3�/���W/��gb*b�'��l�� ��M�()��K�Z��Z]���|;�T6#)M�l�'(��&B)k�-p��������	�o0ISYÖ�@#����qz'Bk�q�K7T��ނ�*2��>v�%�U0�p8}}�eK��T\C��<��~�` ��E ]܌(�u�?��#����b鑅��:�YN�m�yF�P|])
�"����V������$!��p6�J�5ղ�/*�t��h\�?U3��܎�'���W���T��K�x[�l��R���}��4�n��U4����t����|n���͝:e�e�K�Q�A=ͩ���l�0.�]w��{y�tu^㹐M`��s1lp$2��q��>��#�2/=�ǭ?�����Ʌ��Wj�6/�v1��-`��8�#��a�1�v��݋�
�bg'�q��7�E22S����D�:�e�`JXT�kK��!v��k^��,��	_�@9�9�^>��!��;K��Y~���D/p�a�-\�C<gUɱq5"Ѫ�����f��� �1I0R��6h����]"�z�M�KE�VdM����;k���Τ;F'�<|�G`�Q��y4|nch#y�$��r_m�sд���� �K�=�a(`4�&%�r��a�ӧ�
2Nr�Mo�i�"[3�b�tOQBrsN9n�Hl����28:�9�U`b]6VTE>�Z%�_e�)���P�r����Йt3`����D$Bv�M�F����dG��TO���7j��P��.�l�"��9�;��)�_/�+����,��D�L���GO��?��MO����-]�I�ˣJ�(�:��f�[�k�F>^�r)!�F�b5p��ӏ�C+b��jVaJEr�,:p̶z̡
E76iwq2�\c�����#.C��[��ٮ�����~t�Bp�[��D����"�|\"MP3�k�BȞ���w&u���� �{�
v�c�0�[`s,���|	�&%�as�
z�ȭJR����9ݱ�9��;?���늮�����^����1jHK�Y�Z�l�*s�8��"~,�P����YS]�:
���1�;dx󗨷�|)�� �j�v�.3�c�*��1FqH@���tN0"~uMNEz��M����&�|��W���x�sT�&Z�>zij:�!������ �[;(�m�ѐ��}K��&�	wiU�Q޲��])��9��n�(�gM�F���S`x��,�J������v����-'���4�@���Gnu��k�÷�ۓꄂ&@}��F)@�������!���9�(�B훵����%IT��t��O��C��	dΌ����[���k�W�8�䯭�R�щA��Y����}����,i��J�C"G@�������aت*��x����.���F�6��3lѰv�����>���`C65=�Ywo��̣N�� ��n5g)Y(q}��B���Z���ywf�%���%���,�욙�!G#`�Dp�����@�tNG�M����v̖����Of�7��4	:���.d<��i�U�P��?L��d�0ӟ�y��'!Z�]@�����$+��90`#�E��yӝ/@Qʸ�����*�I;/�E�����]u��=��O׫V�y�F5Dٸ��sV��� ��k�JS6H:�oY�!Jw���A���b�{WY��ѹ�KvL�T2���"��`ӝk|o����>.�?;x�Z�l��#�cf � �޼����b�[zo���AP�$�/��4'�D��p�iڝ���B4o'�j;�A��D�>�]J�'U��/�hQ:�$�W��Y)�����0
EG�>K�WUx���a�NX�P�h-�8�f��v:��[��yy�M�Q=j�=}�\�&o(�4+�%<� ~,�������F��Z��i�T?��M�O��S%	��MzB.?�(�������>�Kdo�ׅ����r��!�e`�?N��aO�_�V�Iys.���D��V	�6��'Ũ�u��nد�#�fFGk����n��
�!	O�y���Cw~ԃ����.B�ϡ9�_~\F��}�]�Ce�i��rYՉ�(Ŗ��`��.!B=���'�'�9K���k��5�ē������$�{�J�мԅ�Ŗ�~2�'�N~�
.�D�SP����w�W��̄��Ҫ�d�Yv.���_��?h&�ҳV����ʀ0�s)8�{�ku��o��e�R+�����7�ּ�
3F[[���s��ɡԋ���{�n{�ڸ�g�?l=�mϡr.������E���o'1��%���0(�qr?�q>Q�WX_SW�&e��kS��y�ɶ��3�U�s띷H���4`{Ӑ������7��w�?�=T�̚P��v�����/�Ȝ�a�*z�s��������E�u%���Y���g驵}J|��B;Ї;u�y��M���_���X��t��P����7 =��+��NX�6�V��ʯbG}�������Ie���XMR�-��eK}GKKl�ں��R:�����hy�I*��&��0��V%�QS�?`�P�Y��f׮O[娎�%v�`6^�]�0PJ�m��3����k��L�͵x�t��4's���������w��֚:�����8,u<*�U�3N?z�؆κ��U�W$3e�T��Ɲ;`e�0�[Ɍ:�z�-��2�Y�|��� +�PI4I�^���������T���P)I�����@���=]i��ۯ�#����D����X4�hu�@zO/x�U++�#(�[�)J"hĠ_Y
Z����g jm$���:�c����l��Fr�(W�ٜc��[�h�"�� w��D�M�g����<pNg��?�X�kw�߇*_���W�qx/����zTeM齬l?�z����D�SV�_�ơU�TM��ˏb"��U7�>|F2r�^�Q(�+ͻ���;�M����HG�K�%F�#���*dۙ5Y�3ˤ�-k��[JC�� �z�ff�/d��D� y4u������k߃�c8hM=�ƕ��]Pm�hu6�68]W�ii�+�
C��t�srw�O�Z<�I#�v�n�'�ZOy��u�z�hB_��������>�L8��)��N���0� >a�Vz����L����kK�!�rٹ��}|rdS ���w&P�w�u4��/3
s�z9��')�`3T���1���(B4�\>��]u5�TV�y�w��cJ![t�i�u��V�e�`j�!+<u�]�|Dk�[88-	�%�``��ͣr�����*jA/��b�@���,$��[h���� �̮6���7ä.}�#���-���3�[�W�H�Ȫs�m&":x�x'y�]H��7���+3CA~�Q:	+�H$5�� dT����l�cL�����%i�*.:�O��	���lQ����!)ت�����t=tڀGl�J[KAC������Ֆ+�Z�V����D��v�~>�`P����-�T��'��8�)�σ9D���3Jd�2#,Fԁ�)��]_#;UBړ��Ao�!S���u��P���<"ӏ.��L�e�:�k�/@*���lo�J��Z&�v(�����5�I-�H�ߔa�.�_��F�Ё6TRx��X�|BǷg��Mp���l�,G�fZQ�䭗|��$�r���!#n��	�rm�I$짲0"Ì�| ��TiZ�Z��Kk�\�&�%C0�S��.��25��?��� L^\�~Z�=$���'�kX���[}�s.3F#�S=
�������D�ĽGi�y�n�N�MC4H���B�����D����D�F��NP����u���n\�"���C,�9P��i+��V�2{���(ƂyߐW�R�Đ���U��]�M��h��k1�JWG!#-�ٰ�P��k�kC�~��q�?�UDښ�XdJ2��	l�f��5��gъ���e�-��S?����K�@��o@�ZH�`�r�':~Z)_4@'̎�E}�foL(9�~��{��f�j:����_�;��� p�����P"�Է3���I��,����ᴁ\��Ap�Q�P&ܤ�������Z��`�tJ'TX�L�}��D �"���
���!xvJ�qX�j�[I�1�R6��O,�Zp�@%.nVE=�S����v �i�
���s�-��
���%��JSo���6�� )	���Lx��>'����.ث/��ŭ)�/q ���e@�/;��f��7�!��}���X(�B}fP�����?4֜＂���@�e����[i���t�%���8�-��!���f�j���]��lo�L��'�Y���%��+�<�0E�t�H��`�nŮ�v����((+�cf	� ILZ�D};=�r�3��f��x�~|�/��|���x�齣	I$RJ=�&��[�lf4��L��-|���q�T���j ��8#�s�EU8����Q�G ���������ߌи����7 ;"�{Ckb�&�啙ZOo��LlX�o�L�r7V#���QߟN����$�?������Ӌ͚o�p��]d��G�D� m�%rF��h�U���lǼ֛,^̬��H���+��A��^ʊ �#x�Xvm����-�iގ�pWl�Q��Cxe��	�?�n^��v �k�b=�c2��M����GJs �9��`NR�N�r
')!`�+˹ �BCu�Lov��K'/��
�C�p�����d��h���e�v��0����m2�70�7���k@����)���n�/�H��2��O�=0��ܭ&u`)��vq�:�aY)�i0;��p��&�z� �]�z""a��/\����} 򠐋��©��b�
�0�'��]�Vmh���_c�As���ZQ� �H��3/n���P6B�ˀ~B�7m؅,`�2P�v��(ZV'�����2%:�l���0N�x�/]��xr���x��g�_�H���Ւ̜I�7�2Ƅ;����I�d�o� C>K�t_%��c���|���Ųs�s=����JA�I�?���h��ٍ��,\���\���ϝ���ܙ�՚��F��"���
o(R��]�'G���6
,�qZL�OSs��G$�l���z��Z5�
��8@��RQ�V�rf
�LH����q�� ����Ju�M����s���z��Y�×��W��]��0�YʘBG�Fp,�HZТ���'����}�d�m[X*�R�ו\��|e>���5��t��d}*��#m)6���@�]�4�d�������=�v�adb���3Q��<^(�2�_O�8����2��Y�>�<��ӚSv�T�b���hcR;o����M�����|���-4�z;&8��;�$�>o|;!A�����@G�����E�f�׺�y�m�s���^6@9�<͓�wE�!k������D�?H~&n`���x���[��y*�@����X�j��^���f$D:d�42`1�"m}�PS�%9@2�v�;Nw��.���:w>�P<�,ۗ]S��=��*^!�^�a'U���%ORD67��%�j��Z�U)M=���B�)g���A�E>�Ә�-��)X�{�x����e�֛��ъV&q�x�g��,�(~�{p�}O��f�{�`���bs�<��#�n^�g�ʽ����Ll��[H~g�g�Y�#րJ��ɐә�ʎ��U�Ϝ។�p4VW����]K.���̘��}: ��|`����Jk�Y6@ Ӆ?|����T>M;�[����Tl�jr���s)1���j��V�B�^{��'*�3���^l5�Y�$z�Eܼ���}���7;�%��p��:s6�.��m�#wِ������T�dr%� ���C�}C��챏������+@���y�Doj��<�v����Z���qZ�*a�+ϟ
�\�<_��ž�
�=cuҪf�	3����P���^���R�����'��s�Uq�T;@���m��K�G�O�N���~��m��Rkx�c�4s��=%����YE���l�L�O��$��#/�*�������:=�5����
�4`�	�N�z,jK	zH	�i��A�L��������#YX��~�����iX&�x��\��bL^y�a�q.��[S���;����bu��,u�#x'�p���`�V�	�{T`�Rp��$BUw���z`�3���+��n�S��p�$�9����U�g�&7\̍�<�j>6�tV��������+�c�	�2��ڪ�2c������nv=N�)�7�	�ɹ)Q	�"��O\�a��M8��K����[W�X5Z/�����R�}���!4���٣n��j��;�h>e$:c<n%GD��y,F>�d�!�#�6a��^���^�c����
	R_/F���G�H���%�,�d�9Gȡ��Ŀ��c���	Tn3Dd�`�A���k�[N�6 N�f��͆�쌈̈́Z?D�����CF�"~�f����˼Ka.�����w(�����CG�S�-zh�s�U��lq
E����o|�L4ā���m�'ڡ��_�����A\i��v�mf�q�|ՠ|�Õ-�A_��������gX4���?G�T}}���Y����;�Y��v�JL�����������!�f�p+��x����VxV�Z�����u��͊B���	��2�v�D5r�4��t����QPdz���t����
r���Ly�J�ʗ%��HLɮ8�9P1�����LLj�������
I,y��R*Y,� �ʡ�3s���b&�����Ih�_��H�=ћA�-����zw/��X,O5�.!V�HNi΁`�m��h��}eH�SCUL���&�**��B���zd���[���Ug(�Nǝ=���ʹ���Ѯ1��g�WF��͹�@/��K���	ӝV^�_��=�뽲S^�Y�?�. �%� �TE[7u�w|
M;N�@u�������/C���� ����]Z�y��`ع�o�Rr�͖���P��D#
j�����O�A��^��<21����g��@���+�p�b�lO�P�(��c�s&s�lh�FZ#�Af�	.�q���z؅�g�[��Ty�b�{�IL̅�$J��3�_��S�O{�drY {35Σ�~Z1�F��z�t2T8���.��  �`~�F���kը"��o7���=����y�{"�5��8���by5�_��~��W�@��1��i�qG�Z�l%�Q�7�H�జ����'XY�S�{�; YkzqH-Q�gߌ����v�酇��,�8����/5p�Y�n�[f��Y���Zd���Bb��Z�����Vq41�>i/@�O��Yz'���>�3~r�H�Ý2��
��yQ�N.W*�G��JP�QR���_o�7Ű�k���Oy;�K� ��b�U�NtQ7Ƙ�o�eD\;i���_�9�'��]�S�7j�(���@�������0_ٟ���1J�foH#(�O���2������d��f��.SdA���v���2t�B^�ZX�t�z�����|�k��A_�D��._4�v5<��x�~�ge�@b9E*O���o��[_��3.
������֡�ب�,Q߸\�JX����훣�͞@w�*���\r�$�ѡo��2}���ş�P݈9���|e$����D��TⰟ�����QW(���̰(�/��іp���@$
��`!���\(�H��͇ ����\���U����������%�sa_h?b�U��[j�+�l���Oٰ�]j�= 촅Iy�l�>ћ��h��[R���GЫ��4�aA�Ƒ[�$&��i�#���ͮ�-s(���O����T��%�g
6	��;f�]�nRcd&6}�\����RT�2����W��vxl�%|?RG�f��^���vQT�-m�n��3h�T�jŷ�<�깸%���.I��Lrx���FqF󋖯n�ԗ/��o�Q�)�N{V7�/ڸv#�Ǿ}�)a���u�`A������.����!J�bD�	�i?ʝ)��1�Ja�qXĖ##/�7�3�+Zqt��_�O� w �{CB����z���m4�~p�?Ú�H�ϫ�wo欇ǯ�:{h谭�>7�g���լ5u"Z^����}�z���D��(��#�c�!����e��~�[�A_�*a�p��<*ɝ�+E�J{�NZH.���P�S�S�t蕼���S���v+�*�td�D��>�/�%Z���<�F��.�"�H��d����([?��Ac=%ntag���{$FL3}��1���,�o�,��y9�73Gp���"�o��?��|N�U:�)�x�([ K1�X�;�(��m�|^e�ul���.�'9�B�̪���w������I�k,ƣ�)���tZ�s"�1�&c�bi�/ �_r�^�����Ҵ������ݻ��>׼`Y9N�f]����a���h�R�m@"�C�.�<#$/�k�En=c-��e��Ζ+�"Az�=��d��"k�>�b?B��6���Ӎ�u��r�u�Cp�ފ�e�ųX��A����b�!:��]�=�=h@G{l#�p��x����6�рFRՀd�lG��tx[ގ�,���T�	pE���8E��48�Km}@DNℰ�S�\J�|�����A�����ޱ>�[u�D�������$��m����ce4��tM�����ѓ�>��Ah}�o|�'�~�|km�\s�t�����C��8uR�b�ՒΪxՅ��M���k��xٍ���~�U� ��$��q`hBY�S��^�]俪��e�6pe�R Y����*2c��g��z$ũ����<V�q�t?Nt��e�N>%�|
�}Z�8�~&��U�Mp�m����ԅAϵȽx���63�1�_�ָ��������!�Y��2��� a ��8
���ۼ섥�ƙ0��fi�p�/d�<QFq����ΐ�^YyIx�P��P���)�/��JH���F҉�+j�F���2���>=Գ��ި����0���vaa���="ε�?[�*�[;�#������Saw��*�ۮ0$�F�v���l*����,U�����8�Y���e]d����`nh�U�l)�h���W�e��3��W�}��@^�aI�}���r�' ��9>vo���2�:j���t�A�"�.��T2F�e���@�Z��C��^���/������f�vP�yi� �@�����w�P��p�H�!�TI�$���jt�"�R	z}u��Z�M�Ԛ�9X�uZ��ɏ��l�KP4B:Z^N�)��;���%� �����uæ���_����PLd
W�w��r�<��n*��ͪ��{�Q�sR9p�#X�s������}:+1��9Ś�H�$D�3�{��M�D��=������ X�hX3��\���w�09Ļ(��L�]|�|���FJ�� L���zۭ����A�c�e(��i�꿟 5z���`�w�%����S��QAk�s n3�ϷV�~ c�`��hF}��4 �;n����ᣃ[����rj���O��w��`���	TwPR3{��3L�'~<�<��Òl�M�CA˟ު��6�e��Ĕ������U�O�����E�p�]ν��l$ PB城L���k�dO��[W�>�v��D!h��4��ك:�O�d�����'��O���$���U]�N�7DRi��ąf>�(��`�o�סOr&���҃%�1��I�������RJ�y���_�^��������(O����gO��jL�`������%+V9��W�#��H��~Wl�A9�������<W�}�=�%�Y�.A ��ˆ,�lVA%��7���0�"{<��fc����x��ϓ�ڒ��{���2�k���T$��Q�G��N��O�g 1��ȋV���y5�׳�����H��צ-�����f��x��c8XQ���P�!����Y��E�9���>_�-q�V�����q�C�����&U�7ws�!h�{E4����UcF^e���;�o���e��B���,���}Ԇ���ʼz���Hjz�GaS9@RQ���LZ2g��FU+��T��IE�	�*��W��S�tr�߇gZ�� O��=�kI��pzAD5�9e��x�]Q���`��u׌ܟaX�m`���p����~q�_���H`>�.�#A�1�q?�͓�з)i��7bnn�5�7�b`�˙M�o��{��R�ʬ��h4|yBl|�5��30�7��I������}h��e�ƋN�M���P������̱�DВ�e�VsBPkLH!�VՎ���({�D���z�S�g?���+�7��^H�sFA=�:�i��\�z7{�fty�ʂQA��F�r��Ï
C���Lt��R�(�TC�������1%٠c���Ǆت�&,��#� �]u��#��f���ϳ���5��f�eLUrmui�9�|Q5���5�����1�J�N�e	��r^^�/��]����X�y|�r9�G0Ŕl�]���%±`V[ֺ4��Y�S٤���8�M8!gWt���B�D���{\�_�D6��Ģ?�<K��/�>}9��!�B���J%,�F�F�v�����l��+�Jc���@>���.�>�D!"�Q��C���P��u�S"��"z�NPj4(;.f@����D4@�ı�0bH>&�
1�..�x-6�D��	��(��}�����-��3���\AZ$���ͻ�i�W*6|)mI��_�o����	�8lT�]����]l�}v!R
���'Tџ�s9\��1#�d�����o��5�>q.��,7X��_�jCE�~ -��:�FiI׎'!'1�5�=[+���o�	����]5��(��2�]�7�2s�L�Z��M��d���I8dz�K5�4*(� ۑ�ʏ�sx���}i��Eo�����L]ɗz!��]i���3����ܱV㜉p�%�?��㔎�-�OK�U1��y��L,�A&�忟<�A*ͤS���:R|�t�zK�Ia�1y�9Ը>�t�"�ֿ+�JY	���fP�q���/�F0��e��P�tlQ���ƿ�|/*Gqwn�&�C%Ő�cՁA������h�S�O��T������ϲ�ȹ�%D�ɋ���q��r�V�*q/5�������Sz��X���$%΂<Eb�5��fFM���4*3�Bf���L,���)��3���ݙs���j�.�a����oA�����Ŗ���^���y�A���4��n������q����i~���S_ި^=q`C�����Xx>q��沄���uv�PƊ��M؂�&����;y����aƙȩ������e�����I��fP�T���"��Lb�*�Za[�[�`8��ыb�GNħZ|��՝���};#4m8��j�*Ɉ9J�N`�i���%sg�	F,ҽ��qQ]� ��yJk;�M�M��!�����\d�tvN�cKI
V����L�A  9�*�6�W���K1C�����$ԕ!h�A'�K�;��#�2�a�U,�����0�Y�=�꧍��! S��)־��{���\���s�p���H�t�jY���$�-�4�	 ���C���d4@V���h��ɪ>u_8̷ҪN��7ً�n7F��Ӿl��H�à��ۉb��܄�?�����ځ�:��b�F_�L/��">�O����N�
��-̬��p��z�2V�⢒��QD=�zF*��f���h��^d{�o��X�X�6��7[��@8�!6�
0�gT�����6�"؝i�l�w�h�ud!�h�}$q�3�>�d�Lк~*��������m�n��,#�4~�p@r���LqZJ1f!�6f�?���&���NXC�ד��W=��@����"0C������-t�H�pc�s��$�=bC���7v����[��N�?�6�y��d����#2�	X~�Ϭ?�9�nыR0Kގ1�ȋ6���!��_���l�cv��j.y�W��s��#���=�[U��Z��c�ַ�2�r�������us,��Ձ���"��?,�t�X�ۨ�䪗�熶�<(�dO���b��j0����BM��C�{z��6p2�51_��ŇC&~LI���Z�WR>�-������	�az����5ZɖPC�Pɢ��xZf��ʌ�Ϯ�=Ts��B9�� �yC�8���I�9�?�ub��\~�p(R�~�����R!}INm�|f��N�D-��b�q1��Wp���-��� |�[&����b��W]0Ov- �ꥶ�T�Ў����:�#G�1�w��km&W>��Q���Y��S��2��V����X��;Piu��ʆ��ᖐ4��ҭ��7�J4�����x���/�UhZ���Lm�Pz��.�q��m��.fx��vڨ�$Q���$Uy���ۻ�/�7�D�]�J��|ta)]����M�k�|
�?��/��&S��<d�0�f�G�3���I��w���ܠ�A7>|�Q��TBU�~ء�U'��x��[6�}X+��+=�s&�������
�C<tH�4��%4QX:X��{�,
����,-( G��7��naIol�2�\�VQ��r�4�M�����f�����z{ӵ�B���d'�cZu��dW���'�G��\���"�A�)��"J�/Bր�Ǟ1��B*��<�	DM2V��c��.!go��9�Ks��뾞A�/�/�YE����,�`w�ǯb�CG}�f���q�XŘ��*�(6~ϒ�Y���ra�rW0'C�*�ǅ3M��V�%�M��W���w���Q�j3|���]ݸk�p>0h��@- ]�قطp`���y��n����r�-���� ފ��	�``�B�xל� ��1�"yWˬ���q��������p�a	��:��?R:1/��w� ���e�V��b�obA�u?he~p� ʽ�l�.�N�V�(�Ȏ_fT�l�xc����2B\�h�n�%)�Ek������=>9�"^�G^�C�L@�Rp$�9@��aA�=s��� H�Ј%�įӆ���~W���@�)y#d��/���s��&��u�UtO��R�{��s�.������m(S���mE&�6r_/^��k��|�\����K4��)"���L狚��
�[���~!���n����9w���Q,x]WQkZ�n���sF���Q1���]�<｠�{Wj��`\f^ķ�B\�^����+#��ת�ծMhXmx9�awͭ\Ꮕ��N�q��TD]%.r���q;�;x���W�3�e_��� J_�u�G@��uJ]o��D̃v��x�}J1G
����B��'�?��C�H"_����.B+�fݫ${�!z~X1�qR�%9�f���K7���?K?!:���,�&������.����6�F�&�>�~(�H� �n/L�ާ]�&[�U@kX=Ks�����"s� �6�n�P�|����'\�vku}ƽ��&��z�(����m1�0��0�Uߙ�^�s-�T�b=ݑ\�m��M׹ �m���Z)�=+��y�;�����tuR���;��Ē������0���М
���i���ߐ	��.59��Aְ'�g�MXz�߸�C��J�ű\��kNc��cZ�lh����	-9jEש�{TÉ������d������R�wb��DE7���9�l���D��UK���}*��ѭ�[�lW���rL��A�R��!<��Q�{F�9��А �5)�1���?�Α5Dc�K�H�Lٛ�$��YË+4�>�t4��$�J���*W�s-�+�O�}2SEu��̃LT1Ⱦ4~��L��kL����hY��7�N賎�N�?�k��c��������k]
�����{�J(C��t�?���5f�m������8���M�͡�k�"�q�����A ��C	[�y�4K�U��h0�D�=�
�fOѺ����9�wB�|�QPo�{)�|m�o�0�<��3����H{�	�e��GE�{��:R- �$�5���ѵ�%�.[a(HL�?@��n��ۇ��J)�?o؅)���N���A6d�\�p�	gm���ieR��Ԁ.>S+*���^[ ��-������;�-�r���a�V_T/cGZ��_o���Ǻ��)��˧b�dc����.�Z�I��yG�rw2	����s~R�"l\�����>���WS�V�_�u��Hj"5��tu0dG7Ϊ2���Ǌ��zx�P`vʵ4�ntF�t��L���C�5��p�3¥؟[y��ڣ�
-)"��}�dX�ѱ��̡��s�{������

j������t�~l����%I�:~��} ��'�I/�5�s�?�_�J� U?\�I�d�K:��=a\�l ����ؗg��6�{o�l�P��$}��;��M��a|�*%j0�C�.�}yd&��@O`Պ�l[���ܓ�|id�o�� }�2qޙ5���ؽg��7�z�uk���
#�Fn`V[S�w�s�p�p�M�^�������;�7!%�o�@F���q��#q@�v�r�u{�;�����C�~xu����AK�'$�3�,[ـ�h��J)#�gN���k�+���;�<������*}j����Y_��?�@I��O*uh���2k9��5����
"GZ�G�b��aͿ��n*��p��0X��l��d=��������%\j_A����e�18\�D�L�T�rE�#O!��e�>�/�r[e8�?�$`P���ի��#�pQ��\"�ؼj�8O2y�#r�x[E�Ό��T�i2�mT�����i
E���6y!ܭo��1�/����~}���G� ֗Pz/L��^�-p�w�E	@�R�F}��	�n`|�D?D���P"E���Q��|��4 �4�f�]�F��
�Mct�gͩ�3����e��o��E���}r=[$�(^���,����x��1d��B�5��Wց7ŀ�6��y[�J+C�Ry��
@_#�KF�C萺k��Þ��SR�د�����W�NO����7b}^d�b�e�9Փ���EՈ!��E*0c|��2;��)�����y'�uB�.��GG�}k�����*�{��nKe�e!Wg��iEۓf��
��W�u�8 ���
y�n�P����+��f�t�P���d��F����ОH+��ǯ�s���8S��n��T����?X>��շ���Oʐ�E�[���"�gā��>�}Z���Ji�}����uYH�du�Ȗ2��}�n���j�;�ٌR��lD�g��]Fc昔}v����ρMp6+%
������И54�Dx�����'N;���4��i0N�<����d(�ރ��qv?�n�lB��~lU�����I'ѐbMqod�B�z���|�I��
p�cⳞ�9ӛ�@��y��������"����n�q*C�ڗ��D�Kw�R<��+��5"1zmr��ϊ��+-?�D${T�e(�,>W�7�B.ϛ�U�5���(�s��F-?���E�s�'L[9.cs8*�eJ�� @&������V�e���j�u�A���g��\���<㮸�VT���xD�+�������
�v��!�Bp�0���.�!;�dଫ�Yy�͠�v����aa��椋��iu� �>�Y��8�UǪt^��.� ���h�1�᝕bSLZ�n����K��\�G$�P4����f��~f@�m��~	P�]J��c2H�Qɞ��~�9����1B`�Qn����풵�_G����)q^��,lΏ|���J��)3��`q3���8�<��,�U�� υ9���ִ_9Ē��Q���&�nȝ�N�L;���gI0Ph����<����IO���@Q��f)���X�0����Y.�&ؚ#�eU��ad\��� 1���r����֢X���7WZu�=�>ڄ$�î�@�ʏ4>n��w�S��{	��4N��#�.EY �$:N��9�j�A�𡫗A�i�I��M���r�Q~Ȁ�$Dy��j��	���}º�y�z�Hآ���p�ڦ �fT�Ddw}�3�Kj�tw�	Hoƶ�(��(������U�:������2g�+�v�zE��>)|0���I77T�R�����aˑX�}����.�h�KJ� �{� g��%��0��㞁`�~�ZY�w��	�Pw7��X�`E�
l�[��P.�K%��A�&��MK��ӆL+<]��<a��)sʋAXQSR��-�ņ����OW�~6e]N�0�m����_�	Q����[`���'J)�Qg��S���x���O�TʾMi!�T�T򄡭���� �?���uR�{�ԥ'�HFH(���L�V��8<[�%tPvib]iK-' ���}��x�/���/�`�c������X.����џ@�E���q=+
��k�V�s�JNӽH�	�|e��Ptg~�J�v@,��EH\[�i�b���<��B!�:�����'���M�@��DRj���w�5DÍ"z��b�?C
x����n;u�M�1Qh=9ڝ��F��Ĩ-w�,��g㧒2�T��Q��)Y�}���8��(�'N�%�r}��ɧW�i&���T,邀+�o�Rq�T�Ǥ(Z�'���)�Oх���t�m�6L�"����,�{e2)��x��{�q��m4��o��G�s�\�k���"����x�2���BY@Lb��Q�j���k�wj�LE�t)�+hv�^��V�
���X����d�|�cb=$M�LmL���җǎ<�^-f���t�<�^�����W�F���uX4Ƚ�H�� �2���ݥ#O*�C���"_�N�'�V�xw�Kh}\�h����qb٧p%<d�X���!���ܪ�����|6$T4m0��+��X[�;[�F�7X.� I(�O�z��~Ǝ�Qy���"e��{�u�hu�];�
�h��F[�(^J�J�a&�,�e)�*<Ύ��E2(�p�H�5|��\A�m�|��M�%~ȭ���{�B32�]]ÄrՏe������x,��&ۍ�7�����݂�ϡ�N�!Z/bZ��N�)ɤ]���l�ѱZ�&�lA��AE^��\�xkeC^�F�و���(�o}��pF�	k���OV mFdH��R.i�D�p��?0`^B6>0`CS��_�r� K��It&���{��<8D3񆖰�C�t���<�����c�� �Y��@Y#[���9S����3���;B�k�c�J����S*3�5U�!��<�+U�:�1�������\�����F�Q�M�bA��Mn�=���YY�?S5���>�D�bZ@�K���לj8����m?r<f^�u	�ړC �N�0������r`d���Re�iXw�m�U�eG+�\�4�n4%�bB>е�R��)�1��	O�^�v.w�R��[��"!Ȁ?��sA�Vnj�H�����҃*�&w�aMs�q��S⫵F��r��$�b�ls�n滥u��Sӛ�m@��D9�ة=.����Fs�O,]���g`���tm*���8�KUNa������C=��x$Za����\�u�L��X��%n��ʛ��s{�,j�W�7{!�^���t�T~��xk+�������7z��j��@u���ȕNMx�
�_��t��Д~3�p7�Qm��M9�Ͳ9z^�x�~_}f�ȑK-�`��װ��Ô�W������yc�S��)�0��>���y�s ��b�+�Ȑ��t�����a�A�a�<�F	�ƥ�[?����{��}���@����\���ʋG�C�Bs"G�67�܆KO�m+���X��] ��4�[pW�����w���Y$"z�4����A��K������1����݅�b-��d����Op������Q�>i"��!�1�(i��bn5��>� �2?[�ã�݊�?׽�o��S~�!��-Q.�j�ms�����W�yr����)lD��y�<}BSD!D�s!����V��q��9�O?|^Jnj��Z����>1s�.�>����eyН(���K>P��Q�K-�����Bͳ�l��r*���R�;�V�m��Ģ҄fg�DV2�OTl���Ⱥ�?�S�t���D�նKO,f���'*��5�:��+r�Ӭy1pm�~x�&��hQ:I��"32�����߬�DK���k�t�F�����=���n˥hm�f#�Fv��<��(�Q�3�W������i��**�&�(\[/�Z#.bu��_��߹\��lMnz�x�$؎����w�e@(X�R�ٴ�'a�JhL��ƹ�C�|�h�u��Od}�4&����g�?<���	��� �������ⱅ|�&
9��5�&'���-��[>�Q���Ft����?�%�qV:`Q�G]�����ۣ��^�[4��pҠڐ���)ȡ������a�:�~)�ݏ�R;:g��p+��F 4�)YĤ��\H��"5��^~��]��C��n�N$c��+�W��v8��$&!�.�\C�v�
���n(�0S{*��E
����*s�@F��,��!T
8���ӌ�q .��� ��)��D�}��	�m��S^l�*:��(,IO�ϡ9�<�VV��x�(�R_�?e�rY,aT�X�:Z��E�ť��2���N�(|�7���1I���mg �>3|��5�ް�R �oel�(����Q�F�Bk)��	�C�=$�5sS����oBn�1����)�v�LaoG���ú�E�4�u�?K(�E��ߵ��l޵)��7}VD>5�GB̐�~���ȣ��\�oo`��r�QtC��2��K��eٷ�q����m5��r_**�?���Y,R����ġP:շ��@�3r���z(����������[���R[W6%���,�F�OڪSC$^B�x9���;u��BQmJ'�! @$�&zs4Y����0������g�K0��L��>e9�d>��y� �$N���q���,͗%Yh�]�%6*�MSf��006j�ZP�(���vv��ǃ�Q�~!:��m��J�k'�\(y&���L*�Rn���z��J�w2֧ % ��̓hEV��6ˋ�@��D���]�Phr�c�9y��!��M!������p�)K�ieb�r�.�1wIQ�ۈ��H%���zd��Inm�b�s���`V;Ϋ@D�?�+���<��:(;;0�T�����:�f�?d�����}HK��G�M)������|{�����k����Ϥ3 R�nf�L~&iL��EA�-@J�/s�A}��mI��#G��)E�O�g�FN�V�af�5��`�o�P?p؟�Do����G��ma�N[��؉�����iԼl���Q�����Wy�h���6�Q�_�3�tb��߬p����^�E�^fʫ�dHD�E�<�j0��v��"���T�wѫT蚚yo�����V���Ltϴ]�Q�v�*t)�o��{S��Q��ˑ(m_�M��P�n��L,K!��fs�Mu�į��`߷�(��(�(����c�N�UU����Ȕ��cb|;���ײeuu�E���m��,˜��+ωvWK��p�8ܶ��6�ɮIc����z����vr��~�u���|����*C ��=��BO ���H���������`l<�����F��/C�c�M�d��n�P�ǅʐ1����̂|�N��2k<r���&j��=��P]�Jy��_�+KS'�G���=�|�-=:�� �N�,y�}��]�����N���\�mp�p{2�a��%�-�R����Vx ��0�Z.`�9փqÃ�� �t�`�7�i����E����9tL{ݦ�-�4��5Z'���Cn�^�?��k��:��P5�(�����aCCpS�ϰ��c첶I�YI�n8nk�����ְ��$�5Y!��p��gΏ`��}�`R�ifց����8.�r��4>Tċx� D�ʖڼv)-'��RB�%9���_j"W��m��6[R+��tS١F�7�濛]��,n`YD��Ic��B��>���ݾ�4�X�
��LF��^�����>wb�]�!� s$�d'�'�s��5���tϗ��x*���N��~Y�}^�/��*2�KZ�n\�"6y,��< ���$�Ï%:�O���_HΜ�8aMM��Z[?9������=�wp!u�h]��,rx3���_ɝ���:c�Ӛ���׈��B�b�E���KÚ{�����x�����B�^@��တO>�)7�l�m� \<��Zk�cj�Ģ�!䳩�Y��A�W�Ip�x?:����@y0FyP+��N�qV�P⎤?`Kh*��~�z�OV\J*8��.v���H���F��F�-�lRez�n��+�Nz���l�m%mD�=eV/��!u�K%�z�����j���y��_��'o�@ym��N��5]�-Ϟ��@�l���Ibd&�3t�d�����]UR~ߕ�L�e�5�H5-w���f4X!�Aִ�]�e^g� �I`��]�P��#���S�.�N����S)�L���
��2Ƀ��Ҟ���8el��.,s&��%C�ͣ�̀HC80���)���l!�y/�XFXȮQu���V���,��YF��Ȓ.K�K7A�S�k�+$B:�Y-}�S�W�t�?xu	 jܢ�&C�h���!�
�|��%N�4@ٻ�/���A�e������=�#�����V9�eO0��L1#Y�R�X_�-S?l��1����L|�vu��Ҟ?�����������T�*�).�b�L4:���[G0J�y'q���� ��y�(�bg��;,�!B�՝��Z�b�CE��-kl���:;�ßHm1�?��K��h={{�O�8dR|
!�u����qT�K���9̑��	n�r��P:%y;V��C Y��&1�%_J:�Ҫ�ڋ����`G��^�ƍ���dy�Y'˾���&o����e�� J)?�>d��DZ�]���*ayC/͒��@��]�ݐ=81������b$gt��8@��$��
���'�
���z�\ c����3���d�<	ڸ�1C�|�D���	�V|iuL���ɨW��JZ-@�&	]ņ �eh
'�D���?�ap����K�Hpޠ�eau�^��G�VI�c{t+v>x^oΈ��M®����!���Lt�U2����h��r����f�!"����f�)m�YD��"�+�Z�vn�������Q���H��M3�]W�m~�.�Җ��0�@���9���\��Ѿb��T�x�b�����鐗EV������߀�M��Z�ʵX��M]Ϊ��.X�_t!����Fw��qڪ$�w뉺��ꪪ��c2J�B�9mP���e��)gMd U�oI>*"�꠿K�Y�OL�LW�������b�x��#���:*�@L�#bLm� �>V�04f,���8t+����V��a��z�f#d���c{�Z��`S�'�9���}$�i�G�d|BJbX���ӣ�����з1 !�hU�~B�$5�V�}�d)����O��E�r9o��oǱ09
O%�����6"�E�D����45 _fv	E����k��D]�ȫ��K���Al]���]��y\E\��I�$�sz�&���qA"o����$��n'�����>X޹af�]�M��q
<���2Τ�^�����'=+%�-�<�uwUѾ	yet�ێ1 �n*̼ǜ_���PB���5����d�yBmL�AZ֔	�f���>�v�]v9	��E2	�Q��5$�]�im. ��0p?�ͼ$J�c��{	r��k|M�ER�����B`�9G��e�w�,[�m��.L?Ao�.�ݭ��od�_��o�R��TV�>XM�`��֭?)�����SkJy�wߥ�����Y~s������85� ��~X��7D��(NH����l������FC�X��f��M��{�p#��3�,:o�� ��F2�^;w5Q�!�������Z�M�������>�K��7ڢi�v5A�uN^���ڟnL�s�[�	����_���I�;����9pͿ�7OR/�E^%���P�&6��d���8��A
�g��?,��`.V�b�\8퓬���F	��y��W�ϕ�j���������Bb���D��Տ�SD���Y�Y{�me�|+��O��2��a+�$G�690\��K���G�\^Y1%�H77���rwL5L��Ƅ���F�ýe��;���x?w�[?ٽ?<�k�7 ����s׵O��`�1K�&�3����ʑ���Ћ�ى�I֚o�&�+L�a-A�XmC]�j��/� �C4B��U�����}ഽ��pE8�k6\��c`��j��"N�")��2G�%��Ɲ��q�j���_��x9����$:L��H*(���(GbD�d0?`���/��[��	����(�*S��4�J�uW��W5Q� ������j����b�(�1T�3�*gK9=�=��i���lڰ������W��8,��
i�_z�<_�z�+L��t��/��b�+b��А�c:{<O��V÷��ΰ5�He�.Z��QF���벐�
���Y�g�&���V��_����x]x?�������u�!��ѥ+Ϲ�u�a!&ќ���|���9�PɁPPQKr�����M"��S/Ԏ�ɛq{��h!n��7�_~*L�څ 5gNk�.�"�����F��稦�1���e/9��?u�e"o8�[�U��Q{�[Y��uV��黡�bԃ��C O�Z�X�U�B]�]q�z'��s��v/_.�,�+��&��/��'�C�PY�L�B�=M�F���w(��g���w��J�%";��{0���-#>���R�����o|���8S��>�5j�0���5q2����_/<+'�m��_��4��_�.��}̠wyo`g�3r�@ts^���8~�����߅>�����ү�i��>z�H��7���T��S��o~����(ʑ�h�.cI���"= ���6��B��q/�N�%�L��U�]j?_-^��3ay�ʹk���N�pT�?�נ5�M77w=�c���<�c�����uf�p��= /-�׆�N��W%ҔM���Ɗ��R�{e�ɠ^���%��{>�@MW���;��-1�P!>xw���{��~�~'�<
O"��-)�S�5�~���	%o$�[��	�y���4�>��p��B~�W�S��%Z�����%�U&��\u!�D�g6-��CУ��dC�V?��/4�ju����ɢ��/�/+d/fC�	c9���h?H��ŏ2%��U2w�g�~W�8����U�����Wi8�i�����Z̟](6`�/?{=���	�y n��$�����u�
���T��M�M��4*�u;�3�����"י�b҄6#�P�S���<�O�av>�0����ԞLAA<N�zT)�����j�I��6�6���!�hf�U������ �㘆@���O�a���
��2R��?�� ��Ƀ�Q��X�2o_q�y)窶VBv8*
����Bk7Z;��?�	H]iZ�m�u!�6;��G�A��}��g,�"U��M��X�/��6P#� ����&��)�k�R͖�FYV�)K�{fY���I�/\s3���#7�y������ ̂���-�T�c/�w��C_�@*�L��P��..'A�O���7�]ӭ��%5�8�V��6v���F}�2��.��u����JF��}��_��,Pi�m���'�I�}v�v��.�!>�0��C?�G��Z����s*����,n�(��!s�ѱyb�s�_fc_�-�'hi�>;U\�����3ߪo#�D�B�O��������ɗ�* �+�8��pW��&3�+��W� Y�b?��	�Q��F4g�\�e9�~|�1m�l��4��p O�����p7�8:I�S .0+�aF�ښ`:�-`�-����p =��o�4}p1��BX�B��he�P����ws�r�F���sG�O3	��'�Y[k͓F�����[Q�0�sA,ߺ�z���{DX�KX:b��Kی�x~ͪ��M�(�"����[�2n�F�l{�z����|]�����!� ��iG3,��5?��`M}�a��Fo+{67��AC�������-��},a��w��c�p7Nc�?�$�z�3]e�`�\d}���ȏ�3���[�C��0����'�$i���U?Np6�V#ڶ��!9V�� ����T��VHK��/HŸ��Hge㈽J�����:w���mNb��&/�d�����7���$�����&g���N��� �]b$�n�x�f�~�G�Y�L\	$W���#���s�D��0�]�T+)=�JEDE�#4ٵf�Q`���(�<��vhӔM\4�����ɨ���G�ߎ�_��,�<�%@�-6��a�x'�k�Ÿ�w�8�"����t�0�kNo��!L�V�M�q�6��ѳd�����]�6-C�GSj>/w��%~�Z@�#���{�h���Lʞ�*�h{���x]��������� \P�Ƿ�c�xPLׅ�ҫdh��*�P���{i�퉭�#O���)�t�fs�aI���wV~��o���i.&��A�+�
�GMK��l�T:R�u�c����B���d��dG��&�+4$r�t*C�#�Q�{��Z�Iz�up�*'�,[^��Z�;��E�E�I�B�RVYs<�d�s2���&���Oۇ?)���-`��L^�O-R�m�k¬Qq[�9��UwÑ����Ș���6j%-k�c�$S�8�M%/[�v�j{7g2��#�Zf�[��	���$h��[>�b��]PV�T0k�Z��`�H��1���,Bهw��e$Ҧ�D�ca��c�Os~��
�j7�~�TM+t륷�C7�\�$>Qv>	���ӡ�#�)Qyq��	�饛/��}�ϫP�_��G3'��: +�Xya�E6l�����x��-:S����f���;3�$`ב"!"!��{+g���]���4Y;l�y�IM팉tY�tǈ�48iG�@`���c�a��<�*��pԴӗ>[��K���� ��� �d"�ȏ}� ��~i�`���x3L%����fo�?5)HL��r�`~u��(�,Ȍ
o��>�'.��`ð��W���ÌH����}h�vM�(��E�+~����u��L�$��wW��T�񹇊z$̔�s��vX,�,�k��eF�pE.*�5O��ǗZO�$��w2HŌ=ia>���c�o�K�z�oHE�G��@��v1�n	���*���tV��%*�eD���:�@ ߍK��p��^W�E��P�֘�I)@��t�~� �(Լx�  y�0�Q�#�ׅ�BO(��c�mkT����Gw� ���A��ʳ�S���{�`��V㇜x"���7�]����q%�<��yپz���G�I�2.T����oK/�Щ�@h*�vb�f��;>���Z��&mZ��\a�K0˝���G1�Q5����=������p�7���^�fac$B�I��8GN	�.<����j!��M�e�ذhr~ ��.M�5�]���������z��U\y�N�sXҡ���~,�uYU�m���
�}X�Y�m�n�U�1�E����f��V��ų��E�R�-Z�H�4,~�T�	���<�[6�|�����w{����X;ł_Ϲ���b�acur56>X�6Z�$ n�m����h����O�7�s�E��t�	T �p5���6��V�ٸ/�B�B������2ܟY\	��!���OV#0�������2$�ժ7o�JZ{��1 �q	�W!F��X�glh���z}NoPE���reѕJS5C?8�מ��]����q�ͱ-^͎zs�~Y�+CN���U�`ߐ���EOb��u���Y{L�(����Lmz�hU��[�W&���e�H��l��"Iy��m�eR�
Q�?V����u��M4ҭ4�$l�`?ߟ�������W�u�$�#��INs��t��Sn���\ y`�T�$kPYK��۳��Gcm��.��/�� �`��gK����}D�6~�R�Ô��t��d6��9����v�":DG�k{8tb�f�����-N�J�I5~�%���/Y"���ef�������M���ђ���������;oOY���t�e�l�{�\�1������ Ӗ��3�`����ֺ�B�>�����/�̟>�$G�s�C���r��%ݢ=��KlNn)R�w���GD㷝�F�N�Y�/T<��&�)���^��5pBف��[��0U�*��-K�۶�����>�������z�\p�pD�L�Ŏwӥ��b�&���g���;��=F�3�50����2�@�Àg;09�V'����796<f�j����ATg#,��{�d��졯:�R?_��h>N�Qh��NX���?oH�����B^"<_O�kxLG���ػU��N�S���#�qʃdR4�	���B/��Qac��w�Y,���O�)��K����Ĵs1�P)����O}s�� ��	/��c8����Z���b�B��6��x�um���iP���>�B�Jp�W�>?���x7�c�����{��蒌�OLS�i�"��_�A�f�iy ���\�OX7�W�N{M!�*o���j�cN.u@���,&�J_(͸�,1~g�|p
Ȑi�DR:FG�zoO����ˀ�n���z5�a�}}����5��;�$��bM�x4K_El�S��e��!o?�w���xM��e��ĕ��8��?�k����:ҋ�gr��>�4� b�
����w|���_�����S�@��q�P�?�iki����	�"h١��N�b���O;yX�C�x��3*���\r��N����gG3+慝\�`A@�1X�Q�<-�n~��[��Z�.��z�@(`���"���T�	��A�ܨ31Vǋ�	V$]��h�-O3H~֜~�=���t��I��m���A�ɇ�����#C�X9�w"�>��w#����:Yˮç��3�R�K{E;���Q��YȊN�R��C_;2�=@��v�<�̲�Z+�N���#
���|������ge�)j�4o��� CQ\K�%9�}{?��V�Ҥ�)�$�Nn�]�Հ<�8����ы)~�dl�3O��(8�OL�5|tTw�~���Beݲ�ĵ�����B��?i@|���;��!�!>��I���߀�������"���d���0�j����fJ���(F>LSɷ�V�[�CP��z]d�����l:� �E+u�� �^�"���8�A40���3��G-�Tp� E��:���x{o�]��Ib`�E���j�M8m�?̈H�ê,?�$쥀D>0�A�����yf��|?�	i	~ys�(s/�B��"l�=�Z�
�z�/�O@��?y�-=q��9<eq�o��><���]��KZۑ�hk��9b�q(}��M<�� ^�%�p�!o'}2�@����ԎBd&?�7��߫O[-�z(���[Q�w�L��:��Ăw����hiPg�o�L�E�gg*(OC����=�c�ns�}.�ٳ���[b���JC�Y����D�]�*k��шXRg����Ŗ���BO��"k'b�$�J��v$��cCG�5�Á�I�2
���R0k�4CP�����Ty|&i�
z����-�?B}�Ex �P��e��,^Ɨ8��yUǽ�����K�L�1�g�~!�kP`��;�.���+Ź�N�F�M�39��0/�:��G$M���_�'�l�䩸���C�M�T=�t�f�m��M����E�̔���h�G�;Y�!0'�X��F|v���UT�����QC��`��&"/ܜX�C��z��Oq��'�O"�t/q�����U��$��}�x�baC3���=&*=X�do���R{|j1O�>a�R�U�Tb���6w�.���F��´�ܯ_��[E����)p6:WꀿlF�Xj�_���ś&L�����Ά6��a�>���|s�v�g�ڼ�DJ��d	M>qY������#�	"�Ϊl,p�C�@���c���6M���*['oR|�CH��'N)ƍ�]�*�[<iw�����i��W��sN�W�3�޼��c�S�+�#:eFV�TH���I��6H"Z�Χ���(Q�f_H�)���`:;�g^j�M�i��BZ���%V�_����M��1H�lR�J�:�_��<��>��.c"5RDOs��֜�M������[�R0�|�y�WUH;��bL������P21���+�#�G��<߀"����l���[
,B���?�5ʪ��Ի|,�-M"�����|w�^_����󜚨�O�c�&rR�\���2ȇ������tP��/��f7��󦑗��0AZLF���R)���������M�}�z�ĺ8�s�؄�s� �2��B��^��?�zyX���]K�1�^"/8�Қ�z2��j�6��oMGM:��E��I���+�t��������m&:z"�-�T/�yPEAOOK��#Igi�D���{��X�uy�l�G��~� J��q�Q��ѕ���^���)Sմ|������#��mϯ�}H{����iex$[�+3	�g�ШnOA�T��C%���!��� �(R_1ɸ��z�Y<���7�|��ffV-	s2�Q�g5��əB"GU�W���T����-�'��>�1�,7�� �?����#��V'� }_e�n%Hw�����:��?U�.�$�i�w���h���]��2�P�Pj}��J�e�QI�V�{�+X��(BQ��i����'ת���j��gW��Ƀ@]�ܿH;�i��-A���IC�j��IXg���L����_�=A�Ŋ5N�Z#�I(ۅ��/�;�y��7H�<c�a�<!�*�0ޗ�Ԩ��>�K�*�s����l.?	�Z���c���Kƽ��)ޖS���� ����#�8G�ŏ�m�U[%Hw�{�г˔`z�X5/a ���!nIO��:����� ����{=�qZ����V��>	��
�KI~:�|{�.�c1�6�h��g�VL�>�H��1H�iy�|_�ʀ)u�g5�푥��+h��|J��eZl�!�=c�k��jeɿ�G�X콑t*q��7e�w�U�����B����=���;x�kj㬅���W�&��U�
������e���=U'����OnX�ǅS`�	���
�Q��8ܹ�ĸ�E!U�i��{�v�R���X������J?�5���b�CT)7R��775y��ɿ�Wbc[���G,�)���W?ۼ[Wk?����vQ/���n;�9���β�"{�ѕj<�0K���;�7E#�p�#��m;t�	�Α(�Xm���.em�(���+��SuY��fe��h!l1�]�F�c+�T�WZ����HѭL�����B�^�ϋ^����=�ʙJ%�t)�,����`�
�#��ϛ{T68�^Ni�Ǥ�"�|�R\5T	Bѫ�`�?��B�MY�	Y_��8�{����V�#l=�����y_%�]ޮ5���4@w��]'�M{�8�h��oVu����n>���{����![�d��8��*n�7$p���4I(ވ�g��@fW�vϫjQC�u:3ν��ZM�K��R����a�����^�Gϗa���Ko^���x3��O�Ƽ�d�mc���4����#��֛�;o�[�!.-@�R]3U$��(�	��	��S�݆zH��9��s���d�Q�3�G
y���7۶�2le�AJ��C���Q]�i v�%�Tݚ���5'��ʑ�=��lbۈM��u6
�Y	���{�B���`��瞸��k��_P�NlWq���V��X���q�7܋�K�H
,`{`���	�+�0�.��p��u�����W�����z��EBL��+�V����[B��pV6�	k$u��\<;w��a2bZ���\��]q x@��l[-�����_AO��<{Q����r�p��.1K�}��0+����/Me1�C�'��dʘ�;�#�Mg����#�mzm�0��eg�5���X!@#i�X���ͩ�ԙΈ�����<ϭ�6�i��cj�V=��(�p !{���+�����K�.d��������@�A��I����ʳ�Z����@d�ct��6������%]�sMY�N�^D���|á�ۻF��͋T$0�?�b�(�>k����� �b:�$�u�HQ5z�|%Lg�e�3�����q�!&m~���,E�߰9%�j(�*3��	b�a�,�;N�Ix�w5��z�����5G��=���P����M{y��s�M	��9KI@h���*��{!��?�1o�idt�?�L �1}Ds9x���耧�IUd,/LEOF��F����	q�A��F���a}�׌�Ɵ'�Gw0��`hc�$J�7�Ec����W��n6�&��Yת'�u+D��c�X>�O�'�<�E��Lw�=`�� iy��l?\�[p�?YS�ٖW�s�Ǟ-�'x�<�9��G#Y!�d���:�5!6W���+g���k	�ݨr��zA��:�k�]�t?�L1<�9N���9Ch�X�$-j�̌�J� �oxϸ�5�OZ�!u�y�����L`>�FC��-�l�qG@�FOY�n�C�~����vq�����A++H������6����7(߈���=.����z�h$'�̻M����Ȋp����wݨyz;oN��Ŗ���:���3d懐:�:qz�Oh�ӝu�����>.j�t�9�;��:�t:ſ$޽�M)�����Z���Q:O����
����@��FԃϷΩ�qLS��B�]��B���+w-�@��p:�zk��W�
#�,_y��:k��	O���I�l��c^J#�˃���)�&�T�
�,�:fI�/ u!W%��s�s����0r|ި��QI�MMUV\���/]��9r���Ą���Z�-�T��L.��D��Q�]l���I���3}��B�AULz��b�(C�w�√�d�w����p,�3�69̃k:�7Pwx{�g�"Isd��|h�fޞz�B�0�@��]W8	�g���ZE�{4� ����p ���NA����i6-Br>U�+.&��*�s<��o��{���m'�k��2U|�N�Y�;�����B��gB�-�8��q`&uI;�ʑ~:�l��v4n���kO~��e-_J4c�P�(�O��Wt0o���R��8�����^�E�`��p��)�,���h�ȣ5Tk�������Φ,��0��8��3����[�UV �e�h�n&5���j"��)L��R]���9��Ѣ竎���K-q�b�Hev���p�X
T�E���jx����F+�X;��o�gJ�_�5H�H�4�N�Z*��0��0��0F���-]�w�7Y`��)�N;G\�X������^�9M�x���.�j�^ÂI� y��a�4z�oͧ##�6��M���J�nT5w���[��������r����l?
�5=g�R�A�'<O�oL��8�甉Ѯ�U='�<�RU�/l幺�s�B�kMe_	_fR����T�O����F��*���sܟ�_�"�J�4C���`�N�lq�e�c�=���ӻT��
����c�`Dd}ۼ+��i��(#Ό5(R�|��S�]4�ݲ�DE~�4aMT�3�g�Ú��xf��׼�|��&~�R{��ti�E1��F�+�zd�xO�p�y�~�̤�<�nLr�I����3��*	��q��]��1�L~B�,��?�R���z�ү���'�#�
6�if�y9y+X�a��ymL'^Xf{�u��{%V\�[1��vϣ�l@�(ҏ���ە@]ݶ>���P���K�lص�9�����wcU �D�
z'Z��X���f0v�MGj�߼[�'�#�(����[3(D�m��r��b���&A��]+&�N��y �q��r�c�=�t<z̘�"4Ep�C+��>4sa]]�V Ă�9�hEw��T�읨��\:JC!T]�k4� O`�r�?v-��$Ƭm3�$G�7��>(�9��� ܻOQ7�-�M��r�.u&��:d�Bo��:t�)x����vZ������d��ڼ���'���N8�v��WB�E�?�A�S,e��r�4�����Bxi�T�s����%�*���e'��U4Q��.mԉ��Gm��?��*=��0<���o��
���&��`�A]��;#t�\������\��|��ܿtgǑ*K�����U%	�hC��"�
S�5n�Ş��i����Rۺ�:���zM.�,	,�|�L�f�2�]�yAOb/u.����`x�W�m&øї�&���G+��Y J�\��A�A��7^� �b�h�Col᷶�nR>�� `v��uk��ȖD&��#XW�h=��\�E�V~L1�@�0�ι�fr\��^���'ɒ� U'�^enM[+����z'S�!<(pPdǑ{�p�<o	������m������~ۭ����[�� <<��46@��(�����[��pdG����]En�%����V�]�5�$S�|�PU��-y�����Y����l�h'�0���J��4	N4�wh�M0�P<��F���ZPY3�o�	�nz>�OT���������Y2,�Xs�����哺��9��fۻ���E)��P�DՀ������G�6�QN��FI+sTXRo�<fl�[����-@ۦ9���9*�:aW��'���Oʱ1r��8���J�R���&	�b����L�˜�'GF&��Yya�Wd��B��"~q�?�q�C}d��
�١~j�0�N$r�@�g����]+�<>��d�J������t���oeY��2�;�z�
��8�c�?��^GV�[����!y!�*�1k`�.�6�`o�����۸����]�Z0�����C%�6L�j�(�����)�<5{8:�"7^F=����m�@5VMVMp�Y
6�Ng(��p�}I��*�Gȷ�8M�TX���\]n|1�d���@��Q� ``޴�(���0����^����R� ��v|�m	�L%�\�xw�<6|DB��8hNׇ�'"x��O�1o���란A�Z�N��DR�[ڧ@0[l�$<��V}��-{'$�J}�� ��d��U������1�8����Է��y��>��)�9�z�^Zi�efs�2�/,���� U��kD�����"9����D��LP-l��:�b4�ov�j	x���sm���C>ќX�Q�Ӄ�zƏJ�+u�ľB2���:c�8
��Hr�e�{Ś =%�DrU��V��I�B�(#��-� U������Sc��ۄT8_��x%�� 2! ������k�O�P��Rǘ_,�p+(���^�d(��d2@M�������L{��o���,��[�H�`�P��p%b!{j)�n�Ce�%B�%ղ�>���h���kC9}R��4z���xwt:�<�\�;F]l��~5^���baw7�W~���
��� �r���/�Ă����D�gG����2��
#�P��g�0��D�Ii�0S�dƞ�잔Uc��%Z�~]*O�+ƕċ�S��Hu|{�G|P�H���]Z�k�jn
o���`�����j��oU��w�!�4��g�?�;x���_�X��D*��\�r?���㡡VM�-D0�
�nS5�M�+�-s��$��dJ�Z߼�up�'�^�g�N��B�����=���9�8>��HC��8�a�:���)CN��Z�jF�p�Z�i}uz�OS+��έrB x�ř�$HW�#�, ��+�����)S.�~Q����I���-h���J�\P1���9{n0ǈ�[D5�D�%�A��(7�=�6b�o� �2[ ;�eE����2FH�ώ�y;�;���EB�~Ior��N��5!���b��M�үmG�,4�ۿ��(�eu�ٷYm+���X��@�ZL�U�(~�����D��|z������p�����	�9�M�*I�:r��{T�[`�pX��gχ,"����Y�(EWL�O����;��h�� ��+r��Hn �g�@�?{��_w!R6B��#@:�&T��v�jJ�u��d��_F�u,0�~G��5oU�=�������Z_�g�.���
d��dGQ�D��^�P��x%>�\g��o�AQ�}�C��<��n9TtڃjR�
��e�-��:gP_�7�ŉ��A��'�R����y��7ܛWP��+�k	�䃣`S�[%y�Zj�ن4Z������
�
]��d^��݁��$8�����W��o�-�r&S�+��y�^�����C�,��@�%���� .JA����4E�F�Akآ����4�Yػm�B�<�!}oŒ����~�?��п?#N~8~H���Q���a��km�$V�3�k�����c��iI��ggze�l���X�2)>r��T���bC�<Ǫ�^������i'Q��;�T ���#&h#���ҝw��W��Nǈ�,�u��N5���I�~�zu�A�����ʋt�8K��_ 3?Ok8K.��o����\/RP��'�q��N�-v�1dYSn�g���V��� z"h6���9�Ĺ� ���m����Id�����$�+@Ȅ����� �$"zy�zV����y�d~۟�j���_l;P��D�ƥ�`��1��ߙ���� �*���J�uS°E�ZPL��H��._Vj�p5�d���L`�B��z�i��� ��%T�(+z=e����F�yD�Owk��л�$��d�C!@� ����Q�3[�{t�qbW}�"�O���u�G�ʞFȠ�k	z&�ĥ�YK�^�<�� i���T.B�%���(U�+)z��y�>W�w�R���j!��q�*\ '�Tǣ	9B�������&�hl�!�a;��������
$	���t�~��:->s����K;F��)s�I�,|�K ��ߙSK}�Kj��i�P�9�?�ho�F��z�N�Z��a�e���'�^��L���/�"�x&l�TO�7���V���t��&���,.}�M����W��ee$�V"a�b60M��Z�LuM��X�f7.� U'���kR肭\=cv�v�+�臹qW�$-����	3b3��RT�+
T!1�]��>��r�w,O_�<��X�ǈn�W�(�Cc) Ʉ�w��$��3Ǔʙ�3��E��^�!����s���ɯ��n>�4VMع־���͌k�(Xr��#�i��x�c� ��"�!��+���1=3��_Z��d��hE�A|����'U4�eBU�0�����D��0߫����/���[R��*r���S��E��d�s��b.w\a7ɕu��HA��Q}A��$q�͕���zJ�L#c�L��Xcf>Ry��B`�Q�v�њ)�oj��������"�뤒��O������]&������	`͎/�جHG��d̅E�tT��-�5v:�+��V%u>n.(�=�'%��)�G�r�@��ƨ~��BBbҕmy����9�߭�rR�k��S���ͿQ�~#`XKȸ����.̥��3�R�x ��}��D[�8�7�6`���|]�dzk�29;=��!m��0\}���b4�RR�I��:.��#D����8F;��%%s/@sc����Y���Y��n�����"&V��z'y��YM�y��m%�Bc;Oh���%�-��Z|��Tnﶩ>���=�+��J6+�����5VH�pa�;ﻅ��?an��C��>�*<~7s������}#��K�9E��^�r���2��`��f��h'�0�\T�ͧ��86���i�NO�����z����K[������aMUM"f�5Q~`K�G��*N�P.���)ֈE�����ǂ$l�#���Oo�"s;��-�&�3R�
%�16p ;C $�v.fq��*ו3ݹY2=NR���(_�����Ј02*;��]߄P�(�Uݏü�L.j`ocP{r�յKj���:�5�N�s	ꢩ}�f� ��y.:��G�I��z��Zm5���BI}K㨮�ؘ�>��x$~�G���_Z�� ��]3�I��n�W��R�L�_�P�1d� v�,�/0��#J앨�<�©�!�j�k~�YQR~0ӆRy�d�.9��%��e��c�hpB�����t��'���6ƨI|�g�l���4��UF��VʄF��T j7%��I��z����W��_�n���\��Ah\���-i�{�������q�{����cPCLJJ��]��K�oZ��MI$��R~�T��G�>ӭ����Q,�W��8{y����<[�S�כ�0(�H	������++�aB��s��\ ��Y�^`��?�Q���G`Qt�o&d)f�=	=��/�=��ܻ���Q$M��+Эy��a��Y��_���NsM�h��)U+��)�溴�^qo���uq���a�	�"�<���@j���§�J��,��p�))0#���o��X}Pz]���E?���Y���Ɩ{p��HS-Kx��ٞ��8Ԫ��Ƣu5�Qπ~���g-=��X��d��2��0��#���\}�Мi��8��n�4�w�ˆ��;��$͕9v� � �/,b`*4�a�аCll��kmf����7[u��%wQ��K4�^���BǞx��St5��{�n9��o[@ݟ����sh꓂ϵ���_� �S==�S�������A�������A���X
���;X;#{%�!�_%q�X
�H�":�R��ɞ1(�F%�9���Y��j�lc<D[����S��+�/�l�G}{;"FSCW�(�5�;Q
j����%r�ee\"�K�_֖1��.��i��*��A��sa~��!�-��jV�a��\D�7��a���|w�5r��m9f2��ߺ����o�h#A"R;�F+�8 �k�墳�J}O�ne!��m[	�B0����I��c= �A��vE(FȂ����x�� h�3 ���|��
W,͒�f�c-ЛO�q�Z��8F��X�r�M�oG�H�Sdڥ�����h	؅P��z����8}S|�c�G�!������)�qtCw��VT��KA�X$j́�St��w����2���Wyq"HI�4' 'UxNӢX�9P�̠�o�kop&j�̙:��cO[�4�o�2T(-�C;E�UN(�����*\Җ��YI"`�����Z��@�y*|�'od�`��S��3�u����`����v��ٿJ<�<���~JP�"Qy��]��x��c�!��o
���x.��C���h��p���W�0,�UIЇ�T��y2R�׻�%�OyI�.�c�^�&f�6ϔ��a�P�(L�1_��Yg'f����Y����.I�t��8�on�餬P�2�ه�Dx�8)�0��^Z�<�J������~��/JS����5��+�
��(������8ɼi�l��	���[m^*��7#n=���|P���y[�֩�hE�J��ˇ{�}���+y��g��+��ʨ�K����Ta+���HV�7�Ɉ$)�H��-R_R�d �մ�hO�gq��.���w`�/��;���;J���#|Hx�A�}4�٨g&���5��}n����,�����X��.�1t������d@��2W��ڀ�8���ֻ�*)�\���z'9�qM�ܯ=!9�By�@N���%����|ʞ��V�N�_!HS�z��ȗVPA{~���� M���I���^p^�34Ո'Yz7[���aQ�t�B��gY�]��M�w���#����~p��m���`����#����][���l��*+Jڨ���&�l~κD"P%��*y�����S8�����J���r��Ԕ ��pQKۑ��fĆ��+!��xS�m9�
D�Ɲ�`A�&�o'@� ��kC���?7s�!
V�t����dk&�QÚ�J_^�)Y���e��1Ip.qO@r���TrB�y��+�ƞg��l�7$$��.D�P��y�ɠ4�(5��<sx�o���Z�,`_�b�z�:��x0b!:��~מ�M�(��	�8��H�'QV]�Y~iz�خ�L���J��� T[v&L��G�����r(�Ԃ)�gG1VZ�/�I�;E�{���/�L�M�cu�)�9�i��Rv$v��Y�����B��Î��xbU�y�}�8(������g��"���Z}�4�n|_�z��A��g��ịb%���L �H�f���4�uD�p�~{�fp�L�=Z5�?!#T�k5��g�a����6Y���h��8��HxR�>�AE>��b%����Ҫ�cB5���^��"����S�ɳ�61�+mus����}�+�����I��A��� T��w�fQ_���K��vtv�"kq����9!rd5�0M���*,���zB�T4��o;��se�i�mn}y��pN�ݢZd��Z�K��͵�5��ĵ�<�02q3i�8`+��%�B-Y��r�3�kT��}�x��1�*����Iv�L{�{Վ�`��CY�@o�.��H�H�i܄��{�B���tg,�L
޾M��Z�D����&������j�O���If�)��eRC{8Te\��峻5� �&pd3��ث�-|��_�~xq�t]�ԙ[s3��,�i���E��Ghy��4�&wm8���	�7˩��B2M(�EJ�ac���9p��,�f'���b`yU\�H"�����	�p�T�fVZ�`�F{K��p��R�0d>2h����X�*��g��=���HN�Ƒ�b���߷/��E2�����?T��i ��� �:ս >�
�aiPN��e!f(����|��*����e��(�g��.��a�����R1�" ��gJ+��Lm:4ՂQI������ށ�P�z[�(��e�p�N5္��nߴ`.���uS��*h�,|�o	�"�-�c�����4֚�`f��Z~�#M@IC��M(�+�iyFy�s	�k#8	T~8�X2�վ�UI��Χ3�	�"�5{]���\��$NG0�M�
^J&��[d̢+�v����;A�g~,?��<I�ߪgE�Q.�bf��߾�%*}�i#�3mgk,�;��`���1�6	1K�h�>ڧ���{���z�=	Z�{�q��e�Ǔ)D�K�	�@�ei\�U�_s�^F���DXL��<��R���;��WPƱ<sp��,�Ԉ�:
�k�����|K��h�Ү/���Y�:���$5�&�R?SJB�e=a������g���U�ɝǠC7�C$k���x�0Q�h���O�~����SP�6�����qC��9nI���lc������p��(1�D��2�52��S�7���%F)��MQ�N�k���o������\Ǐ�6NQ+
<����I�CպF�B��g�v^٦K��W'�q��sOs��ر�f�*��h"x�m�cȺ�/�
��+Ƶ����-S�Т��@�<����K(�N���G�1Ř�����5;�J�rz�20`��Շ�	��A��1 7}��,��vFI����CY�^R�E�`�-�6�|�_�Y�Kv1��?��W�8��XE�R�1�>,1��-N&!�ڡ�x�Ƕ�����Ij�9��|W��4�f��|�ʻHHa����䤾KtI"��Ѥ�h��� mJx��}/5|���V���ԉ�m�ЖG�I0k;.�b�j�}:q�ӯ�UCrʹe*p�,1f����] (R�֩�:�8����|�5�^�|d�V�<�)�ɺ��.{�{y��~�9l��6:5s2K�!1�n�I�������vl��R� ��]�n�گ����Cdt;1&Px(#�TT�#�r؇�Wo���Ol�|an�c��Ϝ�����V���1jZ�2�TS�g�� �iW��O�lFv�/���Y�'��y�J1E�{'���5(���o�D�w���;���ކ�4�ʭ�uV��X�x�MH��	�7�H���+.N�J_SL��i��w#k��0mN�~�l\R����<�ָ�fRJz�0z��&���g���j�>�_I�9�Cle�R2��D��zb2Su���X�?����7���Q�J����drc����#(#�'/�S
j�>~��/��O���c&;�9�;�h �k$���1̩���9��T��jd�(���U��c
�d#�F��*pX�C���HTq�@��1�� ��\�W��~�� M��E����Ui9np�l�l�2no��Ѱk.��L
) ��{�z�f2�L���MT�XM/�	2���ٺ31wd�v��z��)*iە&��r�E ���	�R�l��S����*�O��&����ly�$�dYwג�����E��DX��<+*���� ���u �qAX��"\��*N;y�z��pi�ζ�a7ҵ�=*�4A v��Q�d���)��3�@���0�� ��e6���Y�K#�_͋汦D���.�S�{���
D��A%�����ͷ�3<.��Z�mʂ���ҭ/zԄd�j�}Pn���G6�`��Ql���a}�i�F/ b��\,]X��F4��JT�$������	�U�����[�����2+RPP8�~E'��ʕPB'/ɍ�*��� e����\����Uz�ӕrFvg�1.��> �����,��(4WP�a�]��[#6��XV7UR6y`��	�c�y/�$֎�)0][��=	"���`pR���l��ե�A���Ji����y�b 3���=��x�����K�)�2_n�k4��U:�)
ш�(?�Fː�y��]J�L�] �³�w7���� N�/�W)M2�]��e^7C��(�}C�F�Y�W�y����v�*g�����i�S�'�u^߸��I���ݛ��k��=3�����Ck?�4D��P�(;P���~�Q��(	�]��!�˨��=XFXm���`�/ZJh^s�������!."A���e�Y]�_�FOK��D�{�(&'2ٝ��ˣl͋��[�`� {���j6�X�{��Z�zG�h��n�^rͬ�U	���Q�Y�TR����U3]| b�����"f����*d��?�7�݈~C�x�'5)�2N&m�ȹF'r2����eзo)5$��m�*�>�}V������j�2��u��Lz��yT����T/9BG��-1�Np]��0�1"��'��Y>��-$a�a�Nן��C`z�e~�h��7C���>`HڜmF����N��:��U�f�%cH�-�d�,�[q�_�,$��Ix�J��abbO:e���s�DFZ匃�ɒL��N�h�hƠY�[vI�[D&���BȎ�@��wp^��7�g��tyd�A�*�y�O�*���r����z�B���x���"��_&�V�Cw�������`)����=�A�j� ��Pp&�������w΄].R�6�4�"ۑC w�@�=��ӷmnS��۝I4�"̆QlQB�֗Ja�3`*��wW��q�'O>h�:�v��� �	X����zQ�ġZY���~��:��H��z�������b�aYu���c�U�tuy�W���Z��f~>)^_?3�(n�{��D�V�����j�E��(<�$긁s�f��Br����0c��aL��׏��ʐKz4��	�k��HL$���]M{��j"B�sJד�����b���At)��|��S�������PC0>�Lhm��#eg풊NeMF�6nw�*��E�mV��WX9�&���CF�0�B`�E�.+.&�#�An:z���E�|y��X�%��B"'�G��D�W{�v�]dL�kU9O��<*�^�r0JȪuµ΅��Mh��N
�ros��]^�E$#��U��|Ԋܻ����tK�u����<�Cƕ��
	���D��o-y��r��NyLFf�2�x���d�*��"�3��ҙe̖��
R�{�a?Z���n@���F�Z�c���V�R���|=u�C 4"������^)��ͷ�R����H@�̅9��@l��:g�.�S_.4κ�H�����令�Z�Ң�j�gp�P�P���*f�<4��)���o�w*|�3�ا2GDrL����(�v4�TVhB�1=�bA.���"p��B�|K��
�_�S���n���T7���:;���Ta
aR��l��`��O_i0�_�ap��H.�a�[����b�D�n��|i4���=���)�������L�����k��B��cS���qsG���q��pǵ���U�KF�>�!�RL�
v\��Mީ���ǧ��m��I�`�U~�_}�y���!�N����fLI�����j�M��]g��Ф%�Á~�a3�ig�N2��1�����r劅����lv��k;�@ߌ��,ay����()J�8'�a�u�f��O3 ��8`�s�w�֏��$$������5��.c�I�K�P�]�Y���y��Tf����q�0�yM*�� i2�)��ոce�z�q e C>o����fIA���J���"_*�0��	C��&m�!j\9�g���_��88D�r=�(
eF�fr�um�e.�ZÈ	���p�<���.��ʱ�^wEtnt5]2�:�&C�\��u �)��E�����{��e:�5�C�)P��o�-��[2�*�ƣ�*������q��B�31*{�]_%��!tm�)���d|n߶�<��\��{�� �j*1����,�Y?l�p\�\�^�.�,ӓ8i>Ԣ2a��˷j��9�b�/Aҿ����u�©�(X���M+C��k�F]Zy<��q=�tܴx�v#�l#6��!�N}�ZH��M0����w���G��$�\���r���o�G��C@:��$&��6F88s�sHa�t_���פ$��k���c�р7�s:O5GmϾ?@Di�̸�L2IӌfV��l�6�6��
�/J��p����SQ�ʒU�V[��e�ۭ��ex�Oe�g��R]�v���_A����J�6�I��gRsެ~y��'�A���M�^�Ǘ�rr��kg�D`jCJ�{1:�Fx�37�C`%k��j��zo6�[�T8p��Sz� �jk�.���"w6��NBMK?|D"���8ĝ����w�>�W�H&���t^@��T�Q0S����F��*d2���,�;�ۅ�?�)�S���;������1L�~����N�e���(3V\�5V]��Z�)i����Q������5&r���[��kU���/���G/>���Q��En.��*o��l(�˕m)��R����`�� �r�s���P�S�>hBkWFV����[bTѓ8�:"~�bL�Ѩ�۱��P�=��1^
��7o�p6�h�y0�Uw�c�% ߘQ�V��)>� J@W3��>��7�/���/$g]����S���ѡ�;�%�)���bD�cõzZ�Gz����Xv�uύL�O��ӧf\���v����Ӹ����:l��|����g��I�D���!h���xf��)&�IB�t}(rly���Tƹ��������nN�*�sw�N[Z���(�����V���h�U��uhԡ����(#W��!���vt{{�܎V)�U����^��9���6��+LD(1>ֹ�5d�k�r�VB���7eo�oY� c�� �QlaHhNj����@g�]A4=��Y����H�Q �N��̱�o�8���`���� �t9"7���|,x�|�o-%�n�Z	d��B��$����I��]�͇���Ä	�T���+���4mg��f�|O�!5(����ŭL��Y��u��u�]�<�y1ꖗ`�)e�h�X�~n�J�N� ׅ��������!�X(��'+Z@�Ȫ�
��!r�^J�Ӵ�;�����6��zK-։/"��H{�殊!-+GH����[����<�?���)[K�+�@r�]�����?U���z�g�z~śv{���>ב����n�@ݎB:mV���l�,|&��A�?ˬׂZ�Ұ��GV�7ziJ��9$�E�[*(�A�OI��=Gjߑ9����\�6��Un��B������O�����F�l��u�&[<��Ʊ��u��umD�O�[ܓ�;/���'�����B�Q���U_L�k_L��Z��O���qh��=(bF�p��Dk�|��ɍ���Qp����'c�e
di1a�5Z��A�4�v�3)�O���f�w�kP����3�ӳ�P�M�3����Ϲ�ݐ.?X�B�N�9a�P�{>�� 8E[�<K�܊�,��!n2� �h�������}E���LB��&Wm��U�D���x�
�if|G���.���d-ir�~����?�K�%�A=o������`.�ɑkC�:�߆P�_x���1j��C����Iǁ�vt��>���ї��[fX^�R煬�L�ay��,��_(��QP�!����q6ȷz�����)�,�� 7�W����i���1��S��=�����B�+�U��A��<VXna�1����TL;����ŧ܏Lk(�=B	0�I��������.��=����g�ob5s+elȍ6DP\��u�[E�&���d�F��U�6�� S�
֕��>t��B,�	�"*�B:o�Ȓ�߶�i��������?|U��.�U�:���"��u�͛������G�p!	7R^$�tt̆3&[�88���<%���(������"��[�m e*D g����5����5����;r��i���x����y?��M��N�y �Ko ����=
%���,�ׇ��]W;U�S�uhѷ;H���o��$`@�V�:�K ����KYp_<+�J���(�F�%�+Y3���#��VV�tmK=�8����[jЕ� hm�1�5��#���MzE�~	~w���!��?a�#W��C�KOۄ���_�>&
���5��2%��Ͼ��0r���t���%�M��$p�\�t5�7/\אk?4JDZt��y�.h�����@m 2Z!���觉��C�~�xlyլϠ��$�JZã�i�f	}^r?�q^D`y	��l&����h�����j���j�D@	}uC/��?J&S���T۰Wa����ę(���%�����R��!E�g��;��?����kc����t�,!0K�JGnWv�Q��Q��#�wd��.>I
:�3����oUb���C����X���`�bU2�[!F*�}�c&�/��]�-X���Ĕ�o��r��IS%�r�)�F��F�l?T���N8L$���w֛SS�D�١yp��UK;�ԁ;BPz�@�XO_*��O�ᄡs&��1Vt�W�Aw�BTu�
�F��!�B
�h�f�p��u��!Cwtۋt?�*��B��C�e.]�(Zq�K+4MM}Yf��|FP�0\<ng:�qH2qe-y���]/n��+�������y�Ѫ��q��WLG)��)$�8����n�qכ�Cȳ�۳��ˌ �
®��Y����
Ri	�K!�/*���j�>�T[�f�IJD�2U���L:*����
�^y�����P{^��WГn��f]T��!{�^�x�Ϙ$��pO��S��/�ٓ	;H�Ӳ�l�����<i����`\f���r�CR���ڝT�_���Q�j5� 8�o4�|2��%������0�ƿ���0�hbU���(q��]�8��f����䄮1l+dd���*��5��*F�t�7Ő��f
JH�zў��z��ϵ�g���x��w�b�v���%δR��&��d�K�Ϙ��W�zcj���Tq$c�}վ}ͤ���	rtS��Fe���I���h��1ڌ�h�!��������F�޷��3������Z�0^ط��������=�x/�[W%�m��1�8�'@�!���pj��X
�'�tz�J��M�ۗ���m�r�x��J7]c�P�T���c󨝺�fP���f���@a�m��̈́��*��9�mv�����1٫W��		K̊�=̌�Hɴ-�����H���Y̞������(�/ׁK�m6DbԼ�'p�Àl�\_����N�"H��(58+��)7���&�z!����K裑
N*{�'�r3��3A��!�m�m�W��+�E��������	� a�_�<�|$�E��6�֪@ұNݽ]���C�n�]3$�17�^�q�:x�BA�-<ʼQW��
�l��YY M��P�B%��T��g{��{�kz�p64�)���ѽ����]j�S���bt���%z�g���|N�Yb�q+���)+��"�W���艭�)��^��'.rj�������$"U%�ZPLo9p��5]@v#�.�Us5#φ �zu ��/�r��"D`������=|0s���\�i܇�ė~��2��P�+��ߢ�X���"�����3��Z�:���ow�Z�6�]�%ĝhr�]��\DA�]j�zu���2�	�~�ۜ-�{��KK�� ����	`��{���/J�L�"�^�MGCWK����^ ��6'��0�����=Q��zт�	�,��W�9�.�Q<� "���EA=���
��!o|(J��=5|������Ct�{��������y�O�Zfm�G�L��&H���)��iY��;�f7�ݖ�U��/�tm���2l�`�Qڒ�?�FI�2R��l���m��<�=X��.�R�irl� [Ԁ���+�~o:��OS��,!q�1��E��YN�����%��cI=�`T��5���_ř�?1��̤p�i)i��^%�Ϡ�((�E4���)7=�[:.��vS�$��!�U�}��n`5kZ*2�� H��<��b+$v_��e����L���M<�P٫�y��xisTd�6��5~S�4�#!��VD?1�Pp#�I�R�&�����&"*��>(���y�K^wʀ���/ #s�	S~\f ;Ӡ�S����"���L�)n�9�fA�"-i<��pW��R����t=.S��M}��Q��)'k�?�
(?6�|��0Z�3���6�m�
�X���Su���r�
�iu�$��nm���u1
�� ���Z���~��K�]��ͧ!d2�Du�>)���\�f[ '�F�[ǍH�Y���M̀���l��p�z��@�y���$�'Θ�" �wL�`7Uq9y��D֟r���@���W��w�$���U����/��\?Nɉ�;��{��G�E(,Y��&��<�������hb'*��&
��q�c��vH���a��_��u���R;������{b��L+��J�F?[X������	{r}��l�N0�d��3��&�O�%¾�Bh��1Aq�@#Oe��<�B[���
����D@4b�YUฦ����\,�(�I�K7���i+�}��r=�zHi�$�4��H��s��#��e]5���4ĕ���'�`	䠂ID)+��\y��C�Ч�x�+�H���4Ք�iz4�����?`Qz�?�$X�r�(�o����(���&�y1���A����eŨL<�,ab�;�qYw�PYG��\ �=�Z�y���@�n~�\[4%X��ͯL툳�	�̊_�HM�T�g+�J�S-xg\JOtWj�9E��x��ԓ��҂�py&8@M��q�A[p�z���R��)����Ĵ�h#k#7�A2�O��#&4�_��#����A�Ee���1@�[����|��cU-��>M������vw�]+H9g�S霓*�g1��S���ei�e[�Kn�x�?j�*}Ɇ�'x��6!&�tH���(�����
������=�y8��vg)�P�!�y"�g�N�_��5����-M ��KFv�e�F��焱�|gF�?9W�\�tG������|�ψ����!\��d�,"��%q��L�:F�I����-T���l���;:�Ym6;Fa�z��/����!�{`�U#�������/~�8V(q��F������ܜ��S�Q���sko2Ba��v�r�h.�.ǃ*�������'Ob�S�?_�.��_�ܗk�MP��5,��zZ�v������b�-e��2K���IQ�����i�}�nPnOl�C�\T�?2^��b|қޡ�K�os�������/�u��??=4yj��B�m�&0�
	}��n��"��U�|/���y�B�����r�{��7Ka�x)Tii�Zd��W>*'IV�n4 JI����ii-��^3&+Fc�*w������O��~8�nɛyr	�Ʉ��� ��,'S�s��Z㋁T��6cR�<yU�}ZG��ZQFJZ� VS6���(�-!�7_�9�r,�c�پ�3c��gȆ��_�e�Bysd���a'���^>0���j�J���lH���Pl��<GZ�a��j�32� �PcC�M��ď��+�[��7&3�׾�_�� ��5'�W�w�9AR�^�Wf��Qe������}�- y��0�_E�'Su=��JZ m�u�w]����4|g��	����Ҡh}�u���L�ճ��?d�Z�--�lHT�Z@_>�F��^m�	�����X���[~lՅA �72��+n����i�>�I���A/ĸ����rx1��t��@��~�,����%2�M�M��J�s���^�C]g7�%��f���.�/�Ԙ�%N<������wH ����c$u������rf�`��v�^"�!�R��ٞ��I����)v1m�ѿ��	6�j$��p2�1��W�}�Y��r����S�����l�Ϳ�L]͏�ɦA5��a��,D4ae�ڵ|8�*���	�گ~�@��SCE	?��J��1w������8�'Ʃ7��,���$U�u�G�o���pn0��gj���������Y�ʱȏ���][U��ލQ���G�Cf�
��`��w5��@R��B�m<��H^)%�r��%9�+Ǎ3��eઽ�H5��[:O;E�Qo�~�!(��BiU�3V�^맻�b�-s�U�sJ?�')fR�%������Ł=E[�����lő	�bz�y�Izg�� ú��� ��<{�j�&*kr�C�F�#�VF��ĝ�G�����:b�y�{"7+�,R�s��*��f�剴�Co�9�<,a�H�/������%���5^ߣ��;�m"d�'#̱:ŉE���[n��{5{���kI����B��%�Ieҷ��考��MU�Ab���R�>(ڷ�,��Y��Dޖ�T�GIDO�t;u����
�#��C�ooW�X�`ͧE?^��.N��Ф���]#�l�T�ڨ]��˴�3Y1=O� \dt�R�
�'�ڥq���y6�Q��P���7^<��$�S��ʠ2x��CZ�k,�a�A����[f��x���׬�CE�C+h�5:�A� ��L"a��(Բ�ꉠ����;&�5-5;�����Nz�o���
�X�Z3Ѝ�J.��J�K��)�]��ꐓ!��5ċ'������Cs�ٝ���y4v�~i^,D���n��;�9՟�?� ��\�U3P�O��KG�KىQ�ʲ֩z{��]%��4�zv�S�uh �\m���������R�.'�Iك��;L��zy`?���O/�� _`o��r���N��`ߕ�xyn�έ�PH�!��ߢB�r7��)�2��)ws|�`,��卛�5���yT���*�䧐n	���>j�+��l�	r�yq6����Q�U((�g=�!6�h������Z՟�l�/��)��V`:[F:������䩯"�Ɇ�?��>�����Y��$H��Ѷ��mrU��ذ���v�ι��_��b�h�ep�s;tz�c�rK��jW���
�k�t.m�"h���qh-����Kh��ԯϟL���*�)]ņM���y�z�x�[r�QhT[WW���aQUI��yط����,y"^��$w$޹��l��mN2��-�J`��Nԓ�s���Vyd���p^���gl:>_��Uhš�]�9����`��G���Z��|]]V\���}�n����l�C�<��d��a���Zl��avyYo�o�j�+�v�:�MQ[S����NB�ƃ.8.Y�k2ظ��0^6ɰ�$�7r��h�K,�S�vQvi��Ƒ�Λxm�Z6��t��T v=��Z���RX��x5���I�u�8��C{�uJS�1���S����אU1�����2�N��b� ���4���@v��3��F�q�@C��h��!U�7��j��t��;%�b29����l�!�:~�6�v�v|x�T�K2,QϦ.�ZM����8�ŵ�X�o���M��������ܫrN�Y������jF���%p�T�QMJH�?|��6��4b@K�z��-b�,}ՃϳƇ���ӌ��'6��U++�`O�E����`���O��{���������!"b�5.$V���� �M� 6:�
�9� �����0a�5�
u^�+o���A��������y�oq��p�c�����Y�ٻ����(�Ϧ�sN���fYZ�u������L��?�x�L������k���pȕ���P���}e�ٗ<�����O�yH ���V+'~���a���hYh�Ǝ�f�m����1u1�o���U�\�,Z쿫ˤ�����a9zѭW����˛�G0C$ǃ5�\r�[2ʘ��	�~X���3e�Y>��G>�ĺ���2������i�E�+2:=�,!��P��5�H��Ĺ�����x:�Xq�(��z�Yk��2s��6�$��Ϫ�KaT�cىj�C%�B��TT��̼?p�q"Y��{"DT����TQ.[Ox���meM���Q0��9��h��*��mŅO�U(��S��a�.�~�	�y;��u��Ӄ���� s��^H2�Ka~Ci��3ˎQ����=�5{���/v��!uI��o�&��8�~�=qP�TC�γxT_��
���e��"��0����B���y��e[a!x��Gl�4,���l��ǮBc�}^��`8��0	�O0�[R
x����IC�z0~��#���0�Hb��qA(�~ R����V<�X	�9���{��4��M�2`RI(-s���A��0�EkqI���3���k6��|����@u5��A���.�=~��^d�P��p�,�B����	&<����^�wy�d!���l(���L%_s=��v��%o����tzë7�Ӈ����wNك���3|��ՠ�wx�Q1�t�U/�f
�3W�#�se��w�j��[���ϑ�/����l��AԿ.�%Ę��W�p�R�͞�[�����\4E���p��޾����sHb����e�������)��Γbbc���.Bz�3ɏ��j�V��b�J�� �'�i[��Η��U�<��#��ЌX��ݽ����^���K���7i��~��=E@aP��C���l��'��o6�{��;6u��.C�އ�sB�F�e=���p��p.`�.�^ ��^v:�
�n��ؓssI?�(������sT�e� ��-B�"oԔ�X�~9>�"��7.
�V+��_O_��,�Ku���Y��^{OB�;�N>\N�
^`�8h�7�>D��∠��DB�w�&����N�hE5�S
�zF���$?���3)�VfI��ZA|5��1}���}�%��!Y�<K�ů�j�1 �] �?���������MJ��@�>wj>.�v��+�
��$����i{��ŏ��c̾p1�O^D�v��_4�U��usާ��:4�,���O����ڡT�Q֚B_��<��>E�'��g�".*�nF�õBw��pfvx �
!��$���ly�z�2�pQ&��د��#|\�������?��R��T2�� �~�1J�|�#���R�E]��@*p��k��[i�6_�1���� m�j��ƛ�8��C�~�(��EA���Rk�Z�b>˟>u�5Á�����7D��DLT�v��؃#Ƶ�%���aA�p��=4�/~L%d/��U��d g�EIM���Y3�<h|�Zh��k�U9��*]t�x"-�9Y���������H*9�_K3H"N*`�#���;�01S{|Ʒ�_{(_Y�C�R�	�,�In�k�E2偁Av�V�B��%�|57�ivsP�zVKɍ�q©���˔��{�S�C�P��@R.��.Ν�� ��m��儷@�2��Euc�U��-�䴌y�S����{8��Vˣ.x�*+1{����ȡx��#B��[�!��;�s*�Q9�^�VI᝹�$�rpCUw-g�8�<����Yg*F��l��W���%$�k�u ޽���G��Cd $��^���*3����!'�7�V���i=����p��0g$
?��CU�L���1(��Hs��� ���I����$�g
�?��pL(JaX��n�X$��!�˺���Z�MhGm3��u'Q���د�8g_�" RmXU@Lw�� ��̃%�r؏6�i�ԫH��"w%]� ��*��A��xj5���o2��Ѫw�,b��Ӣ	��x>J]��m����#��.�=�$�}W�ɻwG�(���ʺ�!�պ����ݜ����
}����:�y[�v�s����J�v!HG*F���_�-�{��g�`�p=�Py�\�!H�فYj8��Bt>�NFQ;�ǩiʾ�H]����<젻GG_��ϓ�� z�s�x�>
�*n*K
̈́���5��MG�����o���fYK%O7S� m�K"Nl���"�EV��4�|A��ށ���H�Q#��W��X�Ad�g������\��;6�6���)�������w�?�X_[��Oڶ�D#hE�������6�$���qs0�V�CG�Ч�gT���H��G���d�/��#߽{K��J<v(pR 4�\�r��/;wG��S���YM%Dя�4߸�0P�R%�$�8���?�}c��a�l��e����/Di���P�V���e�sI��v�E��Oaorq��pU�C)�Vc�4������\HzT�9� x��?�۫�@΀P�����X��4�M�4Ζ(G���{�������瞡�� ����Y���α+�?��5�5���p���|���������`����M�۸�����[���_K�Of��)���]U��QKƂ�7x��>pTV���:��ܢZ�l+.�ߊ��K,�)M|�I������n����j�;(�S���U�
[�n��S@,s�7�Q�t��$���`
%v�\�-7�	,eN۸����f��R;]7h �kioIvl�G�5�²�w�u���|(��x����ʽ����N�3�k{�!*/إ�D�F[k���$2x����A��� n4��P�eLJ��:��kp��v���z�C�WjcQ�#6�j�(K#�?��c��D0j--W.��s�>0��:C�m�B�S�Y�;:.��a)�Č���cC�v�r��V�2����SuQ�`D;���0�6Ǉ�2�)��{ZFq`fi+~N�N�v�&[ސ�B�(1Ĉ9��0���]s����o٨hl8�z���C�$����ԑ�FQ�e驐��4��,�!�l������H����[w�;�%:�F���P�]�Pa~s�Q_o]\*AT���I"_��"U}��i��Z� �8��Z�w2ՅG�O	��3>�m�����r^k�!ē�/�℧�J�T������y)%��%����4þ艟}��΂��^ھ9a�,��$%O��1�##=C�b\�A.N#D/�=�y+�G�[D�ҝ��ߐ�7��w�'��Lr���J�q��J����O;�d���@��j�xjM�'Ŧ��q�gO�ŰMɚ�p�j���I�TAϘc��~͖�Y�uS�W�����\	��^�cg9�K��8m��7�0r/�~��X�æE��L�Pq�QQ$oh�/�ˇ���#�䊳�L���t�k��.=M|�� @�G���ѫl%w*�M��}��c$��O���HV����D����OM��<�jK����*���� ��#�9���2UǶ�����mL��rW]���v�����R�<PAbf����G6�r���aQ� �WPU�`�3��ƳJ��="���'mJ�f1t(|�_u#���^B��D5��u�p�"=l{QexhAw��U<�{�P�0<�c�* ������q	X��=$��V���JV,����	^�|dr�ǿ�5�],@B%�q�ń�.���7n����4@R��#~����|dZ.ε]�F%'U3Y{��mE���qv�\���<P#6��6��"AW��ea]^�#�W!O��)e��:m�9ݽ�g��}L蕔w54��g���"���d�"��kU���)��&�|v='O���<?Q\�i�j�u}úV?饓$�Y�}#>�e����5��r�T��/|���!��629'S� �$���#���jC��:��V�dz-�vxK(d��^���3�O��Jzs��2il�ܓ�4�

��>��$�3w������v�	gx����̰��A�F9+k[7�������3��+��mX���Z-�t`A2���2�lk5�J�.�ͦ���J�t���b�}�+Yj�� }�r	�a_���E��8o����`m�`���$�8�J��	��Ew��u���s�����0ԧ�d��q~�W�d��`Ľߐ[]���w��aW���[�QI$��h������x�M_N�����S��8z��S��˓���}h;0H�b[�]� Xf�'��4�a�ѳ �ſ!͕>N���x=;�W�A>�7��WjJ���99�{��M������u�%�+���� AIj�(3J���y�)�9�k�ulZ
�p�*=���+�~�Ӡ�ie�b�<�L1���ƛ�AoAt::f� �Ԍ��
=¶��һO ���?t>܆}=p��u&q�d+�2f�J�djW�_�����$��<���q��;H�H��7� �����&�F,�Q5�9�v��������z��p3�T�p��sl��T���h��N�������Y9��6zey��
���oD�.ࢍ��5�j��0���M���@��Q�	�s�oq��*�I���ɮUA��-Uc��G�~�Γ�}SP�]'��t�ž�8Š����AtE|�^�<���[;���j�Ի,�uڀ)��ls�86��D�[�r�lAS�#~�V3���˿ni,6H�74����d��lZ�I�me�y�ns�&�ዋ=�׊!�zأ�������.c����G2�;J�|�vֿ�qv�lo��y
a�^L�ƭ����z�@��/-���7m�.����?9E�	�E���a^r	C`<l�;җ�?�V�b�c��t�9DR̥�{�7G/Rϧ�aK�%�m���λ�WZ����i��|�u���.Ӽl���nut1�AM�I��j��*L@���&���A�2�#y��J���|а�a�AIa3�^�k�Ң�#(����2<�{O���nrb�!��*u�q����?�a�9ߕ���s��g�g�N�4T��w���=����\eƾI2�ȠL�"�%�����.E�!q�4�(�tb�w�Ji9?6;򮒳�� i|�� <�
������s�{d�|�sm���_�c�VCD���X"k��.D���~w̶wP�O�A���dLFW����J�7M�^�3Ա_O���mv�H�\yGF0��W4�!aqh�tr����O�H]*7ڊw�h�)���ʝdbqѨ:$�����i��+S�n�V1�X����+c��� �/B3>�WE�T��X�u?�Cm��_�vW �2Zǵ�߻���&ʙ:���!��	ǲ6쪣�-�㭵��֯�;Z�k�թ�bz4�xS�O��%���u7��	QR;0��CU��°�U��ĜW�����Z5��S���G�o/_�L�����2ϝ�먂��(�ŵy�܄�~�S�~��t�_��$�^bo� !����+F@���2������k^�p�B��#GX�Ii֚e�.�a"���3 m��-R@d��_eV�,[�"n��Ǩ�X�L��ݎ܆*y�����:V�L)]�[��Һ�
���M�g}8��9`�a�3�Rp醾uT�6^�ا�5W=�p��Q:G���3��I%��E7 �
�����Z|�E3p@(�ҋ���b�L�w$�\��~V��ܾm|���aݸOi��q)�xLD�i@�"�엾ɷ/q���[���U�/;��~�����\U2jN������^�3dO_���#֋r��ϭ���Ye�m������a�q���1�2�/>d�GR�B4�u	�E�P�y)=��#�A-'d��8�FX�4�F�1�%$`�N����X��'�%����J�����Q
�$��B�q4�. wm������yc 	����cvvR<fs�cm������YFt&L�C����gĂ�9)�A󉑱4?:�<֛6,p(���[��V��?������д�9��P��Y�������/�f���/#>}�^籕��z	�@K%A��4@�Ef��۶�[UI����l[#�Q>�
�@��nA������H���RDF���E=K*
��%y7�?`�W~��1HĮ��6�T���UkP�=�??�3����i��k	�kqU���3y���<��.�q��������5���͐���44�q����<����P����ޖY)���}��=jg����U�*Ou�X���U���(w�R�w��3g�ɭ@��_�j��=4��z
���#��SR�mgz�˦$/�{;RQW�Y�.�2I��´(ֆ�kQ5��&�М�L�J
�+B'�+?:VΑ�L�^�8z�,�W�Yo��|=p��~t?��p�\G��<Y�G�\I뻄W֝Q{Ve���j�$ ��1i�#u�oF��pZ�}0�&iM ���g���&YY߃����}%'�ϙ�#৹���t�?��d�Ki(O6)��^ �8�m�/��Y
��ߋГ�4���kD}�t�ŵή@�Q��r�p�gO�#��Hx K������S����$��Z8���y�%����4�0�k�4Flz���@io@�e�Z=�v�8�O�����Xx0�lVt���$4WR��35$�X��B���~��V\��4G�4[�m`G��:xw�2�*s���I�Q���CL�
�T�E;���F6���>i�	�i:~Vp���Y���k+bL�n���
V�G"B�v
����5SwigkHO��K�s�Z��ɑ:�do���H�������B/��S4Bre����9�v��0�ya���
�V~�����ܟҍ�7��|T�.��c���e�i�`��s#��
��}��S�bX�>zv.>���G E99��`�-�r�SU���)tc|O"�l�aP�ٮ��ӖRJ�|�睧��&����M���-c���s&�)�O`��WRW��m�?*lgr~~os�j]��J�Q(]�͡�5� Y@'V4�~~{�*�W"�����������'�8�m,�<���)���}�pB�R��ߗ��gǶ�Nb>�:�h���:L��{�B0w�25Q���0�.�ZI5]�ą��1�5���8f� 3�ov�������OW�\�APYp��'��f��Or�6:���S�M������ =�����/� ���
���f�YS
���L�LL�˰w�r�>ͳ�(\q	9�&N&!X㹗��媩����	,e	�Ŝ�d�Q��a�g���(0�0���į<��ֵna���"�����C�BT|�Q�q68y�D�dCZ� ��SP
����nֺ��~n�{X�ly;�<�~3�����L�2h�7�͂K�~�K�lȜ�pʜ2{�xd<2~����=Jaũ�l淋6�̟�qC�M)�g��	����+<�t��F�&��]Z�`�{�mg�KT��Ar79�5�|�nuڅ���O]}S3қ�����Z�߇����|��q�Ty2cޡe�u���O��[!+�O�T���+�֘s�{���pROx�-X�_��e�Dã�SFBbPP��f�c ;��bTx��p\A�+�<��'�*��wP+f:�r\:� �ɀ���/�ȇ�C� �MHn�$�m�-�� _��vF!^g�X���O,py$�6Q·-���#��C>v\������L��qJt>>�Ť�̙�J�Y`��0��J�����_|񮲷�H �����_�c����-��Ђ�){�;��a��}���'5�͜ ����14 +���{�2q��n�&LDx�uK|��բ�R>�k��\

����*w�M	��	F���ߕZ��V�Ʋ%n����^����S�s̿'�Y�m�j���~�A�ԧ�\��.o�Ǔ�'��S���LW|����Ao�Kk������q:��4Fd/��GB,�<ov�}�K�qk�����1.��P���ff�V�V�	-J
(��b>d�Ϣ�7��2L���y\F�����џC;�]�����7�?Q|\0"`��D5	U�bO��Sip=��t9�#�>:�#������+�_>zXrޔ���� �R�÷�s"�gHq-���ۊ�Z[�Z����{n���3#w���֥��O]洂��8ۇ�'���B~�1�up����R�K�9���{�f�>Q�j8���Bh)s�x�"b������7�Q�?��~[ww��|ŦZ7ef&E������9�XI�:l7�(z�5�WWk,w�[;����,_G�t�jķƩE_z�ڡ.��Cņ�AI_�P���ᑼN��v|�U�v������[as���`9�������t$t�x�0�6�n��ǐ�ޟs�Ìq��\��#uti��HПl�6M�����.E�ʲ/�q���t�p4��}� p���0�:�hK ��9w��!@��Jz?� ��& t/fS�7�1�lV^��7VeKE�Rօ0�����>��2�� �컾6F��6v����%��O�.Qo$B��b��DW���ڤ��* D[ZT�@!�rTz�s��.ږ<�qU��S���@-]+�Qq���s&�\1쇳jל��G~&ӡo��D�����r�놧��s�vщÅ�O&gS~�B����^�	թ�GN0�!����6w�
L�u�qN"[�"���i����z�j�^"��9��w�γ1cR���J�35���>���8��D����-;%�����Ch:��l���Eð��8`����GR`,,\��##�
�-��,�_�sH��!�"������+4��ݤ̂���O�g��RV�A��� .-#����o&뮬�wK��+p"�|V�Ι�����lҴSS5�`�G��Q�%i��9Ol��>�(�j>�	�.��#�m+����^F�����9�>�䮱u2N9�V�T�6��	rƹ �_ �γ��/�p4aa)%�zdQ:���G�+Ho�䋱q*��UC.�?L��?1�e��?�=n��-��%�j�Rz��} ���Pճf�������B{Aa��`	���Z�e��s9�W�* ��nĺL�u��_d�_l8P��hRo�Z�q��@H���-����,�\P�>��f�b��4^O�����;�����<�D��Ӗ�^�d:q]�w� ��:�H ���%Zȣ}�C��8pV��P����і�r�A/HTrlF��W�x�n"�5'�?\�\��& �~r�23���Ԗ�z�.t���>g��
�"$1��M���A���Ħ=]��m��k����GK��Ee��-��"����ω'2�b�1��c�<	F�F�ܩI�����Ģ"��/
����Ĳ����e��S>7D0�i�Z��3�:{XNc1�.�ڢ���jJ>%2�v�{�������z��^��� d��{�02����'�q���\
��ݸE�(2����ǌ���;�<�>�`�6ծ�#���RM"�ت#u�/���A��蔜 n��J�曨}�����9�'�n��㫋M=/�|�h`�<��W�Q��Z(h���p��VނҌ�?������������F��Ы��a|�M�������ɪC#$t�MAim���� �{-o�����ۅ�:�k�DЇ��.�ĠV����Ѷ��Ywe��/�\�,aw�]/B[8���q PX�(̅oQߙH�m�������AH��Dy�\w��
��1�!0�{�|��v��!��:py�d�HcCPv�ތ�	�`���U���S���s�����F����$º/�W�qp7�݊����+�F:a)SE�q,v�e�З�8�&�:����k�y�ͻ��ԙ8�ƨ��*���t�.Y�$�)�7����Z�=�k^5ˢq"=��m囓��%���1d�5��L��y.���㯘R{cr��	A!ެ��_b4�@s`��F˽<�װ�U�4<�m�C��[Z�ԩ��l��hx� �}ݶ�}w�y�ã�4�;iQ �y�n�U�W����X;@�Y��E�~�
�p9�w��=GK`���{��xG�����7�6�{��Kp�%2c�l-��~�P�u��0��d��p�.��0ME�H_��T��0�6�AM��]I
���la��GW/HA.E�p'�{�0����	�n
گ ���Xs��ۈ5�6��)gY��p�Ix)�@��*~T�1��t�D9���m��'k�����a���W��4��R�n���� ��(���KG=T@��ť�]���,*.�v��9pB٫v��Ӕ�q��@z`X(i��R��0U)��~�
�Y5����1��j��;���~;Y��U�G;G|'���	�o=2=A�5> ��ش�Ѭ�$o�4\�z�҃0�ʍ!>J��)N��ٸ?����N�2W�M����B��p��g@֭'Dy�4]������
3$��Q��545���æ��LS�Apu����#w���Z����5���?Ȼ�� 3�.��IiӂHyF�C�?o�l(�U����+_w<�)��z:�(����BU@3��%���B�Qԕs����2�+.9��oVK�'f��Z��<��6]ҋ�g)���Ԍi/%�(����x�*<Z ��HT[a���T
�LBWߎ����[�J ��������m�X��;�b�5�������q�_��סP��Z,2��Q<�Nj�/��䨥���^����<���s� Lޚ�� w����Z�wV����UN������Kpl��'d��W�nE��nFnL���j�[�~j�%�MbP��A��e���̦��ÿg�/GU.�����ʽ���C������,�b��j���6��<�/c�V���U��]y]��e���2��`���F�9���
���a���s�"ğ�}%�=�F�������c���KmyK�,�) ��,����i���zĺ�-��?}V
q$�vٝ��;�l�VWQ�!��צ�Z,LF�Ka�"�]�X!����K���j��ƃǊv� M�����ˡ
�7�M���T�R��=x�%�?�����Wi%`�sV�
UO{7��5��r�i,�~0CGMc��y0�^��ȝnJH ��j*�|ܮ�iDca�׆�BQLD���1��[���q��s�iKҐ��,y8
���\	sH:�zje�v=M1��7<� ��A�t�2%S�����ʲ"Đ�!�K#��q�>ҝ����ũ���ęe��0������j����Q��ԯW�&�[4�D+��{��F:���qpB\nl�'���8p���x�9��t�A��6{���xx�_*�d��u�	�HQ~:W���FV��&��w5Z���옎�!��ƫ���aI�u:�y �0�� ��ZF6�A�gk�$W�n욪6f�>�)Em������{���uM_'d�\�.S%W�r�w��� S<���J�Po��i
���}j���~����e0Q����pj���/L�ĥ��Gt�h̼$k�dSԋe�ψ�F�9�C���G��Į���q����<��{�s���-u����4�Dt���Q����,�K��I�a2an'pm�J��d�23�O���V�/��B�]EdiDO}���0����/���#˩C�' A��#� H��t�����7��"�4��8�`
@�0����~ͤ)��h��S����Yhƺ����}n3�T��e���� ��A�{q�W>(6RZ����sܟp��k��ƞ;��ՙ	i�>_px��W��Y�x	�q���c��؃��}����dQʫH��o��VF��J��A������s'�X�7�:
S)S����@C�GVLG{��%��s��ِf�s�|�;rqq�*!�~s$Y�7��p_��zF���
��OJZ��;�*�Վ���ã�e���#��&!�ވ�u��˹�p�b���6�
;/w�ĎaFx�Gϧ�ʐ�(	%����8�ɽ��
��0�]�[���Ji6�S	��qLg��,��:�ڌh��Y��/a��]������4�c�|��{q�E�a��R0��%��e�i�P%iº� Y������/�y�(�Y+pV��y�&��:c$G֩���Y�6&��p	��@Հ����C�"�����9x`�˵
�c�	�Q�8�X�~������J��1�s�܉��\��E�˥���U��������ćK=��;�ϩ�i#�T�ƥ���*jr`o��J���t���eD`?�8_���"�����Y!!���dnE�{���6H�3|�t��1E�d�}h�S�c\�fz���������C��ߵ���i�:�p7{���0��e(8K
��[I��@?�V!���J1�;y;D����5C�i��T��P��Lǀ������_�j@cSs�>�b��gf�T�Z��~��}�`狑��V��߀�����秽���n���+� �4�s�e�v�����T�0q�9��W�aIxi��}]M-2��/��0v��3}_�����>*�O^�m�g|��!�N�!o׷s#H��@h[�	4�z��] ���?,����?L"��T��N�FY�cj83�4\�L���
P��  ���P/����ƛ�ƺ����H���.2U�v0&C�Gʼ |���c������t��[�,x��Ԗ�q�~�����:=��N�_6H�h�feR�JZz���<���D��x<�>��@RU�V|�$E�b\��y����᭠F��9���q|�'yp��[��/�(��-��QP�!K�x�H�!�s0s�_���71���Ґ�l8Qv�:�$p#�W���.����Ȃu&�%�z�@PhB��d��=S�N�|T�f�J��y�4G�DJ�������%I]�D�KԸ��1�LG�kuL��V��(�%�xi��o��DD�������)��.��
���%���?�����B�^�R~?U��+���09�o�
O3�E1�Yc}�#�|�XVxb�mArs^!��*Y�܆"V֕Z ���ZPEgMW'�q�|���G*�KL��������]��^KC�Z�C�)~�Y� ��ʣx�^�r�MRx��&c�'��Y(~���19�[ �xt�-�5��	vP4�ŵX��r���j)��G��c��6��no�A�c��=�ٜ�!�l�k���`A��l���ƚ�b��5�h��3��F��e��<J��c��Lҝς����Y�z �nYwh� �x��9'�������k4�Ӳ��n�o�X�/NV���l>���i9��V�k��������Ы�����|������Nq�j�r�A�X��*��u<�6�՞R晛�\3*�b١�WL8Rhǭ���5��3���y��Y-��F��o���t���N�ۘ�+$�����l�l��,.a��ӕ/�%;:�KI�8�0�욏�£n�{	�1�',Ti�`��d��q����p�'�o�n���߇u�-`��W��@Jo�\��W�W�������nb�/�����T�ӅAMTu
�5'ҍ����#���O96+{�[$üU���K
C ��&d.����pj`�~��	��!k�].G�A��D���ֽ�B.��OR�ɰ �ǹ�"���3Ḟ'{�|����Q��� U$��m*?0�����4d)�z'l�H��J�(�H2>bس=�c�F��򶼺e��4�Z�h�W�r��3/T�x{u�
}M&��e�U4	�����	������L��$ؤ�V�Mr��1H4�L��c�@y�'͋��`=�3U�^��
hF�/..]ʌP�����.�ƪ�=S[Nb0��\0�c�����v���@���b������'�j�j��se|Q�P+z�@y�������pv�?�J�)	��d��bGʌ�ʸ��G�6�#J9*�`H���6��"���'�n���p���/�b~�e *FB����W�~��]����-�!Eٮؿf������jX���=����"r6�b���R ��y7&�u����Ոt���nӆ�u6�`EJ�W8?R���������2�	��I�!9���<�y�W��U��GQ��+�����#�*�luA��4/\��/�Z�_��g_e�$Kϻ�ݒ�~�Ԕ�{�5v,)��v4�s��t�N�Sn����(q���ϙ�)�WIwir6��f
��!�aR	@$e��>�$�m3 ��������&�>Yu\u��\�.�&�fU9�gs��op[�.C#���jUA�=*�0
�Z�UV�\�O!;]�i�)	P_�^c��!��ָ���!���P�Hw�G��S+��L��'��E�5]��,�0�g^H��ä�cY'�+�1w@���H ��Z��dei�%��B���0��D�8D�z�l֢���'�F��\k>�� v�C|U�������F�3=\u���7
b1�-�E2kJy�->(]n�`38�����/A��A����������w;�; {�x�i��<�v��w�n�GM~�q��Ny� ��r���!�Й�X�{��P0>����4�_iy�4�$޽s�B��C�m�L�,K��0�٧?E?��&�ê���|�,'��N�Cx�&�Ot(/���ؒ�`�]TVP���fI�K�P���jh{�E)���G��F��:���c+�<Rw@&#�?8��?X@MΓ�P�k���h����\���;���g�CM��@X�ص�懀O �ytd�@��׼v>�E t�k��Eg������GVx��N�m�D���:���<V�\QD��$�W�b6�P)�C[�$���$Zy�9�����l�݌|�'��������2z��8U� �N�c�I՜2�"����"�R��G �c����e��Gܔ*-rF�`D9��Q�kb!��^�HKm��)i��
ޤ�Ӳ��`�K�hZ�Gr��>��	��0�-"�v�49Lq�1W��#���BRo;=1x������m�Y���ӱ϶ �q0�}1������\�́�L�NW�P/�>��spa���o�#H�81)L�Nʭ5s�����eE9l �ڿ��%�b`�S���tk��{UQ�o���k$��5�I^W���}18��.��F����g� ��U]���-�h�K��O�m�6ܥ]�!�-:Q���KS3�>����賳6��-��#ɗJ=�f�j�G,�<�z^����6RЈ���".k�w�V���n�7���W�f}A���uf_���
n�~^�4!�Q\��z�Xo�YW(��G���B��JF����m�
����a:��Kq�#�u��\��hڔ��M�{����I��T���[�W�����e�+�O`� ������P�o���u���WG>W��%���`@ D�&�N<�Vc��L ����S�cF��v��L�cTG�[2j��N��d�����[n'�586�������KN��S���\�z�wV �et�V3騏�-e^IZ�H�O�I�W���e"�</T�wPT����+N*��2�O����r��1���+Go�w��o޻�U"���r����!�6��s�1F����ټ=�+�R��c$�-*�v�Ժ۟+(��p�t G�~JM,�<��4
�����W��%a90ڂ�3�?�$9B�����b�\���m�|1� O�� �-KI>��fZV�~�u��.{��$�'wXJ�8ʿd�ر�?|r�� `�='����}#2�"�KO�,�5�+a���u��f?7bԞ�:㓎ɤ�*+!��kNQ:]F	���s�gZ��kP�Vi���\�W����0(��ޝ��/~�.���(�HK���ȍhvp�n_�NXd�O�G��97��ۏ�\�Èyi1 tMke�MW,�h�X����^�(W�d�7&��� C��iH�<iQ��б��u������$/�\�qn����b�qgt��ZOћji�nI��8E����V�ʈN�a�d���ڸ�f��!��ő�nܾ2��#B�^�/�2q�4׃F���ʎ�m�W���+|�b�],�w���i%����e�Q&���{t����ʦvE���J�~e��{r���b������Hv��h��$�Y���[2a�'hn�i���v�S��Q��T�iǫP~��5���x݆"�ާQ NG��D)��DJ��톬��1��t���:�-�,��AI �$t(�(c�̷�54-zծ��і�O�#�T(�h:#g��Wa^(ؑ�Zʰ�%��^b���O�fH$���9�^��&Q7o��˛�]�*T�޶#?O4q&�kv�[�q�� /A��K��@m\�Ϫ�\B7��e���M'��������K9�R-�����m^eW=1}!����S��������$i^p)�\�rԹ�&zW\����)�5�u��u���d@pT�>�����/�<�%�Jr"��L����3���%]'S��:�.����Ol�ᙕMG��N2.�+��|��>��]��h�/���W,.�킋K��
y�ĹI,�U�0ԧ߯��2V��L�uH�z� !�hQ�����Q�39���8U;����\�Bi�7<�C
���۹�@��c�yh�>���F�P�pm95��/�s��4����B��a0�������(�(�.�iOp�>���_��L�le~�M�-�X��ET|eP�� ��<�ٗ�j3
�6��̼b�'i��2���Ekw�D���b%�/�����a�q\t�yc���ߥL�F%��X��cL�s�)玸��X�B��g��j�O>81 �����?N>�J��AE��9����"�P4���F�Ι�;k�[��'�b�}�;���
�p*ē�;�56��J�Tߛ%�&f@6��&�?�p&`�ݷ~�����3����}�I��]*SW�����EQj{P�FŐ[�4��Ǚ��n�*8�^K�	8bt$6x�W(�4�¥��X�[J��C�y�o����7�-��TK�T�D�f�|V�J����}"2to��J+����IXj,k3v>y�	P�Q��j�T�0�D�E��Ff�.�#&�PdX���<Km�S%�N��N���N�Wmn�
��ܑMt�%LI줳�/���՗��,��:?��kFzi�x��<�ݗ�{I�	��FUq�L5a&�Wc��� � }jP��%��2� ���Z�D�J�잾��MId�`o�Qo��+�c�r�Z.8�~ ���
�+����q.)q�F�N��ں͜[�<:��J�x���� ��s�M"Q�-2/YvF��[�d��^:�������p]��͉h��ڨU֐z����+���tND�Z5��(���}�<���<��J�sb��i�@�Ĳs��BY���N��Y�c%��\�-��X�Qo|�zW��iX@7���ό���4����ٻ%:N��;����G`H����,{�UZ�c���R)Q�ZbT��5�VЦE��)п f��V��ܩ�w�����R
�;����)%;d��<Y'g�(�^�@g����m��Cp������I�hV���^���u�W���F�"٨9t˫ �yπ����wmC��n�1�@�|���A��O,sfu���5+P��KU�w]��:8�q�>F�pv#�M��8t��A����F"Ey3��8�ʊ
#Lɲv�j�<��2�g�'^���q��S� U� ��Y�4��t�Cp�J�/!њxT:�dGQ�J%6�*�<�Lg۟K�Ѡ_p�����Q�H}q���1f�c�u1>��jC�mwљ�0��v!c]FX�d�j-m��CX��S�<E�P�B�p��	/ٳ�a
 �֎N�?ŧSGb�<����S���q9lE������P�mq���ٟÓMLg5���euju��F�ы�v��ա�h��Mw����d&��7;���_ğ�PV�ˑz�9�ZL���g*��ib�|��u��H�u��/)�#�W�Ґ�Q_�M��1Ʌa�zhJ�n8hD<�o�_3�/����fO렱���O��;n�'����P�]�?`G����xi�T�D��>���t��H2�,$��}�SO�CR��#R�n@������I30..y�6y� �4�	VC	��G@	���lN�!��U���eC>;��L�RXXy����U*���%�����aJ2��-s�iLkQ��OZ����t�����@�ށ$mo�l �v�w��[�L����e��W�~r�":wQ:�|��^p{ܾ4sJ/1���.�v�)�n�����3F��%7�;��oq=�t��GjK��`6��턿��l�j��D�9�ޭ��@L��6�_(<.0�}+���r"�o���A�p ���<�?��ǼRK���.�H��Dg�X��bd�&����R�qN�ķ�P	2AL�;�L�d���������]�|�o!c��oY���ͭ��w�4Sd�VdȢ�ţ����~���m�_�QBy u[^��I������!��T�GĨ��ΐ��Үҭ�d"��g�Zsbs= ����	�:��T� �.�My��8��C�-�Ь����w�Ʀ�B��[ڠhY��D`��陣!��"�[eF4	�8����B6���,P�����uP0sM~@ �?bqW�:��� 7�&�i��C}T봘�*Į#jҿ���0�����d����A�{|���
��|(/|C�珸�/;pC\$Ӌ�\Ƈ\��zf�H��A3C���e��Z��;v��N=�컿Wa#L�|�O�Yuzx�/�f񜏥m��JC�{���ܫ"!�Q�q`w���4�'É@A��Xib�(�,�8��W�9k���?��j�E�Tp�!�Y�%i��)ŷ�����Yε�"����GOW�v�����>�Ok+ǣ�RQ�3���;��$�Ha��
k�e7�SP����Q�<$��k���]���t��P�?��/������s����Ҩ
��R�X� �v����@����	1 ��ԍ�&�ȹ�n��x�\����R��Ϙ����5��y��L6Gso�s'j�AkjL&�A�KoZ�4��K���[t@�;�*�;צٔ���OK��i�H�Ma*�ѓ�R���FP�n��w^o`��`�������c��H�i���������ӡ6Aө�D7'�ݗF���F�������P�e��<�qY�����ҷ����G��FMtI����1��n%o;�܅�X:L�b���9���'q�I�@Y��VvO������/�	�u�g���7�)O�:�=@c�:�av�i`�MC�hk�
�b?��4�GC�W�E�6/(/�d�����,:tv���2�:��I����s�q@�a������X\ˏt[��q}N	k\[�{�T�����'o�3%6�
����cA���{;*&^��/Q��^��E���w��mt��B0q�PNUx `��� �����^_:�����k�?|+C�QT\W����(�1� �_�n��7.{�nT�?��pLF�ll5;>"`&v2�ZS�=��\�J�kN*�6E�e��W݈���@�7@VA��X�δ��e�#�rf�S�7iNRo1_����F_�5KrΞ`,:�H�qk�u?-����J�ZT�R��
e��j�{SSh�(M�ɣ)������{�l���	|r���P�_�b3xY� Q"֕�����D�y'���N.��.2[���c9������o�|���?�b�#���<�ga�)�Eu�Ϧn��Ȫ%nAt(;����*m�g�	�F����i��K݄�������ځcE�<0Mu>��`+ �8-��)y{��<y����(W�9y�V0 �?���k���F=�����s	)MYVp�YT�3ƣ�hP9l6 X˧�?�U��j����Zv?ci���\��q���0,=Y��l��N� \N��>�xu\�N&�Y6л�ܴ=9���2��b�'z���[������PA�M}d�H*� N�-���'��!��i1^��
D������6�E��65ԧ!�S��K�4���^}�T����R�3����X0���N��.�T(������)Ӊ���L�Ԓ�߈�,3�ģ�T�-#�hĹLVX�z�^�q�������:�2���4����	������Qdރ D�3Fﰩ��d��G�Ŝjb���5�g����/4̻�"��[���+�=7�S�ޣ��:�p!ͫd�~�  ݳ�8�V�����Z�l"�/1��V�
����x٪L�C�<�.&�B���Ͷl�Ӎ�n�T��l�dS[[?���.�i��m�\9�� P/�e�֙��R����5 ě�WDee?!-����X<H����J�ǲ�2C�ֈ�Bƈ�[s֥�DR�y�s��	�� [Yև���?�j�/��k�g;�*������;o�hsB��.Z͏�Y������o�BxtE���@��
R
SY
��M4��X�{���Bac)�vuhl��ԲK�N��,�4�|w��F'����t�E���j�u5M��ΎV!+[��A	F&���p�~!{s,O/�P;I��[��Y�|R.t\����֣���NBS�4��D\O�$�Hޥ��5,�-T�y�����{��2?Z���;q���� #�J{ۄ7�E���s�����+pLz���t�|����N�1�k�<�09_�n������دE���E#�(.O�1��	H������><��v�� 2cH�����c\�DU�9����6�8@
w�5��4�#��{��@ޮMƔlK�+{�����t������[� kA�4Q���wVw���ap��B�C0/�h4�tl^�<Pxb� ��D�!�yo�By�
Sj:؍X��]��G�P���\޾!I3$U7+ϥi|(;38Z�++yl��s&U�#'�ޮ/sf�����͹I�+��G,��]�����L�a((RM��Bǈ$#��d��|"�l����^,�>����kTh�#16p�.�7��o�tg]q�z�́"��&7��y�O]_�̊�����H�,p��q���G����+N(�Ɇ �`3��F~2�r˲�FM�XbAD���u��,�5o,�i�,��=�9 F9$����� h��f5�"N���`.����W1��p�Uc6¿B&�I!�Z|h<����bU�'W��h��T%�Z�����5�0y��V��ߛW6jn1�X6��^�?T��ke�uv#�2�?nG��lR�#�3��@TG�8uB�s`�6ط^AhZ��`E��o/�2���QO����6K>>�W�h�A��z�CQz�D���/Rr�E�C�a�F�=�F�gb�*�hp	�t/;,%��s�b=?�;*lí2�%x^ �����)�GƫߛSþ#a�7i�W7ޙ��5�6�>����f2�!��>��5T����g����-��u%Ue�q<!�����O�f�d<��`lH&w(�E��4tO$��@o�5#h�b��ؠkv�쩌o%:C1�Px`�|jAD���B7RHrT�+���`��^�B���P��ˇ�˺L����<i̝҄�%97�I͙��G�4���p�{�Z3T��I��-p��v
m�s ��Ձ���i ���r�hf��,������9}a����X!����s��fv�<�48-�;vO���9煜s�闕0�ɂݞ���!��H+�@���U(��C�i_�*����`��tosV
n�1�V3~H��0r�ֱ���'RIE���j�:�-���ԣ��'�n/�}�c�p��e�P�f��A ��=��݂!*��M	K�J�L�1��D�vT!��0v'[q8l�wI>�Jٝ��x���9���J{��i|��&��7���wc}�%�����Q��]���N��x�t5J��fOlwr�R.}u���O�dlЗy�"oi�f�cˍN�*q���M�B����Ę}��T��>�qe�g���m`�����0g�nb��~��n��
+��%�бÂ�@]�6��PV�8�J`��I��m���I�*���!��-��[�p�.��Z�"�Ӎ
~H��4
e8�*�v�K<�����qEFN�;ʈ���XZ�S���w�d�x�����T�����~n�m}����d_j^�s��:�~Z]⋦�\!~��Q�e}�M[���[�n4����n��>����s�S��7�r�W�[8��/�Gj ~_�̘ؠQM�{��0F�F�r_������%�2aV��K�.� (�aTb���1��'i�Ȑ̈[�hY�����Y?u�`\C����=,�H�f5tM��I�5�2S/p�h�<h���ݠz@j`އ�t�tT�c���7�n&�����_�-��*��m��h��#��*��W���1����t��OVZ�2���*� �M�.���Po��Rq*)%�p���D	�WK�V8�d�Ћ���ֶ2�%�R�L�o���]��%����e:��^� ��5-%���*�Y��0��hl9��e}���P����f�RfP����Ck�����gx�N7y�F��`%�n�����|�ә�`���Z*�`-Y�S�N��F�#�c�B8��C�o�)Q�x�������ӲqVܓ���s��۪Ծ�XR��D7�qpQ�
��kI��D2��!��3+o
�u���8Pd��%��[o8rz�x�:�ƹ�~-�'-���r�<.�i�w���B�q�f��`3�k�7��r����-\�
�X�o�t�?��~(���. *V2��ލ>��O�%��~Y�<d�t�6;
4Z��x�K�s�/&������B�xd#eQ���J4@�_
�ǧ��XԒ`����	@�m��\I�T.n�-���\��z湩>4�8�ʅt�d�5�����m+��z�Ly�As;����|��Jz���"E'/�{U̊[-�C�;q�3�Ι?	�Ĉ��e�hr�u`��Q����G��}C��kYW�_��f�_��H|꼥��h>�����\CwP�/&]f6��DO���I�2 �A	۠��j��e��R�a8=lw�p��7<S�R��h��~]�}3P�ݼj'�?wa�x2��cJH������ ��3�����=֣�l@�^��~8�
�Ʉ��8&M�$����@�"/�X8'���r���i�<��������m�-�I�G@��/XԖޖ�8I�7& ]S�j��=����ċ�u�7�
�]d$�V�������r�	��G�r-	����
��1Y(��,Sz���,�~5�Qͧ}����I�v��`RJ�*g�����.H��hvV^֦G͐Я-1��7g��=3�Th�6��.ބ�n��7�NR�5!�'6
;��)���~�VG/GX���+H�J���V��[�5+�j;�Ɋ�;a[zE=^� �bv}�px��R
B���>���?����}����Ml���v��"YTFT;u�F 0�6��%���NB�i��buI���͞�;��h�O����@$���Ze(�/�؁)q[p�D!���kM�߷�����gy�R����!��xCp�`�ϟ�,��&�\�-�����1�2|J�L��&��\NX�ﷸ&�z����zIp(��X��溚���Ձ^�� Y@��`���U�<y��%5�wc������K���$�Qj��֪}Yo�l�	��^�6"​F�ʊ�?�"U�uǠ�P��M�nҐ|�V�G�ߡ�wǻ��E����C̒���Ѝ�ú�@@�O�qP���M���$�tV�������įA?j�D��l������T�
�9�<i�''���^0��TG���m�a]�M��E�P�*��H�PT|�[6&�l?�t�4!�3�\J�T��R\����>�)��k��-��5�}�E��yy0�;�,��Y�8c�eZ��J���՝�m�F����s$*6k(g�$M�?�5C�jt������l?=����(��j��#�# ���\�I�ȝ8q(�Sw�޷;@M��ҍof�J�(�ٴ&ȏ�%v���� �g�%�"C���iج����t1���Tg����b,��&��<��Hn�
֣���Y#�uc�d�N����K�x���4����WC1�� P~e��z@m+Uintý�����/�O�)�'&��<(��y��>��z��| ���'y�s�z<o��6Ǜ�%�\���p��X�u!q�X���r��A�d/�����?jw���0&~s�X���h�	.@by�eI�ܹv�8Q�Ƿ)�i���嘠Lw 2@�UkN}Qcu�Cѻ;#2����C ���<��T�C�V�{c���,�F��ro��/2���2f	cs��g=�_�,b.Nmt����.�v�9��MU��R"��kBV!f����U�����WΆS���,^���RT�m&5W0��a�C�tc�T�i8½�9�BK�пJ�`�|t:�]�xˢ��ͳ)3�P�&P���t�d�N�]n�~�h?@2@�!{P������ڱ�p��f�cǜ�̥�9q� 5Pd�q�LKlAԙ�������ܱ���L:��D�]�b�Q	��uՖp��.�!,�h��)/��i<�u�BfoC^8��S"ϼž���>���29��D�x+F�E�rf�Fe6,���ㆅ�+"��dzU�=9�r��+ cE؃VP�)�!�9��Օ��@�W�GR������i�y

�顕Aݧ�߱N>�\H�U�n�-s�h$�c�5�|�wi<��8�}+rmm���aS-�r��τ?�z��$��
qsל�4�<76��~�ۻV��8u��L�9G��i������՛��s���2DEbY(X*r�O�wOg8��<���hX���a��h8���qf�^e�41x�ï/��g��"�%���>�8�#����]���}S�2Jf��'��s�� �`6�k�L:�QN���P��g��	hTZ��
�-��VJ��E#����)�PS�؄;�1+���?����5'sB�W�_�Ņ��	d8�^qc�ײWb�!�p�|v��N�R��#�Z,^+��8�����d��[�V"�a B����0۹��K	?fG��n�Y��z�-�Ml�S�5.h�;Im+�k�^�ഠ��6gb%�&���LN��n��4��$��ÇXS̥C�o]Ϻ|>��P6)��w=:�#�zơ#�ԟb��߯�﷓���R���=	� ��퓃���B��?q���)��f|�	�]�͇�*k�ߜ_iA��c������!���I#_`�62l�;~�Jֵ; ���͔TB�� X�w��鞾�fұ8tJ�m���d"G����F/�.h+�M��=[� I�R]٦\�|�g��49-���d1��c\	oO�%����E�~5j=��.���O7�����s�J��W��}uܕ_a
; oKݛ<(�$7Z�o7���C7��qǻ{>�z'40`ì�Z)M��8JGH��ˡ	����H\g6"D X�mmX@���7�k�D���I�gU���Xq��q[W�ƏB���dg�W,OHC_eUb[�I��t` ���޸�/]��2-p6�Hٖzxr������%oM��S@a|: z���	J1GZ6^�gS�����n���yГ� 	k~8,2�E-�Q&�? ��|[&b�)�\�Ir��i�����+y:�L
%~�˄�������L6�;��:Bb'x�%N�w���N�'P�+��P��	]�"�~�O�^E��^�tmeݡO�~.�S��$O;�1��3�����x#2��,)�:x�iNϿL���?(-��q:�E8ASBKB���5�'��]`7��G�lah]s�"(�M��/�o��z�W*F��X=@W(�/�(>C$(��;�TG��uW�d���+����/�J�J��$U,��c��o8��/�U�4e�a�v�瑨5҄IJ>��R�)�Sre�S�\����B��D_�֞yV���A���(��>]�i麽:l��o�eӳ��
y+���/>����iL�C�ٜH����y�L⚯��%�N�w���Gpz���CT�Eֱ�1�a4)����]��y�D����[i��	yLQ9�\hU��.�VE)�}	#�ͱ���鹸A�~2WC�^��r{<�
 ����l�^�T��zl;�������bD��]�Uј�j�G�٥l�B:�,(x�}�j��bPs_��x�#e���2��u��b`X�&���h� ��p�ā�J�Z>�b8m�i嵰wS�9�y���ٝK�*�1trwq�����BܰykvN�����:Q5��2���D����ᱝj�b��>�W��|���Y���c�f��Wq�N�Z#��ív�kJB�'�����e���f� �G������(}�A5e�2�D
��e�5��&dU��S�q�]�1zl(%��ɇ;�V)fK�B Xɠf&D�������#��J�w^T��|ڹ�,LvM+��2�*�QU����N��aG�h��[`QK&mb�q��P��J�ڴ��؇*��C^�	�N�G��O�?���J�u�"�]����[x|��JL����P'Y_+音t���^�$�;� ���=k��	,p�*9����w�'�AtꘒC��6��q]��6�r���K$��cl�Y#Dp�Kԅ7*=���1�祷��!�f�Do�H��Y�����_y�W�Y���݀.��F��XH�Ni���h�n&YPv����~�����KP@��\"bC�J > z�\<}釓�6�V��vկ�����' t���<):s�HΞ����-ϥ�k�q�-R=p�#u�\��r��{~���[�|X�W��<YCR�PΤ'K��]	0� Xc���S&,�}���ѷ^��cp�u�+-�ۺ2�jJ��Ǽ{;+�w$y���NJ������b�~#a��
9�8jv���fd>�P���A��]�'����m1a�f%u�n��ô�(S[~�w(`M�w\�29��
������|[ŬN>ڿ�2�@�݈��h���>`
�����}�=�6�JG�,�������N% ��s/�|�ow��=�-��k�ʠ	��u��>�Q"�A7b|O`���^�D6�$T�OE�U�㘓�WH3�E������'(v�2
�����3�h=X�d>qW+hVW8�Tz�ӝ-:	���/	�}���8��
���j{���C�U��Áz�m��@G��Rs��H���ӕP��f��ˍ�^��Ԣ��$�)H^&�&tt�̈Jj�����J��������S�^17n
�N*��S��S3��a�.c�8�gPh=�����EP��	���{�%dfNP�h�н@[\?z=n�Ϣ���@�����:�`�o�����b�W��7{*V�[0o�/7|,���ڐ��gP��N���w̻���;'Un:���ƹI�M/��i�{
{"����Ȧ��*�����
���FRE%�k� �(%ėx���-R�p_��@��x{���K���_^ɩ�
FS��Pd6=�z"�c�X�/� ���Z���&2���~���_�w&��H\��,�����O�g�4f�3R���M���D��ƐT+�l���Zϖ+]�f��:�⎰'ޤ��U��cB���c8?ɮ����8!X�~�d->��r�jd��P5�[���̣����wr��`���.%�Jb	|�lcM���{h��qS�Dg�T��ka���Jp�������.�\GY�&�Ҧ�ɢ�f�|�6��n��W[��J�.~L�[襛�N'�r�������	�Oa~���d׷ǂ�4b��a8`��_c	��V�H֥��T�|��1?EN���_,�%�^���񫏤�9S�
	�� j�Uڡ�nA<��K�;w���ym��qM:E�i@�n^e���)��E7\���y���fEה�!��M�P��$�	9�3!fchB�6,p;e��:���u����S��%+��@UW�	/�w�� ���&!S�8��f�kD�I��X6��`ރ��������#��~��A4G�;�>+�O����2a{��Ad�v�ގ
B�KX�.�3�N�!��Ң ���2�$�KT�Fuf�&l�/�jw�����V�k�x����~]�b��0G)o�X⣫ңh�a��]�Z "�q�3݀P\��,�Ho���q��ԇ�=�edA-���v{m��Y��y*+����
||�n=X�9��t@�#��&a��-O�BG��c���j���S��M��H��uu�hv.Fο,�][Z4�Bc�rz0�$��,�d�C~C
�5h!Uc�-���j�a=�]޻��j�n�L�:���P5G[%�8韶y�J��t�TQ3��$ZX�J� %�\���$��S�G�W�n�0����\���p�� w� 쭥�Ta����6)�
�u��>�r��Jނ���US>R����aE1`�g�ɀ�S��崎�m�6�6�v8y��R�D�u�m�צ`T*�� w�,n����a�ζ�F%&:���@�t�ur����-�0;m@���+��H"��Ѻ� �8���+�a�-kZ`e�؝�b�^��z�|�����sՊ'�Ҹ�n�!��wcϨO]>
�Y?$�����Ig X5��t_��=w�.Y˹X��eCڀ��^E�j�Nv��omC�����:�p,�FLʈ4ɓI S�����O/��x
�\��Q�q���L>��^c(���E��f{�t���i���H;� )�5�~,��Vy`������<r"��9�ϯ�E���R�y��VM5d���k��ǆ�$\�[.�p�^M���mM�=��ѭwۚ������]�xT+��b�Kj�tC=D��mQ0�-�+B��'F�ө�U ��}��f�6���4h��V�sN����2Nf�_��]G �mg�L��*���tY
�Њ�{� 
ƐE}i���82�&�ʹH��.��҇�I���ں�9�#:?����[�C�p@H���صy?}*���F�"

{27L�Y�M�ծşH� S@��{�5�wDp�ͻ�D�)UVwHL��]��(��
��:8B6����W��A��~�N�O3�%�.���aI����WV�ܙ��(�fq*���4h�^��:b^��7��cu��!VEiz�Ap$�_g���CM�����
Ӧ��\�g��}�ri����PL^s��]�Z=ΰ*�E����*�k����Y�&�H,"|���m�����L��$��?9�(�Ơ�'<������ՔTϦ�'d��h�����L��+�- �B�Rd���U�+�yԷ4�+��;-�~Vķ�A��\+e���n���I B�����}�R"4J�Tx[�3=�,���$��,��}t�O_c���+)��'��Ϸ�/�Q��� ~�>�����㻇�RRm^�2�ƿ���L-
#�:+Td�42k|S�ܙ��߅�듪� ����0�XZ���Ė� ��>�o�VZ�lXs�c�q_T�&/H.
��5MI�tK�:�Z�69 }�+�}G�Ӛ��Gi��>HVY�`$I}�V3A�?I�n�w�EHn}*�J:PА`���s����RV@%�cl�vKI��6uH~���c�$>���x;I��@>�}*Ǚ߬U����O����S����GF�B_�11���FH5yC6���n4i�O�?�� 4&�u5����l���Z�;ys�L�aZ�h>VV���Ѳ����9A�I�V�A�BjO��ΐ����"'=��s������/_1�zC��L�S�rd`H��aU3'�2�� ��ܵ'J�W���6a�:ʪ3�+��Lx��׽b_V��ְ��������A�Uն��V?�w�f���l/`��O<�*Lq�Kq�>c��m��T �7pU�7�n�d0��'�K-�IS���WD�O��&�Ln��u�]�L�%���f��,
�D�Lh��2
��7@2�Ѵ`Ȟnn'hU�d�}x⻁5�9�:���D��H���9��@"������b9�n���j��o��|�Ľ��/�nPٌnGs��N��E�������&�tp�긩��n�}����a���8lf×E�c��[�.$��y�Ep��U���AI#�ɝ	!'˷���;�N%uh[f
�l�$�,�����u�gRШ�������_h��j������A���9�;@���;�N�)l����@�B�K=�!l%�AkG+&�-n�3�Ԭ]-�B0��mf�S)M� ��~����{�,�SA�݇D,�A����	.*���-�H݌�0C��hW�C�����6������V���%Y�����U���7.� �u��)���5:��Y'�<�b�h�Q�N�ȸ-�, ��՝��V4��RPLסC���=��*z�T4|�T��tP.�0�z0-�ݫ%E�&	��0PXr�К0%k pLw5@�Yґ/��1���x�uf��@O�ď�8���٘�Q��R@�CF�� ��&��vF&����HgJd�o#��8G�ư��nMԟ�V0j���%����5p�Mce���{�$�z�����+hi!F�@�H�ܚ$��1-����ˁ��kq���sE�Bh��iV�;]eC��PWRg�]�#(U����;�3�y���6�""wL��4yV�ӧ����)��o�,Y-Z�GE�W^�*��=V�D*v�\Zo�d+(��)D�9��b�W:���}/����e���5S�/��8����0}|�9�m=�d6W�a��]ihJ��->ۅT@���g�Q�ڼ��Y���	�ѣ�a�ʜ��]jy��9\ȸ$�,�?�Lh��ƭ�@��F7�mI|~i�����v�x4a�Q���
�(x��d����j��^��W�}ҩ�Mp4/CNS�\cZlV�ZNb'��[f�dpS�P�����|�jF����e�e�dx%KYp߯�(�p�؇S+�9'�p�"�w�t�s��I����b�L��Oڔ�NC��Dw��4Y���O��t?�#��Ɯ��d�z�l?۞�R��&E�B�'�J��I�X�M������P���pS� �ne��q<a���:֣�h�f$�Li����P��� _�bY�h7b�2o�Biujk�H �g�B�̼2x�V"�0��2�sR���K�m7����T�} �*���hz �H���1`CN5I�X���3z�DK�Y��h`�#̝2fSfq�ڢ��O3�����i�͹�k���� ���!�U��(�����ž��F��-��#�\�T�l����@���K=	9(�\1T
�r�sc�XAs�j��g=v�w���kL>�R��f�<fR���zxr�x!=��\(�R�����N�B�Bm`�R���;�����#݊cjTK�@ ��������Ta��gK.���S�	���S�� l�q{=�����~`j�2��Ǵ���&�ۅp^`�9��c�Ӈ�1z��t䥖h��l���K�K�ij��=�R��r�j H�yB�_�H���|�F�/�*�4�Vy�]�e�9�i�֥KU�-��ƳWj����v0Ϸ�w-�Y��ƥ!_�$���#�����g��M4�]ɮ�<�v^��� |xK���p�{��y	�83��}��<�=� �r�m�W��]A46Zd	�aY=~VS&t�Ϝ� �3�vO���)�Zb���	F�B�\���h�=�ҕ'O�v����`���|t�tc��L����a�K����q�$��6�hf�1,۟Ma"|u.)4=��L�C���>��o��{���l�ȺR#^��3�xl��)�1�tv�A���؟���6p���}9ٴ�fm/f��*\7@D����OIԥ�P��wI=�c�{���F��c�K^�e�q�E�N�`/3�����A��u��S2�l<�U��{-���<�H��k�<Pd�j߫�<�+�S�R���E
]ZX.�m�Ǖ�d���2c:�y��,I۾t�1rlV�p�%h�RQա�hl�YIl���$�Z����� �Ft�7�2��2:9��'!��붻��K��~�	%fO]��l��F�OpN��U?&[H�J��W���+|�fKpBJ�OS�S���0��JY4uׇd�
L*��}�}���rt@�ܟ��՚~u9`�������E�z��7i��<�%��B�l^�鴝aō�8��ώ��s��d9��u<��{����K�5���kG����r%�o�n6����{�;8�
��Ky^�hB8��͛@�P���Z����͋�E� &��yG�Ð� �׿����~_[@~�}l�.j��Lu�`�R��s��L^6�7ޮ��>;Ty��5�'��r��w�|:0�6 r�g2�(���c���Nn�f{6F���ړiߝ+/4C��Ȕ�tuG����G%0�hy�m���g�+��!�0��Mj��Y�R�}��8��ԧ�`y�.i,���k22�7
P-�?�)��+@O�݉�f� ;��-��, w�>�tm����e�8-=�3\oTj>��+k2wjPm ��I�Ϯ�"���c[%��ĵcqp�/�W�	�����s�T�����K�E�#�tY�|����-Bu+�9F6��\�:؄�k�Cj���_N��K�ӕ�0�z
�f����P�읡��oz�u.��/ePt��N��ۻ�%Ā�T�6��ܴ
E:�E|��U�X')~��4�_j�=�J���ƅ7#s��u�i��W8Q��� �pm�rs�B��ag��kbM�Ϩ{��r)�� ��o��
ҽG����*��ߩ�r�\=	���GEm©�OEi�X��u9bɕ�z��ޙ���~&��\�"�}��oR�̩��2
6_���ôD�B��	5�#qR��#L�#�o�Cp=>u��Gh����`�R�o��|A��d�LE�ʼWUUM�d�*��u�5h����n/v�֩�H����ƾ�z�5d>����!����0�.��^
d1�޶Ӹ�����o��V���*
�E��J��FjS�y;ۿ2�ǫc�=o�/ݢ��59�셿�pƋԋ���<�.⤫���y®�9Y��B%�w� �5���o�g`��w`X?;x.�G�G��-��X�F��H��*[W�$P��(A>��{Dr��8��g�9M���N �~l�n�a���MXޔ���E�Z�ߑĀ*y��p�cs�v��T?kp,Ww^ț)z�3+z�Ƕ��UĀ��MgК�9�֨��	M�;;3�����6�8��b�q>Oi�P�	��z��8E�癱hV�4�% Ě0_9A��|�)��W�Y��ē���쁐}�3�'o i������Au�);��	��G����M��Z��X_��{J�9�����^�2��~W�-��n,b"�_h��C���qe1q��8*R�d��.}k�>-���AV�k�|Ȩ߈_����N�����8y��J�Ya���{L�@�.A~xzG�V&V�o��xXF��j�7#r���y#C��%@ |�d��2� )�,A\[�X�}�s@����c��r�Q�M�pE�t,�,��n��1b�y֞`�mE��,�d��Q���]�E��� L�OzXD�Q�y@�r�6��R�6�h�0�/(ͩT�:c{G��h�5���u�bps5H�>V֟�b���?���~�lZU���,�5���'W'#��E�u�:��wԚA'+���@z���
B^�	ϊ$xt����Ѱ�\A@6����$%,��5��U^*��}�_��p�0��4���3���CX`����x�K�[����l�����"[��M:�/U�}���*�P<4&I�k1�}�(j�8\)�H���x�ܺ��/h�{��^`T����Y��n\�Ă�r(z�Y_���䭴S:��m'�b� �	�
����홈׊�`�η�2Jc��z�X��z��剒�M�&�,��A�@%&j���;��?�K�v-7=.޿����C�3̓+*��Q��R@���[�iM�ϒ�`��(�����r���	��mi�f��'~�̬���N��%�!�~����N/����y� A�o�h����>�{���S�ۉVn�K��>c�u�����+�MV:��Ru˻����I.k�W�	�SF��*���q�2ɶ�"Q�XD���4�������9����Վ������	)A�����b�f$�I��O��L<j��t�]�$KV����,�����~#��{���5J�13�0|��Ԝ�]����fE]����)��"�
1���/$��qIͽ���M"I���@�AA����V��w��ǀi��؀��IQ��������9쒋�YH�Kܐ�nV>�*=VWF����z���8������XZ{/0���~&f{V���#ϰ�p��U��尘O�������1��TV���}�dÎ��&�����vou�m	ېA�,U}
��� ��:c���t�cq�f��֊�8���$bl��<W-Ck0n��Y"�dg�8�)^�,��D��Ճ%���F���s��#ֈԶ-#tp?=�tRGp�'@�3P�g�ڋ��c9��������9��(/f������6�AXi���n�?���+���ɻj/���0���w���|��҈��m�L�����{8�!D9Q�ζ�_�L5v�dY��PG1��d&6|k����r��}��K��QJaoj�!۾�Cv|���x�b(�w/2����P��I��{�	�o������z����6��b��B��34�t�����;�����6=T��=7��yPI��,������a�Ls�,�յ�Vo�~,	h{��N�0�c�u*�oL�̸�p>�z�:�9'��}]��_����w8�?��D���Bm����E%��
�X+��\9�u��4mi�z7��36p\�}��I|�	�q�U��S�韧�C��_6<��Fu�Yx�0Žߧ��ޢ|�����+^2�M�@���+�Z��"i\ƕ֯Ō�v�������_%o@�X%�Rg���������rf�]^�6Pq�fբ5��Tb�ܤ�O���lv���K��ަ�X�٘w��S6<8k&�qr3-6��҇��|$�g�[�@i��p��0[�s��b4^���VSp�����z�p��5�j���'Mpe�,iȡ(N76I�-�BuH�F�1�����`�Q��\c��U�y`�u>�1��(-��)�����Y��4b������.X����	BUr7�lP�Ѧw���f�X=/D@9e�o]9y'��a��?s��}.�Lv��K΢d��;d+���I����+�-�^BT�E:�la��P� �����Aʤ~�v��-8l-��Qx�W���#�u�̧�rU`m����\vO�~]!Ҽ�� ȅ�)�� �Ƨ�s==��Sw���D�j�`.L��DK��Ac� ���xFߍF�9�!���;�2!V�^K:���2��(w2_�(F����9��0����\��F���.�DM>���E^0�����%�A��8s�?9k��ߊ��B����r����O[��36�%"�էi����^y-g�O�d=̧6���V����̿�E���M��ɮĶi�����]�i:,}�X@�b�
��H���*1�4>&N�
ݢ3x*|'�2��
f4��b�L�^�D��� �s��Ya�/b����yK]���p&�5�;���5��\�<�[C���?�2g�y��y�/`��{y�T�{zДS���d�qI�J��&����k��+6���Ю�J袍���Ƴ����p7i�D�];��  ړ:���߁<-�1YHoV�9�����!��n(<���c��N�t��l����Ȍw��T#9��;�����3������#�������9�)V!��/���A�PCPgz� �zaG�9r�9=8��G[���Qc��^��E�W?R��MH���@�ӺC\�C��W����	h�Vz���kރ$�F�!�7��f��K��\y�8� ���r�	�U�J��I/0����鮬�ň/����P��/�۫��2��2a���M���"߈/&'�OZ��B�95D�߳ף��ۚ��\��0��%�ක�~J��I���	�"U(4T��A���P��T���RǛ"X�i�w��8aH5, �]�� ¾Hf��Q.x��)�V�x��6���������9;��o@~N_3MOtu�{u�Q�{nL#�I���A3f�h��b;������&�*uk�>  y�(�V�cO�S�19pvt�hJ*L,�eҶ���+ez�x���ĸ��joL��'qtP6j�}�^��w����1T��,�½���Ƕ`)���k����C����LaZ�����Q���	�Wi�P�sUK�zՊ[��ޣ�+y��V��ViG��
�I����"ɭj�f�>$��3���u�E�@��"�^p�!V:�D�m�eL���v�g���҇�[
���VU��A�B��/�)���%��s����5�d�q(�L%`�!��/"�X���x���u�}:x�+&y�z�#��#Wv�Y�ׄ��V
�����6���&�r���r$Eh2��/���?�39�UWuW�QZ2\hX��oY���J�Ң���<����އ��yJ@@���)�3zb\G���[ļ�Ej�!������� ��R���ޛ�vD�jGt"��`|���.JT�} �8�9N7�ay����qH�g��ˊ�\��+� �vɤi�׬2���(�J,��e��uTE�?g�I��TVqW��i8���-��3���{T���Z@*�L>H��eNv'ڹ닛8�G�s��4�տ��l��'�]$�~��u������V����~��eU���B��@dp(�1��j��QHL"h�-:
k�gw�`m���Xos1iH��q�B�@���/e�� EzvcR�hW��%�y���hU�$����Q�
/��$/{o�Rh�%���`�eonNf�� �*n]�"�;��`�_t��t�,������)���56x �x�<���z�p�kU<���t&N
�>�|�'Z��@0r�i���N݀���?��J�j��_^:��~�(܁H�rU��h2R9���:����l�r_��8��q0�^�R'��E��\�l���&yN��ėǆ}��11��}�c1�Yo�F���Y9$�|�c��X��7����6�~wR}v4�[��"�y�6�R������Ǧ��t�p|NN��$�JE`�\��j!� R��<	v��pYZ�]O�x��1���@:7׫ ����;�i�u�t���y8|��21�^��f�U zwR���V@��� ����4ɘ�1�̦��FX_��A��᧸����u����5g��Z��K�F�h;�	>j��T�������1�� �h�ͦIΫ����`���L��)��Wdq��%����E�� "��/0~�tD�a8�7�.`d��)9�⋧��,zV����h�Xȸ�����%z��j�>�F�b�b�Aӝ�KД1De�<(Y�w�b5��(�����䔵�nIje�e��AԎ���-���(��O��h��G1�#�g��72b�Y�V��~����5���W��7:{)�J�	�@��6�;{���@��ܶ��\$DVg��4e{��M��CR�N��o��5l��daIjK���a�6����ҟ�q^��/���>=�'[�)^4k�������d��p;�Ib�3����z(ɝ�e�B��9���X���ņ�[C�Y��7�Ӕ&C
g�\|����W���- q+ ���z�l.�l��2W8Gܘ�%7]�`;= �`b:�-�ƌ(��DO�^fX�5xZG&due�0�>SV^w����0�S��>ONΦ��ɢ 4T6���`�`�E)"?#*g�9'���ܚ4P�)&]Gl�s
��#U�3N��>�NUV;�G'�PB!� " ��ΉpR{�2O�gΠܑ��+Ag^�(]�$|����:ʡ���q��ܭ�	]� �����*7���zjA���d	���˜���qg������X��}����X�Ń�9��e�5m"rG;����	%=q`,�+17b������@ƽ�̲�X�=�IМ�Ha)��q_&��sFm�%����� ����Z��j����b� ÐK��%ދ)�{�.�_rFy�����Z�ӯٚ��|l���R��j���8
���x��doA�(���n�CJ��co}�iヿ��yB��t��\��e�}� �:���d�,c�Ţ��"�{`z�K. ��e�������+N�
����$�f��������Q]/`�K�������7����ƪ��G�/2�:t4ش/����{�S�t�󧓸`
hp��Ҕн)�c-�ɱx\�wP.�<��c�5s4$v]7�m����0�Rbk�7�-�p�g&��'���67Rk�&���s�����s��>�0CT�~f�y:�aج_Gۖ�Ҍ"U���`�9L��-Z&�7�����iYz�,{��6>(��[�Mn�,�㾐k����a�T��9���F�a�@��#y/�NM�!��K�U��l{�cw��� �[��z3ѨXX"�u��>J/�wY#q��qK[��3(���B���*��}ۘ�GD�m���8�Ĝ���r�T<-�e��|��,�X	�c<�����p��S����Y�wTV��[���Cz��KD�M��X�[^O��qL��� �$ߧ���L��aH��y����,n2W��@�C��ܾh	�0��A�"WᶩX����f��Rz�� lޅ���b��X1�h?�S��$��S~����ޤ��D�Yv/^Q@�w�۟�!TRd>z�Z���+V��cTZ��Cs��ε��G������oɸҩlL7'�&y3l�Ƥ��j���g����]9@�]\��T<��&�d>q�x�Α�ҜUm-@t�_4�-���HS��jݧR��0,�;��9��`�Qt"d��v��}ǵ��Z�_�t�Fg�װ�%u���Q�v�k������eb���Id��e��q 2���5�^I�4�,�.�hxͷ����,#gǚ2v����$1���Iw�WܽX��{�"P@�� Fᵘ� N�>uK$v6�Хɟ���C���G�^-NI��@�a��S>�?��{�=|���<��9�Ҍ�6t�H-�~��sI�f��j�.=��8s��l���G:;��x-A�O���p��Ѝ+u-�7��,f��β�2½�'��2P���Jr����bv�vK��ŉC�љ#1֒>B:�)�3ih/�	���.��~�\���!��lN��Tg-�Rx�[��|aZ:Th8�<�.D���V��y6ia�9��E�F3��|�@q�[����:��۶���h՗�64�3����6mX��a�,��}����ieF�yq9��>�X���"T[.IzBA�q�V;������Ӎ+���J�̸�q��gU�'����G�t�Ǝ�U��]J�a�̍k�)�"5��|E��eъoV+g�fz�λ�������oRG>����1�y�s��K~�E�������;�JV��IGTHfHΏ��]~��\����$fT)��8_�m���t&5¹*&������i`Wk���FD:Z��q�l�������K�
�>.o��eu���-���c,����8�r;`��3K�T��ς*� 	�y�'Mr�n!r�
�CϙϽ��֗sl�'��z������岁�����F�,8;���[��=��H��YB�w�Ē%؇���ɲ�X<>�AR����fa�RA-
�Y�hn�N�ј�Q�A���JP��70��jk71��Zk�ҁ����[A���V��yl�m�_	�*;�3�R}=���8�>���Ŵ�� ���ڜ�+��>uR��&jx�l��YSt<�0��Dk�+�I[��֞���~wX�w V��HO��+Z`a����܈mep�ﮌZ�b�9u�������<��=��ÊQ�D_��F��}Sܵ�#�3�hF�ެ��DR��j���p�c�wV�|�BX9/&H��A��2��D�*��;�U��?e�P�*���\�&�V�m�y"C��7x�f]8Xk��x7�{_p�9�2a�V�o�j���v�x�٣���tp��Y�s��)_k�P��'�\�p��=�ϳXc���Z���38�pt<k��;E1Q���Y��v�n�߷M6{m�2�(<IIs�<W�����D�u�<�iJ0�vR�H���cd�6I�����a��R�JF��v�����h��J��aG@UPj��y�᳒����}�.&6�"ϧD��XP*`��ђ����V�y��r�~o�R�وΝe�9����1�[������!S��x�?�M^��c�m\�,�@����q��àDűB=Tu�ES��M`�cCKZͪRK<Y�?1�ibI���kc���_�Ts'0E�a��$���l�n�0�n�U�d�p��
��t�G�0ݾA1Kc�G"}S3�Ko�`�@�QZ�@uFWx%]�a�a/��u�9��zt���{��R�"�nR� z�.JGq(g��ѹO3>���ST*E<G�+�JE�T!ʯU$�������d�W�OJ�x:����gozc{�&*�A�z>X�����v?4�j�]�S~ ����V�D���a���a�/9���!�d��x�b(���"s�M����r����k�	Ak����!IZc�4hk��_�V��r����6eҞaVѺǔ!ߍd��V��?%�M��S
+s��\|a��<E�D���Ʌt�is%�ф��X@"������^��^%Q%{S��S���$-�ڠjrH��6�W��)�9Q�f��W+i N\�(����<a���_�=��ڵ֌s�ƫ�RF�>��NB�ß���!��R�=��W#�@��L�9"1��f�4ٝ�'-|��{=@֮ 1����b�?�3;1KNw�u��&t������}l��>\
H��~f�kW#��IEV�\~~ٷ!d�����������Iक़��/{V(�(VL��LV��_Q��&ÿ?f�����!}1��)�3����ӔɭIj�Z#(�E��9�^&u*�ɰ�z���?蟑���Q��y��[����la�`�	&�0���C#����	�����P �}�o����v����Y�-T�$��*O]���H���G�F�����:��]�ha7����&�gV:pOjb��K�N���
h|���xS*��<Ŧ�~=7=��27m�QS���!�bk��.�"�r��Ŧ�?��;�ũ���!:.�l>g�=Vn�"��v�(%�mO,�-�fsI*�����읜�$R��1�B��C(��	�8]��Ht�a�~���:�z{��uk�V�1��������v��c����ZƋ�[���:Α|F1��b��Z3��<i{����t�
ؘ�u��H�+�8�|��׎�m�������X��p&j�t�g%G��W��/��@�3-���m�4�k�K)��_�E�5�}D���D?<�>�ΞN�;��'$�2�Ӿ��P H�h{�mf�+��ZΒ�f�����":�[/�������$��K�C����;�2�KI�?��*2�;�rjT��mvݠ4Ӿ�������W�<���Vf�<h�c/�@+,5_�BY�E&�䬫�Y�����ur��Ē�;�b�����s�s9��m�cci��U��Ll��eO~����1K��>n�y�ۋӎ�G�.G�t�Y�
h��v�jz�xes��q�����H�u�a[˿! �<�Um{�Ձ_�U`�@B�_ߌ-̺�	��2��S�li����}��RB>l�N��}�z�'���bH �!w�>�RZYɬ�+ޠK�)�
�� %"c3�$�ص�A5砨�IB�3�Wɤ�~�zaS95]�
\eH��J��v^����D6H�`���R�[l��ZUP�.F��=[Vű �[�M{u{���T�0�n<P���!,�}٩�/|���B�@3pEZ��~��o|�a��8~n�a(���R�
��.ӄ���}�dug{J����\
3��Ȫz�%hL�\�Y\\�����z�'J�ֿ�85�ő�p�5����
Wm/���~ˀ�\��"���2>����S��ye�.�PU�F�p"ܴ���=�����G[]QO��2��¯�i4/Gy{�!��C�pm���]i��%��ᑣh�I��W*����l֒R$��|�������V`�d"<r(/Jn&���+�w��K�f%���-UNЛх*DH�n#/}�*���6�����&��s��:	��h��e�jn�X�a@N8��^�� t7*�}�;�}���emZ`6x+��$��ڡ��׺k�1��iql7;�@Yf0��{��Ŏs,�uE�)�ϻ
�T�;��CGI�U�>@��T®��n։�E @�[����������j�'�~p���M��5��rb"�l��zw��G˦�����#��"�S;��i#���ޫ,7j�[����$ ���1ܳ�q��� Ɂ��8OB�����8����0+5�'_�r��F��S=�ޱP�<>W�	��q�����w:qh_`B����������@I.�`#!��	_\�Z����60鷸��7X��-*^h��S��^���v�W�j��A��J����������Ԧ=ew���6\��6N�r�1��ϰ��M>�L2s�D,��2z流3ho�@��Dݧt;/�#��U.̬��� m���q F���P_F��ܐ6�h�= ��D}�]Ҿ?���Րs7�f������y�n��W���D�*�\��S."���,lŘ�7ʐ��@����I�:za!���ٰ���S�`NDY;����D��X��hU`��A���[p�ɄN���[=�ImD(6��n��7����6z�	���c��4��[,Mvq&�$))nPt�;��$���S&�K���VAT:+S���HnQx5;��U������������@�8�fF�-��C�����\1�(�d�A(�_��Ǥ�3�ć�0�- a�m9ە�0@	��%�P�:T�V���R��Ȭ�'����%`�!L���6�	���_����~��3���wK/FCi���J���S��]�v^�>;��${��$��l	��&ˁ��4�'�]�/�}��$�+�n6i��=��EB/��{O�Q)@�
�R]�C�����90���l� �9!i�2�ri�uq����C�#n*�C�8���@��d��3�����ٺ�Y���	�̑��.�QUr�atg�� ��.�ܳ� /�5YRd��Q���Yc��1��l"Lf�s��)W*��ic��H��t�"�.��IM6�IW�5'c/X��S�� Va���&cRi�އ}F����w������b	tMޜ頼� ���/��8&o�?�Z���J�X����D����Wl�SŊAs&���l�q��R��:��/�p=pj"W�6�_P׈��Z��SH��;�����d�S{cs�w�qG@m�c��h��T��\nP6_2�����N�������`S�� ԈYS��5t~�`UL�	�9�n�k�z��PpWi�ʗ �!/���7�~������ձZͧ7�!0e�#ۇ)8���U�߿�_X܀s7��4��t���dEˏ�9�\%��s$�p#g�*1%@�j��&�\�H w~��(C	'����aџ��`u Y�n��~�l{羷��"������G��8�/�X�S�jt�" gt��^����z��x�5Yz��$�Z\ʝ'�6�r��N���%.�;0��.v���P�厅������D ��0���=��+{���M������
��̾쎶��o�^��C��	� ;p<�5	d� 1oo-7vA�י{�[*�'��~'�%ǂLa���$�2� ȇ9��%iY�i��}o���ܽ���P�un���'Ə�)�~+2���`:���J�
2�%w��P>M�Ws��18�
����1�Z�2��l%�;�*|�h��%���=��1��!P��i�;P)>0�Y.�*ےl|V"/���7�ՅpC��5�a�u@����oP���$n�:[޻<Es$nqn��tZ5�Y�i����� [�6w�2�g"Lk(yzי����0������N�S�s?]"wPm�Io�0K�n��{|YL�T��4��Bw	��~����-E%�C�,��)�cP#g\��oM)�a��b�y��n���6�LZ	�P�їH��B��|�-h��X�e��ĸ}Kt��%Ȋ��p,����X�տ&X���Є�g�Ì�-/2�^�C���Ȣ�P��S<BS4��F����k�O�)YJ���'+{�<��p��ȧ���?N�.�`(�f98Xh� ��ɏ�E��E���ϙC6�� �d�rR�m�L�1_X��1㶁G�����x�b���e����X{6���4[�_��$�	~�>B)q�u0s�H��v��P �����I,F�.{@_R�V�_ׇ
^�6>BW"���:+$��.�va��Hc<L3n_�D'��ɖ"�7��r?�VKj�����-	$$��tir��nP��;�ʻ�)��a<1v�<�9o���5�x ��]s!�\c&Q{j�H7a�#��Yj��)� [��n��:`r��ߤE	~� ���lh_�Cɬ�˴>{�"����N)�������-�"rۯ��|8����j�/��5�q��P.Vx���4��(���B}� �ȅja�Y�5[�Y�_[k<���Kϲ)C����$�?��Yx[�v���g.�wX���|!�) ����,����_��	/N�v��qc��r��^��,=+�����b�˯�z7��(Y�Ƃ���)��5�uM�&EA�A��z. �G����c�
�s���n.��1�Ŗ�Q�` ߌ�f~Xc�ngz�&��C���j����E�(
�(T)���>L��Kz �D��,P:��2�\-���'�Ԯ8�GB���EJԇ�ʆҾ���o���$!�&&�z�fJ�*��vN�o�Bb�J�G#�.&|-�<��aj��1�
�#�?���YV��*��Qʕ�C�W�{�H�����;�U�9��h,��ѓ���r�Z��؂|ϗ�&7� u�o�ȇ)�CWB>(�*2�-kgɅ j��`����GN'2p�_S�zee��?qĥv7@]R�U��`�^��U6��p�R��,K6�m��B����3$�0�j��͙&�]N�N#޽	J�)��X�h����ڠ(�3m�O	 *��Ϣ��deU2ln�D
��k{�t�4򊙟άE��l�E�"�`�*�5� ��������ab�Ug�W����n,��J���z�8lɎRn	4��K�J����jbrZq.�Ռ����O���0[�F�&�;�r� ]A��/T��ZӴ�Y�\�d�d��V�h���4�a�a��RB03��'?h9���E���~i�5��B_VIꒂ譛�!�`�y����܌d/��3B��m�ʋ�'
�Ը������ �;JN��OH	bc�
H������Uz(�� �J�09�خh
�~f$�?I]d|k���	�{F�<#��vf>�/e� �q�k�/v>�iu뻏���mc��`��O��D��Td:�@B�NR�"�ZW���<g��X�}@�1��7��'��/�̍��ԁ[�ܤ��0��ʌ��1��䞟�ly�����w�	��I�Bܦ+�-�L�?���So�b��b`��C��w-kbhf��Rڝ��?X<�Q����Q�IGf�i��BB	˿��`���h���NZʅcQ��g\�
ү|�V�,f������+�G5p������P�1�f��}_�P��e8��ujɳ.E��W�d��$�\D �P�%z������V����(v���+f��c���~G��oj�R�$;m��9����� -lY�-�J��:�؎lk��fj5|�z��&v�
＃�Y@i���H�����*�k�9��#X4�X����Q���$4{�Xv#j`�D�ҫ�����Xf�z.^|^���xQ�u������d��v�,�h����|Tw��E�AF>�~����i7m���$u���3 F����k��3#����s.^Tºgʷ�m� �SbJG �f#We���6/5��X\��;M���X��_�/�1��t��:'� ��5�t�j���u��(2~'i;x��1:)Y�Q�"PE�B��C��;�3%n��Ҟ��3о���ola�f��q�px�l?��}@�ao���[�����O�P��e���ް!�˱�4wsxf���Q=��ԑ�WP�`����p��p��1�O�[�{�8�����|h��$4g� �FW�r�T��`�Uo��oV��c��ص��!,I��Y��޽h$�P\�&F�[�o3VP̭�X�m����M���RsM�Q9h!�o�������0�B�΅��ꮈ`�J�48�������<����ͬ�O��E�%�	"�3���u��iT��(O�	��P �U�,�Q�8��Q�Dړɥ3�B�s��%氃��A��o��hɁ�۲l��w���*K��%�l}(�	��Ho�X[���I�i�SD2���(qJ�.R~G��}�s�)wz#pp�l�p�e��=jW�3M�R�h�u�-��b��Z�s�m����T-��Hg�
=�mPdŹ�7�]����g�,܈8Yvf{֘�+�aRu��K>�+J��ܤ���4=a�9����(B~
����T��\���A=9�PՌ����5�n:3#Y�{:y��l�_����q�9bg������OJ��)���,��'�?GO[7k���N#�H���S?Ī�����.y�d~mܖNL� IƒEQ����B���}*�k;�2����d�w"X�ǖPO��B�E�H�@@%���8T���%`����=m�bB����R�H�?�U	�w��C N6X�@3Q��^�|p�������x��(�~��逜�/S�#�\�3�5����=*��	o����8O�p-��0R�,N����=�Y�]:��'w��(�{��5��C�~q�
o��ndi�d;��,�|	����:�V��	��b����SP���y�� sȏ>8���^"���-�4M_w���t�Y�w`?�d�	���|�n�d��˦e�)���8���9]����WAde |Q���A-HB���b`sC}��"�Vg��]�̪���O�&��/^���n��*��3������������)�b�T;�E(L'�U}"�cY�Rt���@���y��aj��(�fLoߗʚ��ퟛ�瘟YPG��Sa����t��r)�-Q�"&�٩�Xb�<�V�:�q+���rP�
0Zf_SRml8��J-�;��fc�$ }a!�Yp��_����m����F� >�}��h!��d���akޢ>����d��D��#�J,$���ۻ O�b��`ݡ�V;����S'� ʺ��o�'�7H�������E��(�J�:�d����<���2'ꧦ��DY@�e��֘@��JuQ�M,*?9hX\���AF�j
bo�@��o_4U�]�p��9�����C���e;�(�lⴁ�r��%�߹�(�@�
L)�!4�¼CA��CoAd��]�*b�;<jk�䨖op�A� }c�����%�T��3=0	uP!������hRq��U��#[~Zh��f������fʈg($��e�w<�N�Xp!�v~�@�N����$�3Re�,��#��U�};K��ѨdQ�
�<	b��n���,�Wnmo�]��'.�FXi��6 ���2�e��C>�ꐟ5�<������@��*Z����'
U-�!4��ۙB(�R�6�Vm���몑9ů�������{ܮ�m��I���1�A���mϺ}�٣��cɌ�ڨ0:֖����X�lQG���*<�ץq��\�:�����dWC,�J�t�����O�Pa'���&��������IWG]q,��<��q��.r�ՐͿ���n�;�� %qP:tOե8�E�'j�GWm#	��%����r�:r��^�W~C���7T���w@���S�ɪ6;�{���w�����Nk庲uO�&��D,u���n��/�?ZZ��fw�jT"n%�B�R�����,�����(3H�<��'j�Α���3
d����'�VVC�g\�H�#go8g�x�i�P)Lկv�����L�vk����&OV����M,�+�YTf�����v�d�������;��c'�Ip��m���Yo��Q[x�E�x��������Ky��b�A\�>Ѯ�$0O��s�Y��kN��'��"��+H&`n3�P�-ԧ��Ծ4XE�}֥�/�ؾLW2I�������Q��R���g��������M���D�h4��'c����nޤ�I��J���y�4�z\�r�Dbw[�z���f*i��*��U�FLvHT����m3Q�gK5�F��xC���!C�I4tͶ�~�8%�z�3~������ϱ]&�f.,KEv�^�a��Y������nYl�ݰ3�A�7!z�*���ɽ�	W6�|��h����SD_ڋ%�����%
R���nV��C�<��M%kc��l
�5����{�]�v�]�����)�A&4[r�j�5;d�@x��v��޳j�:����vrf2����:��3:��oD��U��+ݓeZR7�L�؏c��1��bx���U�hW<#ͧ��7���_�U������^I�(�iI��o+Z�~4\�Kh~;�Jm���G�^L�VI��)�.��IU�CjW���{�l��ԉz
j�jl�6țMKC�ƃΉ?�����Q�B����F�.����ڧ���!|q!kQ+������:�d;�����j���9�ƎD��u��N9�7oA�}��x⺷������EO�g@�Qʲ"ى:���	�ǧP��|�����+���k�{�O_��	��:Ze cz��ޏ��|�!�6�p��K��a�%�dl��������9�w(���"���ufU�Y�AcD��"�f5a�G��"ƠyRU��P�B�ڲE}mF��y3{�6-��	��?m��^����vV����$��D��������er��S4�(3��u�D\ɣ���6ƍ{�Hٻ�Q�=l��+}�|���؋�~Inj��ST�wo�n?8�n� ���t�7w�%\X�m��Y5������ޏ%I�ۑ����C�<�E{� i���[M�lj4�ԶҴ)�-ʽ��L�J�RS�I\O<�Z�4��Q^��Bq.S=�m^7�/=�G�1�xy�d�r���^G���Y�JF�������fe��M.Nо7���y����K7�o�x�#JmG��k�'���L#m$j�&3�5*f��O����.��pD��� A��IF�4I�i.U�'<���^G��n3yh��-/�V�Iښ��/n��Xg�Ni�x����tMk�3��>��\Q��gTs�Y�	�2�-��d׸���mR��R���|�������������hL������J2.bv�Hٍ�[��b�1��n�N����hx���!�S(ykw2(�yd��1�d���N��<O<hχ�9����c�2m�q)}��-	%��N�錆�Q����R�$������:|��Vs�~�"m�MS���X9{��Lc��^}"�ξ�!9��27l[i[��{}Fw��4�S��x}�Lӎ�E�Q�Es��U�ij�;�q��L '�����X��![q���ڣ��oa���q����������A�f���[��]��I�U�^�-�T�^���w_�����Y����v̫ɜd1�F�`d0�-/�5��'3�w��5�߅��u�Aĸ���Mp�nk�?P��r��(�O��t
W���:�+�!s�<a���^��~p�� �tz�f�}�ђ���A��K����Q���e�D��V��np��g�6��G�{�g���[�� �*���͕��_E�D[�)�n���$�_��YoϒAS �O���Nb'����\�$8߅���V��jU7z��D�
�*�Q�cDÀ�I�-n+�^v��`�t�B���U�a[���]�%l�L#�[���&��	�_s����
�(WNkK�g����j װJ(	�;�zO� ,�P1c�c�e�����|e�C���o�,���*�/�����'�(��K�D��/'�˚�����AL�z��%x^D	j��;�BF�u�ȉ���4�Hƣ�F3,hʋa�e��9Z2��0�lt��H��T�zmF��9��[�6�1�y��=�ƾe�ݢ����	�����i�n*��v~��z:�,�)eM�L��/Q�P~l ���f�Ż�g꽂�}���
���e��J5�YE�{3�{�$ɞRc�������ڣ���.6��d�^"����p���&�! �x�����OV5ߩ��t;�c���V8�	+)�2�b���>�Gk���F����PƼ�Uy)�9�%�n�p�q!y�����*Ә�8���hl$C�D����-P�B�?�j�P����^�Zu�'����@�u�L�A�Ǽ<��e�/c}�t.n��]�Hi���#�D(X *��k�8>g���4��	��;-���Ă���=��e��럧jj�"���^�{c^`���L�	 ƭ���m��h!�͔I!�S���,e��F�d�遙��$�v��+2���Y絏��m��
,/L��4NeaR�p8�3Ѥ��Jc!GEvu�p��
'58XA�I��+ ����1n�T�q�2�'8��S*ck�	��G��.���Q�$�O�\?�ƹ��~�-C��x���p�`�dI��+i
�P�����@	��u� ��>+K0�Ǝ��(d�R
L^�^9��t<�j�G�R|
ѥ�䫧]wYK�O�����vZ|5�$S��\�a� #�"0��*�L�s���+�ʱ))�yd�+��l@���#�z�S+�R���T��F��� ���|dGi�Z��Ѱ����eB��U%�ؒ�*�!98U,�kE&��TP�sD���ޢ���S�%+�009���u���ߛW�u\�'u��% B�S��]a��Ɖ��T7��s�w�[�ԙ��IS�����v�r��o>�]�
v@b���X_�V1�-g93�WἯGl�C���Q��ƞ`�m����ZE��/,��ݒI�$u�-R��r��U�s��2���B~j��D�PDN�ao���TN�Gu)�T1{{�E�j���(�Eς!�5#�F��^��p��~Jg;fiӅc����מ��!X2��p'=���!@6+��yT>��jW�j�w��4��>���>�Kg��4t���׭_З���Ъ�K��R���gM����(R���}�i35]c���~Ơ����J�:��j!�_���
n��}�a�,�9�ؘ/f9u}wк����dPZwu���&��٧�1��y��Ʃ=�Sf�m()��=Đ��}�$|�+Ww�w(�ӧp^�YE-Mz�O��CA^[����>a%ԧKƍ��;�Z8>I:Ӈ�uD=7���d��-�XG`�,J��T>ԝ�'���:c�ŢH�ЏmfK�`x�|{��ƻn 7MO�����O�iym���g����*�v�S��u4F�>�T�h2��q��N�=�#�w�X�ʤ�;��)�a{^��ɘ?NX:�����D@�$�1��R'J* ��1<�����V�yG�v �Fn{;
�����|$}Aٵ���=/ً�ϥ�j�u��,5S�R��"�f3k��)%�+vp��[/�G@���밽{\S.z�6G萛��*ˏ��ȈB+{|�
9����Y�>D_�"�
��Q��c�[�H0��99ٰM��� �LJ�̠���3�|�^��tg��*��2�]�W�����P�S�l�c� m!h���N�x��T�<�Ū��8ܚ�LCl��\�ރ���
��g�VN6�Qve_���[z����J{m^Q!p����^��}��bޘ�I���v�is�݀�vB.v�{�?E�uJA>�I˦8�� v�p��P�{]��oa�Zy���b+��ނV�����T�f�/m�}�:�[�F0��W���q�t귪��|������R��)�6ˇ��HZd�IM�J9F*]ͤ�L����&�D$z�܀��(�&�Z�� hK�R4:������ߥX)7�^�t��zT���UU,�f���`�{=��� �-)�������x�)���j�V�!�}����.���9�>�̆U����
��������ea�|�]�g̜��1o"�A��pIY�٠'�R��xۂ�%��C�*�Í�P�������:��� ��z-A��%��������?W���ݨ�_y z:_HH;��Qa������ze2X�
�Hq0�����H�Ų;0�I�Tt`V��Z�2���_
�Ei��f��.��0W`��~K[��#/�7D���:�"uJySߦĮ�a��p���DFi��l�k"~(>��;.�*wF�����nf�y$�Ug-�bJA vhR��Z��@���k5Qqe���ռ�ܻ׍���H�u�%�X
~Ԣf׶KGvJ ,���ߞ�	C�$�J%8�#�� ������~�����i�[�R_o�hn�b�aw�)6o�����_ݶ��s ڲ�?N3-����Dy���z�V�w{�IP]d��E\Q$0��;S��ru;�$Y�*���m��3�+�@20���l�f�d��f�I.� ���dGO�s�?_KO�	f)ݑ���Rq����'"��'Z���;t�sU ������ �m�\����kz����خy�]Z��(��?{��[|�̲Y@���g`�<�^l�'�u�qq	�D5I�	�n|,��׹���Ĕ#�[Ry�j�g��܂�/����֋�ۯ�Weq�{�x}̒1i�@�o�r�ԏ���fU����Ӊǥ���^����a�X��BUz��%�x�M�h6T�(ya	j��0z� �^�����T/��Զ�)\�U�Ě6�o�Vq.^�JM��̆��E��@%wt�2����"��a7�k�8����B�.4�9�����#(q��?��n��Ԣ{M�p���wýE.��o֪�2��ޘ�����.��kT�$����gc!�;{R통6^��������ɍ-~|��?��y��=y�����g���:�AaБ����k(v�!�Y?l�*����-K�O�Q��Py�on_9�ҹSg��G��_���㊙���P��_9��}@G��gǆ�Vj�q��?�;�T���@t*�х`ړ���b_��ã#�����O�)���ՀG�;ᶍn���$����\5��TRO%�M#ʮ�]�՟߯f �T{�U����� �^k��N��>@����8�9��oǓ%V;AÌaX��)� ^�ֽl�\�|�5�M*z��U��M����Bi�M��,��0%���k�r���h�o�6�}���2q��8� g	�S�~��ﬢD�sy�������1�ܭw��/�����ﺜ�!�,��t�¬T�+/��X���T�� �ԧ~M�`��ç4�]�X��Hn�Fvu���= "�<i�������JmŬ	g��8���������^�{��Ϲv�R6�as��ڄ�21i�ɵ�Zh��S����^	���Y�M��H��M�;1�cV?��&����Õ�+.G0�ކJN��m�$�FAHFUd���q�qI�U퉽(��v	��aW�b�l�{avS��&�m���^~
gK%����d������K猶�$r�Kzߎ�z4#3��E�7]�+W>�f�&���9�R��zҗ{���T���@�Pua�g��J��7�m�c����^;�I_������Ub�O�	PO�]�Q��Ir�����>
v���I����}A��B�Ի�$��=��XX�	4�O�G0����l�Q�ǴAۏ���\]� �����y.D���wZ'�X�1ULX�(á�V��Oz'���x���؅Z��;-�q��s2����6�-�N,ո�_+߭�p�S�3Y�(X�|��cz�s��2��B��ޚ4§��֭���7�Z�o��`���������*���"�q
�l�N�Y��Ϥ�����PG|u��0�&xh����m�)�3��Y���!��~8���s�{�8���\6���4�����X��2������2 g��	G���o�z�}<L1χˍe]?��@9��m�BPq��e󠯼?�lA�^�dn��r"\�[)��ia/�"�!7L�k�v���gNY�&.��,M�ڒ*?���^�s	��m\T�D�n7�Q2�
T"ɍ�K���C��S* b�B�p�,ǜPϡ��T�o�\��OM��ﾊ".���7O�����@������[��@R�x#��{�d5���FX�������q���M	��,�J����n�{ۮ�	��L�M�L����~d�[���^1�3f�ox?���&�x$5g�β�H�)q�l	g��W����C_c�2�~��G.랤��)[&��]����-(��5�$;�(�p���<�Ug�@D��ĺ�����87�O�d!��6����I�[�� D��0�+�\�Q�}y.�tZ�}���-9L̘"�K�b�>pIѣ�{O�=J�0W-���6����2��<U��~�a+$6���=�%��H���?�8�������f5� ۚ:�ΆI���q\���������CI`03���` ]��\Ў���*4��(J*������ŭ�G��_�ʖ)D"6�.�qR���^YQ���U:�ۂģ�����#R[-DUqU(P���Bv�h�t����O�oY|�?BᎤ�㼊�c΋���]r��w��e�	�w6�[摞{E���]�m�U�ʛ^\��y��86�CY��E

+��G���qN�\G�[ ����2�	�N��A�t��� ��`�s!�iK������'U2��\�W�6�$��T�f�i";�GMH�DV_�[P㽊�T���O�K�M� �65p_Vdl<Kv�#��{ܴx���Y�SF�%�Ox�{m��T��цr�"�D�v���|�#���$O���2��W���NSY��z�M�I|��B�f�}\-��VH�-tD��뱠ܣ
��{�E?����>d�&F���|�9�GT���3_e[�[
?��B�����xp�V7����^O*����\_�]�]s���̒��#�s]�?�Mn�������.���?!�愱l��|�����$c�!b��*JCz��[�����d�C`�
VV
�͗ˀo���?����1=�Sֲ��2'�_�Ӻɽ�������Ve��� ������8|�2����7��O�.����E��_�H��(
B�)�g���v�/�4�J�x`���_M����j��ۮD�F�g�f�1�s/���hc(b��m��ao�����t�x��׳����L"����G�UR�#'^ ѧ�X�n&pK�/C~���O���07å|gOY�"
�q�� `���y�}5D4�o��
:q��8�i3�ic�Y�[*c���`לm� %wV��j:�����J!k��)D	H�����`N&j��c��!�^�,�� �Q_�rP����\
�����ڷ8�` v�z#��`�5�	�tY�:%5Z+�h;����˃n���K�q��.v�`/��hDYN�ėf8읬�h3Zf	�?�-�����I���	O��� ����N�q;�+�L���k=���Ha��i���
|(Օ[�-\�$2nD�A��$4�(�~�RoD���?i���a����m���qy��\N�
ֲ.���fbɟ/$(�Gh��~�y}��HūȓB &�����⿁��H)����O�O��(x�,5��1�!�[o�g�o�l�
�S
�TY_ZSP�ڊk?pZ3��N>�(��Ea[�A�-X4�)�	��<�%���ť�X�6ŶcG�~zr@258T�,����\n1NOH7�v,0.E1��.���=�'��١�Cp�Y�ᙣN�_��]��T�Q��m���4�}/c#4�B��P��V��l����dޫZ���4���7�����ak �f����!-�+6��g�l�̏�&r�1����"�@��,�1B�8j��3;�{��"��0�:X�0�i�ýyH:�+�+,t����,��|gf��H��S����x;�_~��*�ư|&w�����QH�Ӆ��g�l�$PA�/ps�p|z��
̄>XuI~|����)'M$	W��v
�n�i�(���$�>wA������N�-@
�׾_�m���ǓB�3E�:j�R����������
�h77���8� ��uMf�Z�[L<Ր,9pG��L�p�dE�8�!n�H������hIl�L+��av~V�� �%s�}g�ʾ#ڀ�+/W�!J �X� ��۔7�"�/)��G׺8Zt���#u�phJ�ע(P*�H���۬ER���9�&�2k���Ik��e�R��m��ߘ��ޯ�Ȅ/8�LzQ(��B��"�w'&K}u�|���ܕ�7�\Uo�_Rjr0o��NOA�n�J{s��q��S�8���t��=w�I��<���5���y1q�C���9�V��ξh��آ=�I�5F���k��:4���,`i:��������G�^�������p���#xg�xX1>c/H������r/���Bӄ��f#lgsY؛�F���l��V�+���<���Ql��E�z�uL1��R��׆Պ��!��V�Q�j�/Z�3n�԰FR�I���M�/�r�":�p*�R�AN�D��� ���`��Ա�Nk��4��E���W������T�b��S���´�g�3l�/���꘏�0��P�鼔�@%�;�/����	8�ʈ���u/���`觯A����,�-��褖1�fĬ�{�n��[��%�%���}��weh�=��B|��~k���a-��p�PxO�M�P"5 r�
G�t0k �Ǐ[]������c�4���n���W�i0�����i�}0�d�0�L�R��tҞ�U*ܹ���*<��K����c���@���g(I[;j�u4�����dX��G�,�xj&8j�K)Hܯ>(��G;��ló��Y�Jl��h.Fgk�P�Tm�]��3�nZu7�jU��?t��[|ʆh���FI!B�IFd�J���Ӌ7�D-��k��9Ң���<�oq��z/,sL.Wq�%�G��&��O��7�p��*n�J�����������{ζ~z��p��?����������jw��AR?�X�RJ ��� �a$2�������<�T5
�@��=���RT���^��Аx���!��(gef�$�~mBO���0���y�u�y@�ŕp~�vL�	�����D?��*a����QE���s>��Ђ��[�)A������8Lc}}��@m��˫�Wr���b3�Lq�4��
��_F>^ȧnhBJ;As��Г��7(Zfm�^
�����#������  �i���������*��k�)�G�p�ShPt��w�l�!��7�Nx�W{���~!�jZ%���ڡ=��>����\IM�o��8��,=G�.��T�� @Ez��pV$��� �l㐮O�{�=�B1��C�kb�a���a���/�ىR���WF���I��\|֨%
�\��ۥx���b
�׷�(����6`n�*���\�/�c���;�s�zJ�Ƈb��JZD!��r��3�+绰���Sc�bژ���������|9}2��n�S�0�b�^���6�K�O�L�])�x�En�yr(�&O���2e�-�J���F���Q��0� �X[f���&�%YnD�m��|Q'G����]q�������$ɝ�����F�����ҍ
����Xp�� SE�ʷC�	G�o�d�NbUT�?֞���n��Up@�,���AD�����_����4�2ѧE��º�]	��\�jr84r�{L��Kӄ2��Όv�4.�HJ��Y��"��KV^������P��C�5qN��� ��pY�Pj��LK�;��`:\�Cb�EIJN���N���[d�~�b˗LL]W�`��(�
D��q)�����Q�$����ទ���JM�H�B���*�ϲ}׌}�g��S*0 wf��p��ҫj��#B�Wء\�B�G�-�u
�.8���/I�v����y�+�;E.5~=�uքh��l����
�p�Ln���!\�����z	�{8Ĵ%I�HZv�Q�5��c�|��#�:���e�w��:�#�
�T-Bc7O�4S�̕x���s��"hʸ��N��v/��χXqT���9��,ާc]��@���[�
�����)�'��܈#d��W�{+�R�}�mEh
	����ࢸ��e���O�>�f��ID���vm�l�˜8K�PJ�2g�NUg�#Xp�q�,�6Z�?}��
z�_��e��l-^�u��û�#�o�ƹ9n�Z/� n�R���I� !��zn)��=}�����aY��/�א��t�g����\��Mic��m�}i:�R�o��YG��I��H��e���Pk�bA�Ԛ³�TEYd�����ۘ�<_1�K���,E� -Vn9H�t���Nʫ�������$C�r��pI=R��3�J0+G1�^���F�-�1�X7�����yg�XID�g��<cG@�rpٹؔNձZTҎ]d³����u#��_�Z�h�;�xO'������Y��kv&��h��v��tno�E-�"�6���8����7�.���$]+ C� 9�3 ��l��hv���Qf|�zp3o/��l	��%����~k�٧���/X��H_I��:�D���z�̯������M��REg{FH���
�����& )r���$0�P�◾@�@�5��4ag�h� �:u"��Z}ʣ{9��) �ݍ�Xs׎��Ƒ�8"��i���j���\Ay1嘖􇥚(b=L��ה�	tubN����]ogx:��S������"��ڶY�y�����,�YĭڿB��3yݴ�syq"\���z�B�V������$_�d{w��{¿c�nE�5�˃h��%.\�\��1ipt�+q���s�O�7�Em/ɣ��W�lERK�FىS�'����<�H��mi�+�j���x���V�V/���3Ǝ�,��i���v��8����Dl��@��6[�^c[�z�|�w�<βC�6y�M�I�Nd���s{��!zHl ��|^��U���O�Skm�%hT��37�/I��ҕ����jϲ|�6�U��Jj���HR=b��Srj�"[!��]���(!�UI�C_�
]®��*��0���m��za�;�ë�"*M����n5�L�D��t�ց�/wC�ް�,�2�A77��/]V�w��i����'-���;qƾ� ����Z2z�:J�����foE�[;�X<�S��g V#��{à�a��3|3�=g�X}�lBg9�-1�G¤�>v��:��b��SQ��;����%���˩���A��ھ�.*�4��e�% a^��l��ge[U���ڈ�S/��t�iA���^�}]Z�1�X�g����F���p-@x�\/��|�����w��h�����?nJ�t�2Kzb���t��@�W�ߺ �O�Bm���煰�#���u��u|��>PXa�Z�='����P��^�"���������� "w吏O�������X�R �f�g�˹||��)e^�6�_�:��7sP��j����,w4�?�Z=Kɨt{u߾�ٶ��|Y#GYf�e����վ���}k}U��*	k�ִ5a\Ǽ�0�N�*���sⱺcooI�'_mQ`;xt��weK����J3�"�&}Ux<wS	C!����g�H��X�U���h�M��+�'oń�%8���ȡj� 7[��- n	�(�c�Z�i���Ӯf��]DL�/c�����F$����0x�l����3�{!��YJz�R�� ���N2D�5��s�aj=d��/)&4V�������F���l����'�C�7c��BO�ќ�>�a��Zg9���nG��?0�,�pP��?���� ���)�В��m1���@֓��v�{�s��]X/��
�?n��V"5�1�AgHUM<Ƶ��>}y�=$�$�_İ���%��dN)͔�mT�ӑ�?�R�j�CF��zO�2�|~��KL�dR:��[���JC% �B��@�M�}>��QxIS�<Jw�@T�h�����w�Z ;zf!qSMgּ{���U����N��x}���s�%�����9&?F������_���ٚ�ƟM�c�o�> C:W+��������'NqMdx}�?� Ƴn���ֽ���^A��:n����}��*;u7N�֗��e�3d��`���m�2��D�f��l�E)q�����"}rs"�P����s�.$�`�3�uq�#v�T� ���锕�1N�#Rs_i:H1j�E����2��pwg�f�����{�5r�4����|]W|� ����BCW9QǶx�<����9������4�������u��(n���fUqt� -]l��=8'*b|�cj��SE/�����Ґ�?�w��I�4Ŋ��(�L��)�~��p�+c�Ӏ@~�,{�LYG1."f�Sٷ�І`@�`.-[�����Â�z�Ç����`��ddf�7���;�;�����)������X M��ֺD�����������B���`� C�:E�$�҄�
��9��\q��#��Țk_74*bj��\����I9$m���`p�c�{uv#�>C��:y�i����h~/�E��\r�	���@��l�^�h���	����jf�#��ɡy �e�o�g��-#&p�%��C��J{��Za���o�+��C%մ�@\����!�L�w��$�d���݀���É��Ls�KT��)
���H�܍J�#��5Kv�'���E5p�hn1�z�2_�+�o3���Z�W5��b�;��g�"�u�/�O���P��ɿ�������R-~9���=˚��q��s��&=SNY�X��� �l�2x��#h����R�����3p�:F�Z]xN�"`�H�C�����mZMA���n���i�[ƘX�+_\}����8��#�4���;�L�܋�F�~��{y�;��|�� �H*��nt�(�2�:4�OY�L�L���ӄ�%f9�Jf�>P`��u�
Q��5��;`���Y}i�ƓږX�8F���p4���B�?�x�o�/%��&�y-	���*[i*qZs�aӕ���0��A�R�7�[�^����pE���\�&���1��kær{T���%�e�ٳ����Z��65�fL���#\�q�a��㸭�u�������
�l<��`���u;���bz&F���P�
w3 �h���*��	�<;����Y�F dS-dd���;&���'�9?e>�'�;���綗 P.&0��n&Jvv�zm7+cf�W��j��F'�!����Ŭ��)��A��^&�5k����E���Dt��D�TgP�Дe+8��b�����HvJ�~+���xP@���ۍ����j���%���6@�7�+���*�
��IZA�7_�Ќ���2����h�x��@�V�x�uu��S��n� ��l7�����R0�`:������ry�*sł�5Γ�9�xè��eM�?���0̽�!���~���:i�±�����ǹ)Qe�쾒iJ,K��J��E�9G�_���|E�r3I`	c?�%���E+^V�GWz�	eQ���VVe�I���ԑ̢��=Cu?`D��/ކP�9<����r�u S��t&��f�(l����pf)ʟ;�w�J,S�}j\Z��M
e�t��De�S:3sCbn+�Ks+=lQV�M�L�3��Y�
c��8��:r+�e�ڑD�HWgE��G�ˠ=O�/����L$Cv�DԗC&�sSN/�Ay�p:�D���Sre_6��i>��[3�e���͵Y�O���`���C:~Hk��L�X�b6��� ,���Z��	��(���9ٻ	S�TS�Ka�K%���p��Y��˥�n$�.~��ֵ��9B��'�W/�8"*�m��%-/�7��Iqn3�힆u�a9AqZ�^�:K�?�b�P���� �H�ؚE�A���[Yl�B�����"C�����tRW���QԿ�i�k�B�l%�yfS���V����-ct���W�I!ef�P���jč��L|qw�H�C���s�z����5���GIM��?Z�YS�� |�˥���N@4�c#"��p`�����1����:���F��V�'Ӟ�,��P'�wݛï#�O�I/(���%_V�w�_�s|�k���b�BT����BkG��{O7
H�������vV\[1N�����2WƟ�-�*���j��@����P�2-+�mq��ϵK
-_�玅\���(�_��%,U��UL������i^��>�)
r��2�0�PQ:.�4b*6�wuJ��!�i��̝/K܇�C<C��>og���f�wC����$KV矌����=�#���)x��f��3&5�@����p�c-Z�x���h=��G�@��+U�WǠżV��IIx-���.e�����H/�6ӊёG�1|C��-��T�����U�V:E����Q��S��v���6g�̈́H�l�Ulͼ�pT�r�e~�h�*���W7���#su\!^�r�BN-K���Z�w�0s�~�i,�R_��u�|�� #zO�5!r��dU�'`K��M��"��dM0I9��Z�Q�-f���!��B��k�q��N.�7G�°�����$��ܩ��������.�:��+��l=�1Y:ƽTj���_S��-t 94q�5*G'�4T"nZ�*��h��Ƴ���$���@�Л;?��i�s��=!t<�}�5���eG8Y���~n����eQX7�����OϨ"y5 ZN�PD/�pz��ػ�'���J�mٰ)y��Q��7�L ���o#����	D�����5��s�M�"I�^[$1�z�@���j�F;�8��������&f�O/�H#m��!e��`:�y�Y"E�>�0�����O�dE��j	r�o|T"b<u0ח�뽭$$�&�G�pFJ���n(�\~$��#r����&�"�v!˭PoJ�u�v����Ǒ�GZr�(�P
�'2�7�ɥ�H�͑g�2Zv' ㇃O����P٫�W^^�@�,�m���aF��/��It��v���kr֬^O�^!]F�$C,j��~=�6m��rOL��h�E��"p��,Ъ��DC�E�,�Yɒ䃐�UkW�}݊�]y�W��܌JH�������ٶ��M�^�aߖ����p�M��L�r�>Y�����y�͌�R������zp}���@��d➼Ȇh���짗Vp��kW>Lٽ�L��&��fM�뱅߬57�0N�mN���������$mm���CL �7ܽ���Y���ˑ����|�㮼�?���$G��呀��|�"�;�W|O���J���+��>����&&�{m�v��+^:&9WvP'�K
���!�J)��&F����	XpE��>g����� ���ת �{^%�*�n�A"��8���2$6E�MDdCFU�f����"�����.�e�i�tTs������WMO�JY����CE�K�[�!P��e�Q�ӗn� �>�K	b(۱��;0�V}vWT;��|�Bε��TC��k0�=*&�}���X�2N󰷅����l�w"���+ȴޚ��x��_p�ʪ�\g�o�7����������?���z� p��=����v���'���0~V��rB]ZU/dJ�/1��|n2�`�d��b!�Fk|�3S{�nl�E6�%n�O��H�S&�9vٮw�b�,�){�X�z.�h�����EiҺ�A��Th% �!�B��i�D�m�[.��#�Q�)�C
"��I#���Z^~\�e����K�C�!�T��&QY����3�9�6et����ՠW�Yj�! #�n(K�2[t���5W:�,N ;��A�2��<���
E��6�R_�11օQ�l�oh�����$��@��A���E�Du�ΚSJ�Pi��m���-�<�7�#�ť���|<#�8Jw�EĬI�(�B���� �/�L����S:ۚ*1=fqG�U��n���@8j�+�≟	�2k����݌��Tw�%o�e���D��E���8$[��C�f$���-3���l�+I�x_
eCN������a�d��#]Z��O�����M�O_2����X�v��[i 9&TZ+��2��cFUEC��J���Kk�xIo
�a�R$G�9��;��#�G4ZR*����S5���M@��AV���ɓ�H������4V#_u��]��>t�Zw����IZ�Ԛ�<&��2��E�S%�<��,v䀀�0�\��W�)��1�.�[We�p)�����?u@vDP��S��Ĕ�[��H��|�}9r+A�ܿU�.�k�3�"�uu�d}9p�c�A�Z$=�Ρ�H��Z`��ϊ;�z���.����?:�ŋ&tO�
ƣf��G�^�V�~@Ϙ��L�=�aR?�*y^-G}�Dէ�M[��/.��sW!�������
����{EF�KhB������Λ�43�O���S	�N�{�m1�R�;l�S�Ԫ|�\����4��'w�]KV��0oG�������� ���{��J�A��H6�1%z�N7���E�f������Ӻ�w�����QEG���u������s�2�tk�4�Z������.A�j����oоH�z$�]���}9�<�b�~�q4p�Ew����sks����x�9�#^M&J-�u�[�@}]��He���`Z��"%ޣ�$�w���t�R�$�{n��.L'L~����n�ś��_�4���δ�������3C�e�a��>��Xp!��qЕ�Ԉ� ������	��; %ֶv�NPs]��`��3��k���I9lH���HO�^0���eYy��u	���))N>��L���L���Z��!���^_�M�����ac���M�o�7��'�4�B���J��a8¹�-�Bi<���d����_XW�H�C�tC��T��}sȹ|.�9��.���	fp�<�R��(?X��W����/$j��d�3d���vg|���e¿�;PxΖi��wk���4�{�4��w
U���dަ�AFS?��C<�m��6@ptQ�U��Z��}��}U��t��"�-47��:~
��63;C��t���$�۫������Q0��#�T��`���LHz��'��^��I���+�^k�����b<��4q��v�$r�Eg��t�^4�� ��N�B<�b@�{AQ:?�o�����;�{���Qaf|p:�YMV(��D	訅�&R9,4˳�r�%�OʣZ�ၩ�p���K�Tr��W���\��׸��v�xtVvҧU;3����N���dC��!2 wl2�:TU��B�V"'�Y����wD�l�>AMHI� ��p��_x��a�Ѷ�;BV���)D1r�iZo���"P����>W�Gƀ�1���ds4ow��G�yET���Cq������c9^-�m��ep�����; ��c������%
U%�.�p�5U�Gu�⹺��]�>$G�Ww����3� �PP��� "1.s��X�00��M����ț�u'��_��̢e���[���O#y�2���^�K[L�P���!2~�rX�+m�-̮��}�7f҄Vu��}����%�b������	�k���߾�0����9j�*A��a�ݷB�% {?J��$ʊV|�Y��)��O��MxA�R�_��2����\��Vn��s���-Q�g锩l���WO�&U�T�g���R�ah�����O�Do�[\�v[�ܺ���!?ɑ��F�c`@��Λ�&�>s4��KQB�C�W�h�`�oC93+q�A{9u��N�1w���m�&r�Y�B�=�g�N���E��!Y�@�ѐ<�/T����	�����Fܹ��j��߹�{	AE�t;Ӂ?}V+��.���
!�1�~~�/H9���_E�j�zs�:���J���!��BI��2�v��þd��05�w1g���^e���kil_ej��9��n�!�L����fmz5�G��l��c����(f�0�Mp���퐲�S�N�-6�}���_h�Ū�g?�Q�+u��]͟Ԅ�Wߜ�I���nꪆs�^���}]�8H��z(��t`5���:���:_s���4�ʦu�}^|��T��Ag��H����D���~	�#A��:m��������at�A�he�G�#B�^�\I�*�o>ӷUUB����ņ�	� .m��o@7(tF��h����V�	�ܘ$uۍ8f�ob���OM�9Au4(:��Y.�Aٔ21UΣ�aQy~�v��2W�#j�����6_���p���O6J��VΠ?!���������I�*K2�8�����?�r��"Kӻ"��]�n�<d��."�Sĉ���
�H$O��<�N��z��_o�J<�{�k|�S6VSq��7�@��ɣ���EH�^o�C�H��!c��W���z^�����/��򚕤�k�W� ��z�n����l���z�2��5U�|��_���)Q�R�o��f���!d�n�K�Fs��d!���o^��d� ��y�/��T!����WzI!���(,x u{������
C��U%�Cݫ*�d�]�a|m�ɋpY@�C�W�S�
�Z�������e�ʥc%5̑� �G�����D��m�7 8w+�;�۱���>� skQ�FA`Ϭ/�N0�qՙ)�˜�	U�;�Y��ɑ�u�B�R�U*M�
-�r�$c�J�{d^����ՠ�1�rR����|���7�Ԍ�x���]���L���	��R��׽�����>e��7,Ė���|/~z�Q1Q�.0!:���i��͢ɛ�̓sY���>��.O�����۟����ģ ��w�o��	.Χ����d�ouE#�w&�[I�$$�UM����ڨ�T} �e�Rɀ���[��'�t�s�5�2���4f�{�R�������ݦ��2�gmH��xP�ҼK�Xk�7_��3� �
��"5�T���D���R;�[[�/͵|#o��-v������D��C�Z�]2e�bP!8Nv"�Yi�A�,C	��ccK{���|t��
�$ɍL=��,0��f�]� ��b> ���4��k7��=�)ݍD�c�f��O�о^5M=�2OX��RH>�d���;�&9�2����|�i��<�neJ��9���Z"�f���O�¦�B�H�`߁��,o�������k��.G��9x�f� V�kU��x�{7]���ȕDp�P�8ٙ�|��Z��,���5�V��T>��F�n�z��st�5("��'���CA1,�b93�����@G��p��˖��D�1/z��}IsQ��a�	�f�U��	,�t߮��)a̶���Va�Y-$��N5��8~JNT�2��K	>e9l�wJ�̞/Egc�pr��z� ��"�..6��!����m�2	O ψSo�t�L\4㐢���{�C�.<�팴��)��x��2���>�	̦������5�4s���SQ2Q�����Ir
��4���\]f(�o޽�$�Hp߲��"��0���J�gc39�[��$������/�M���G)v��T�țA�=��L�Y��+b�v\��{��L�'�I����h��_��+rM��;���&��T��,��*��5���PBl?�&���|o:������I�����M���OC3Uɶ�i|�R��YqңI��H��i{��*m_��D��π	��<l�P��DG����/��Z��}�WH�.��ۂl�4�V�jqCd��~���2o������#�	h���.�>F�|w0EX�&֘�s �'鱍}Ђ4.�	���'�<�YY����c�?�ӕ���Du��c%���d�5�PQ}l8�_8��$8��n�"1*���?@�L���jʁ~A8�Ē��>sS�ȵ����:���D�k�9�]h���x��w���_A{��F���:/�]�=5�u]hM��SM9�0\��G��^޺~�ZY���Z�0�|ojL��l~��y�~mӓl��u�(�< �܍����1��g�_�]k�WU��%T�:���K��n��a�k{�y���G��ە9�A�&3b_ƶVQs�T������� �Q%<��o��m�C*� �>��\6�l�����-��3ER����u�t`�Yh�e��8R��(�Rw<&#����fQ�p��>��8ߙ~��IY�B��[Ľ뺲k�j6q�=mfl�Q��Dg��*���N��t�%��g��~\�q8YC�I���R	������ji�LC�n�=8�h�7?d�b����+�P�={�#3�RH�s`MZ�IN���0r&+R��K�ȏ�h��Ro/j+��+�x���EBF���,�uT�X|���!��uI[Ņ��ݣ�U��N����B�52�H ]������^���Ȳ���
��o�5�3�����)�4c�A�*�a*�*�+2=�2`S��/O��tuK7������;79��A�A�_���;Z!�,�<�I�]i�������l��K�ז2���p�6�pՄ�Ӕ�ݦ��.2̱?�N�y������ �w�=H����Cq��R G������j	7��>���H!����X:�YQ���?	`��VbyRF�X%y��Ԫ�
H<�c�Cj�cW��5�N,�g�ޥQJ�E3(fB#��m�y�%q�J��E:�{1����ҋ��mA�}Ll�+<^�<Fi�������ǏL���!W+�	�4��TAK�s�R��:�0l�k�~@B�0��+���r���*���υb�r�4u8�M��!-� �����%���V9v7����Ns�@>N*���?�&p���f�QBqGzP]j�JJ�� �?����� �ؗr�@�$XdglSTvFS(0>t7C�%�JY�Ɇ��z"^���@�)��*�Jw.o�`�@vrba��`��и"x�� PE�+�(���[��G&����?�f;	B�x�������ڔ>_�U�Mg�����>��by�L�~ʹ��ަ?W��@>�2h��a��O� "3� .�J)�|Ls��=!��K�80�������0��L��zR �jj�a���W�t�F����j�p��KFuW�ɍ W�1���:�[��>k�BU����6�*��'�!![�I�9u|�a�[���͹	�`�� �Ce��ڔ@���
�8٢�����G��9*�(@��QKHk�)!�?m@]���-@@�L(��MH$S��B̐�dB@�hP�d'Xg���o:,���F�# @�C���RX���m�)w�hb�H��\��kЋ��qt�Z�l
�e����YB:h�D�����z�	���έ��ukk���f�b|�+�T;H7-�S�*��>` �C�
���}���� y**������S/{�bs`aL4�ވ�#�:`��(a`�X&����}���|�؎�ӏ�'�#�5��@���2�(+�(~Ǒ+o�o9�ßW���HK��b'4�-F�^�_,�2@�"����k2?6��'8�=�
sϩ�cG���+���4�\t9��N��6����l_o���o�������o�Bo�geq���Jx<��']���g�.�ر�e��>R���ri��f1O����=M�������ĥ1^W�vZ봯����9�/��~<�+�C:��t���􄦙�����>�b��;��'�a�bq���s���W��q�k�z���W�����#�7,C��]K�
d���S����9�Bi/١��
Y�����5~��:�W������-�W�P����.tD��&	����m<�=���~^C2�&{���B��#B��'|Β
�"�f1�<A��u
@X�d��=Ceߪ�wrT����eJ���b۵�?�a'�\q�~� �����ad���kps9{aW���7����n����Y��,�ƿD�e������rJ���{�FN �4?���o+f��4:C�&i>>՛��fp�[�1G��#j�Y��V�c��s�`��يEY�ie���Q:!�l��>4�r5�⑮��.����������j���5[��Y�:�*�,B������V�u������r�&�5�+��NZk�H�I�q�fUDt��4��Zu@M�E~�Ђ�x?���C<(���6�\Q{eW�S}/w��Xz�'�Z�Co�.	��ۨrq�X�A���&�Zo~�}��"+�q2	����'������m㘽�v1[���)�}������7u���l&'�Iý,�E��K�}�#�]�+�=u���^ǋ��c˥����X�6��#�|�& qr�J{�3Jb������9>]x��9;w���
%��~
��Iћh�r�L��c�x�� J
�˩�<��EE�m~GOk�U�Xv�Y~�i行A4�5"Cӫ�J(.�#um��nn�.o
���g���!��k���>_�Ť��3��澁�J����:M{!��6� �FY��n��߃2#q�P!]�p���bF���.��NKڡrĉ��KiR�u�=�w��p�R���IF�HIv]۹!�
�-`�?;_+�ĐJ�5O=�m�g�%�ٰ���8wu�p]���&CD�	4�.���e�ՙB#���أ��C�l5=yFa�s0��ڦ~S�6A��������%B�$��,��v�>t�����|t��"F�ԛ�G���;I�@���	�\��;���s��ڀ���L
dd�ږ]KP�;�RG��3.z1�2�� I�@	+�hi ���M��`h3�z,�0� Z`�D�'��6���t�!h�xFG��~9#��1�����:�}�"���0��-B����y36bX/+O e�/ )�Q��E�[�����aɝ�e+�2�);��YRD��:����.<���'1�+mu7�����k�ƥg� xx��
YZ��(���fKΣ<E�4�N�m���g�u�S)"gH�9�:���X!q�?f�ׇ�x�ı�a�:�������D�~4��P�b�����2D'A���3����Hˍh�8x�2�����W�;tB����o��*=s�C)B�k��1 �[K���'?�����O��D�;HOU�I:tR2�NL^L��0��h�!��9B�� ��{�� �]���82��to��ѫKt�/˽μ�
8k;-�� 7�X�D�8Į#�Ï,<���̄�Ԛ��`��|7���tIxgOx���` ['uy�M�&����`Y�N�RU���I�F��2/�6T�
��@�%\�����L�����tg��݌S�7���sz]�d���T�#��M��y� ��Z��C�c<�~|��U".U6k #7�<䧅�vǹ8G�*�W�̭��b.��0����$D�G���T�9�X������i�2�P��\pZ|&�BVv0�^�j`?��0�:�.=E�ʡ�jo�O�k�n~�g� ��~�l�q�m�{q�;:�M�0">y��"��Ek�k�g���,dYs[��Y�|�#�&�%�c'���4PC*�q�������  Pv���H�qfc�ݒ�Gp�w,b���{��g����@�:F���!�$P>:��<�`	�������w���	F�$��l��D�?z�@�k�χxo�����PX�M��:��d�5�$VI�"� s2r��θz}���!ˬ��1�jR�k�
�&ܒ�.��̴�_�>`_�Z�!�9h�KEM��h��;>�R�5^��ާ�߷�r�o�q�T,�B����~������۽؋= 4Ol�1�n���)F��}T" ���m�\�<�;�T���7v��At�ڡ<��d��"���l.�	?���5G	hr>="<�_o`[=(�-�9G/$�A��ǖ��~��5R��d��t�rl��������wCa�w�g$���D(����̈́���b��ս9�����L�	��_�D����n������0�,"���j�}�X�{U��]Zd��:?F�G�n�$�ھ�6��FGw,���V�����;��L�5i�#���6�I~�)���6γ��b��B�(�!>��8ͻD0��5�)n!��;�U�M#�$�r|<�8+yt �b��Ҧ0`kCv+��MGԐub�K�XѥQ_��`��]J���i�oaN9`߅.6�~��M�%=S�'�d�Z6�M���j��?�=L�|�n$�>u��i�#��H �a{�<��V��FW�)-�-�����缍F�$���7��y���D�2O�N��5O1fȲ�Q����Z����q+:�O��́����S��q�'y9��%+�M�l���j+m��~�m=�ِ�R�@B]S�T��-"�����R��%�$���+��umL(���ENSS-�g[bbCg��ث�W��.��V_��m�>����:�MWJ���9��5.�H�#�,�S��;�hz�bXSV�@��k�A��z��2��=%�ԣ)z����-)ׯ9ߑ[��K�P)��^�_���Sr7��Ɣ>l�LGu9��E��וMA�i�y ��	&ݢ�-���8�M�/����<�����C���͋j�㤽<�oC���!k4�EQ.r�)�,7Z�1��ݦ��k;ݖY){=���S#�S"�:A�R-�Q0�p~������`�g�--?8��1y5����!d~�$���V;O����$=B�E�dŰbR�Ҝ) ��a��J���ǯnqr�u�Ȼ}�f�W�� �	�P-�g���N\IP;��Q�,@��4�>����8�:Z��/jF%M�!�՜mи�� �ʣ �������bp��g���znnl�2�W�4�"�{)'�N�2��tj� �GU*Aь1n�硃��Fn��[�a�]�ɗ[}:�CG+L{�4-�'ޔ���=��p�<�����w� �j��[�Z֥���L���v����l�w�g���ki��#t��L���n�����'CP�*�J] ��<�,��k|�EP�)j��A�i*`S�ĕ����`։�k$Ht�1�L������f5��~����j�O���v�Qq3)�ʿ�7�Ճ���/��砠V_P�͌�.=(�]�F�&�o�@�N�;�WjE�ff�L���st�Ӏ~��eM϶ �����z���EM�3�4�CEbʀw1m ���Pi��O��|O�P;q��}��T���<n�+S�ϛ��؏֭��w�bԂ������8����ϊi�5;����	�u}Mu�Q�L���Դ�����"�s- e#�g!�	$�Qn��c1T�t2�9�1��_�c8s�x`�	����{�+J,��$��ȉTV��R�nh�*�d[� ���������K��/�^��}�����x���aPK�A��*�%]�)�VS��(�7�� \��͆�0���RD�;�0_7��Q���CU����6�9��S
�`ɻ�w�[tXLp��qNj����XD1v�D`Ƽ�ab=��B$�n6����%�l��9G�E}U�썷�ԟu'P� 	��0$��S��Q�L��#��;��p���
��� 4��x7	9�T?3��x�װ�gD[�Ҕgd�z�������w9���鴅�`������궥V��d�Y����	��xX�jXv���~ {���}ü
.�p+J���S��`kE9Iw'�Xkas���y@�G[�	��,���җZ���VGVW&�������h*�* �4��}�q���/E>�� �r8��53` �߂#�u`�>���Ae�LE_��N��QLU�p�tcĄ�����ɿ�j�G����3i�8A�b�������
!�V��7��'9,3}��(O^1Dٙ�{%!T�z��Xf�H0븡M�k@P����B�m�M������E�(�n`��D��-;PsN�X�N���hS�Z��\���K�)��E~�v���ĳ���n({�j+A-o�]4&���1�S�܎b�ؔb_���/��	�ʊ�h�z׮�׌ݰ-EaL�zn|t�Ib�Ñ�m>�H\�,�mWj\�)�^V�?��Aj��4Q�nvVY�Z�/Us;� ���pg�K�?ڬ�f�d�dJ�w��]^Lh����NR�����&E�L|���$�I��]�4r&t߹n`�c���I$�=���<Nq�v-�BS���#�q~����;�J��d���$Zm��xr�jY��Q��4��Y� �<R�5L��;P�IL��B�5�oG���=��~�&lkZZh@�@S��K�X����������&(r�w�
Q	���M�.�d�S�g�uR?
�3��y�&�\�
��� =wI��9͕�ܾ�o�d�����S��b��%3�7��&���2'D2 ���Y%�����p��{?�S��W ���/o�C�A���?Y���?ґݸqO��y�M1S{��M����>8�}�ߏ��f��i��˯�#؋�6�+�.�м񅾫_�*�2�w`����R+1���i����١{���I�5%Z��`�2��.u�+
W����]�ٽ���<������/X���I���_qs���s���/m�������2"�j>ӌ*<��M�����GN�QR��u�����#���ʉ$�_�C>�f��h\��q7�ʲ��(P�V�>2z=n�d����i��{Gn�M(�Z4D~���	��ک���T�:�`�g�����ێ6T�Sj�-x���Ʃ�C�����=�qW�#Um�W�������.��ؼ�Oå;`�e�Y�)�gԈZH�K��h%�͂�2��H��c�*$��b��
Dk�;�����W�$����ah?��� �;�X��WGi�7+B=�1),f�-�4����N����'��]�w��_#~�4�jp��1��������:D�z�������C<b������.�.�?܏4���˹�>>=�7�r�*���|���T�U<�p*Y�v��*Mh���*��e�4��"S��л<q�X����]|
:ڍ'��ņ��?H#���(�s���5n��0l�����S`��T�t�)l�����H�W�-}YV��G�6��W�!����{*���g��M��{���>х���D�9�xh&�瘵��=8˽ݓ�'�=���gd��)��|��b-Џm�Hݡ|\�_ȉB�z���@���Z�ߕW�TySE��x�4�q��8�
�(�z�Y�_�� _E�^�'�`I	�s=���-��V/4��(�Ǘ�T��DZ�u�疿�B��Z���ߚ<������a���#kT���ʽ�a7��C����θ���L��o�Й�,)�o��}�&��9�3��bL;0�x��
��"�%X�L�������=�'6e��9�/2C��Ǒ�Y\�1�`�����J��b��-#�Z2ּ��G������}�:��Te3v��v�6�����l`�gj��n�H�RHz����L8Bu�ժ��u��M>���F�j�-Q>V��X]))9�]�ϲf��(юq_{��{2�4tʮ.��j���5a��t��*EW�Hb�K'%Eh�A���@�@��fٴԻ��u�>�i sw���UHz�n]s�������a�a�V�Y�F-/-Ʃo�ǔ�>	�`�/dWh�����!nF��剑0|n&��v��Q�S�^��v(��Ӣi�+s�~���Y�3�����
ߕg3c|��2oa{��8�[�Ms`�<%��[�9z�a/�u��l7[��H�5$��EK����{@��;�1r�/�8�d}"\�F�
91�N�����O�
����6j�my��f�ڑEJ�:�(hg1C~�6�u�����Mש����ܮ�1��8����S}�n��t^U���i��
nX�:=�M�|Q�i�EwN�:���I?F�ۃ�O�ɐTo�j�]A����p�a��(3hE�<�g�E��d�Q(��_�>p��O^����v�u{}��n��Q��̆g����j�Q��\�~�G�p�p@D�P�m^��:�;OWv��&�fJ��}�#)�-��g]�F �-`��fs A,�1i%z�?�Ag� �m�0��xz	��-�C���<�����9�]E��gRm�:KW�a�1����Uy�Xh��ۉ�������$	�����+k���8�b��sԽ�*E1���0�/�a�;Em��53��z��� 
�Y6��
G'@J�՗�Zj LzPG��#�t���;�[8�9kJ2�&��S�hD��6��Kn:��yܔ���@~�al�5^���1!��x0�.V-�B����1	q���ycD��P̊dh��Ah��pu�b��Ԗ���˨:�ˇl�:uk��z�s�FmC�"(��1������.��C꒓�}�(:�3�2v~�`,����X��3H3^����T������<�ihbw��:�ߢ�d����[?��h�9&6��P��4���kÜ6b���9ΰ��F�	39���9�jo�*� ��`�i?��sz\��h
�"���������V���;ǻ���v�i�^�V��BI �(D%HB��c�Q�j� �~��-��ԕ�*Ɉ�k%�l}c�G݂�[_s�����7�(�Yn�j:��b��V�!U~��=Z����k�ȇ�;�=5��\=T�0��)ɕ1v��J�@T����^C��*(%��������k{���.-����N����!�z(�I�2�	F��tj�B(�(��q��#Ȏ0��r�X���"�c�����-��X��zJrz�hjU\t���A��J$5l	��u=ӳ¨zg�%��I�/'~Fj3�f�<.<����2*U|w��{<��D)�H�/j����_�& -�'tJ%X�pP�dX~\�͐�A�_r��uK�Nw�Y`�!�3�Ht=���E���]p���Av��i�o]��HJO*z��h2�$�dT�7�#0���Ⱦ�\Ae����(�8���}���Lfw�����Ǜ��h�� Қ��'%z"<�.ႝ�Qռ(2덯���ٞ�d���os>R�T"N�ƝCO����G�/<�J]��aZa����=E�4A�������ص����ҿb��{�.m~�����Nn�T�Ņ;�|!hnE:6��qqWc�;$�t<{���4�-��g/(�%d\��r��F;�Y������U�<�{2"��$h��Oy��Z諥v�ޕtS^���8.%��=i��pB��u���V��ƭu��J�-��]Tr�y��M�?��W?\?|�B#������>��I1�O(��"g(#�2�XP���^��F��U��)��3��-6�w.ذ�<`B�k����TpEan�Ԯ^�لu/.5�W���y�	��H��Y��IRQ�gfW�$��6꘭03]��c@��F<�*^�u��3x?8��j�@@{ə���|�h��:-�p����X�|���D�����������q�j��ܒ����@�A�M�y���Mل���2A��w��dXE���.X�y���;ev�-s�!|X{=���f���D��2���q&4��֒�1�����&[]�[E���g�|&)\
��Že�i�qeǝ���DM�e�.p�0-�X���Y ޞ<�����r��~i0���+E��ӑ�-D)�b6kn��õ:%e 1"���;�-��Ox(�o��f�Y�Xk��ή���t	Y��Ŭ�䢪�߼X�a��I$#��7m4�*i����f���s͗A�W~ o�"SmW�D�r�e�5������:?�9���v��~ve`+�h"�f_ϔ�D���WO�r['�P7��@��5�$&���"�uܾ	=�5��.�΀��4�k�r���%A���qn_��Zw�%�b'RZۨK�Р���Y�� �f��@m�\
&�$�cz�N�C��3���n�(����#r����&)4��8�ڷ�|	|\��o���������
� �[1٢����c8U�Y�b4h��U�f�.JX�p�p�	!�A! lX/��9�D��|L� `U�c�Y1$T���C��% I�Z:��%G�u� ��o��Q����c��pͲ�N���|KXPK����\X�Oh%WE�:O�H?�ط�z�Y�����">���D�,Y����C��.�OUU=e��Idʔ�
P��)�I@������n-L�m�&֚q� l��b��Ȃס�G	��p."��PE��BhC���r�������:f\Q��X9�gK���`_u��&����lБ)����nհ�
p|�A�]@���IW������7�z~:i��5�Ѳ���V���d�	�J�c��;}�P)Kdl ���FOɾ:��H%m� <�}�0����]#��Ia�����7�1��_5{+���'�<�h�QfZ�(*�K��#�g`=��Q9`!�4�5֭w{�nQ�Y`#Ep_l�"c|"k��8�c�T�w�B���]��y����%A��'�2.c��(��4:�<���n�CM����
��v�H�M�\� [9��g�Al�׷e!IP? ��ql���,�>��#"�@�")��Z�}+&�a<�:�%���\�}	c�������߹
�ax�`��!����s�A��9+��P�u��8b�S7��t�at(��p�)߁�~wJ�X�U�xa�R5e'��K�B'��Dhv���`������CD軙STc.�{+����'<��p=�ɼ�y����$>(��b�P�ġ��4��痧Q��6�@K�@�Ѭ�! ������u5)��J���`Zg<ٮt�?��G�cs2�$�h#[ߥ���(h��:N�/D4�lO�ޗ���j+��5Xa(�������[�E씰4�2��Ќmt#5����0���%�����X���)h�U�D֎������Kn7n"�|��+V�#�U���Q���pm��{�xʇ9,e��G�ٌ���[$?����af����������Bk���;u���n��_h��="n�<ՓCT~�Kkt�;�1�(�]�9Um�x�v;��^��10_�lx�����S�|X4B�^�v͞���X��_�����T{;`s®�k�C]x9o�⿸"����GE�=��N�'�ބ�~�H7+=�[E�7#x�a[N�����J����E��;�	r�%rg���H�p�Rk؋���b�N��-a����%�����J��n���f!>wD:zq��MfM5�h�!�h�AǮ���i�H��Ь�]�u٩���*�ɘn%c�2��>f���
GO�h��9�0�̨*�K�e���w��\n���,YS	E��h���� �|T"�$�.�G�<�]�������A�[7���ߝ����p�絭R���^:#a�0Takta���.)a�L���ʬx!>�	�g�_U?�*ވ�EO�N�� NQ�k4���?i⛭�^:��#S!� �+�'��tM��]>��ɖ��� �
�r�o��K��?vG�G�c��tjW�����|���p�W���C��f���c�&}� 1�ّ����K7E7��r�������x4 �����;"?������Ew\%��1�s���@����l��9Ă�r	o��$&�Ax|ڟi���&�灉����Q���Pm
 P*�Q���|i�r�_�u���lGOBH�&H���=A}������e՟���$_qҩ3�j(%�;�֤�|��J�Lo��l�Ѭ>����|���[}^~$��?��D'p�`#�vR��N�	��	P3�"�Y�+f\�eGu�|�0��{��!�RfD�q���a���v� �`D�[���qe�nP�m�k���.�A]&J��b��t�E;"��<#��$�s����`�8��PIZ�b5cm���R.H_��Tt4V�b�w��kR�c-/|Cu�L007�fj\r�5P��bl�{0ūym4
�#���ê차+Zk��N���s�\�|��5���-�"ھ���҇�ʼ�㍛����R�����+S|��tVE	��ju�(M&
`��U6
Es�_҉.D�T9��%�b�]�^�?8����bJ��l1�_��]a�n������P��^�#�6�w������1t���H!����'�TD#��o��R��n��w���b�V����oۚ[�Ėҗ`@�xdt��XI�:��n;Iq��x��'�o���>�Y���U��	_���5��������Ko&�`"�S��6�Nt��x`�y��R�BG�}�ګQ�~u��6\?0;��w�E6ɍT8kڜz� ����^�w��e����2� ��g�	;�ƿ�`��7����FV�
��x��qT����y  ]��p�-�K�0�-�'�0x�5�r�4�U�x����"�~�q��t���W�-��{8�,�Ϫ�80���S����];E �~<\��7�T;,nNg��}ʣV��-�r6�F�x+�����Edp^�� �}����5��a���Ij_Z���	R����*�;"�U�5hR�e�ԝ.p���gJ��n��e|1u��1U
�#v���B�/a.�j`�J�ApD�d�q��O�6bBt��BWwI:����h���4Z�&�`�=���>���H�R]{�j�k��������G6"�bl�{#����1(�%�{ǘ����A[/xD��8;�y�J�^��H�B�$�F>�{\$�	��= ���5ϥ��W><ow�$K�}-�b
WN3� �yA��$-�Ϗ~P!ނ�2�`�1z�cF ��V�R`|{I�3=�>�����}����3WQ��JK���`ȅ�0���u��ʯFk��J�s3̋[F���l唇06D~���Ѡ2x�N���P��wBo$�~%�j����ub��K>ƈ>��34�hE�}	���^dDwj�M�S���#<
��˭��5b�Z�]��R�\�e�~���ʟq�L���)wخ��iGvw7.-Lxȕv� ks��2��M@�܅ ��r	*�U�.D�<U.��3�V���j��k�ٍ$Pq-�F� ��S>Ϳ�j��	����A�o���
�]�N�c8e��,,��M�2���M�cx�E����� �t ��J��� .>�H!^���K�Ɠ���ӟۥ+2=X&��\���D�$TL#��3�"� z	�s��ǡdbo�����H'�-��eƟJ��3S�5����Q3��j���2(�����x.I����Ӿ���	)�n��C9	fovI�Q������.+�du����9
����d�)R�Q��#|�:S�"��l����V0�4�F��k垆a�D��#x��s�~Di��X+�Mo��Y�
�9q� �*j�p�J��x�ġS��h�7a�k�T�Q�bF���#N�A��`�	��K���Hz��J?T����J��-�������CӚU�82n�7=���Fq��}�����V?��7��<̽�#J�d�������A��b�Kc6�����pov
8��fG��i���gѩ),�l�{�ʥwz�u��$Z�t��|�]��4�ǩ4ōl�����tkhhO���2��
�z��@ڟ\�;��R���Y/r>Hο6d�l��sj�Ƅ��'�������J��A��A�k���˧t櫯K�c"&��s�fd%a�*m�=�\1v�A�`��E�ϻ�n�0eg���[�[�Lk�<7�"DP��3Bc�r�kOx���u���hx&s�v���Q�C�--}�]� �U��N��2;�\�z�ܐO��u�8>!����][���vU*(�K���4��@\�w����o���� U8쪂WMi95�G����Č�6����:
�� L�P��R��Ï��(�s"w�en�-�f��(kbz�ڢh�(-a<�b��J�uD *`�|����J�\� ���>��*�,��s��h\��j��ڻ�VT_�E�7�fJg#��𐘑ssPg�>�5I��k�M�JĎCwX���+d7�vM�R�>�A���:ګ��OR5U�2bh^���L������eW�&�Q�S�eN5[���)�bX�YBaj������1��f�c!ƙ���rez�} ��Ɨ]m��RPo��A�R�_~;��)I�/p�$vP:�{]��(��N����!!�\�X��A��[Y���0��0�����h���Έ�q@Uh�"l� �1N>�I�Yh�0�C�`�Q��xD����Pu|hk<r(��3�k�<`������8���N��}t��k�f;�gMz�ԏ{��y'�����֊�tZ�Kw_��('�#�h��n%\Gkʳ:�i#��?���s���Z915<��k�{~��pj^��|�p���Yi8��1��ϻ7J$�&0��Z��@���o��'l='�	K���Ȁm�@h��>�����g���������������V�}t�&@��Z����{Ń�F
^�0�"K�������u!���8���ow�����S�Xm�7��i��0e��d�_t�BHѸ-���8����-\+��o�0�
����d�`W��5H��đ�zy>= - ����N8��{6�������m�^���:\���a�m�G��N�$a箱�x��Ҵ�Ea�X��)b��ce��Ve�3Ä�Lk�׉K���{��m�n�<_-�Z)����C�b�\�A����vح��5d�[LƂ�='��%4�0+����ӑ*�2���"� ��v�8N�G�B:�s�����K>:%�z��1bǾ�[f��q��E�Z��}� �`T[F��K!D�'���w?F��J�w��0��*�UqLl�k`���X�A���3ÀmM6�f�#3)�c��}_'Ψ"X����pφH[��`�nf��K�8X�L���A}W��u֢�c9�[�H�ۿ�6Z�ak1��IP�pF���5��vx�xB���_<f	��7,���j�z��5��X�^(�J����}�=2�d1^�����g�M'/'��C�m��)y<�/C7u��Eç~R5��QF.0�`v{�id1��R�[R��u��(�{Z3�j3�rH7���%�+y�� ���.+�3��jT��)�����9����h�e���`�a�>a�o��
>����/��k�VuL��2υ`&���T|G��0D���}�����"�r!Iw0@�DM_Ն@$��J�[O�#Ǹ,
��L�����̘>O不�܄��Eh�~.���Z��l�����j���Fl��>D���؇���F�W�L��C��(n�1!GRU[ᶭ�}r^�`�Tn��MϺ�֓��#�30��ռ1�*2;�>4Y8�e�_�ǿ5���&$�Ry)��?N O>r�L�.�z?n���Zuj(�<��7CNM{�u�Bnv�b�t���Z����o��o3c�O�p��(�Z��#ӫ.Z3̛��u�'�����Sp��߆�T��a
�~Y�����?ҋ�������Y@P�Nai%pT��,���Ί��SI��͌��2FY(����ϭ	�!O�����?m��l0�� ��g�9����b[d����;��x��'×��ׄ����[h ��s��N��
ȁ���1Ce�A�^~N��WGZ��fŶX t]�U��ٺ������Ӓ{�E�Ye���Vfiz7&�2��ƘBCY���\�'W��QS�m�Y���j��'=H���LVAe��jX��?Q�rJ�i�7r8�ˤze\TZs[M��R|�A^:�����������K�i8 ޵���b�@q�/a_�P`ҷ�%����F:��[�"IA3F�l�Mb��X8q��j�3<Ȏ�wЩl��,�'�}�&J�d,Y�d|��c%^M��q�A����(�㯰���#*n�W�!��ܪ`�}_�/�%b��U�7�F��&�����D�����f����v���i:��n8�������`�'�(���vt���.wl�L����0�wY�Q��)ϛOI�Zٕ.��|�c#�u�9^?��Dm�P��{̒��({��"\ ���u)�<���i��9:�w�Q�}�*SaON���
��tš�/���h�!�t8����:N�<���sH$��7��t�X�{o��>���w]xSx ��=뉭#ín��7�М�m=!��]�H�͌J���!�@K=���6w~ӜX����nm�	�VP���#�8�7~��;��Ԩ'S��}|�>�\�Hk����
�@�F�A���>��SX$=���H�gT���6�敞���CL�l%�`�l��&E��x���'"c�%��=�d%,ySS���b�>z�l>"c�2��B?���c�ӏ�)y�`���M�Q@������F1�N����>Н�ٺ��,�l8|� +���7�Ȝ�v_��M%��)R��� d�,�*�Qo'���Z¨c��{�z��!�#^�,&qF�|��ؖ$6��ħ�Ў~d2��	��>�N��Yp�Z��i��&��>k���h]k��(oPl��oܡ���׎yŞ�>���?e�`�*�k�:�+nl�P�������)�=ֺ���o���n�a//!k+�V��zߎ ���`6�����Vl�~Db7;�3����%�1�8	#�#�n�m%/��>��;* OC�A,�<�L�������AQI��N��U�J��#m+�W_��߯��)6q�~o|�v��.������ӱy|䕳X�׉@Z����^��׸�(���b40���vK	�n[���oǀ�V�e�����)e�LHn�u}Ҭxzx%��;e!'�}^�@�M�{ (���)(u?%=���e�/���[׆���8]wZ�lp��������.e��k� �$�0��;���
�Lغ� �ׄ������w�_��e�b`T\W4|��d���`�G��0+�Xu�WD�j�8Q��V�;e�,,�Mz����߃Z����/B��EE�F:ѿ���,�����0��,K���%�9)"L4�_��5�d�_+�M�m�<^�-q�(�g���Y}
�n��GԖ#�:p�-a~�`��O�ĬX���t9�j��ÚK�,�Ζn���8��QRǘ���n1y��Fb��2�	��"Ȏӟ��?�V��ˌ�"�Nv㠚��4t���1W�>a�C�8�3��D���U������09��t�������]j$kb��>	��HTR`�G[���ˢ�DJ叧�b�w���A���l��(��]�u{����4��/��i.�T�9��7`�h��^��
��|�l�����6�E|J](�����غ�n=*KW-�H y-�c0w�V!s9�Gp/h�N�7N-'�aL�BKl�;]�v������)7_v���;!"y_܋�^I��X�R�ٌ9�)gܮcs�\/+j�5�9//p�)!%(��w���veƐ5�� .�B�l�@[c�qD%��+J�'������d!��J�ڐ��O�d����UhY�%w�{k������QEi�ȽQFa9���Ne��.�h���>���%��2��7���7wMƽ�v�_
Ur:s����Y7:��x�xJp6�e	���u��I����f��	@�8�����Ȓ�"��Z�V(	����n3���y���D��s� ���-3q��8���5J[U���r���w��P��߱����>�S L�܀Е�=3����u{���)�+J�n�\��E���z^-T��!Ϲ�{�`�}`��p�B��J�=Z&8��<fyJL���T,D?|Z��஛�ڞ�MS�����Rg�.�Z
M� �V,��꩘�˿�'�����v�	Ζ0�	!|[�-O�|��L�@��\��WN���u_:��uT�Z��R���i-������f{���>#j����Zq>}į��	y�Y{����K�G�q�뭺�*M|)�E�N�_C��g~��/<@;-�\�Th#��s�*�y�G��%"�v�} :�1X�%+mȓ�e���q��K�zP�i�V���W:B( EG|�e�!Wu�KՃ���NBZ��0��TYY�,�V�~�����${0G�b���.�*�7�?�z���P˜튅���^�q Y'��Pt��>�4�%�4����W����K�`�o��Ψ�
tz�	o{�2�H{&���A����]U��*��e�\��p�V{x�px��>�;y=�{��C��:�=V˽��l��pDpOV�`������^F|
�:~워{�Of|rR�Kιh5R�3�ޞn�A��V�F����rh�m%([���t�f�Ō�`�H��^�n�'~6��
�ZS���$��
���S���O�H���Q�5�;Z���n�|���I�*�m9�w�S�gf�R��GcY[�^n�͹��S~�C�|���aŚ���R�2�u�&����	��a��n�P�䒜�\�xI?�s6�T�̀�����������M��7ǁ���G�[��0|� R��4�r�f_�[����6.Ġ���
��
A���[Ë8s�P�0�*�����Ao� �5�]r�t�PH�-X�� ��g��i�S�8	���Ӑ���MxS��>ư+1�ҫ)�s���$U~n	f�«�m� Q)ʺ���UH��	/�{���:�o#�yݽ7p�X�8�~�Ʀ�T�;�Y��׃��hR� 1�����\ɱ�!{����	S��HlO�C)��(L_���e���"JF��n��賮r�}��2���t�����ٍM��2���H�-��i:jm�rz�[z��d[�"���5��g�����KL��k�P<5$��}W�mQ5�Bh��It��������#N�<��D)�)� �Q�䶎z���BɌ$t!��!�Ii�b���v8�s0���a�oA،����^>�����Vt�h�<�7�F��'��C�a�X�;*Ǩx��a��O�ǬԱYj֨��(n�f�yz7�-�ߏ��n�k#C�}v���X8b����뺪�`�2�� �Z���pV�PE����hQ���L6\4���]r#+3�q4��}������J.�jw� J�Q�pͣ��"��V���[nm���B�ԲG�ߝƥC�aK�B�KT4�2mD6N���t9�⳯E�ןؠE�����A��a��.�ޏ�v�4uAT���z!������d.b���'(�_���Gݷ){3�7����pJ�j;Y��t��!��F�N���Y2�x���U8H��G���G �W'6ۋ�+�|`�\fޛr)��Ap��'d)Bis�2!iP�B� 2��
]���} ����o���+-�li���6��T�xO��EF����;�S�{����O���k�|ac�mv�E�o$`]�k�����07T�jz��=��]��=�]wF�Ġ1F4�I�";֤t���k'J�\B��S�Q���c��3�<�[<�a��R��O�E%��1ڳ���G�y��<#�.����Z��@�3)��"oKh2�*���~�}*���I�8!hx�+7�Ry=+4kkG���T4DJ	�:�tB\Ը�O9FiA�c�"0g�k����<Y��I�P6���5�/��C�Y�Ê�D-w�S����x������~W�D�3�͆�&s�-�bx<�{%d~Q�b�.�e�8�;���7ԃ�S k��e����Jq���Ȇ!yj~%9U��f�����ۀ�%�z��{���'p3,D��+�����h�_�3��'	Ώ�5��&��|t�G�BߖY危]<Zp�V��l�.� �R�!�Z�e���n�pE�V�Ll����^x��O��/F���yk�G* �`M���,��2�}+��IuU���=@��f}Q���U+40�P���C��<d�I��j������
!<q� �0�_�+�B`M.r�>O³3M�7��� b�-�^q��I�w=��g�4�޸0�*0K ������-����J��+^�%�8Μ{��Ep�$�������U�}�Zp{|��C�U�H	l���%���4v�d�ZB� ���K̊�
�&r�����_�=��8]`�t��l-���u�a��;�hpI^/��ѝ�e��W�o۷$��1��W���vga�y��{/f���^_3S���L�;��t�d��]8�K�d��t�Z�
\�NmA����F�e��X�x�Y���E��6�W�cK-+�pF�0��H�L��V']jli�;�p˙��Y�^o�[�*��&W�����' �`d�G"d�zw��:)BA{���+%.8N%�!,�DL�s���=���Z�,���Yn/�`9x%�d����'ېD�h&��DM~\?ק�����,�O�:�[���8Y�/y�ncj�`��F�'ढG#	�Ӹ��$�s�䓸�k�ߒ��AXh5�ڏ��E��y ����i�xM�fi]���6&���f��d" }2���'zn4P_�j��S=����[Ak��Y��@�[sܙe�ɹ��T��O�ٮ$)0�v7s\����&^ƖY5vPb�&����5��L>܄-���C�XgY��q�]����+���+i�?�.].\�I!|���Q96��x�UYd|_@���u-�h��QĲ�Ȋ��լ �OQ��Ғ�F�u��pḋ"����"�g�dM@���ж��9���A�e���IO��1Rƿ	ě\�]�݃��DV���m�ĢmV�`�
ig��=�Ex��O�[����
ff��b�H�FE�4�Y��@��(>/�L ���V�S�+c��� ��_�)����(�,&Br�r�rR�t����A#��R@L��[M�*fx���JF� R��g�h[@dY0��a�QJ �M�.sb�����ɀ�;0yH�½EK��~(��lE��2���S�C8.4�{d)H�ڂ�.FT�����!�#6)��/��r��l��A���<��Ԡڐ<1$��ck���Q�O�9��_��BХk�nV8��i�gp��f�X{��S����j�]�C�Kƌ�e���b2o[{21$C����?-wQ�C3���ѩ��c�~H��Y4O��Q�7�v�w�V��wuwW���'�W��J�yDu��M��g-ܥ��p>X9T��u�q�$i֥Rj�@���#�I}�Y��A���n[�gA4i��֧��
)1�\�C���ԊHG{�S1��=�.���aO+������x��f�dU!������	���%+7k�Ѓ�2h�� �9+4�lMFN˭ݲ�r�Ab���q#q|�z��� �fs�C՛0Ϛ�i5>�,�� V�ܿ�ǝ��*P��<�{%���(�]� K�S/�5�(��c-��{Ex�e�s�����8=[�f�4�o���1c�|�mMD��;ڂ]��H�|~[�@���)����_C��h���\LUj�@�.�	�ydm���'�E�m����r;x���� ���̥�3�[O��J_�b�}���u�~�V2tԵ!{5�|�O�p�W2	�i���A��r������s ��:�?r�B�R��8���n�!5uK�������W~�TF�c��K�8��+�>CE��we������@e�yOv`	���ͫ-t���D�m�I/:�\3��j�<�5�/K#6��+�$��'0���@�_M�\߅������n6���W�{�b;LԸ$�L�S�0T�Ϲ�u�>��!r������)a\φ��T�'���+Ĺ��#�n����s�f����e���d���HU�5��#���$��g�Ǵ�C�ÖV���K�nX�
�e�u0�7�'��jV����۪�ZG����8���P��W���T�(3�%�Q��q��˯$��P5�l#i��!w�p�'��Կ��@�)=�eE�'4�\�B]J�k�T$8A��-Kɣ�GvdF�q�	��T���*����cc���mh�j��s�A�e}�}�*p%
���fu�0}M�pP����&{��v��~�A����\9B���ە4 ��o�TЏ2ms���i�'�ȃ��*���hⴆ�v��	�ٓ��) `�ׅ��DM�]#���_����_�M�V
E�g�N�{�0@q;k˱�6�@�.-����2�tg���xj����Qk� c�)x�5k�b4r6�����_�����T�]�,+�LQ�3g���3#ȃ�6I�U���G��e�/-��܆�\!�P�>�Cas`�19xl�"X�#}�V�IpG��ۊ���K��ԗ��z�B�}�����ճs��t]M&`Xur'%2�J�OH�䇳-6�Q]��
����-��jw�����^��8�?֕!5�s�>��i�V7�w��pUu7�v��İ��Y��>���2���̄��N~�:2�����9��4����`7}�0oJ�e��&"d߷�R�%��(�7yg
ߓ��?��b`$��&���~,�!����Hک�v=�"<1�μz�2Z3٥i��z�xL�����'�PXP���D�1�Y3��X��F�4�S��,G"(�f?���~ ���G/r����1%�(J@+�2��xY�Ț�&�̺y�p�$���s��m�8G�s�$.�Qı����l	��c�hm����ê%	��(�ϸ�Xg�R4��Lܓ���%�K��� 
��Ƞ$�'$�I�����z�N��O,���W ���!�Q����|��6<n����X�G3��)�!��9n��o�36N1J��r$�Z�h�>p q��d}��&���`Wڂ*-z+mf����Kt!j8~�C��J,=�Or�����z�`��%���a��J�UN��nL�2����=r��\��u���̔-.�KE(?��:�V'dx!�>ܩSv��36���y峨����M�Y�^��9����ѝ"�o2]���xzn�P.�b��!���,�Z��-���J�vl��@��:!�dB��+h�L|�Ng�8O����.!^�É�@����	�q�gME�Y�Sk^�A��owa�ω!D���ڟݼ�l��D�o�M�mﺜ��h�l�	��+^'�p>NS�Р^�/~F��i������0EYm^�؅]� )�{��SF,��R�iC�z��v%�l���iP�i��\���&>�چp��r8�<��ќ;���IDY`��£]�����	��;�G��&��NA}��ކNV���TD�<��N������iң|�Z����ve��f�R㾇Ѣ�g&0�^#DgEdmp�[t��4��|7���1FR- 	8�������>���nN�j��c*�D����<6�KZ��I��sFb�=��5���ր.������h����#���l{8H���!;#�v��Dy�
_N�6�j[W׷�)0҄[M���9�=Y��W���o~:�6^�z[U*��Y� ��)��.��>��r*-��լ��.8��0�KV���p��c�q̩�:�l�� �1(��d]�̏�O"�%��5/1�rҔ呡<��x}���ra��#=��[l!Y��w��Y�8'j��/�"#�$��LZ��F�4��Gw���kw.�!}�SͫR�����R�|�G�������0y$�XH�lk��݊��J��{�������Dl�� uVxǋt|���&<�A�.�|��!l��)��N&�T�,�F{��443^�f9Y��I0�@P)ęe�+LO� ��?��g�=���o�j��U�5�m���~eP����l�������~m�C(��I�G�����0s�ã��scs�:X��H�/m�t��9�Lyz�xo�ȓ'�^�ZӜ�m�	9�3t�dM�?�k4i�v�f��c�E��S"X��ܡ��q]��d%A�C(�Ǌ0@��k$�α?��)˼�nA�u�S�1 �+���w�1���>+Ggy*N����Q	�iB�Wа6X޾BO����W�q��k���/^�pd��C�l�RY<؆f�rk��ӕ��N��h8`e7�C��5��W�	D{����U�M;o��2����|'����r��,�7
�������׭[}{_Ba�Qq��=�.Nn�Ø|��Ơ��� �7�!^ߐ�� J��y>�up���ȬWT�ȏW(�p�+���3YY��7�| q޾�5��}�^%rxu*�ބ�T��]<�.l�܊�5�-f����Hx,�t����g� ��nt]����Rˤؗ�=!�2Idң�nC��f�����6z^j�)�v}^�J�l���G�+.:���K��7��6�h�^&�Dfy���އn2�ͻP�o�~�ǦYX?p���Lq�+B�����F6"SG��V
�>NaJ2>�:�軩�׿��}Y&>���iN��2A;L����3� V��W4tΆt���+=r�tz�!�Ăuu��/)b�y.�gK��Ɇ�*1A����MR�ӈ����	20�[����p�P��)��,̍~��b-���ހ�����>�奀Sc�����dS�?�f�wj��~����h�)�����JaQmA�n��
�0�E�R($ٌ?��0�H��9��@i�0��R���/&��k}n������ז�f`�[o�ŵjZ����FL����B�A ��`�ܭ~��RV�z�y{��RT4�vk���E��~���;Z�Po�.&㷺4��4�bZd�׌J�If�W���qѵ���j��)K��*�&I�{��e:����]jH�^��Ju�� ��~X(��Y5�c���%�����GO��{%T�f��ZJ�D��5�Ȭ�Ea�pU,R;֑��8�=�t�[ƒ��c]tH_��*.�>$X��EZ�!	.�M���J�MN*����m��|�ZjV)�������7p��!�n,�h�i=�񪢌���݃Bu’m��2�%j0���g���z�����(��ҕ�#��|ׅD�䷊�QWU!v�v���e1
��e�N�1�g5��~�j��4e2-�9��z�p3��8�PF�R1�>A��xR[(V����o}H@Ym�h��:��Ȣ�����/e�We!�@�}@��'O�5�)�=��+��c�	\�+�^ˤ�_0Ά��VR���JF!<�'�aW3��)����K }xVE1*k�V6�q��0���G�\�FB�f�*�<�]Ax��R�d�QZ��`47��)x�� ��Y�f�v] ���"�Mޮ��y$����؃�V�/�B[m\4�����ŀ��#Ȃ�`Q�0����#��l��$[�K�inh�v�,ņ �=o���8Qݧ^��Z�>�< T@X�7���2K0�H�C"U�]��6IvF�7l�|L��O;b�
Z۲��W�a�ʾ�?��Zp������$}!�K���齜f��7nFD|�~��Y�E�����'gup��"��,�˝
Y֯x��R����x��rq�uP�.����%�Ip@�>}��J��%V�U9묨���.��E���[I]�@vG!!�؁,F�uXn(��z&<�}���R[��7^ܞ˘�]Mо�tE�Y�c �j�X�U��eo��o_��Z<p����'��������8�![+�A��1��*�4�ad���~�ޔ�M*���o{�����L��x<�������x5������eP�}Ǯ:��������E2�^��#�����A��ȷ���W�e&3��!��fת�b�d�8�zYm�#���z�n��M	GJ�;W,fF�8և�s��L�)�|w�gdfA�C��EذhK/��Q*#aʋFw���{�i��J*��I'��NO�s�F������$��@����n VPɽ���9���|���%�5��^������[��΅�X�j�����;�`ݩ%�$��r���VZ��鮹
ϣ�����(��4��#�Ry�qS�
��໺�/#�� �!��Ǩ�r�'���Z��'5o�T�}A�f,:��Q;�d�����[EY`l�~��O:�v9�4`�Ԟ��ϩZb���|��Q�g(V]�@��p�v$�¡��2>Gq�ENv�J��wЛ
5���<���dBb�D]0}R��!|�M��_�Y�,�F����A����/����|v\�ˍ���~)�v��o��ⶾ�ֻ˧0R��wd
ˋ��lFd�n�E*c��=���O������1�ABӵk޺�5�/����xI��/����.B��{*�P.Y	��W��E�����s��|���/�ۻ�|��#����±u�Y��ǹ����d�a9��o���G�)?U�Oz�#��E�p	��qR��u�
)!�CN���u���dû�-xX�n�ֱ�H ��7���77�2B��~���!�^c��^<�%ç->
�n�����ߨ��0a*�zwQ�"5�;��gZ�����wzu9��v���[.Ǣ'���}�;-_n�4$Ƭڐb)��F��
�8�h�+�{a�=Q���H�	&�H��J
ؚ���:�`��`���� �P>��́��"�?�����y�%T8e����j�&=Pv�W4�C�sgM9������nSp�'K3�8��Q����`S������.{\��o\)�2AӦ�m�|E�1�h�~zD�O�dٝXU�턳f��{<Gg~��,�+��Y;��w�3I��\�j�.��,FK���9m͍�Rf��h�/�`�ҽ��R�,h�@�x�|�͛�QӚ�d�y����|T�"�"o��e'Πej�& VJ�x�e���F�	��<�˴�Kl���bP��(�=[���x {>�� ���Sr�V���C�O�j�j��N�t���Ġl�Y�m��sWJk��Yh(�m�(�	��>;2���յY
j�v׀ջiK�I´R��ړ���TTR�k�D�P�ْ��� �"�,��ō}�]*�j΄�N�{d�\4����ş�Ǎ�0?�+z4&�i,}��0��x�RR��AK�"�/��'!}��y��?� j�qRPL����K)㟉ݶ�|u���M������.�\�x�;pb�Pa+�a� J���3@��t��'�Z�ZS�/�^�Ԫ�)��H(�P��ߝG0�ۯ)�������m��3mn;Yֽ�։���^��T��+���W��zc��Y��X(uAy��j�σ��������|�(;�.e�����B
�z�n�Yȩk�ʸE@��%�|��r;<�L�Wl�c����8:=Zt��{a�r��ő��ttd������ʏZ8�*S+,%r�A��Z�t_���@�	��/�A��%����S(�C�&*n�Z4ޤ�p��a��|3x2�+�
@5�i���o��[�Lkz)
��?C��=�����Nw������<f�6B�V�	iȽ��G
��}N	�t�Um�k�F�b���3<����#u2��zd��uB��!�YNN��M	a�����D:�{ڊ�����|�.���E�t���\�)�7�	�dp���>
��,�4'[�%����Cm� N��Ў*��3Qn���D��oҍ]x�,_��̅� ���	^>�=�&����I���A��`�H^��G�ۛт�n&����s�Di���p�dϙ�[2�\�,�a$%����O��6h���
`b\
I:����&�/"�s\��p}<	=�o�L����fв��ˑ�W�J���������{��1�i'u o4���d&s�P�F�(
f�~��s�u&5��[��R]���=L��lZV�e�����,)b�H���9��A��ă"w]9  f�o�#��I�x��!]���O���ޕO6XoHr�%��@��·�bE&cqAb�EV�[�����ܡ�J�;S��m��M�{�T&t��'�:DeQ-�'�H�X��>�e��X�/j�[ � Lh|�
��L�������xZ_��t�˖Z�Kv�'?��2h�G�<�cJ�5,%�:��>5`��FG0�*���3T��bWPX[6��������ȶ�M"<xG��o1�<�ݠ��]+(003����f�on�Z�oB$��볿��R��U�>�db4e��btÕ�F�e���)>�$����Й�Edz.�U�lح�ɬ.ʒ��ݷ��&&���;���cH��]��g�F�Ѧ y�˼T����ֳ���>��n���Lkg��z�y�Q�P4��xfk�Q\����K܍ow|\��-���~;*�@��b�`������~�Yn�mRb)"��P���!5��O�]���5n��55����=v��}��=�/B:��S�3����4�XN��"�C��n����{����4V:m�l��zBo�.,�ک�7��2Y{)��Z�+�6�nk3?�ܥV���|3M���	>V������݀�%��Q?�b�%b�*�eZ�X�U�����@a�޶����� Blkl�=Xsk�{�=qC2c�]	�T)Ps�J&�ӃY�j���c�ϡ�p�%�3��TT��;2�$�Uߤf;۵�f����w�ۊ�N?e��v�y��O����L�5�W�(>+JR
 ��
���D1LbQsWl�A2U��S���B�j�V�#�.𡌤�;p��5~�2�i���M޸�QK�V7�7��5�E�_ٍ��CH�eh��]�KG	}�`�A2��<�A�7���S��b-}��k����
���3)��(�>=�S��Z0;>>Ԃ)i:oo��W�_&3�U2���T|^{��X�i^��q5���Fז�����rK�	��a ���)��*̽r�G��< ��1E�� u�V�%%�C�ݿ�TME���Z9�������|�rA(�L�
'�!::D5« F��Hn�7|TJ�GDDπ7��+�ɜ"%&E��S��}$���&k��vކbg�w`��=i
���/7�W�;>7��)�����&��1��'%¤�ia�Q���K٘��!|J���W���I�F=|���*_`[hz���$z�U[�9�����r5�8�-��X�G�L��#H%�U�=���r�Г�]u�k[�^�@X#*hn��^��GpZ��F,w�&x�B��-��e0kL X��uG-n{��n�:��a����B��o�_����?�r���aD�wف�'d��
\�.��SB��f�iW`2M�Mv�2Feoo`�-`�%���$a|�ijAV,�%��x�o$�U�1��-ߙ���E��� 뛋��s��ο���!)�v���̏7�G"���wc0!]\�gՁ&� �˟S���[����`���E��,��^B�`a�d�V�'��F��6��W_���l;���R�W�:� =�NHmv;c��&�A��EjdT�u��E���o�o4���+�*|X�C�p�z���K0�?�㘠��w�!]܊�b��U�����=�ϡ�tm�N��xT+�«�^<���ؒ��[�ۆ�;N���1�\A�u�m�B *�,R|Z�!�=g��s��H���n�W��������(�U�6|v>���;ͯ�d��6�F��7-0�>���F2���"9�c�xL-&M����҈�|�Dl�G���e�m7��;	(�ƈ�H�}T4�"<�����2���iV�,<�w��:������/B_�7��D�0�������r̩�Syx�gW�5
���}+�d�������iy�p�[��M�t���?"Y�|,��Sd��Dm>�����\J'\��0�x���5,=��;a�Ü��s-6 �c��G&^ұ�n
���4��0"�1�:ȰU��{�������IQ�gދϖ�|�X(T"���qk�^���O������2�l������U�,�xr赙5bF�#���7ȾJ>Oi�E��bC&��e��W��u��ޒK�I� ��yZYk,�h6b�ջ'Za�M�� �����\vr��Z9�B3u�`������w��.f ���l��aoW�m򲵲�vg}�VH��(���:��ב\�mJ���E]��LǏ¯�0:��V+ ��R�Nt[�@mn@R5 �P~~'���:�dy��8� N�.����4��ܨgJ�&
�lF"(]� �@Ek/9�ך6s���̕:t/�.`�����SZ:q�����(�Aa���gM;���oM�,�,^��c�[��"$`g�+�ZÑ&C�'�F��M}͙#uaL;�@>&�%5gm�I�(��8���<7�����>��6*G���IKv1����k�$��U���Gh�AE�Ռ�;���$פ���p��'��pS�2�kvn�X^�z�@��b�ڵ��?�z����	�����44>����r~vI� ����;	:/�&<�S>A�Yd��r�_�!����@d3Ĕw��1N8|�l�*��c�z�[ay	_ƽ�_(��8���[��0���أ(��ԇ�	X��Q�'�p�~γBR�`/g2	r��ծ�^zG�c��g�/:������=֎ L�a\���{���#��GI"�bBR� �J�� ��CCM6�8n_Ģ����S�xt��?؛�¦�(L��v=�s�rE/��|k!�⨃ժ�l/I���B�Y@dS�S2S��z�ب�*�ˢ���ט�w�V�����.�E9�����)m�������oȮr���QL�`KC�+n����A���t]4I�#fɨk�=/��݉��$���n��օRv�/@e�4-�C�����M,7X��cE���
/�K�}z�{W�
I�x�'���7�k+N�Q*	B0h:5|u�y!;x/�\a�)宺�'L4�:&���׈s�'���{@���I�}�y�_ q:e�M숝���� p���7k��*B
����J�;�������{P�xN���ƿwz�-̩���9~Pq�"]$�+b��Rw}�B���P3���}�@R�=y�"8W-��Y��V��|ğ"kCG`-b�ET!������r
�`l������~C�����T����
�0lrt���p�As%�q{�B�Ԗ_����w�KI�E1�wLo�mM�E79�e�Ƴ��6R�@��y�	�d��qL�������uǒ�D`���ڣ;��_U�r�[$N|��2V�)��l-z�pΤ����}�r�?�^�����GF���Ǳ�UP)"Rؘ�z�C�r��\����Iw5Q��u�λ�q5��=�(���^pe�4>b�Ӑ�]\�p�P5oZ���g��W�V���ٖjw7�͏�A0d&��'|��D�\�B�pZ8^rʺw����!��zgӠ�T4��R�E�(Ulzݠ��� V1ٮ�#)������������a�	���Xb7��x���N�H��Z|3���'�ӣhڤ|��Y��a;�S��j�J]�-�+���@b�!B�`��\�N�e!�"fh�����uv���I��~9/�%3�o�*NJq�+�t(���s���o�L2��V�,m�\ƛ�'�R��{'W��١����oD�l&��K��c{w،����@��y��Z�l�/��*'t��SM|"�%_)��T퀿�q)ܪ��V�W���X^�"z�q��r�;V�|v`����&G�y�G>O_�Up��Ȥ+�	�!9��(�[���j�]�8e�jB��&� �{� q@�S�vR�f��s��,��VeNu2��O��X�ho�d ��#O;!?y��ڧO�q3���|a�1�FN�WƱ{�~Uu6*�Y���H�1h�R�d�s76��x;�ʉ9e�y���t�  �����J;qR���O��2���jKH<�R�}�y�@Pl�M��,D��O^�):�{fY��KS!�.F��l��m��JM���m9h�X�K�8
?h�����y�V�D\fdt �	���FvS�������&�&�vZ{�l2-[g�@���G�ua2�����.�;�=O\��m�^�gV�B��
C�z�y$ϣKF<��:�V�m!�:W�w�nc�&��9[�G��2��k϶?�����3�%f-����d�<t	�{(s��������i�1й��cp#X��;�Ε��H�@��ϱ��V#N%맳����%���[gs�+iY�B�S���d�!$K��]~R��4���W8�IZb�q2�t�.5�0�����v�W��ލ��oK�� �Ybt%m�D ��+�hд3 �M����]ٸ�5s��Sal��c�wf}�� v���A�i���.3,���xφw��Yu����A�b#^4�)|���%�z����s�����;Hz�6�B����p��`�k�oi�b�����������
D�Zn�'�/�P����;�z����>��3��GX�,Dxz�L�^�Z���3��fE_۱�ܲ����Ȫ:��-������$������װJİ:��c9߫\�����S�*o&,������x�̻��n
��C~2��"B�w@��t�S�D"��$e����2ظ��)�g�i�N�c�-\5j_��e�.4�褜I s�1������Y��EQ�%O�M*�10U������S�bY�0K�@$���i�5S�v��yӌ���"����~a�طZ j�o��J�h>�M���jݜ�ٔ'��7$T��ՔJ��_�*����0�Zv:���&vA�*��6�q�cG�.��A�ñh 
���cqX��Z�k3۞1r�8a/3ZS&ף�;�iV�,�Bn!-6$����q;�;��	�f���^��jd��\!���qdձ,���`�7��Š*^6���D ��`�7�Z�|�s�V��.�JxdV�Q�&�!�9��lC#�o���2�7*��r�7+W@��'��n�}���\g��[��K�Z}r�#&`�N�쳮�`�g��M2B@`�"�ڝ쵃c����*���TX��mxu_|�7�̠�M��b�^Y� ��S���Ԙ��%�ȹmun;�]]heW[c�	����׬p��a�S����_J�>U\y3���[��>$t$���"��'LR�����d*��èm��T$�G��|GU
a��N��{9$�1�k�H+Xe���$Z\;���d�ļ]��C0n��QLB4B��u�{s��eC#Pe'T'R}�f��»��|mIgAf"�iɳ��J洬Nr�s$���!�	�@��Yd��n[���bŌJ�f�C�,�}�+�2@pwPL�� aK��Dz����D�O�]ל!�T�%K�	pTꬕy��]�7:��_�1�}#��Jt	��Bil�#�>�����]І�rT&U�^j��$��aQ��ל�8�Ng��P�2Q�z�$Nt�%����b����c3;�kH��ꎚ�94��.�E$য়��V'<!�m�Q��Q��;��[�y�A�$���k�ƶkxR�X�ś�jf$L�*k�K|�b�"���`�R�r� �^�@� ;a��M����a�n!�#AX���hώ�F#�Q�k�2b��Ax�H�8����*� o���,����;�w�XY�6�wZ�X �j����}�f�
+�)]�bI�x���Y�1����C���h���|�M��.�?�<��"�����ݯ�0BT����I�H��D?��qҨϮ�pkW��� �؅�t`;�
k������f�G�O�YG����K�"����]��jx�JM�y��c�{��a��3���c�\f���~�'p���ݭW�Р+��HXD�����w�]zE�ݫ�c�Y<o��#Vc��n	��-�e�BQj�E��Zp�;�b[�TLshM�A|������E�wB��v�H��&�n�2�n�+Q�P��QqL>�Ұ�_g�%kjnc�s��ZU�[�1�����՜�xj��̚'�~j巑�7��~�e�I��o(C��[~��80�SQs'kU'��U)�w�4�68��5uq�9�>	ygr�w3������ f��'�+I��8� =0*�si��J'/٬�j�U1!]-�9^�w���`'�}>c���O���q�f�\r�S@�n��`r��3B�s#֢�wUtGO���"}�&|��:Qݖ�5�S�c�hѰ:����X�4���+q2%v�av�5z�~�B:��k�cjxr��s˙���M��NV�Pv�}��M�YkJ�^T]��ɑE����Uo��ZF��gB���e�)a*��7��=�?�1���L!��t�$�X��C/��k90��u2�h-�i���xT��+ ۤ8��{w�" a�P�ZU�)1���c�R����6�(�pٛv�sy�Uȷ�rY��P>��tJ�d�su�f�3���nI�R�N��Bc��������l�rΫ_x����Xg%�ƶ��ϕ6���9� H��9� 7�����K��z�|LQ�e����x�y8%.@����<�Q�ɹ ��R�9�.A6%t�*��_i�1+1����]c�#k�b�Ӥ}Υ>|�r�p�k�WY��)8�$cM���C�^u
�|!�Ɨ��A3X�7~=*�!,�B{ZXr�[hL��W�##Kg VCY����r���
�d{-(�B���u���s��y������qm�0������*S/^y�'���+�}��f:m~}`�����Ԧ�����0��%buʡ� Ҋ�W_ �����%����B&��]��'H�+��c}f���K��_w/\2-�y���vb��
j�v���� �$K�h�/h��w�}�v@� ���dT��ck�X���>(a�"��RP�<�5���D�C�"�;�RH�kc�BHo+�%P��|V)���jt0>�v_����� �2��-Ę�������n�c�U�!N�f." ����Z&�L�_���v�ձh P�h\?3UӼ/@W��V�	�,�}t��ȧͽ�X;��N���3�_b��܋�r�p����B0N��b����$�K�.. Fa��P<��um$���a��j���P��{	z�J�A=��2��T��$H.� )���*�Ń�ó�8�e��Y _`�/r�3ʵH���H��U��8��#�hk��@V����������р[�����ȱ�nU6�W���2v�v3����C��f������6a�][VU�s8���(#�N �9���X�z��q�Ͷm�^a��M�a���\R����7;�=�F�)�����'e�#sg�}'�beȧ�@�ݎ��.h�J���@4�ܚ�Η��c�: 8��y����c��hW���M��Kp���E�������i� "c�Ҟ����qg����򇱱}P�8��C�T��xD� A)��@?�ž���1TL]+t~�����79,�XЊ�B�c��,U�?Y�j�;�4�e�j����"�@���bYBT�d)i��u�D+U�$��a��1�'�˜r���kr�V ���ӽ��Bܿ%#O�K;�1����J��S`c�ڢ��[�d�k�ҿn�)����5�9��;Iv��rm*����Q��P�p٘S����| ��bb�E�Q�뼦-
T��jM�T�]�(�#���>�c�p���c*E�1���1�B�#E-��.c0&��Jg�L�6���*C�t�B���툤Э���f���B��vͧ���J�B���q��V>f�Z䕶�}�vF㹔�m����0]�
�g������;�l�ٰ"�v�"S�ۥS5\�-Z�+lm�`���7��n�����L.ΟV������+��]1���UqzЅ����eʙ�vBc�LGsB4�Z�Ϩ׭�~2�3L��|�����./k��Q�:�k�ܯÜ1�,��6j�&���7��#��g�9r��T�a-+N�{��W���}�ô���'�.�\o�I;5�QN�?�/C�G�.�̭��C�� �*��؂���fp�W�f]%^o�O>@�:'�NNCFt�x�s�?�v�R�2��{�1i�AWĸ@[����X�>�t�M���!�0���kW�Sf�N,$�<$�=W��W��� ��ˇ��Q�4|����1dƮx�W�;�P@}I?�n\��e�p�6����g��g�[��<�E�Mn�-��`)��६�����P��������!��B/�
����;��`ob�Hj�y�)�	�7	Bt��:��D[p�([�����ݠ(�@�5g������h�����w���ȗ��-�#�gD���fL��+'���B��yď�>��Ȉ�"�S5����6��E�!Q���K�t��+���s�����?��mkz�1�C�3`��p�^pk;n�'��i�xܫH7��+ڴ'�mW�D&d�}�E�S�1��͢�vܭ�1\�&=���-��PX�|�6T�-D,$v?܍��/9��Pw��#%妟�ԣ_+�AX�p��$�yZ���ǙÞ���k.r��N[�����ם��=�D���4�ނx��\���
!2^T2�i�ȭ^"J^�2)�F�O��/��0��k��쵄>��Fh�ɨ����,���	�B��$6�"��Jgn������K�ŉ!�j�W+��oga ��v�X����PY��TY�~�]�;b�.ɯ�qE�_ɰ�/�X�R�T }��6'j�ɳd*e��>��@{��QR?�L��W��Z|�-U�6���'���,Lv���k>���߭%d(�hZMH4��Jc�*#�=�s޼���#�`.�к�2^���D���-�}ogZR6��\cB���zt�f���u��۱.�ӗ��F���q>�fn�	�?�ԓ��q����(
�ۖV	�f�o3��WڪK&=ֈ�;%�
�	Z�nРsR�UV8�$Xh��*���
�C�bW�8N�@X &�6�qHZ�=�Ku��|H����muɽ�b����M��!� ��͚Л�n��)�P���\��0��^���|��\B�O�j���K᧤�0n�*����xe�o/1��z��|�х���)��VUBk�����mx�iH.��n 7r� ���vh�y9ڼDTF͆��'�^�s~�k2��%/�X���SȌtT��F��#��W���^�l�v�<���fDy�M���K15f�0p���GN�G�
4���Bi������G���Ǖ���ť#��dd �y��>�1(��<�S�9u��_o-�b�	���5��
F��nDŊq� S����M<P)c}Ս���3[�t����YAa��L"OEH�Rg�����y}jG	7E��8w��Ɔ��I��I�H�v}���X��b�TNHdaJI�^���`W j���;1\ڮ&a/�2����O&,��s7"N�wr:��8�v#7���z�i\u-n�=���)�ȃe�g��� ��ʦ���n
����hēM��I�l�cu��D�vF�Hv�U(��P�F"��8P�:�\�!,��I�sЍ\��eTq)"H_Z6kMOz���qe���'(��үun��/�.�%Y������M�~�Һ �j����8A �y�:IF�m���� �����TP<���^@�wAqd 9 ���M��W/sl����]^w-��L,����KJ6�[<\�D���5�FW��ʸ����Lp�}gg߹��$�-C�����?l��@xɐ��h��@4��R���%�poe}��k� �K�X�oõ�ws&��\	�p�c�V����L�s����f����k���^-����e����n��W��ω
v|����Q3"��~�ۤ������G�}H�/\�oC�.gr��G,C>�%2�h�m��r�����Kn9�":2��y.��!� �E��_.�r��
>O#��^S��+ËX@^݄P��k�-��C	ͷ�ٺ7�&"A6]ebE |��xҙ%N�h}��,�_��Ǯ�H�]B��4V|��������n����H;�/O�I4���ø4��È�^�H�nj�[�#�F�/��IĤXdz@!"_��_���8C���mrpv�ԗ���Վhz�Q��zN�8X�4}�J�n����6�P3`+|��Ճ�ߐK���ʈ�s�t/)ɰ����=�j�$k��wR9v��-\�}�W�!����c_�7�w��Iى�UQ�����!�H&��J�|4�2�hm)�rv!*|�]i��i��sq��4Muণ`�(�nkr�A�1����,�8e�5P�S��R�*:P���1縵�{s����D�"�[+�Ћ,��(�I�;ꈝ����*��Yr�dMxك��0�(-<٦V��}�-�/xF����ٟb��M����!E6��2T�<���x�i h�#�V�1���3��̅���2���%j�{�@~f5	�"
��G�NP4B���K_Q�@�g0�B�|��k& �Y�Uo29$�����V:���q0���ѻt^��\P����G�	$�N�CE����+ó���\#��J����v4���tS<�[3�hB������xM�hS�<�ԅ�F�w�9xQ}�Cfh�É���~�_^�Fˆƴ1
j�<����؜���gP���T��(�I�dӗ؛��%��%����$�!�Ʃ|~s9��o��F~$�@�$�H�]t�ֽ��f�o��cc|��S������<��U���������	�@X����&8�7�?{��sk�j��!��9j�'q���W^���t��x۬��דjM=lu�{���4� 
��mVu�P���x���v���?������~`]F���>%���iC�Į!S�*���.rT�Ξ,$��1�=]�BviF��=�.���͗����\����c�0���㥾�$��73��"���i������̰���}��������e��A��u�MJ�t1���R.W���_�H6�Q'į����^����z9�^�
���aϼ�J�g���͞})XS����Ez0(�c����Ru~������G�?.r�P���t+0���������N$���T���K~`���^��Ŗ����9~]�&An]�W�^��l�xl�h�]��V���6��Tr΄�O7O3���#^`�"��
U�8�F�r)�1��{�9W1MG�����6:S�3��|���`a|9��x��쯎�\����C����w���Y?%ֳ�aX>i����L�?��B!6���$c'�z�����k}(/>$$��I^W7�*�����ܒPɌX�&$�W����5yu(��И����#6j15*&�<zP����UyGh*�ԘUQ:�b#��?��//o�!Իj�~���&;FS��) ����Z�=j!o�rmR�T����nC�<�x<i�,�,�{�=s�Yqx��p�ۣ�@��P�g�9A����T�!��}�P߻�C ?�c�4B���Q�?o���;�d��..gPw����bl���@S}��(�c8��א���~�I�DA��>Hj�o�oo��^�y�~hf�~�฀��Xoh�V�QYzw�1�m&���4�AX�^`������� ��	�Rl�<�H<w��7d5�V ��SV��<}dG�Ť�Z@�+� >9���ǎV�ĥ����c�^sF�c3�\�x���]���mί�[g��(�K��_�OCI�2�oZ=;�)�E��V�X�w 3�i5g.��vX��ے��c��b_�����Vn�i�З��L��R�}�l���!��m��}�k���UF�<����;�V�܊<T�.��3go ж3����X��]P~��@��8�������ָbZyD��PОl$����� &}!�h)�ql���ގ�6d��"��գ��ɽ$juvF�TE����Q*3���Ӌ�N4�\�2��Zu���"�����0 ��5��~d14�9�=I`��R�u ���Ձ��w	'y����v�]#'��k|S����1N�Dw�at�q�u֫O�`���	����^Z���$<U0�W�t��)?΍��Ekd�x�f�����5pHCFă=�>�fx ɾ{�	�z�1`�_������E�9
�;5^c3���� |@q�p�8%Tq�N��I'-U�x�v����lȟhN�����f���ug�Ɖ�k/�I��PE���tv)�ө�Z�]���^E��M䀜�,M���̪��P�E ��>˫.��q!��Z���e��3gh�9���h�I`bY�����B.��Rfy����;�s�^�s9��Z�X�62���l�t~�PrhA��^�+`�,��?����w���Ȕ]�Ko� �V�i{���/�	�հ���I�� �������?��xU@�3�,�(��9������"!�������SsM���[_:&i��-�b:��R���J�U��%�!῏������MmI]��&J2F��H��Re��Ǒ��ڳ|�`�(�� ��!��r��Nyf�M�����̼+jr̛�����)�/��|;���[|�~N��X+w����Z<�ǒ�?p� �e~��n`hV�*=�KΜ���g�0��x�I!�]�=7ZC�q+vt���ҍO��v���Q���qs�p�f��K����?�g����֐����u@�,Eۯ��%����SA5/�;^��kxGF�-�s��Ƈ*�9M���]w�L0+'��q\*��q�&�}P����uvǅ ���<n�x0�a�������|I�d0-��Qy�Ԍ�IV����QQ��_���������.0����PhC�%#	�����/������U~('3ۃ*�/#����4�]|��-��}U��� �~�;�(�e�sJL&^_0۴�s'� 
��
7������^A�����u�����j�Q픿F��-�q���&m���&j�Z='=+��6�)\tUs�4rb���/����*(�ŭb��y�	ߛ�
�h���}��%�91�&�,#�	�r�wO%�PŹ�9m� w��(�-�i�`ͅ�b�jPB��Ym֎�A�8@9r~��(%�����茽P\fsG��ݐ$�}�T��{�H��Ζ�I�5���W�M���9D�^�öeu-	�+S�6r��7�t&��(�O8]��e�Ȼwʷ.�qw��Ƽ)����C�O��ɜ*����_T���<U�+a$!�zy׈j��m�r
 �و{s��ւu�q+���ݾ��y�m�	#��G�	�B%�)�l)��Sg�d���\\7�	�Y���4�F�w'��p���r]��%�=��s��Y�
��m�b,���G/����b�5����	g�\�$�(jsr	ߌ1�S�d�`Qr#�R�%,Us���S5����)�I�`t�-_�����Z#�z�㵛<쏬b��>ce���E����)�i������E>��c��$��,�2�O1�Jގ먊������݅v�)�'R%��e3Ɂ.�("��x(��0���_�bĖ_�7hU�ikh��z'qO9�U���3�>��<wcA�c+Y�+�̨�AC�a����H�4RH)(x�]/q=�k����S��\��tZ���T����H������q)[<�8��Q���Z�{�2�����X%�kv ��@�(��ڜ�i��y��#ys��'g�,��dew����C%���\�\=��`�u�$�%�S����w���;����1r�}��{�� �&�u��@���o���`�7���n���W���X�o��'ɞR?#����@�^��@5.���;��O6���8C��d�(�~�8ST�I����N��������R-'#2WC%��7d��-@+�`c@����M����܍�`��&��mej��ă܄$(�ԡ��f_�8�|�R���HMI��:å�S�x@�Dtw�����枝������w)���<���ȕ�Oh��T����*�6�瓦���R�S���Z��AX}h!X�R�>Xn#w��l{���4BJ��hD'r�~��p�
~A'�,S�vY$I�}��e�Q�x��<#�܆Q,�'���{s�����[�1��ic5���)���Q���;�ä�L�ur�:<��S�qk���7C����h������Y��m�`7�g�fԴ���{��~:b�=z��}C:@�s�:�y?&U��N���1TaMoM֧��jLlP�F$ƚ�`����T2^�Yc�(�f�E��d�N�m����,T��1�рѭ�c���Gx��f)������m����Q¶:����;�5ܡÊ�},���y�6�bo�@h׮����pi��Z���������En�P���k�zm�����UV�@��Np^�C��������y�Y��B�7,)���YqAC/�zr��Z���2�$˂s_%;l���s�K켿���@x�#����zY]�wp�E�U�6�n�# \��s߈ԏ�ɭ��`C	��)�����l�z�+��,���w�����ox*���ԑ�AJ�b���z?/r6FE7�GR�y��/�����6P0����$h�Y��+�y3��&���<}�^Eff�(�6"���a(�%A��fY=�.�Ө�� ��������;���W�퐭 ֝���6��[%r��M�s�b���o��Ӽ2:���c��U�o�'�M����v	s���(�O�D���{�n�"��a�0��<����YZ*|�ѳϖ��x�����˃]n�R���!#g[I@����^�����i��L��'Nބ��9eVFƔ����6O�4�D;��ٶ��n�.l�m�_�&F�ڲp��̲c�n�T��k�f'
����ԇ��\�/$���?��"~k= ��� �7�8��2�&�N���+7.
�|	+E�P&���xN>[���k~���m h�3�os��i۫�"N88�A �'C�l��.M�4��Qjuz�����j�D��. �ي�uR��J+.�j����EV�Dl�ƪ��ޏ5t�T����N�͘���uC�z�j�qy��6�V��Do�
=�M��*T�[��z�L�}�]
�!OT{ڭ����/�XfC5�0���*N�p�C��z�����Ѧ�����A^ᯔ��I܌�
_�̠���B>Y�
���cjO��/�|~8�J�ē�Vԣ�����Fh�q�EN�'��Jt�3I:�9�n],�E�]~ٸx#\�����?���L��e��Р��]�����Z�]SU�6��F�(���,�����NA�g<\�YQV�/����`Q���8^�!/ �,t�ح���d���Vq|�6�}e�u��T�N5'`*�_\!�r?��x�D��<
�[��i{"K���Ɗ����U��D�5�÷�"�q�����T��	�
�F0#�c�75��j��e�j̱�.�:8����{,��(�n5iH�)�'gS� M�LB��'�R�r�W�fz�� 9y��l��
8�@��DVN�BR�pS�i��,w�)�b7�v)QASIu����]鋌��*�mb��ۣ��	n�Z��%�� ��y�8�$��~ ���H�[�F|S�U�h���yL��|���5���J��A;��=ZF�bY�!�[z�D�Rz�ϒ���
�-���E��]9zH�Wm���BT����g^&��n;ؽ���#p��琸��޽?�Wp	���3�pr�R^X�r��mN-Cf�c����yqbBH������_��T6��۵+$w�ȭy��aq%K�Xzgf� ��WiS�Mt�OQ���#tX���2���t�".�f���|I�3_c�}��f/�2�:�(Ka"���Q�5��~�/��B�峫F!�k�*�d�~#]еo.�d�`��d��9�>�}$(��'�n�2�O
y�c��g����Mc�|��0�k��2��5�:l5�rm+�{��o�d����P���ǭ��Q����?��օ��i��ܕI"|ς\�w%tA���!6L���_��ZJ|.�����,�nC��� ���g�K1�8~	�jW�u�<Ei�c�A0;+Z�{�ڈ�[ɉ�Hf�>�I�{�p�0�p�*D)Jp1��S1+�[���{�������|r�b�L*����Q.�ɾ�-��%Y��}-Z������89���L�p���=)�کBһ���@��ʍ����QR����PH��{�B8C�&�g����3���
�E+��`��S%�����-2[2P��J?�'���sUh�;��/!�+�y�T�Y�6����Ρ>�x�o�b�5���e(O6�Z�V
�[�ŵ���C�����]IX1�#\���APƖM�I��(L+��ʠ0��2�M�LF���uK���6_�n�����'Ҭ$-Z{ L��P��G���?J7]��+ǀ�������ΨoOY�?�P�d[;�l�3b
[M�����Kx�|�2�u��q�>�i���Lr� ܙ���C��n|��Ӽ�zZ���v�X|c�v+�n�tj�?������:k�G�u�FV$��,��I����ia{�y=��UH�/W�5�5����ƖO%��>D�_o�U�̈́ZRՅR�Zn��Ыr��i���|}ħJ=\��0���I1͂�N��,&Ɔ�ۅ�)rg�n^)Y2�5�� ��t{�x1	(wRYF �F�-7�f�2ߙ`�{h\_�!�/"��
��?�_R��̖8���q@��s7e���g3���+���1Mמ� ��w�J,<5b�q���x݅R��xY`��M_9^Z��m`n𺯘��=�_-nZ�u���%�3=�HPt�B�^bدx����r�2˹���}O�k훕3�t_�:K2ؘl�]E��T�xƗ1��͡jQ]F�UL�¼I`)��HCX�09�\�T+�I��}���M�u�W�Z*zf*	�@�Um�F}�\܊�WE������$�?�������	[t�v�������BRѫ���}�Ы���\h�X!]�"pݼ۾�"z�X31�����>��|��x:��F�8���d{j����oWr���]�\_0+�����ި�N�2���3^Mk��)z ���l��)}'�E{�0�����	��nLϣ�[(�3[�e����AXs�e�����Hq�0茙К��(T��:a��=U����q��׍�ޯ������'�sق=��3��J�d��X4� �[ĕ�?Y��E3�{/FD�4DiE�B@s�h�1�񬿹s7YJ�SeׇB����4g�/z���{y����m�&ΰT'�xY�M-�AW���;W � ��VnY�ü�����Sѿ��Y�Ƚ��eA쭂�ite�ܗ�Q>}��琍P����0�Obb�<���~I�j\�ۑ�XA(��c-2g��զ�����u��y�R�0M�(���W���u�Eme�7�[��~�	�%x��3:����ZGp=��]�hҿ A��㣩;mQ����Ӏ����viUr���_��Ġ���I��j^b�v�!����z-��T�"��A��b��,����_gڝb�
R�8�b�C;č����TtC��fk�e��҈$�0e�#��uG�BH���)�b���?��y���A�?�#R�)�1Z,�4C#@�b�{'��sK�ˬu�����%�]J�&EۅUd�x�Y��9�{������Z|��jR:��~ �[1�їmj&]rNR+ޟ���1<ff��нs�c��&%�����P�a��&s�7���j�"o!�l;�I�Z��" �B� ��e����h �=0�� ���k
A/��X9	�-�c��
y6�4���k:�Y;��޹Ix���4WQd�Ji\F�Җ���U"�7�7�8��1�{z�O�I>�0�s�����.���w�Q#X�͏�R�2S���*m��W��8eV�&o�*i����"s8"�W��@AQ2q;SX��є����F�)#�����I@���UyR"���������1
��P�*l!�疖�U{����4��i�^L�=e4�ĴG�\T۸�*LQ^���ӗ�=�8�2O)k	�UlYꂠ���3������!M���F���j�`m��M&�#,�~)
6YY���J'����ḳE��>��SX����������j��z����
��J��K�FTN���0T�2uC����@r�'C��2�k۟�zm��7hz��QD�/zSk�8+(c[V����r[�� �J�A�36���F���c�Ҵ�v��N���A=�%g��C!�����i�a^?g�/�ʦ��Q햊�V�����'��?�H�Ѡ������fg���U�5�U�x6Dk� �W���zN�ؘ������UY>�}~���K��.��N���p�ފ��;d.1��2�k^���Ch��GO5U*�ʍ�vVI@@
�B����nePSQ��X�2&mY��[�&2I�����zpuxL��y:Y�Zٛ^��=^+�E��]�13�HQ������k)�N��`��dRz�5��<i]A������Ni���*��z	}��1@IJ&ˈ��-V�'
��Ѣס�g-��6Zi#�p���x��n{�^��ֺ�S�ؼ�J��l�s�TСe|��֨Ûs/w	B��fŦ�t�O�Mcul�]�8�]�m��۪:���p:yE�dVՇY��Ǐ��F@J�:�e�z�ɇe	oրq;����B��3*r���5�qiev���]�W�����W�P�?v�~�p���$�
�:�1h&������V1�;|��YXsl�Ƕ��՝4ih	 6��v>5�'��T�Vځ��<n��,\��B�3�����=d�[`d�V�qi2�}R)�P��#W�F��k�^��7!ou*2�*�w5D���n����ID]��˒��Y�"��z�>V�Q�-�H���?_�'��'d�ȶ��������:76({��ja���f�%O���
����y�&7f��N����R7!�Pt�ms����3�M���l���TgC�}g���V���Z����"��8�|=�'k��_�ۗ�w��~����7�H���N�N��>/8�Cb����'���֍����%�܊�z����,�9ѓ�u���1�{�#I��-�V��T��6�ұ�x�(K㓗���ZU��k
ZX�O��0���JW��T�6����1�䬕��&;MY/���.,T�<n�vN ���j՛;�[П�p�/<��ܵ8E��D�!�U�}���/x��!�?أ �u����3����f�\\[L��
���Ƶu9� �gy��%֌��4�����[e��n������V����@-���T*X"�Si��S>J�3��YfB��&ݗ��w3��7E���+h�A����d�z��W+o�GZMfn���I��3�P�V����q�:��m���)��o�k��A��\{�ZBֿ�Z
�>�������2!��F<�X����xUV�K��5�l�����`�N�nf�\�00���f�H�G������+��H��Pu�n�5��5j�q4&~�2�o%
���;����f�І��:�	{��ZS���W� q��,���!���y�4���U_к	��J�k��cM8���ř�P~��Rh6�U>�e��X�l�Ώ�g���.��h�2 �wm�u&E�jf@n�ʨ�J�D�j��0�K�$�
t�q�;�jE%7u��fe�e�����#����ҷՖ.�*����.����>�I,'Rd��b@ɢ���_�iw��Z�A��r����
�"'���Ib2� Y��Z�۬j-�̱ěV�rP�wȱO��/<�y�����
(y����]��ɰ����q��;@X������{!i�4���;�yL�~��(�H&0%��TwU�Ŵ�8&d�CR� xl�s�-��~q����tt �%������\����q�|]nS�)�#�N~��yV��ύ��ȶ����?�# ��ѪA��2��@p�N��en�ǲu��}c"[�!��}��>s�s3F�ΒtJ@�^�k���J�T�>�g�ɺ��մT��dk�b3E�#8xn8ݬ�����5���n�Nvn�����}$;���7t�e~�ǰR��R3��4��˞8g���\CK,`Q��Ĉ�O9���$�����n�A��u����x�Y˥EM��M� DU��j�%��;��L�=��G|��1Ǣ�z�_��5�%�:���.wȀS��X�ܟ�@^�Dџ]!��b~oۧgb1ܳ�jVo�ޅ�C�n����h�&�����h tÒ��1�-4]� m|�V��w�$6���7�7�tI���b�ɬ'	��`�^�"�E3#&�3ΐ���	�˂�}�%b�~��
%�D�;�ʈ�&�M���b�1��jlNL1��,	�]�X�P��a�g�^g�]D������:�>���wd��$�hl��%{VRL�y��=�nMa�W��m�woӫU:n!*AO�nfM��N�]� ɻ��DX7W����,���o�e�7�fD7x�Q���5T4w�f|f꯲0k�Qe@�DYĮ�N&z|E�ç�_eVs��#���c����8,}��}�^�Q��32	y�ǽ.O�[�5}�^�l��0;TY��e�:��b�~_$d�$
�#)�8��;��� �b;�ծ��@*:S\xP3g0#�uav�x�����) a �h�Vԯb��G�����y�+�H��HV�\8��KW"���S�����H@W�r4ޣ�js<�X�Q��Q ?�����u{n�"��nv��6��(,��_6���e����L�[ϴ�p���k��h��2+�^�r�hm�ӷ��	3P�(��rj�%��P$��$�{�Y<R�� �R�-;�:��XN����8��a�K�x���O���#����Е�]g�aO���C�Ե�8�з[�*}\�XT����J��r���Ð�\\��rX�eߋo�X#����C�ް.p3��Ѧ���[�e�$2{;�Z��b?���i��P�M�X��#������<mq����<3�GB�i��	���[mu!%ͧ���%�g�I�Đ�O��@`�!nDP�h���T9HN���P�4Қ]�̷�����V��j6��jCg���5YHS���,��Rd�D��1u���*����y�>��� �z��IUBP;�
�C�c��k�[�C��I		�����,��c9��b�.�lZ8*PK�5��E&A�qL�q��z��\Yү�������% "���.��]$(\R{W�N��mJ��o�@���E�鸺�A���2r�"z�+*�^��ѐ�a
sJThUpa'SFgo�l\6���d���옲o�:�J��g��
7$�Ƣ��͸/H2g�?V���4O �HKm�Zi�}�ͧDZ�V	�l5�`УA�d�A�z�nc�y��xn�_%�0�EJ"3���9\������jI��lp~b(���n2 dz�m`��6�_��ډ��Ϧ�5����Hnjί�,�q䞲�SHm��bᝀg�����8�Ff�ȉ���?%��O�+����j���7r��m������*���Qt��t�tԳb�p��O�K%/��<�b���-XB:�
1���5l���\�êxX3=-��kY����Ւ(0D,��mR��q���Y���I\��)�E�6���Ml�7Yʾ�db��]���� Uk�In���m��$+Ԏ�@�d��Eq峇U(�9Ӓ�t�P�Mˆht;�{���|^i3�ەdLpy�H�Ad����߻����*�(|�ġ&#���I\?�<D������?��c�m��a�C����PM�x�n��=7;͔�U��T�.�U�ta�˞|M�s�AD�Th��hݴ<�Y���n�k��4G��>4@��c��p[Sx��*R���;�:AC���7���П�2�Ԝ�Ig�������]n�à$|؉\;G?S���n��C+!�q�i*1(�h4���'�և3X��l��4 T��<h�4�L��V�)65�?�5�}zֆ�(�{੉Q'���C�!�~ J b��宍nd�����إ��uz|X���M��lH��&}�����~�`�N��Ꝼ���ZSsw/�2��B��h�d���ƨ
V�G�C�VĜY+VI�R�Չ��`6C�:��Po��skm "�<�ἘVd���+Q��b���<������[Û���l��&à�������V�Π��AZ��GE����F��)=��8�ʟ�/|g2�����r�٭W5�RP�uk|J���u�q�X'<ِ���Ha�����[��*Q������xme��D�= �Q1� q�s]�'(�\��mK�l�Y�*E�Ӊ��K�i&�z�ٳF?i}��y���$N�sf6��b�����%ʬ���6��q�r篥��lW��Z���}��t����8{;�C�7Ro1FA�cʦĥr �$��ė)��U������+�?��ͬF�I�x��
��}
�%C��C�P���P>�du��v�
�S�p7����q<^ �
�-�\�@�#u��d38X;���G�~���=?�wQMy�:I	qU�W �AA�X0"�70/Sr5�m�g��t_�)�@3~����q.CG��qts��E	׾�g�&���	l�9y����	L����{��2��^m����6_��"m�3�NT	U�eH�*��mδ�V�K�����G��:j�/��iل���=��a9���<���R����oWoM�g0��<�Ɓ.�}(���0]f�}�N��ǉ���%��+�{r��Ć���zG��y�b���6��WsG������'h�O-{*�'���<{���>�6f���b��q�D��B�?3ǍY"�vn���HC[I��b1��XG�� =��z-����o��D���M�X���^�9OlV����Q��r��u�)1}��(ϴ��"c�2R�T{[9�cƝ��L��"����^%h�}rH���n�j0���͊ż����6_��F��O|�#���C3��}�5�|H1a!
�?G�^��5[��<GXø�A�����Y�����$Lh�]��&��f;�|��^_=�ElrO�DJ��g���<�<[�Z\(���6U�ֶ%R�H��8�Z��	)�a,��Eif��E4��s��@���s�/%j�R�\(W=��ܢ�Y�J2��i�&�$o�lI#wX�6�>�iE���3ƅ]+G.�VX[8�['D�[#rwg�%���g�pԫ�8��&{���2a�ʙ֯Pa�m���I襤��W��j*�!�o�ɛ��M�L��"�攼�O}x!+��1�����iP�>�R�k=�ob�%O��k���yo0�J$3dQ$������q��"��C�7�{+��*���j�FEt_�ޏ6kt�d�\�� ����ԧ	�{ZM�~����m���kQ�پpH�Ʉ��6���:�"gB������x1��)�?�nv�$5�2�;[�u@�V͋����H�G��]9��}Ɨ����c ���I4rKYΆ��rLxA��ɮ磥��L�ky/�	^��e~��ѵL��;��Żh!z#
�qx��>"����l}�[a*V>��8�%hI� cw]�"�Dn��w��$�	Rx:6��$�|�;�T��Ka�@x��q�HϚ���`��ژb��Z�$f̸�uA��"��#��gK�"U#��IQ��3j(��)�� 3U	đ�8�u�B\��j�9�D`�E�Mˀ�Lg��W�O��E��:F�2����L���"N��Y�D�c��0��[��&QX����Ѓ̉�V�&��<�E��yI��1<�z�N���&� e.��U�L�����-�W��mā�����fxV,Ou˙����e3~��oD�&����#�EeVZ�a9�e?�(s��`��z�O?�C;(�BJ�
����)%�y8�x1�.���5���;�.#�Zu
eRC�y�q�d���?o�Z�<ȓ�j�� x���|��'W�zE�����o�2�pk)��r��g?}�A�������wk�.f���w!�z�{�R꘸+Q��#vG�lwW�*�a�ų����$d�}�f�&�I�[trQV&���d'��F�ː��N�x��C2I6�6i^��P�J	}Nv�籘5I�E�"�P����4�=P{���,X$p�`����o��b����U��q�i;�|{ZQ��Ye�UW0
� (���ɲ���,`�h���칪�8�	qto�ODpsG�����檐֎1��8��`�bt���?����D��rh�~��+`&���| �Ѧ
n�F�A�L
�����8����ל��y8�ދ�s�:��?;�1x�Q�WFv�_��6�6h���vչZ��*�U5O	�� �pP��|���&�=ۏw�p?�q#5��_�*U�ڍ7�b�+�Q�>�*E�UU�|+��v��ϺM�~�y�W�K�_!\V5��+8&����~�&�`�+�E�0
���=@���~�7�T�Ag#>�q4gm��E����'� ���Q�ɿQ�$8����������iU��{�H�I~�1�-���,a(�]8�D{d���ǯmWug}�e8�K�rT��ڷ/aGg�|A
��6.��t��|�c��Ǖ�(���r��x%WT8Xm���#r�r%�)z��0ۀR�J�Z�7͒��R�4�Bf#�>�^��%�h�yP�US�?�=�?������t����]�|���y����yg�\�f�X�B^�B��M�)�7QM(-��Un?K���׎�%ͱ����j`�<���`��9��u��j?l�C�� �U,7˝3ȡ[��g�"�_\��1L�w1�$a���B8z�q��j�m��}��7����C��V�6-o�`$O��2����O�j-�T� @A���h	 ,RK�B�Ѿ[�ӝf&#=�c�<Wl���V"{L�Aaiq��J�q1�%+�b�f�)���B{�����d!r���t���I�s0�+�(���y#�%BPg	��K�~��ұ��-1��g����c��!5���/`[ ~�V
�?��a�2~�3�7U�<�T�J&==����<;�7���ǪGC|?�q��Tm����5wU�cdH���[x�P�
Q��o��)�[b��3n�"����b[z�Kx�]�']�	3Wy�q��O��9����}�rry(�����}��V������C��I���B�m(��?�
�x*0���e���)J� Rj����(\�!L��Ϣ8WZU:�3��F���)>R4�>�)��G�{�	^�:+]6+����ӓ��Z�����#����A���i�H�2��4l�D�q��SF(��:�V:$@0������^a^��e�ߏ����	�\�2�ޡ���ݟVOuu�ų���ǾA{Wc1���)�i�z������p�z�Ǽ���xX!��$�9��`Pl��N�x���yT͢/T��G��/��Jwh��K*H�@�c��X�����T��f]
aWr/UmҾ�E���1خ$H��59�˥ń�|D�q`Zn�{�#V߮�{O�8���R�!Xn����+@����hy�x�mh �w����q�t����o��&x�{�v4ť�1X�08�n���Xh̰�ח��:>�"�a�2�U�ޑ�η�:=Zj�6�9}L�3�C���ag@\�<|l#wQ K�K�UC���F4u�R��&5ު���g0Pٖi���[p�[�ԧ�P�2�T��q����zνx04>`ֱ�h?4�A���{��kG��ʁ�9��+۴H]7�,���K��x8�9M��n鯪A;ǰ`i�m��Ģ�L��qz����
J��R�@96�n����41(��]��o����3[PR�GZA�3�!������<$��z�ڇ�;���<�k��u��%iQ�ӔD%N񻦊��S�<(��4iv,��,=�K�O�ʑ�2"�\O�����i�u�x+'߉���aUÛ��X�D�\Qp�H=���}v�n!��".��U8v��)$��"����=;gW�;>&�Etw��/'s5-Uf<#�,P�ٳ.�L�����]j����}�l�6:P`|�:|ѫ�@�g�)��H�E^����D�5f6t`�D�̉E������s% �͠��	�K$�]��x����߿��@�V)*�}��)�u��q�8�Mf�7�~��ܘa���T*��3=ڜ�ma����[�Q ��9!X�'j�c�EK����-`��֮�=uKǗqC$x�7Q4�r�O3�S>	l{�i��Uw���9��Mͣm��u�| xl�~�F���˅g�~>������~�����X�E�	�jO��F�xDZ �_�J��O�
2�����fJ�kU�|���$�ఖ<&+qh��`P�6-��g�W*���q���v�H��di�텏{�����RI�&�!��_��{<d����zV4�꼷4��cY{���tr6��B
ߖ�r1�!��=��(��dm?U򂿎�`�k���!����.��b`�����AL�4��e���A�3���z�, �����j�liѫ�᯴'M�@��U�~�GlU��v�4X�W�4��� ?�ڡ�y�}�fr��`����D�H%�����-��О�cC����h{���G�"��c�oѿO����޲��n#���ZE99;O;OR�[�/�8Z��5�����8�)�>���^����g����ý��=S{ި�j�Fƅ֬p�y4�R��.�-���Լ��>���2GK��}=J"���[�Q�M���]n��0��=4��3�I��p}Ba~I�t�VG?pW�X�&�넵-��5x���h��6�I�g�.�B��F�����>���,_�+8q���uE�����x�	���@�s���,��҄�ݰ�=^�r���n�\N,�nbg��|�=��G�ѥ��% N{���/6W�]H�o�
�_�`�8�>Fz���t��qZc���g>c2���`��q�ʿ����з����U�,�;>/I+�sH��B������Q����NM���ldt�+����q��|�V��g����u,L{����|Z`��;���=����r�/��c_������#7��ߚҞ�q�����!�����\�L�����4)���z�S<hw%���> �[�@��:0}v���͆I�'�Mu���I�~VJz��T��JsD�6AZ}�����{�g"taTD����ǅ
K����y�1�#a�W����O�+�V�m]۷?�Ļ��D����<��pΣ�顭���=��.�/�pY�P%�gqv'����Lbt��u0��O����qQQ�ct� ?�\	��%G��	[�U��xI��	1��Ea:Pm����?2��*�z40���t�����(i�ͥ�n�hĵg�2%j;1�G0�
�o�]乬�3�d��)I��L�9�4�!��DM�#=����;��cg$���/�N�Hd�l�<ĩ�e������� �p����&�j�7p1��̍�j���~��1Ď�VDڇ(((:���U���z��,�M��/'���MEo��"V�"�zWx�j�}9�IY�(��Y�Y���X��?������A^Lb�����c\'%)�=���#d���柟b��<(�'{�ζ��@$����G�l��	��f���S �0�s�T���7����
��*7��&Pè��B�z{2R�^�2��9^�1��cG�5��m˸<�?4��S������Q���D{���]09�u�u��X.A���o�pH�8j3ZK9�婰#�a>��}Z�?�PZ.�jl|��b�;�z�����MR�pJ:5�3ӎ�piK8�݄�����	������8�Q%�J�
�T\�-��qr�����އw3�Tp�����>�[p�Q5�fT���탿�ǿ�	7c�I0�9�Hۭ���X���2傲�A�����4���h��?"�m7��v�C�Y�]�&����%�])����O��p�\���Ɣ��p�AG���|B�Foc?fѻ�(:�!Ң ��2̷�JO��k��Bg�AlO^Ʊǎ��B�>��nT/2FK ��6p&�F��8��+�tR�5e����/C<YV?�Г��� �<U:��_��-�����a�{b�hE�i4�M{���<t�w��-�d��Y"۝�q1�#_���́���c�A<N�������X/߳k���D���VEo`�/�8��?C�
���9z�ǟ	&���&��;Z�@c�_�u���L�j<A��)�/���mŧ�Q���� R�f�ZI���g�gH�E�]~SPm৳��`�q��|���*գ������v��r���V.����)�����N�$���yv:lxw+o���Ͽ����
:(�	\�H��l��.'_���k��tu"�n�xG\�o�� �I.�u���+ҩI���JW��lO�O�p�4�XU������Xy��E��v��m6�EZ=!D��;�|$�n1��Oj���ؾ���U.k�w����$r��{ŬS��C['�Q�ߪAXɼ~�^5��-5h��v�INY�jC�!|����3|�F�VН1<ѐ�1�c&��� _ "�#�Wt�� l�|����i*3�Hm�����]�7hi��� ���1rJ�j\�X|6oXQu$�M#��3��f�xF�y���H����@<�A	����[��,�:�4������i�ʺ�<1�w/�\����YI�t��8��ȧF��Qi�yA��� �
N���&�.P���������Bާ|�M��1죐;�6]<+o8FG�u�K����7��CQyc��i�Y
4�h ��?�����7/�o�} ��Į�A)�������{�$����tG�����blvw��h�:�-{����E��������ޛ$5�t�1:�"��K���}U�QB���9��g��G���|��Q�]D�Y8�h����c���'<�jj�uų�Q\b�����C�$gy3H�����EdVJ*�_UߝZ�L`}��`r���������R���D�KX�S'��L�|�Oq�w=�;����'m��Z+��iM5u��q��]��2��7]�ڹe�}��+���xk���o�R*�#+����PƏ]�&�ڟ�	Zh9$}��j� ��5��ޙ���u��#v�&�Ҡ�E4G�nt� 
����PNt���T�c���HH$tm1C"O��J�����8tJ��If�Co���=fc����x]_J-�do4)Eؐ��ݛk	\0��4�I43R?VM?l�� �/�ߜ�J ������z�<�2l��)��d�m��ˁ��H؟���i��0�Ч�����>-���d]Q��_WX�r`t��[�|�b\ٚц����
	N0J��VDH�D���m��P�)G\�����?���m��U|W�ʭ�����Tq��!S�P� A�"��pN�4m����X�/m���Kx��I-��硂p�'Q��
)(V(�d�,�A��E8��/cXCb�dA�3����aR�9}�7���1��&��:�U�տG��"@�|��n0��l�� �-*�7C�p���βE�$X���\��s�qHtX��D7K����o;&�V�9ISQ�'֫���۹JۢW,����9�T�z����ϡ�+�X�n�A�w��n�����Q����͵V�Y�!�k���ȍ�$�Q�%GN��"�2��hӦ�����f�z�ԫ�∓Ό�UL$����-l�sٚ3^�>
S��J�l���wFsZW�T=����R���rBUĸ^B�bB�� C"9����,�z�ۢ_44���9.�I�tJ�Aq����|���%2�+m�朌�5��N�x���0�Aݗ��4e}j" ��/i�5�)�[�W\LO�i������E�M<Nٔ�CM8��f��#��lM��௙g�À��ܗkk��5�����#_�>��ŨB�(�j�|�R̓��G�?~;ہ���ơC�\9��(1�=kYN(vsf*���hV���Sq���X����Hc$Ot��*�{=�X��{d@��w�<Fd-��Z�.�U��X��F
��Ѹ�e��Q�h�6(�2�H�����p��f<�f�;�	""�4&�/w*�f�]��M��*���\��Rj�hߍF�Hx�+4&�ʎ��:
��X	�n�dZ�J&��bxh� *�5'X�:��b��^����cbtp:$�z��2t�:�o;d�w
;�j>���vN��P0e3��55��!].$uG���e�ψ�v!mý�fRŸsQN���?!�_O����[�� � /O�)>�(���J�@� �no+�d��҄���U/����,�h�C!6 �'�C�4�y���G;ݶn��֨<������в5��zU�*���#4��mֻ�q�G��c��Nm('S�R�:P�"�b�9��C����KL}B���oY�:�ԍT��b8����Q<O]Uf�}�N��Zh�N�4�!����/�������N�֏����Z�ٴi��;�����|�.\ze��c�� ɑ����\�x��##~4��j����_�w�1�G���d��0��0��i%����w��?��^7x��쮶�X|ؓ	1�v�&k;�a���gVO�~��iT�h�%�-UFİjh�{*w�JL���&�y���W�٦t#�G�@w���M=ˈ����CE�Tf�Ȫ�C-7:φ���g�Fы��Y&�仜��G�MDR� ��Â��F7{�Hُ��ɡr�o�T'�Ujl�5za&�b��慚�N�"�츲7�j�#�Nl� p��>z��|�i������Z7S��p���akܰv��#e��h_RwwQg��quo]jr�������S�9���xH���u�3���S欗
�ܕ��Y�]�[�)��HPJ��"�*(�i5��F{s�^�֧[�	��'74@��l�̊��Լ�c��Ĥ 4Ѷ�mH��)	w/�EW�!���Ӣ�Qo�+���!��37WXO��F�Z��;��&%�Z�����h��i��V�n����=��m�O�h �V�
���GF��n�0]�����-$1����4Ɣ�@eG;�Ґ�[����?Y4ke�g��'�D�
0,P�cgfġrhg;�]��fk��Q�4ϲdF�G��Zl�ˑ��L���-���a���b`#[Jju�g6v�zO�����΅@��$�;/�!Gn�yc��Z������H(ɾ b�btcB���A෾����!b̚��Ӎ��֦�#�R��)�~n����*|�qQ^��
��Ѵ�o �0#UG�%�h�vI����}Q��-�-�~�<緉 t?3�޻�.t&��K��sR|�_�����lp%�i��	�d~��uS�l'�7��\' �7W������(_�ېY�t|���ZU0G��T�@>�p"}z�7	.�;�^�}UG��f,��I9��t///�+�s���.����F����~�.�@���53�%g�_H���p2�W�@�$����-TI°D��;�\��׶p|w_�iH' s��b^�kDI(�r��.`��)����˫oj<�)΀�`l}q97`���^��U����%���qɐ/צ9�K�V��RA���3��S_�	��n�-��k$�G1���$���;�;�i�Y�Tz0nZӰ؉j�CEm~�*���� �+��6e�(��W���_����,<��X���C�7���.d�'��|}'�4^v�m�y�3�1��L"�j��|�{+w��VN���v_�Rc�D��
o�f{M���,��/v�"�壐*�p+�u�)M�[#�Q7b��y���nБ�!�.>����K�]>���U�}|�mx�%��α��;^���8t�~#��;���X? E��t��8���* D}E�hE��]l߫���u�ܲ����^˘�� �4 H70���Hk ��yU�����?�s�~����T�I�V��׍�Q��ڸj����B�#͓�|UtU�xbkw��$7�@�.H�����8��E:W�F^���11�> +#�}�~�ƨ�L��;5;)x���-�ݧ�&.�-o�����iF��h=,���t3\���.܍KGjĕ����޳v������=��s�|��KLb`���)�veݦ�x=����L�lk��{�@%4c�g��^�7׼"�%�����e�q���N/��q��1���&�T���<;:���ԇȕ�k��X����&l0�紵M����� �3ȣh��J�)�[�nQޝ��з�O/���S1G�R�+�H'��9�R����)�T���q�48��������F��Ϙ�@s1��p�cN2���	�§�D+^ �@<�PA
*+o�Ľ���}ũ�B�8�z�|N�&�~�gE04���
����(��$�0dx��2 ��'{�q
b���s�j���E�Y��~�O��0�-���^�&J���#��֯���9z�g��5�c)�A�� ��~���-������s1=D��ي`Gm��4�F�X��ʫ�2����*�B�����`0��q�+�����������N_�Z�8/�lt's��Ӻ�.���	DB�+���=�7��r�OM�����*g�	B��_;���4�n<���ffH
ySA�b����ʣV��_:'�6\v��K0��&�=�?��Fa�21���]��>ڕύ�:�lR�;k�\8��<1t�_#�F_�*���U�P}�"�5 w��:���n9W6�C�S�J��,`(��N
9�PU�v
�(6�,~﫺"1`��D��.PmC���²���/l�<%����:͆�ɔ��!b'���qxN�ٸ����ߔ�~��4;�r~���L�@���
�XZ�a`(GE��R(�����sr�A��_&6�9[s��z�p� >�Tu�sj�dJ��>����H�nk*^WPp�������ɡ�Z]�!ߨ����7�q �	hBI|Hv-e=2�y:��5c7~;{7��������Ӣ�1�I�J����Z�]��egi}�&�yN��ݢ?���t��|�N�r�( ~x�R��6ES�8K�HP�:r�cG=i �?�fR�u +�݌]at�x�AI�=���P���0P�ATk����/�Qc�)?M7񄻼�e�׷�R��`-n�Hb��&#n��&�v�^�6@3&HY/N&�7�o���{1&�����B���qxo�ē�k�^/�'��lP:@)2ᱫvjniR��4�w�3.��ty�n��������U�*.�ޞv��|
.��g�B�E�9W�Gy�!B@���^�x��y>���ۃI�?�NS5��(�����gG����퉇o2����,Ef}�W\ck�p?yÍuH�6L�i�H��	
�����@�U��鋇a����Z�4@-	�:�v�!��W;]��%i�HHZ�H,˦�>c:i��9G��!E�g�_p�<�C|A��:f��p��t�%�Ko�='?���Io�e>�S�V�@}#���������vBd���0u���dUIF���&�ڇ�.����e��찖�d��6ԅ�?h��FH�EK��Υ%�߰i�?�@-"�K6ۚ2Z*�8@c0���� �KKo!���P��|�8�slp����dC ���\��p�r�a���LU��%k�
�nv�Q�qJ���7�����@��D�m����D��d�Xɒ�+|�������7"�M��(��vߖ�Se:x[t�j������{dRM���Wvz��\�Ԛ��|L�OX����=�a�M7ʢ��	�L�6m��~AT��drF}� ��:q"@𚣧9����O���k��9����r�`e�ꂺGZx�����>�\-�������1���3Z0aF	!�>���T8cK���"�"#���I�ތ㡲o��!�T-e;�YW��́�ݷ	gl.[r%�V$����2�yk4	����޶>

̈`�����q�᳿QJ*�˭jVD��O� RfÂ�%��	�F����y�::� +�79�`����zD L52kv.u��(eݐɎ4�0���M��̘�=C��G�w_Q�d�22/g�y=
5���~��e���Tca�ǖ�mTed�W�b�UI���.�W�ٓ�ڮ552�:R������jH'3&F� �^i8*���QE�j+����m:������\��Q�<`�S���d��ɶ6y1}�����&�ޗ�ةV�M�L�b\R�#��p�3I:)4�%N�ǝV}����C#���P83��\Ś��Q\�D�/5��<�����Aͻ1�_�'��d!3L��1+��2�Jr�jb����>W�`[�>Z� ��Qkçj�a"�c"��i"շ��B&]�$rn�����7�({.A����ϟ�[ s�FՇ��p�'�i�'�&~���w�,�n�|�9��<Lj�����@���z��z!;e�����v�"F�%��Z` 0�56�[��>�s�!)��A��mh��DW�ݖQ4��Y]ks���H��==hUr���
E���i�v`&�f�� ku����\���G�D@AFľ�P8gZ�{��$'Q¤���_%����9K2���3f�q=�y��
��j�k��N�S�B�Bt�$�h����RF�M����-:Ӱ�G��n���81�q���k�6�=s���L��)���ix$�o1���S�r��~f�@(����n:�@�p>+(�XX0��E	�u0�j�d������ø��qD��V}�l���X?��E�vk�����?c�/�I*��ZY�E�=�ϡ�-�9��;Y 
�pj�9���.��Z����R*D ��ً^Hx�s���8?�m�H��}�A1�����`�%����"l|��#�$��J|g(�9]�*]U��"i�&��xl�-5E�=^�K옏�R.:$:CR8�x�0��ARb�I�s�lr�9M���YV-:2���U%��S�&0U�%��e�x����f��ʉե{��C�Z�j�����Ã�a�Xƈ���m4�/�����7^6x�7:�5��5�=J)<�++48߫�������[�6��4i*�JĎ�o�w���Z}�׽7���I����P!_��to����kޥ��Z�xp�`��Z�>���v����է./&A8>�����L- 3�͇]a���ˬ수[�Zź(�LGp5gN^�ľg�?��F,���x~vo3�U�*��,ė9B۔�Z�x�S�����ѣ�6���n�X���c�L#GG��}A�V����,(�
JL��y=�x�F��΋���	���W���B��Xy�taO�4�Z-)���K���s>��#�jn�����v��7` �'�>SA�ì�t��d���e��j�Y:q.���S�i����?NA�N���$����,h��)7���|���O3�]{#�3K���Y�X��@F��Q� ��y>)���B�5��5F|v����C[^]m%��쓛��dE=��W�Ȏ�(�IV/�PΫ�2!�~]��S4��a�����5	jv�xv��׊�vK/K���z��dq>R�'�DE\L��� ��U�d��Hij�7Ɯ�ı3>Ѫ�M�	�G d*���ӂ�t,��ޤB�"�Y���n}�G���%�%V �B�dJ-����RF���X��Ňw �֌�L�g+f�����>�sH��+�.P�#�)��H&�m�~���g]�&���]�]��{$�����@��0\A��&`�a���B�"(hL�����������\k�$�I�k�>פ���>����21�m���~!�3!��}�,�DD���D��^Ƞ4{����&�
��>c�$����e9V7�w����z���eZ*�ҡPSː�7c�nj:�-n,~w�H�F\\mn��`���F�#�L=l~��d4�j"u���e��ˑ�E'��!��]|[�_,��a����U�|��8u�����tt��^1�^�"(*��9��^�ݶ+�
D2���X���h�^�h9ۦ�.���d���G��q�$�\�~�$���`w�Vͭ���
��Η�?ٰc��{����E��������wR���ÞIY�]���=+ń�3�s�tA�(����Ď��x��ִ��D�ob��i��zV�-%�>�)��4�M#0#�1�h`;+V4��S7V~�\�1ZRo�Ώ{�X���ٵm*�m8��^�O��Hn�88�0�Ƽ?O��q[��I%j^s�9�ozнy��܋��	R�81�Voԟ����?��4��K�$�yw����3_!{>?dh�Y}�2$N�Yz��Mt���8ۃ1����3ނ���(���<��,p0��o��N���$2o� �Lb.X�V�"aB��?�k��� �%����OJdM;���ϔD�jҭH7��0x���\�v�s��c=��R� P�n3��w}�o�_P��H�3�XL���u2T�s3 �U��fz%�2496�ʨ=��-����]�(�y��V��l��G=iȉ����Zm�'����A6w�?�k�q52�-CN����#����v{,`�Sd��d����mV���`<����xq��K��;y$0�H뻽��j�ؤʒf�5�G~�ZA�gr��N�����^~��"�Цp*��G�h����د�y�@�oB�K��1k}�U�~��#lɾP�S3��ʮ�i*OY���o��~{�T�,�w{�� ��lS�\�����B)=�Z�z8��"z+o�ۖ���w�:���}�9��ߑ��pѨ"��n�Ճ�+�=��<=<�����j���]�%�������S����ޓ��%�iDGs�y�	�#�}x��.s���T �~���ua&3�X2/�8�З��i���5�LFz8;���l%�~��o`B*�n�mUzf�r�����Qũ�9lC]��2��91F�rI�����&�5z5)a�����������hK�zi�y�P9g8fxop-$��H�[C�4����?B�-���k;;sewn|����-G;P�7�;�M1 ����ӑ��� DU�h|��H��sN�~��y���R��Q��P�� �Qޥ�����&�m'�Y�!"@��6�mz��B�*&]�(|�@�Ɩ̛2s�J���"��5d���(\��&����������s��e�vO�!�cv��"uڧ"yJ��.�d#q���W��.o��]�Rs�w)$�\_�`&0X�Wcĺh$�w��a��O���[��b(��3s�Q+��)XQ[^�Q]>��W�A�ӓKmʿ�b�#�CZvCC�_����C4e�ҧ[t־\��C��I���~�_�9Kf�ð7ʿ���̱���.
��@�%�n��l�/�eԳ,<�C������So
�"�Ѿ�\��;`��Y�� ��,��#����^��~L�--�_,��ϣ�ou8��\Uffw�iQ7�Yѻa��X^l���1��0@S� � �A�-^�[V�{�Xk���1��V�T���zg�-�L�E�Pp	��k����Ǟ}b�)�r�IU{Оɹ	'^AĤ(ȅ�����U�º��y)�Z�>.kHwAK���E�(��Â���!��K��٘L	`����<y��>-�ܐP�_KF6�1�A�����e|3_쪁��o��2�e[f���8����1Q�
��G��*?E�C 4@���-�-�W���Z`�IQ,�Av��@|�אf��b{��t��M*Q,
�����K��}EO"1|^%o�Ύ�n�<���@h�[NH�Ƶ���佷p)`�9�JbZ*JK�1(>�[?+Z��b6\k�nP�������ee?��Ɛ�-�~�@�o�Y$�+��������^���,��V��J��f�*x	�i�Y����Q3O����ժ:�k�:��oAmr�Z@�����zǆu�;�A�<�4�[�2��D��.ⓞ�]�9;����\�P}=��U�#��o��S)<C bb�4ߑ��=�~�W:�Zr1�������H]ta%�F�Qe,dO<x�`
�-�� �t�����'��P�-y��\^���'1�P����b�a����p�s��ā�x=2R�%LO�x���7%��d��+��.9�$�̺�`ُN!Y��#`�o?���k������9�=#�Z�4^a��U��/6�Glr����������ʭ�A��c�/��Fm�R�����r��xd.����	P���%tP�0)-�^|7�wE/����Tehg���F6��k]�'����̻�S4��vaۄ�����h�'ͬ\*z��}�#�T'j�Ȋb��;uWp����j�"���a��s.�f�U��]�7�P<����9ߣ�- �˧��U�3�\�8(���x"��jX_P\ۍ̙XI�@rj��=�,5u(h�4iٲ8�h�-h@�Y�Į�(��'O4]�-�T���%"~�>�-�BZ��[�,e��D�s���װ}��7K�[^�A2����gfc¬���
�S��,�S��VK3��u�@0��<tٶRL.�`W��JQq����2�W�Xe�@nQA�u��$�r��M�g���d������<���ekr���84�cՉ�ʗR�{��j;Jťp{��t0-��t����R~C�p:��7��x�A����V�h�苒)�[�6|�
�]�慖nXr	�J��<߯�=�D$"��3��Q�R^�*���|��F_�ܩ���@lSQ%�c��G(=�m+gT�����P{1y4򫠨B�ĺ�,�^y��x��Z�3�u*U�����	�`�c@�Kd�5?�o��..���ۘ�T��8/7o�������T:eB��-_����:�|�Z�h�l�I�'Z�p���Y=�ր'z��17@)a��I���ʩ4�_��KĴ
,���aV�4,�OA��B؇�*�p �*k+�����\�w>�D#��1���5>c��Y>��}<�!�֦���3��́cj�P��M)pa�/�V��j�m��TR	��g4v$u�����a����:��2��:9m=`w��A���w���A��~7��f1��*���}jA�|�!_��b������?��1�H��F]Z?�ʹ��\��R(�#�D������&}N�e���W%�؜�
}ho�ƪx}�V�1���=�DU��HÞ�RXSZ�qZ��&�M�K���	0e�|e����0������66���C�\��@�dI`)�D>�yC�<����cKbc	(J��ø��/�{�G�����
Ѳ�z����e�U5ܸ��4�4{X��|�w�0Y��u��ˍJ��ğ_��|a��=c���t1�g���e��TG/�W$����w5��ꎅ�^�c������M�c����6�{)IR�j��[w��쮺ί�7�~�RN��������n*=��(!�u�C@�6�*��M\�W�l*k������Y���\Pf=k���k���(?��8�Ţ) ����s?e5O�г�N�Y,:S��2'�KkkUܓ{����ܚ�h�.���w?���)FvC��v2��\21�*�Y�?�Ke�-�\WD�a��!�� 1���\��*l��L�K��z�"Ќ��K\4�H�T75~�l��֌u�K��l���l��҉���v�aQ�@����Ei<���F�d�w���!��@�t#��#)L �@�����XD)��i�E�xS(��T�	�=����dNh/�R���.I�$��ϺЍֽ-HL�W�ܜ7��X�
K�ڻ���c/�����#v���	�����;M���u7�S͊�E�j~���;K���+�0�'XT�8��q}Y���8d�P����U�9|r쵿 �-b����RZX�ܳ���Ot�̛�]����Ylil�3�Go�(��.�����!�h�ZlS�mf9�Q�$7�^��DGU�6�<t`P�:�Ib�`��+�X��;�(�a	�)k{V �G��`=bl�L�R�p\������@�K�O�`�3��C���EX��P&�>(GMv�+�i���L���ث�(��,T���aK���f�l�^��9TQ�1��]諒Z�S�pԸ�F[�щ;�!Pm�hvz��9+׎��!F|Zz��3)�ĕ��O�:qS���"W�|�������/ `��i�AOR���G%�{�~�v���`�����E-V�R����x��\/�%��K��h]���
�5�Q,kٗ^j�%re7��P��Z݊���]�A�*��D;I�*�%'���?����o�]6�
�q�����7�󎕸/���oy_r�j��*��L���"���r�ī;h������H��K��G�gU��n>�GsWY#�\�p�I�$�Z`lf���N�dL|���@�@u��H����L���$���'�I�4�U�W��b�`��A~^�9�L$���1��PEP���j�#?�����@��ŀ�iR��d�d�����k�y�)���)���m�}u���7��ge��Kg=�_C7X"�#��8�C�t�8?��6�_o�K{�Jޠ��A�m��ε��f�i���Jg�g�0ߘL�5��ɕ�������
p̸ ���A9�O*s����/��<dD!�`��rk\1�o���j��Q��{��U˩%�. @��Ӂ�	��6���B���h*8kW-���/s(K��97����ڨGǐ!�`�ظ��[����	5Z�/Q�s�������H���p;�%U�%�b���b�6��_C�׊�����"����: v�d���@����3?ġ��n�j�wf�~�c#'l�&b�}6�5��R�GRcv����<�;��ޔ�WB2u8��1n>@A1R#Z�>�����欺Q[�%=oV�W�Ɖ���ۨzkؤ]��&��	%�?u� 0H��4�m���C�����x��G�l�*��޻r����  � ���CP���r�"7��lT�CИ�Z49l��$�8!�[9���D��Qv��G=�H�����cCب���o�ݴu��@q�$8'Sh7��	��Sʱ��S��F��#�j�:lU��Dyj8>X�6?[I���Ȟ��,6*i�y�)�v���%���ݳSWN��*���?|��IY �'@HN����H����t0}%�qP[�r4�p�u$���Ĳ��q�aW���gP1�&�#Ɣd1��7c�P
�b!ZI��0��Wj��n;WI>a�W�Tn��0����Dy1���a��� gFˎ!�/;� 8/�;"_�(;�7���p�o��!���x�ǧ��J�"��if1l�,,YxN��A�������FS���JX����ʲ��>�3|�����[lc|�񯸽8%v�V��:`�I� ʤ�$�T�/-m��{�95m_�m��+�=�v>���M�j��~=E��h�;!#*|��ǅp�� ��D��d1]����<��/R�!�H��>�#�?�!gFN��Ҙ���iVҾ���13��n���	�Tʶ.G�#�nJ*�����BX�ε�:�_���k�|N,k`: ��<Hi!$�/�j�-�*��S�+\ck%�I�O��G�\5]J▍:��Y�Bl�D��F(�*ޤ�Q���G:��$��H��)���=iQ3��@j,�5�.f�~�vKD�wH�V7�F�;��������=5��'+���˚7�q��S����ck�dW�2,�����H� ��1�������)3f�缦�@�%I^���,��spW1Z�D������9Vs����)�ᘖQ{l*�qGJ�xRY��9�d��]b:W�|;��2������)M���T�<4/˹���`�Ss�����ƺ}�?�~��pq�lN��?�ԧ�z7�)@'��+k1#
X���P�TU�e~�L��:2�b����(a݋�8���
��`.�5K��@)}�PI/�}Μ
�F���2��sц��[T��C$�tW��� J�N���~P�|�Gٞc �$,O
�ݏ�2H�_\4e)ű.~Ż1XVF� �T��&�H�z�YL�6�H��b'��p�4�ͳ��1�P��Z�p�I���yj�����=�I�-$�ẳl^���݃�� ӏ]��wYXTE�쯥�d��.��ɐ�%8>4�<�~>7�~�O��rA��M5�}.��Ԁ!s�~x��/H��������z���gz&���<#�)��t�7�}<��x�	Ha��>��e�01����) ���+TU���e��F�dYdUl^��O�n�d� y*��G<>�R������H���t_��`ECe�st�6�t�E|�l�v۝�DЉ��J���>}�ֺi�q�V�~�K}1��M�)K�iK�O��<{��r�S�f�:а<�k��+�Μ���7j�b��FeA��Ʋ����
���>p+NAC��j��͛�I�r��(3^���IRmK���ā���i�%i�r��z�ؒO�5.@�jP���&���{`��
���\H�
Y��?Ps��Z����`N0��sW(S�=D�s|���Ձ(���bWt}�^ϟI|����jJ��mؖuX�gCe�~����`c#����rQ�GHX.���_cߤ��%b�@`������6v����Tϻ�+�?�="j�}��@z�]2����Ƽq�/���5��}I���ny�:���+f�?F�3�r��SH��u/N[�c�ā��u��5���*��hK��S�V��S�$�%$��#*�3���R5� �(V���LwE��}�����do!E�o���k�+9oK%׵NW�*\��!/P�r�n��Tb>v�]DI�	C�i]9���/1�9;R�*�����+ǰ�^����-Tś��-Ak�AS.���C:s��f>�f*x5)G�
�
胭������Y�('z�
�Լ���`�y[�@�@zAXБ�&����DǷ1N=����&�'��T,�x�!tr�X��Ҧe��uO~�o�k��8�F9��}$Qs;��A#D��.��^�g�i �=g }����XH Pn�/$�*Q��5��[�{�D1�[� ��)h���B�w��6��X����'x��p�	^�"�#�W��dZ��.l�z�AĬq�X�(�+�|x�p�>�%J�§��\�V\����7�fj�d��EX��6�U��D��_C����g����,t@݇��[m�x�\6�%�6aw}A�	*hu�<��Z�an
��9�<������f�Y�9�S����0c�~B�����~�䅆Y�*(��'�f����z$n�ڽ�w�^�|?����Eh�e�D�m8�+"�7p|��FR'����]�$�N	h��7�fy���t�!�.�$c1A�g��k�YrNg�W��1��H�*^[>�
�$BEN�wfN�2и�j��"��N\߾��
�ߩks��n�I���єh��F�=���v����c��ޢ��pƨ6)�G�1��(8/sѕ��(�+��ɮ��7��<�¡bi�T*�fF�.�m�Ui�"B:���$�eۀ���x�	g�#ڞ'N��*}����w��K��I������_f}Ӽ�ᕇ5h��#;��Z�a�P��4y��$��P��8���	Q<��Ň^�@�u�/��(��C;�a��B;�c��m׆���P�7��0��@i��%ٔ�*�#
^�@�}ֽLo����&o�I�2�K��W�P��=�E5�o���$h�Ԛ�{N�Л 캫�H�ƫ
�4�7�j�D��lT#_���H�,�h���� gO�u����L�%щk\��l�^e��(V�f����î�U���,��w���F�ˀ��� ͷC)����g���͘����z���O�ݬ�9q���%8��Ys�d�����6P�F�\o>��n�����^Tfn��i/M0:��u����H�[n��n�,�]�9��l�d_,ĳ2�f!�9�e��g%(���2���!���@�"�ts��~��)�6^7�ev���77ʏ��D��9y���j-3:cDs����ԛ��QC�j	��d�]ܳS-��?�/��	^���S�=����nw�"jFQ�:�!S.�sK�u�\�FsM9��B��^l͚�1p]��?I�.�_��R1�^�>�E�Q|���D�ŝ-��`0Y��0�3�@	�J�~55�d׉FpuY?��aر� �l�=�o�r0��j@tJo�ˊ� �jA\��ƈ�`�?�����l=R������{T����R�/SaŽq�SQ/Ŏ�'���\K�c�i�#!V\��w��݋��E��#9�B{́d��\��.�}>c���Gm{�1!'���3�����H��VR{/z�F`�Z
���!�u"K��h �a[��c������Z�<9^�+/��@����GK�,�0Ÿ�����$�E&�G���^*���{V�����h�Ej7d�GU>(��r�w�X�_k���JiHd��������se3hfy���9;O�@�'�Fh/�ww����n�Ӕ8�W��s<�4�Z>R�MpoZ���Z�?,t7g�LJ�p��&�UU�4��=�x:�ͲQ�8���u�I�	� �?W�bL�yo�Y�֎}/�R)�"�����H�
^V��g]I/��=bJ��@�YA�QRO��C��Cr��_�N�8����U�W��e�#��,��*����U ;ck��h�E�a��xO�CA�I�h�ǣ͎���c����������o���̝Z�y<���B������ş�;!��tNEccl�i:���Aj*���T���~;ט�>� ��d��w��B������륻��s���\�>=@B�-Q� �H]ぶ��ڳ8�kR���0S�6"�!�;�눖�y,��x���![�E�x9y�&2
h�������D�:ɱc�pS�[�~��Y�&�a�٫��k��Zr�K�(���us��*�f)�F��� ےNH��_ϧW��6�;N�u��p3�P��ZfI����<�榼ee)���=��EӜ]�Hg?t˭�
��>�*��C��4=�,J��C���:�>�Jm/��"��� �uE�gBT���2�*�Y](����T�|��Iu�d.ǻ������q�����o�F�-��Zu��R�p!�A0�{�i�F�X�I%\Any��ʝgCn�7�B��	l�B��'�j.{��j�}��3x��:����k.%Jc���"NV��3-�LĊj��ծ�O�Sk��+C�ҏ��aE;AT|Cb����'��"o�n|�P�;�ʼ���}��fj�{�.]����\�-�`��/���WQp��*^b�\�jͣ�ӂ��K�� �� 
P��x��?�֮Ŷ�wF��1����win�\�$�d!_ˢk��# ��������*V�}9Q��R���|y%BD�N%XB��)5��u�^8�I�pG$�"��qY�2��~�ʂ`n:�ڽ��`x״�q�W<5|����m��gC �����&OX�/��,�7��G�]��ͮ	3���������IC�L3T�U��"�"�^H��h2>�1�4����P�#6��4��@��S;�A���a�F�Z�F�)Aڙ+�+�-�������Md�h��PW昍S�óx�Y��Ԧ�+��j��d�� w�U2�e��N]ﹷ��P?j�$�*�&�1��/].k�4���P=!N�1���%�z)[0Xi�X �k�"���Wq>5��{F��D��"H�-t��7 ��^깻Q��+��T£��)��zה�ލ˭�:`����Z���,��D:4���:�!�̵���%^�� cb���dhH�J�iҬ����P
��W0��x7JN��v#�0�k���\aS��$F���r(�B;l��w��-���a>?w�a�G;�?�����:is���v�R���77�k�&�����c�[�!,�Q7ŀB��m����%� ��)�эC2�k4��q�^W��b�ե^T���D���[|p!s�,��`�ޠFd��ɸƟ���H:��6�Z`Lݗ�#I�X��7�")�U�n���_����5i� �3�Tu��f'Rᒠ�q�Ȟ�ɡ��]���u_\��j��	QA�ܿ����^�/2)\��j�c/��$�$�\5K|t��M�&�5��	��":������"�ys��!�);��K)k���G�
5	Ox��������"�Nߖư<_�vM(j�m���5�i{
�r���hDs��W�q�Y�0��Fci ���g̖*��d��5L����GQ���~L�,�O���$�E@wK�����G/Ub7�B�zԩ"�RKP�i�A��'�AN_��E�IJaY�:���z�_,�u�[ük�W�"=?r_
������rK�G��?�P�ue!?�M�����Bk�M�4 �#��c(��E����ɤ5��u8h%��b�Heeh>{��҉��C�����6���;+�(	#b8NdY����JTs�Y���w�A����±�#��l�~���"w{�N�En�[j$T�oJ�v�DF���&������]���f�^�7�	�4. @�SDKޱ.��sb<�9@j���.k+���w�� A����e����)Y\f|����!�J���ʍ����MEZ1��Y0��������������i���Eo8g	�{=����O�Y����������Z��N���<e�T�p��.�����u1b��0�mC&��"�i����΢�����B`]ٿ���-���#Ǭڸ�����P{HP���s�����t��ǵ���+{��v�A7դz���qm�bf�$�|BArD�S0��}�e��|��d��<��U�=�'=!�5��@�۷�	�-�I���1�%ܤ����$w�ۧER�%WFcor�h�5{�gj��
nEaޘ,f�Aet�Y����t�.���D�����~(���C��(��ĩ���!�O���sTV�<4�b����G���U�5%uF��@	"�@ %����=b�~��{ｇ��ZO�ҋ�33\K�𿤅;~Oun�� a�_����W#=j���iS>��vH*.��ry�7zl���
���j0>}C���,�|]��ވ=�BK��| ���Jؤhӂ!�����5�U8���'p����ױ�ӝ]-���&���l�uhAw�D�j@ɽ����o35�nlO���M�ȕnIeR[�?We�tmv2]2B:s�3P�B&��ٞ�w`ɿrd�M=�M@���s��X������	���eq��=��g�[�������];�I��z�LG�`�̟�q�q���^|�g��ړ��J���| ��D�Mx�)�:Y!R�Ky	S`����[�]������ă��Fa2�@�`�Byd�/�C#�tÉkiup��Kgrm�z��<y�t�Ń6R�Ɛ�k-�y��������s,�8�g�t����kM��1����5Z�ϔ�Ě�K���2�6[	9)��p����_-y)�ر	���{⥊'
�&��%�M�y.�"K� �;S�W (��f�W��-�A,W+�>�D{, x}�6�+~z��\ҫ��GQ��
�Q	Z�8�L�����ymb�u`�����o>���0C�����'�s�܂M@c�����	�|���=+��\D�z7FN�C�����
dV� 4)�J�������I5�l��~�mbF���X�y5\�ϩ��OJ�3�f���H�N��Gri���^��s���J��o����c�j����5X|U��}R"_U!�T���$|�욭�}�l2��,N\��Z�MR������� `���w��.B�&�H���\7r�Ŵ�e�q��]�<�,M�~i�H��x��1f��cH&Y3�*"AUm?+����?3�\�H�Ҧ32R�����uAN(�j��ei����o&�y�MVG�@gv}3i��
��d1��I�p�Կ��BZ�=x�V�sR8'�S��e�l�=(�;��qZ,ɪ���$�*1�L|w�g3Ď�8���L�Tjtʴm5x�.)y,�>Q��
�5�a�k0�u�
o���?����E�Q����CY�V}��e��0�&�X����i��K�_k�:����ɇ^���t�7S����+�?>sܵG�GD��$�+��{��y�AT��Lj��� dm({t��ܿp<��Ţ<vN �fզՙ��� ��}����Ο��.�2��Ta ;A1����su@����Ԣ��2=r��݆�ȇt*j��-S�tn.�D�E���)�I�T�vK뢒'|�]�ֽ��	t��kG���=b�͉">o;+/7L������C�\�W�CHq<W��C�'���cOg2���A��r�t��Ĳ�v��{,����`�>O��>�3��
cyV�*��/Iw-�����I�q���߃Ϗ��3A��p/�Y�3��@�*A����JR� �(�0�mHG���y��)�U��)�"�*���Ng�Ls���C�
'R��Y�uw\����g�J�����"���v��FS�Z'/���Z�Px�Nl�M/#�O���/,�~�`�C�q"eH� �����H*U&e'�q�i[A:��fL(.��%�-ہ�Α���H�
^�p���H6�;l�X�<��������-����$W+�ǩ=�d��p��;�� �3��A
c�2{�6%b!FGT_�k�C狍�������؉�!Bq����K��b2�ۏ�:o�}��B��@Oh��v��:Z���\<T� �XDZ�\�X�rȮ�������ǫ����P^�\���`��">VWx�>���+L��Fr�"n7u�X��d��.��*����
������jD:j]�{�/(��U��2m�BvnlCk�����[����A�4c�M��F `P/I�+A����7n[N��T[[ �Ʊ� ��V�t�Z&%��@�(�t.�+cY;dg	��`=E���u����j��x����賃���j����p���A���]᾽�ew}�X���(Q��-Z�?{*�&Al��T-֯��j���;k-g�6R*�*�����`gB�i�����B;j<����/'�C�N� ɳ�6����Ƥ�l�X�o�d��$L��WJ0���:ė��EyU�vd0�Dp��P�"��7�ul�4NOA_=�\0]���E�+��U�p4����l���8$Vvű!�Ǡc��g�A�B�@�ȍ�;c;�{�J���!����}f1h���f��9�!qc ^�qN��!@�G�!�����6��m��jS{Hp�qN̡�7˛��r�i��"L!"Ӱ�q�O��B�0��������U���0ը�k�!�*@�cow5E.%82�>�������톖V3Ώ�� ������l�S����ݲ�*�G:��Z����k-��p8l���:`w���.OZ~e_�ÂT��uҁ;�$0��]�����?�ms1aD��x��E~�ؗ��>���D6�!���@��|^��&u�J��]ϸ8���Z	���Kvb�G�#ߤɻ���ʔ�3���������>�`���	F���	����x�����b��.����u��#ȩ�v<^%��]�{�=�{�O��}4z�H���1`�0:��������8>��Q���'X���F�'-�wf�|�sڎ���	[�J�d�ә6���7���u.�C`l<�{��!W*���Dz FQ��*X��繀H	����~y��R�|�A8g�rI������'�R��i�����we���TP�e�%1}7BK�@�����,LZ�Ľ��B��>�	{ԟ�e��q�2Ͼ������E��t����1^�f����F)�FDTA.X�6��Y������b�n��[6���Z患c��v��[�E���{�� �i��UY[�o���S,���|��Y�q����.~%-����[o띰������N���¹t \���e#��LF�!��i��V�_�|�Y�Ŏ4A��\"�t�g��O�\�����O�K��x`�1y��uTĝ�l�� ��.��ى�qlu��d[��EZd����i �	�((�-[��EiP��B�·�D�xע����S�4O��P���)�O��<]�|/1I�d��ش	��{z��J	�<A�s����{��z�;��!� �C7�Y�>�c�FB=�gp#M��!E�L�k|�b���͆D����o���?\�W�Q(]2k��N��ګ�lA,�L�S/�7r+�ϗ\�E`wu��ͩ�u1+%kn
J� ��4��5k$D��I�)�Q����wÛ�;���V�Yv��R-���������T�@�q \dN����0p`s���l"�����?�����w�\���0� �k&�]�}v��}��N�3Q�+���p�:���lٶ��^#F����%jk�9E�~�g�J�����)*!�Y����GmkĿ�\	�SY��p�H�k�*vxhX'�{�&V.���ҟo/��"�n��v??S����a!���cF%S�w���z ��C2�����}�?Q�ۭ�~3p���{ޣ�o���8���W�e�ʟ�6��p]�0�2��m�c���T��}~[]f5�?���(�S!Y�=�}Lp�m��,�*��Q4z��R�gmv���wH�g�ddv�c�غ�[&���Ͽ|x��#�>Fm1ů�P���FW.B�k��n�|�^){ .ܱ�L�JN<��*��I��(�G�Й�-�/$�5�-$���Z���N͟��f�\����P����}��z��V����	p���YW#p+�T�����,�ֹ�{�,V��,}��.P�	'�*��|L0	P]�4j����In���1X�x��� �Q��"\w�>$yV٢֤�g��H�B�|��U��Y5S4�v��}����k�ybO�ޮ����B���\��d��m���W�ك;ү+���9}0Ŗ:J蝵�N-#h��\�F��}wD�3G����5��8�{�\-��jM�w�J= �hs)b�tO�y�F"ƹ�q��S�T����dmkq뛝.e2@��:T�	�1�, |���Cx�S�o�ל�.GK�֣G#ͯ:�+��Nn	a �1Q�3�撾wu�>���M0f�$�����:R��v��4�/��a��*�8�RL�L�z2)h���D��I5�녫�_y�t�7-��'��a��8��4�jcL�>�:{ޏ���Z
���G�LR�*�U�RT0��`I�PD�DKW�ݢjc�$�e_�H���,N�!B�&��F!Ų�7��fp��L�@�-mN�����t���AQm��ݼX��L�GVZ:����.����2=xv�h�ٚ[�F��q�z��HC��_S�ȅ
,Q��\3�s^��[�ڡ��{��2P����P��J��ޟ���M���Q74�L-%.��^��� 2��y�W�-�U��H�ީ&Ϝ*>n��]��0�������+��}*����9�`&B��Q8zM��I��j��� ��0�=�
l6��(u�m���	.$%�=!�v�S[���(�f���ހЧb)A�pӼ�ҦN��ڵ���
տ���'���Y%�r7g@�;���k���>��P�l"U���\ly��22��������X)L����wp��$�B�U�O��*[>Z/���)��@�`y�� ��#����W{����3���Z���Jg��k�H���G8W��v܉C�����*�e�&�����P�_ed�t� ��_LN3r��j�t���7�J�5
�_�V�Ue�Ħ��D�#8�F}���JA�kr�$`S��*(�\��M� P����k�x��WD���*^)~��N�!>��c����vc6�OKG͆X dȇ4	ᇭ�	j#�~��d&�5�K�/�y©�� REé�!aS�f�A�A)GZA������~	��E��s���K��Q��,*0��Ŷ�0�A!v�_1��R�nEz��DP��s���Y������~��fr)����4����ӇW�t��)�Q�e �#����P���}�B���HD�c� A�	��6.T�#e����o�5O������e\�o�3zʼ��h;��D)�q[PM���u��5�-uqG?8��wr���i�t�\�������K����Q�rL��})���zh�In��X.�(%����^�%��E�J>?��2���`؞�{��=�ONc����ۉղ���Xm"B=7�.g�����ׁݡl6��~�[!�,�����+��\�Q�9��".X���K�)a�a��?��	�}��J�B����X��,w��]�)�����kZ��Pt���Q�`���!#��46%:�#{�hiJ\������~���SO�Sk���r`}��˶���d��4��KmQ�����%�8�+������SM��L��wW�3��k��
-6d�Oh�Cb4��j[�٧m[_�^��&��e\'�&[��Uc����S΁3��8���"�|3��~q�}O�I��,�����]D����Ge�� `�JU	�0�1r�p��|:?�"66�1b
L�D��`�u�%_��Y�S�C��Z��3;�����ȣ�m�e4m2*�%*�P�}�7bu0N��ɦ?��H�M����k�ޛ��jZ/x�������lW@�"��wa�N�/{���� x���X1��-Z��=8�-�?d�c�2�+��J�L��skQU�G�_k<�:�*��S����Lc`���pw�vk��)v1�߿�]�@�Y�XX:�G{�ώ��5Xa�ώD%����S�9)"l/�غ� �}��P��ֲ^�;����#vrB����	g�a��z�'l�>R>�d%!J��+a��m�H3N�Qs:�1������M��ޑ4�!���U�7Ɉ/z��@Q��%��k��1�ż���$��1DI3�/91�q�J���J����Ұ�q�Q�i�����b=���`�u���¸Y�}')�J0๾��zQ䤧#M #̦*1��/!@q7P�l��T�����>`oׇ���Q�P߽Z��&��$���q�[��~)qe2m���_=�%\�wC�e���z�O ��h����G���Iᴻe����Ij�T�vS ��5���P��/܅�����ɒk��R���jjy������	�A�a�g6��,8W���A�pk|Tl��Ӻ*/m52�[c�I���;%hwAD�x��ȆmD�֦<d́A�0.d
<`�9����)��=�S�dW(ej�~K�a�#�>�O��ȹn�/���@�m�hB 0�������o���������+�
O�x�i(�I��|���		
��O閙���2��ё�*nٮ�Hk��:>7��������2}/M#��×��i>��������#�P���j8^, ]H���]�ȶ�������^ �M�k[��.vB�"�<��/�FJ[�����V1'��1湤uV�HF����D~�-�s��H@avՀu�1���̓h~�A�9�ە$$AG��.��?p!��$��ڴ��d���GV���a�5c��)|��UE|�茗�e����ȹV�<�i����LE �$w�_]�)�ku�����
8P�Z��cԥϧ��������Ji�C�"����W���^w�V`��ʰ�:���a�E^E���Z���N($5з6��b7GéO��N:O�.�DO�>���e-f�
!o�i~_�i���^��_2H�C)�'�*����?ϦG.�N��<q�Q:J����#�r�]�6��2�3�oĽ�ʥ��.�2�w{*��r�9�^|wݝ�9Д`�o�O�Rb�L�UP��Ϗ�����+��Jo>���&����p�·��
OE3��^��-�)JA��e��QI���	%ʃ�=<mG�)��1��&ޕ�"~X�4>%L�X|فy����Ŭ����=I�U4�;zn�/3���v9#?9I@P��gv��K�֋D�`ͨg�<�I�"�&����w�Xv��� Q\��U7��N">?n��=�zr��)�N�$��ϠUrJ#���^68 S�R��;�+#Mz��F��^>�8���
���n�dj���4u��Bg��Lδ'���F�To0�x�%�O��'eO ���g�pP󮷷���:���V�&@=���l��?��"Cm�=�+6�JC�ں����>�\�\X�O���,hӟ���	c�V|��HX'�Y�z�a��*��C�u���'c�0�7o�hs7|0������Ҍ�+��7���7"��k-����8�[ƒ{���2W ���'����ܺ����X��:<�s���![f5F�r|�V����4�����)�>\�	�ӰxoX��G\Z�Nd�W��%�H���k 劐4F��s��l�7��9�ƒd8�"		��u�Q�(�	����j�;!���D�6s���`'p��a���]^x~�A4�I�9�U�1�+�,ݙ6vD��uqUq�U)������J&�њ�����-!<���N�"��@��vA������^�d qH,`V�˨qM~�]+�!�nr�D\�K��=!��T.d�7	M}��V#/��Qq:
���?��ne������}�P0n�ئ�
1��ͳ��@�{��:Ђ�B8w�>��d������_�n �J{��Roj����5�W�����
V\"�������ӺSV2 ~��*�gܹ�y�% �7A�B�9k��Dw)��ԣݴ30Z���n�k��GKE�Mp�`��i����B4b���9�՘3wF�!��z��l[�j�0/1��`��>W<���P{��B1>c�*'F��u��^$�n"���ky������^nb�6ĭBq��I����vQf���%ߖ�B7�C��OǮ�H?�f�.OEP�kb{D��h(A&�Sr!�(��B#�.u����%u�Ц�Y��!��!a�H��R�����Q�u�s��Ƀ��6��g�H��!������Y�h����Mu��<�Ufv�=?��tO�Ή���b�Q��C{��;!g�i���l��x�=瑯�N��5x����:5i�֪lDve���z�E~��)<��t�Wu�y�P�p'��1��9�ZCݧ:C���}��X����Wu�$y�r@mB��ǳ�A~B�<�Q�����[�)S�v���O`rV/�Y�w�lҚ�D����d�R��S���؍�_����3�)q��.˿�0]љ�Q��\�=@0p!%\���`7
w�j�K���-xRv<�j|��8$���N�A�P|d�Dn􈭨��$�Ԣ��EìΤ����r�����b3cV�
s��ɧL��	�>M�n�o�L����>(!�.�˲D(*B�Ã��!�u#]�C��-陲9b������s����D��2ʙ�j,����C��;���92~6�8�쁈��B�R��yf��f�	d��	y�W�(Cp�yq�TQ�(��S(>�k,#U���/���<.��%��M�T�#�i�1Ld���n&I�%ʃ�C�ʔ'���Ҹ=J NcX9\�9�Zg/ �|��}��d�)U�(]-� ?浥ܪZ[�*m0�+x����BޙD�~�XI�c�uXh�a	�̺�m-02���7<	+�/����'T?�W�N���*U�i��G:hq(����,B�+��J&�ӷ�H�?v!�"
�S����E����x� ��lc��4te����?�z��0�x�
�� �'��O_|�F[�c��H�Vi�Dc{�ñ�r�9����|��D�|��d�| ��g8��6�P��d0U:if�����z��M^�3��EB��O�	G����kh�(�G{O{��O��f_�b5����\%h�}�	͹z�I0���69��wCq�u� ��2@g�s������Ì^�R���ˣ�W�@$��w_��s�a��m�
��%�(`����~;q"��n�u�	1�q��j��B�)�w�E"3��+�np�N�����W,�n� ����k�+���t�=��D��9fj�a��A�D|��i]��3Te.7�����}��s��F_g{V���s�tgjjڨB��b��S����7vQ�\�9"�-.��S֎�H����U��a��Jt�� ��o���t^(��3��I?R �=;�VFZs��k}wB7�pǱ�WI�ńS��.H���*�)���� =ש~Z2@�cf�7�[�EQ��)�<�;ݯ��t8�3N����5z�O7m1��,yI���E����}��b�!������H����6vhqܩ`�k��}�E�$���hf�[\���m������F0d�"�B���g��h���̂絞��4+M>C}��q:xK���ۋ�ɊHm�H&j�$K���/��R���dw�gs԰6�{�)� [���V"e����mHmr�j�(�ang��I�G2��i&~�Д���dF��]EB�(�~����;~l��G�y�.x�VR����ؕ��9�CV���[Q�c���~o4;�XJv�IYk���7|!o�U�Ԓ;��j�Y��Pw�� ��,��+pVF�ɼ$�b-ά�ĉ�|�����8	4#Td5���͏"��[��y#0�G�h�Fr�3���/���A�c$��Ԓ��j7�D�Z�D&>��ݥ���yᵻ���u�6�oy�g2�Uy��� ��xX	)���B�	o�9ג
��6�Ef��'����R��q�li(�����[�'uO�ۈ=BdF<�,�VۆH�L�m�N��B�ꋦ�G�)U�+-����;�d��Y�(��ɒj�q�v��AST�h5���o�e;�D`� ��7M�-����pUB�ȩ��#�b��>A�	������Wk�S���G�:��u�ݿE b�D�nuܶ���.�iAz����3nZo9�~ ?��լ̄O�Ǫ*��F�)�c?V�6|��`�%���>�.�s»�S:�2$�Sgq�4��|OZ;�n	R4h�� �f�Y�c�4�|���9���JE21"�Z��@�ص����C�@�O�P�*'���l%�_���(��NתH�h�]}��j�=�-0���.�G�P�8=l)���ஹ.���EL"�l�N�]彃�����Udm]����\�iS�8�%�,��*o��^\�¦��u��֌Q���L��T�su |��oP���\����m�3��R�B9���p�?�w��u�~ 2��:Ee���bHȅr�a\�4$�� �����ښ������/�� ����6ၗ��J �_�co��D��������S��+�& [ 2��D$�t  /�p2iJw�N͘aX+�~���}�Δ�r߆K��0�=��l��F�#�r{���1Fʴ�%[A��g�j1�.rC�׃l#��PC�%�H����ʰe�by��{o�|�e/�E�l�e�S��PBr����m����%b���R�6ˀx*��S�������(��f�������iF`�)�'h�ԯ��y��=Y�@Xp�}�N�1n���v���Ud�y���ێ�~� ��XȪ�$E���!	���W��$��WrP,�p6��"f���b���f3��8FNY0	
�K�W�d��S�#0�,�Q�R���nE��s�^��C]���`l���L⃫Tc��QC�[z����n1��:�=�wص�ަ^�2Zb�b�b�<߅F����;�9O"�1`�s�)*7E�G����zf��h�Ä~7�E[,��<tr�[��o/f�kߘ;H(Km#�n.C��fj+x+�#Ĭ�ցf��FѴz�&����'{��^Z�|�5��x�xX���皍��]�$����	��ߡ�C��JŞ�:����33���ƚ�{mX~Q�W�ϿS�׿:��*��v��d���Z�w2�y�&BQgQ��2�(s�ۀ�!���R�+{~=K�u��OmKX���LǑ������+�����K�/H�J@������	{��$�w�f��	���#�F?��&5ڝ*,8���f�꿭Zщ��	��6�Z �6���U����M�-�������Z&�B�(�qn�7�8��8�h���:�oi��&F�ڜF�Ip�p�G@2��j6�e�di��1�;�]q���,�D(Mv���p����b�3��کl�e����1�j��Sjo]�OX#�'���	��@S%/����V�$��4�>�3 �%O�]q��J�;�*�D̲%-[Uk��dR�/4A������x���GJ�B��%ң0�˹�-y��C����=n�~���5ǌ#��!xzW\lLuJ��Uz*�m�I}ˀ��BG	���n�%(1��j7�Ptq�<���n �E����r�ϋ�I�p1ڕy�x�㣅[�]U� f��Smo���wg���	pc�j����HnȾ�PVoo(^�Z��rbv�}G4��Bޭ4(2Խ�fr�:��~Ϸ$|\�T;~�9��ֳ���wt��1��M�$Ià%�-O=�q*:,�T�~C7�ۏ������x�!��
�t>�%VVM7f�%m:H
�5�U���J`wj>Y!G���E��DC�*��φ3��`�)��M�Ie��5��xp��?5u i�w&Z�ɖ�5k�����u��%p
��� a�g�(��D~\���2+���6z�~=��(��{rz���5VNl ���H2���(=39�.��,M`�X�r��9��)j��iC��'�^y��vw1E��4(CB���6������K �UOiQ*��+g.���Z�c
��G��#�]J���,�,�w��TTBc��r�B�����c!�
x�YEXI���6� O��P�׾�8�Cڠ)� �R��<yZ��֥2U�Y�eaU(߉ȟ� ��V.^𔃋������;�����:�(�;K���h�0�D����=��t�BC������f�ɗ��[�-e��u-�tA���zm)��p8L;BCBtWx�Y�=�>��T gZ4I�Eq�#	w&����=V��I@L�����s�� �l�`�Н�O	��X�]��	�b�{knk'_��`�}Q��M��i��A��������rC1��v!�h,D�e�������^�1�����M�T�W�<�/�Z*�k��o8���4�臿�����A\��ew�Y���������4Q���a����qC{��5�bau����R�u�X���?wث1&-
�w���I�j���U�GL�֛���&��3�0ˌ.˞S)3~L�^����W��%��\2�i�Z�$G��UlO
OVؒH�Ջ��!1*r8��U�͙�X�Mh�o���N�
�z�}8˝�4֗����R+�]�����1� �>��ݘh�"��(5x�iZ,p>#IK���2�� +g���<Juq���
��P��y���la{콺	�u�:
f�FU�^E�H�3��7m��#�6hF���Ǭ���6��E�������G��))�]�F5�%����� k`u/S[U}��W&�>?����9=�p�	^���z�n��J3���Z�,�vP����s�د��P�J����h̒�Bdy*���1uM�:����h��訳6��LQ��!�__��S��C���*�X����)�v2�@���)�>G��؋g��ZF)/L�mp����� �E�i�5�R�Xn-���<��Z�OV���#�����yMx_��|޴FP�b���t�7/�h�^I�R��=yK�5Ԫ���O>����]��*O�6}З��F���}j0�jI�u���qhx�D�l?��U,����'	�助y���g ��E
������EC�>:�ƹ����$c�> @�. ��l44&�~������G��R��bb�އ5�a�T���K4� �ђ�� ���5h�}l��&޷0�2�#,����z�ƒ1�$�ulF5:�V�|����sǺW���mwN�]p�Zj��.x�՘N��
U��B��|����n�ǩob�*|s6�T�(�$��Y��@؂ZQ6y�G�����f����X�sۋ��3NE�����g��ӈੈf�͏���	��W16�m�X�Jv�sR�"w��)���olv��s�ǍaR2��cL��$�9��8�J�;���3�b��E�ҫ�-�kB�I5?L���J��~=Ĺ�`6Bm�'�C;Ycu����i�%��x���W�\
a��bMDHX�e,JY5�t@e���5�����[{h�'�5�^�$���:)��b���58e�t�+S΅{��=��։}Ěl��C�lF�%�l̐f,����F`����MO��+��_�~z��o�p��X~H��(ᮔ�t��l���N��l�k�ӕif6�P�)���`��O�Ћo����o���ߠ�mw�������V���=#V���[[e�M����B�7[�NL���p�0*逴$���BǇ�=je2��.=����6���Xi��,�j6_���X&����x�_��M'��
�>X�q�������F����rw��ck�ay'��T6�A��x >�WVUx��$�LI/�e}Lm�K�gw!�lo�M!y��AV@���4evN&�!���f�~R-��'��C��b��L���s����V�E=�}������x}��GxMęj��B9���! k��ӂ��T��.�:u,Ep�O�4�3 �lI�#^'�8K2�8,꣭]*C��JG|=�)�ġJ���Ւ��jZ�Fm(�YJ���H/��P�[�Q^��'Z#�;j�/5�-1sݙxn����\��Ծr�Ч7�a�|��	 ���M/W�����]4t����)|
v(�kbCd��"��W�1b������������/�,Bllfk��ʘϏni�4l�*���d�W���'����ѝ�����ғ涰���M����ECP ���={EL��N�"����G�-��t)�r��wzo��¿\���K�<��e+��Kf��!P̂�6=S�}�F�����t4�WlG�#$�[�IJf�ڴf���ߒ����%l����!�+�*{���\5���3����Uj׸�
�|��$G�/��$�����+^#�8��r(a?�שo4���Y ��Cd�f��J�����.�H��`��'ܥ�:��7���˹��2j�{:O?��(�C�p��
���?������c��ʫāM(b�a�i5o�ـV�剑<}l������V�l=��@X��*���x�pI�X���{���\uEV��	�Zn��G?�m]����<Z�=Z�Y�h�-���S�  Q�R�<zE�DX�;cm\�0���`��GX�ߔ?f$�Ol������@�q�$+K �1 c�l�n������H��a\'G{؋t��-_�ՊnU더�;a�)]85���8��:�������!C� ��P��cC��.`ZXH1cg(&\k۪��M���z����[��C^�o�7�C�-�fQ���v���I1,	),;��ZV���3���� #^��lX8q[�äq^����L0�f<d�ϯtw��(�*�@6�ޓ|��cR"!�`&S
I��������H��؛"�o����̋�}{\�Zk@�c��5M?x�z��h�'Cf��&?A~@�[[~�%#��n�+|QM��(��^8�B�'��yV~�?ȶO
Q2ǒ����)�rZnh�{�H⾇��)���K��؟�x�O�{�6�IB���n�O��s��PS��6I����&�j�Bu��
��G��ol�s�	�\�u~Y�`�{�zj�4�@H�NOd����)c�a�rܘ�A�fc̙��Y�����课�-��JuL�jY@ �|��뜐�x��(ܘ����Y-lÍ	�I���$�a%�4^� vn������O ��357`�[��5W�TT�tl�˅1g"Y�RG�L��� �?!ջ��<ME��P��ЁPPν�7�N��ym��|��wn���^�Ue5r������;���m=1H��vL�U�KA���j�,�J����.o�ֳW��a�m C�E�'��YUv�y�*�3x�[%8���u"4%�K=D�����<���t`�ho��~���pcu'n�� 3�w���cp�D
<�|	��R'���2~�&cM/��dx�*P����ZCCK<�p:�������":Z�P��ω+�#[POC%ۅmk�y����A�𖵮�)�.J��Kww������ܣ�#� �Z�,����Yᕡ�f3�B�(>�.:)���"N�3�c��x.��z���Y������ �)9=��Iw�����"�;���\����X����{�;u���� Qܡ�R�+�����[����p�S�������b��K�h�����)����>pЩ �3��ǲ�_�\�xT��"��~:��ԁ��]�� D!ڿ>����R3R)7� ��Xw>@��X�^5��X����Vi��<��/�%��e�)k;����`�zf�n���%�}!�gO�C���>��&v�}5���%__	:�rC�W���j����l��^K��~���J����Q�r�\�3r���#�m��f��֔C�8&s	l�%�i0���d��g��X5�y��r���L�G?�����E`,�1�G�����9'Py�Rk5��|�e$��9�d;T�N�I��-�B��������j�i��;��F����	n+1Dec?�K����=عV$�V$��ʦ�q	���`� �Y���{^3�:��#iOr ��H�#�����I\P��X��CT�S��N$9H)-j�`�?v�4g�i*@�l`��u��U�O�� �B$b\�EXC�9�ƕ���t6Yv�:]��ڟK �˗�����ɗ�¼P�1�A���o�:j��U��`Bi�6	���H�bi�u-<�!��[���5 2�N���Kc�U`>bz�7 ���n��?�k��*�����x��FY��՞��rA����:g@�2d�A�}��q�]��$mdC�� t^�j����(	��^  �3q��X�d^�o��lݴ.�gQr�̬:I-�~|���B��f�l�b��d�U#��E�9y~���
*�a�z�})ts�N�<%N:Wm$�5�e='�2�`!�;�{���Pt��u����q|��H�hÓ=A����Ɋ)���f�v*�кYv��d�+,=1��Ip>%)H���aȿ?=,e��M��Y�^*/��,̚�h���j�<�- �d������s�>�U$h3���Y9�'�I��f%3��zV�6՟���%����NMr��x�kw�B!	�������D�S$�����yW�F��,*��v��D^3С�Ջ��V��30�����łT:���0e�˄H��!�!_F9�E,þ���~"�)NT�9Z��X�n��ٵ ��2�V�/��`���AՁS�!�S@�eP@&ץt{��ٕ5>��i-*��f��pnE=?qU���|��A|`7��k�V{h�wN֧�� ϑ���aེ8j����Zǽ��+�bZ|�PJQ�$�;�e��zH�}h���L�/�b3�UH���4V_�oUB��Wf�����|�������c����?�en>'*k�F�Y3�>`���S����z@�X���HՃGF�<^������u��-�v���V Zt�W��H��[ &/�4�Oǥ$%JXe�����5�`O�ՓP�TK%�$S����S�O�
-	���w��$�U�� ��¤g�H�A-z}�=��SP�7_TEd3�q�����-���t�N �"�OV�Еݵ�)H�����D�٫v�����F<(@+����f�\�$���+�fb�?�o^Vab�z!z좜�V�KC�dM��Xr�"Ӊ���]��m=�H_�fh��3y�T�u���E��(n�G
��Q�i�����7�'���yj�0@2��ؐ�FA�"� �8���|�ӥi�k,�/'#i�n����-(�ԫ�v3�];g�V^������|]X��u�tSo���o�X�+,Ͳ��2�-���\K�Z�+:�~�{����_95�����]4�R(�Ntf*�ֵ�����~���Er 'a�Z�#���9b��F�\�[�5���ϓ�YS!�E��u��/O�'���W)*q5�V�4�����}
��5ds r����aFq��@4���BQ^��}u�8�����<ѹ<mΈ�ȩR
n�W	��
��xa(5����'~~Q�PI��u��la��A/�yH$R6�"3/As"M�o�ɤO�f�M�������zjp�X/��|�k��4J�؂���\�㽨d�p�Y��EJ;��l�֞v)�ɵ������.��Sdg�"�On������:ĕy�g*mr[�-HvI^�ʝ���D͗F^�]�~?���g��g@5:�(�B���9��Z2�5�ݢ/�&`y���ӹ��A�.�؎�"#r�� ��	�WO���+��@7���'�������x��S��������h��
�R��[lEE*����#�.(þ�$x�T���a��5 N�7�+��ێWjI��Ae�摚���D��/�b�v���sr:&�7+1Ge��x�*ub"�����P��� �~P���0����#�`��ӿ��;��`X��Yd�G���G��V�k7��z��J����"�Rޭv���vK.�0 V~u�U_S��JͺI� �̡!�m5��ATL�»i�A[��+�
L��7d�k>Fw�Wۂi���x���!�u�������Em,��f��۷F6U�7�	����-e5��,��h��o��]���3hZ����f �,�

��R��R	ΰJ�oC�Aѧm��O�#�[Z��]5
�6K����GJ�s����ۗK��Æ)bh�]蹋q�-�P`A��S=�mv�Q������<�ښ�I&U��2�>��}�#Hs�I2
B��?�c㣖�,!c$�Mg�H�ԫJͧwc�fe��N����_�?�h�_���tiF��#�y���i��=��>�0�o�18w�}��Ws	Dr-5���ʆC8Km2���&�>�	$���dzB�t��ٯ�D���jЅ�"�U��09�_b渽��6$�N.��_$�R�r�78�y\s�E0Px..?j{�;`�W�z5�׭$Z�3oS����x�v�����֍�!f���ƨ���y��nm�`K�A��Ŕ6c,d)�^���3���������X�����ζ�*3�N:L֚ǲ�)N<�.�*���7a��2b�a�=�ɞ(B�!�7:�b�X�JdڣYo2k�o����		sԼ��B ���f�sa��.[����/�_���i�aK�6=��j"b	
,+p_Ռ���MN�ыP�ocj���kw,a�_r]�츎f�-R8(-Ec,vt�!q.z�C�V�~����ڪ�cM��ᜡE�T�1f���NY_Z�G�q���+t��"�}������*�w�Qn���>��s�
����î�ႃ5��#��U$ݙ,�/���P�Vڍ뺷ڹc���#3��i8l��d7�7���l���*��?�ۆ5�^�w��?��	ۡ
%|�-.`D"�V2g�Cq��͵S�Ǔ�YU|� ���}��%R�D�S��֬�FK�#�(�po� ֫z�����ԞG Ǆ�Ж��C�A.�aB'�Cq��#v��`P?�85E�D�+�6�0�0r�@B�k���+0��Se`R�ݟ�K�מ�g�
D��G9��r������(�e�d�I?46������"y�J�ڶ���-sh�L�@hyd�H6t�qq�3'c���
�Rу�����\�{ve@����}��ۦ�wDF1����;�����MAf��FJ}�!��*Wj#m(�q�4~e8������&k��~{�g����U����p)j��|J���7�%�*~ԙ�0����G�U0t�}86�nxF�8kJ�R�r�C�;��r%��5���Q�����w��91�+3�}]̕�\4x��?�$�M��DTr#;���i��[,��\Ԯ`��Y�⥱���|'#o�1_�W���E����qݿ�چ/+�E�56�?��w-�"�oigv+"X<C�l��c�ݸ�gp�}{�yk��*T��+v�/1��6��N��M�C&�&�h�\d	&9���ʙz�uf���>5����#	���]C��F���q�3Qu��mbo�f`��\�`Rǭ���򮺬ޙ�6[�L��\j������\���o*�� T� ;2Rs]����i�?o�M壅��ѝ�w2�|�n���!�â�5�ƃ�(u�o�;�B�
�	�����NO'}��/ׯWEQ�v���9�&+ЖBN�Ot��e�D�pm�^�"G�иW�:���^�V}��I�A�Y3�qV+S�s������Uaz���dԺ0[M�"�To�5�q�|�M>�2m���s03�,�\��[�l���.��-ƨ���A�^N�����#�m1��o�$����B�x"h�� r�H����m�"�#	K��zT��񪵽�"������@��'�E:뻶wI�}�lۿ<;�x���fs��I�_jck�o<������\�����B��r��rZ��Vp��@]��w���l[N5xȯ��,���b��9����A���9o����a�^�7��x�Ǝ<î�!� O ��e�9����C���f�j0�.}��r.QSc��N=My��ac�Ê�iD5TV���N�* �'z�x�5lz�[�bcm��0�V�w����wu2`P%�J������ 9ij���c����ϡ���H�[�E��;�L��q� �:����zch�z�gi��`�����o� ��M�� 6��+��T���1�x���'�K�$�q�Nj�������8�E�d{�c�|Y� h���!y���u:%�����~4�Gs\QU�~�}��K@��RF�Ω[��g*�'*
W��l���@�e�q��H���4��ͮ}����r�' ~O㞷���7�uY��P��<�g��WB�&�ֽ�H;}�b��bT![�DX�Q]������G�^(3{q���2�?����&A"#2Q�@���nD���qԲ��c�V����r?<�����h����ni�DKL}N�x�6NNk����1�|�t����#�����Q2��S��R�6�)�2��ü�1-�ּ�Cq_PE,v6���,�q�Lb�v��R������_{�#�����%h�8����p�+�ir�t�U���I�ur�o��;�)��M���_�o�W����T���ZqL�X<X%�"GVk����;�߉6�uCO�5�R-T�J�t�X6�Jh���X�c��>�F�.�V���߻�$O�ύ9�	5���؛n2�r,n���YB�J�݂W,��W��uD,FJ��oH�"��nl�j��q�
��=+6��q.�H�t�6�MH���r泷O�;�[U�����@��g���#���x1s�;-Tn݅4�!���K�`�ۍL�S|���`�S����C��+zy���+�!��Hx��Sy^�E�����@_c%�?}dC�ޓ�7d�2`޽v5���T+��$�*�_���� ��1�F�r�{!��(��8S�k�{"�uz�u���y��K��!:rqM�!�8�T��Q"(�����@�t�}�(W}�ȏϲ��k�r����n�r��p�Q��T��D��6���=���5��/xjy����T�8{E
���M��7F[8]^^>�3X�S[N�����A�9������_�x��G�kBX�>�o���ֈ��)�>���
���
j��A���կ���-gR��jx^M5�.�W3@�>��h)I���r.S4N�Q�LT��uw%/��3}����|��_1��NGq��S��G�CP5�X���հ���d�!���<�E��9������b0�ŦNLԢe����8��y��|H�2F�W�l�D�kK���N��������%�vh�������i]���ә+��6<u",z����I݈�v���� N����K��Q�R��V�*�U�y�=JY���@g ��d�.$�Ӫn��6�
��v���)�[���쇉���p}��3�������H8z�)�u��z �n&��zտf\��_yY` ��H-���eq��;S�&V�e{� ��sZ�fyF�[W�]�r~*�ܢ�)vG|��]�~_����ڸ��I�?�ٛ.3�{�)e�*]BX1�yAS��\�M��;hj��"�1��%������;IpJ>E��9�R�v�b��`�&�������BN]3��L�S��Yc=�̛��aRٞko$XX��O.�__(�F�j�.��G����t93z��{4ُ�\6�	��=;�_��R����qw��NƜ�oDijV�q".c�9O5;���7�����2��􎫿<*f7��L��͒�\Wt��k�s���%�yK�X4קj��<��c���Na��֔S��S���[f �yU���*�-X@���(��@}f�X��~�^�rثF�|�-�[X%C6P��~����Q!�/.���[���P�H�j��g͐/r�x	xRA��b�� �o�ɝ`�{�s~����F3U����������Y^�f�s7%�E��b�U���MR�ch�3�sf|���&NA���Wq�A�C��%1�<̙�3M(�,jI�8a�����Q�� �G���㩋��&�*JQ�D}��s����p��n�'&���P2 R��eyx�N������6�:�^��1��'��A�c1$Aw��8����3,���NL�]<y�`���俧Ed��)���O.l��MP����A.��H�̗���r�>��ވ�3)E��;��O��-�u�J�D�J+4��UK��D��2���̳Ԥ`�3����Wj�gQهZL�5�<4Og�I�R�~�Ί���<
yI*��[����SƱT�'�c�:O�4d�X��6#�3ū�.��)4nQ��L)_#Y(��w'l0Z�z���L���p���ؑO�)�|×d�>���鵾:w��vt���_Dh�pcy�r�HJ�d������]}���ثU"T��H9��"���@�z�o�DP;)o�Ip�GB��I&��vp�He"Y�&h��3�fP�H4��9����d �d`-kK4���>�zx����q?�����%�����j��'�T8��,�MѿR
H��wQTs��}2?NK�
71��ʤc�1�1:J�6��>��?�Bg8?��dg��l""`���<�>B��Kg�?�w
������˼�kD#���Tw�c[��8��ȳ
�{�Cz�{���c,�{����jl���/GDs}S���o���?��缠���7�O"ݤ{�?n9�U��Ϛ�`�Z�/��?��9.8�<,�}�<�����g/]I?� kb񰔎��Ww/f�����	1AL^�K�ڇP��ʴè0���������s��Xo�������(]������3�[��� �k���R5�o��!fRHo�a�_���|4b��s���uh�7�¦�����&��C�\8=��KЊ���x���P�gv%f|�l~ ��g��^[U�-4R�'�(
?�q���e}��Q�T6t�u�7|j�ǒ��:Fm���u�J�l��itT�X5}k-K��[|�hʇ=$�C���Bqag�M4����,3ӫ�d��ۃ����?�������G^O�U���bs�y�Q�5��/}�"�Ws����&	��,�#�%KB7�{�W(�;F����oj��>����N�<+2������d��e��Q�G;�� v9��pչ:���m	K�;{�a�ig�g�m2��4ޯ~���E�(S76��{��K��z���M�O��X$��'��`��i_�I[P�F�{%�p�k�i��*]�XL�R
hK7�M�QM�iК8ك'��%sZ�Q�����kҒ����d�5M��߹9�q��PQ�fZy1y<3͙(&-����k�&��Q5��V��'���{�dל�E]Y|*3�+@@�Zzη�IfA�I[P~�#М�V\ԫh�����&)�ڭݿA<�#����j8z��OYP�-)��=E<�׻\���R�3�>�{�P�4"F�׏(�׎���P�����-ӷ����%�́ޘ��L���U�\f�L���8�3�/#�����O:YW�8��e�����V��иb���o*R[�`�6�_��i�R���Kډe���1?�K8M5 �-&��r
qoN	��5�7���8����N�q�@˭�z�y���C�x/�T�N���z\�h�$m!nq�Ix�ZV�KBR̄�\��y�w�	�.C@�צc��F�ʻ�	��f��[���C�8��uD�7,� |meD9�}Eޮ�<���*��)ʣX[����*�_���BC�Gd���n��m'?��;�V	\;Nh�����{ku�kE�� 6t����x-b]Å������ף��+���T�X��駛�~@L9�X[�V�,9�o���Uנ�sf��3��$?ei�;���IOk}<( ` ���Z��2�$�?�f����.s�A�]����+�ɪ|���rw���ә�T4�z����Y��������ڣ�C�[u� ���$�ü~���������õ�c���+��nt���#����vDʾ�<U]gw��=����'�'
 �#ӱ\���s�aw>�V)�*kw_һ�"m��Σ�4b�����o�돭#I2I���.0��*n�2L�5�Y��-"/J��X8�D�4�g��:_��4�{���#IV}cƛx'��AV!���?n����R�އ\@����5��;�2�MPb�Q�ç�6��χ�2sk���&��9��>0
�5g8�S�v 8_�+{����͂����ϹQj�ϖ�Q��T�䦨
ISf!C�|��@P ʧ�O2�'���3�iu�8z�&8 >��
�l7��Cp��AKN�	��s���w�x�v��j�0� �P�̻t0I�)Kt�ZQ�������lj����j��ж�����`0ci�V�s���~�f@<���İ��/B�����5���~�t���&O�T�qNs�����Z{?�����E�#� ?���q�q�*�7]R�^w������ä�C�&�a�|uDl[����(��;�N�ƻ� ��߁�(N�����N��7u���B7p�J��$��!�?�t���m�B_��0-P��k�7�-�@�5H���!���F�Eѭ�^�	�+����SL�`SQD-�T��D�&cV�_��_.V�s&P���o"�$���RW���U�t�5����w�
�t��(b7��R���,�,��>qfQ�M��Ik�I	����ԠZ�>�\�>�"���|>򬆧W� ���j@{�#�vu����*��R�W��=��?G��W��P�����&�rO�]��W���fU�G����ad��)��}�n� b9�
,�I�?^�k��:��?� T�p�Z˸쏻/�,�{���q�L�]��W��T������.�jW����'�!�d�"_�L�вUñ���_�;�W2�c��W{7Z�q6hń�i��g�z{�gE�X҅��>fL�o�lO����3�|��l�܍9Rρ=Rܙi]��D����,z�
s  Ry�H�>k�n1�S����ח����TJCP4�CS�������vu��.�#��y�2!%|���gĴ'��%�*B�n��o_4ꋼ6�ͻc9�>X[U��6�r��u�1����;� >H��n[��-vM@ُ2X�B��:oG-���Ύ���M��>��D#��(p��9YG/��whr�/�;H��E��|�̲2�� ��˦~SLƙ]:��/Tp抰�*�&��I�#!�Ȏ��+$/T�ru֔�����J��/���69�;{\X���)A2�<�������fOV����O�rJʄC�D�1�R�.y�l&Z�ϼ�ǡ�i�gEk��R�I�A�=U���S�J p�4iq��� ��\&2�(b�s5��������aoe�>��Ͼ��PLm[ef��:��CR�8�ЪL��f��\��u2L�4�Q�4� �={>�������)��lh\KQA@���IK�mد<lg O�1�o7�;��w��@GV�\��fV��!Tv�3��w���&EPb`��m5��a9R�7��F�MU\/�E"�ע)P/G�3'�F��n�9>���n�������.J�u�(�~.?��!=�+xJ�W�Z�\��M�J�CZy�n7RL��&�n���(j'�����BBw�s��X��P{��~����8��Qsp\��<��?��eu��Vf�Kc�£�
�1�o�JZrh�j5�l�d���E(q��N9D���Ν06�]K�"���7v;cc���=5�� p����.*ӳ{9��L��ǳ/5����T:h�dH��v����Q3��[��ۧť䙹����p=�����>�E7�b�yF�D�!�g7�?� ��ݩ�A�v�DcFJ'E(�V��	#X!���g:�e"t��J�����!�lV�1��<w��~�"Q?��%%��_�Ҝ{�Xx4Q=`G�%��Rt��� �u2ȡ�Ι�����.��U?`V{?��h�aQ3�5��lي�t�G V?q~ǃ����rʶ�]{���Z%���;G�B�H�|B��SA)^����
R�X�Xܞ|��[�e�{Ld�i��}:�a���&8iMCO/R$� 3B�j�uXg��S]�'��)�I�a�W�/B�m(��%�� P��$k�rC+/y�Ŕ3�\�6)��Ro�-�I����!�Q�	�}���cx��53�2IP����tN�W��cE�?����Z�.�\y_9(�[(=� c��S�z�%2{I�9�
;�'&Nӌ�A�"H�4��O���fp$d�{�X�F>��}!�����#^8��fc����4�͔����0�#aߑ���j���
�P�tPa�Mw�+E3"�2ݡص]�7�Y�h��OT�~�����B�R!�T2-��DKN��s&>ʃv���6pWC��S �Q����R�q�?um^ۺl�"V�v��=�L��|�a�����v���'�Ǯq�hlG$c��F/����� �H��A�~/��PF��MAJ%e��1M�ؤQ�����c�n��Rf�p��ߖ���N�e�5��+�E�	��:^J̈��b�Ҟ�E��������q�.�`P��c��RǍG�!�r~��kS4��!*�y�Q����Ȥr���Qϣlm�P*��J�?%(��:���8J�����nT��������x���%}\��A�ʼ�_���F�}�� }#��m�l���VC��ѯ�Q�������d���f/������ۘa�^}`o}��|oR ,�c9�?�A��Ǒ;�I�W��;9,*L{S\B9��>]�dg�]�J0A�M�����؛:�x�m�Z���Hu�Q�T��ڕ'��R�!�P�\�.�;X�Ep�&?x�;_n����jjz�^�����(��<��SoT*3~����ge�W>."ڿ�V�~��.��{�mPߑ�����9f��Au��0֩]�����ۊ�%v0�x&~BZ���9��ؔկ�;��rʞ�>/���%DP�z@ihx��X�6ޠl
���<QP�0~�N'���1�C=�G`��v��z$�����J7Z�O�ҍ���n�'q%�B���o%����
  �F�m�B���#-^×6g�i�z�Y��������@��Ka�WD��&�_�'���a '�/Z�&����N�ȼ{f3p��S��_�����KE�vx�`�w�T�`�1'�]=�_]�j��G2�Tq<�t��5�4I��!��>�\��)N�
{��?o�>Bb?���1����0��ȝ֔���-Ї�UʃmGv��b-�@O8Ҁ;Ld���Τ
8���֭�����sa��
A�#k4���/F�=��E�;/�g����ko5d��>\PL�7
��Lf���COB���ȋ����M�L�Jk`^!e�}a���
���ZFJȝ��XO�s��7n�J�b�����7�5�:�]Ʉh�!����P�;�_ʸ�U��.��-,�����f�_o%G�ǰ��I7�q=���iw4�:x\t��_8�vWy`/�3�<�#�uM�|��
�^�kI{/Z	��{(rc)��$���q�xS�GxOkPMmgQ�|����P� ���wc���ߡ���ŧ�	������~��!5#ǒʊ�9�M'���YU���8��`��K�q�敖�b��B�q�Eu *ɯF����D^��?]����k�Х&BGN���y����{��-��G�b�1�^tb�)Y��D1
W�IGP��d�d���a���M�خw��sq)�b�[E��N �S��~�i�ډ���"��GQ����Ǿ�`�/�
�MP�F���W�ň���;v�$�?��n��A��t�ql6{��U<���[l�zd��c2.���s�'�oA|P^x́�6��6<��mu	D���fO!Ttp~�k\k���l�~<G+�#�&p���)�~c�~4X>�P/�l���m��U�,�(1R�^�R�c>�Z踋�"�N����K���g_FE���$$v�|��k�]F�L�������K�1#���z,�?��C	4!�ߊ[R0��/��.;B�?��������3Mn���epEt��Iz$��̈e�Ց"��3t�5	�El�,�#���֜)�_ʠ��*�#��:���$Q��к�[����[����¾JN�[����w�'�M�lBegR��tl����B"� �Ar���7 ���x(mYV~��:(b�_���K�p(�)�~v�]���8��}�",��U2�g ��z���׈GC�"s�>��M�(S�Ԧ��� �	�!�0�O�}8�ά��sSCaG��|'�V>� 7nL��eJ0��\�I�7,m�%bu&��{S��`��6t����׌�V��ǚ���)ܔ爔�[�ϛ�٩����`�>盄�r�&���b�J�F��t��p�/�ѭ����6i�Ē��g�)'��߈�]M%g�C���l�)�Z�C������"��ҹ���vU�������uߵ�r�C�W��l��v�������y��4�v�۔�� �#�6-ӡ`�y��a���6=��_ڊ��eU�����Ľ��p97I��R�i����*������:h>��k��5_�AEɄ�P��'�!�E靷�����y�nG�\�c�,iot��X7#W����ʮʹ6O�N���
��A�
�����-�Ռ�-!��@�� 4��3�_�R�,�t����m������%K�M��2JN_q�}��n�9t��R@�n�fNp��'��v3�،��Rg�̈́�t�~Bn�@,��{��$M୹�J���Q'D���g47X�^�wY�%�:?K)d5�R��A�b��}���踮�c�j+�WF+�@V���vr�@��FҜ�v�'��K3?�m^Z9�$wM�����	���F'd�Fq�VA;���){v٣/��4���چI�w�-Y̼DT��ć=�.�(PķK�8�H�����(�'��%2*����S��֗ЏM-0�v�\	�JRZ'��H4�Qy����?O4�V7@��'9�kȐ@��pmX��/I�{8���?�H���E�z����%գ'g8�ӭ�Y�ޫ��F��˖jڼQ�R;�V�x���WWj�I~��1�[nl񧩥�23'���f��������N�����D�!�ȃ�.s/QMN����Re�:h��iiT��!�i���zQ�&�k��|Q��X0+�i�υ�-1�0�v��Ha1 ��1�����%~�c�Ym����%6G82����"Y�OPBɁ�U99�*�ũƚu��8��	=�?���p�?rW@F6��2����#����k|_@��V���/0؋�݋\K�i`��k���NBT:��[���w�A�PɄbt�=��P�_&Z��-:��[���VZ������z���rl!����=]l��R������+��l��){P��� u\�se
@A��.��@��^�3�^�w�=q�� &��M��L6��>1���!���� ���s��6��1s�l���\�F~��˙��9E#"���;������F�����کV	���?����X�B�Op Ą j�d�m{���C�WKק�LbA�ɼ��E
�YA6��>��������3T����Wg��5��>%�S -�F?e�w��0zA��������)]C�"�̈gnG�f�����ю��'~�2B�=\�Rh�����0!� #d�{�l��8�9O[z�qƓ��9ɟҳ�Cm��S v�'�='%o�y1��v9Ţ�>��f�,Zs�8X��
r�����.��5r3� ��7Ѥ��k����m	+��&a�A���"�k���}2��~&��QB����tp:��@��P�H�a���1	���:<���8: Y�����t	[���t�G���$���!.4ϥzN��Ň��c��g7췀o��b� c;���:z��i�͕��d�i22��zQN�(�����2�]u��Yh=��5�m+��Ǧ��f]���NN��L�H���
z��dV�/e`1X�7������o�p�ˉT��Nq��{�AG��Y���vgL�^ ��1���H��o����Ch�8���'ɤ`��؍�A��#��g�)em[�(}x��zY��qZ,-ϐ���pQ���7�U�	tES��Ƴ�&F��(�[ŏ%ӭ�A��1��eR�Y�8�Au�jMj�9p���m��j�@��?DNC�a�����X���ט���̡rw�p�]K��w�,k
m:�8���<D?0X����� C ������/�h�B8���넍8���_HmH�"�<�H�.�f��P�H��R2H�}�)����	�q��A��	{���šƸv���C��O���R<x���	��UaE-�׵�{�7����ծ s �^{�n��z�ъ���� ����,�2���閐�����e)�&�Q��A�nT�ۯ���[ ���H/�qg�'W��Q��5t��n�z?�dփ��8Z
[�ఴ�ݒ�IL�}6U��p-vZ ��4�
� 4 ��D���6X��~�Y+Ս*��*���&Ď�F�������%�5���+V�*�	g�?I	��b��!7R��s�̉�Al&����ҿ���f��/Ȯ Mp$e�?��:�%���W&QA��:�KU���q���B�zd+٣߆f�G̴D��W���o5/�`=v\�P��L��uJ�)����~�p"xF�3?����㑕;ڤ=֧*���C�"��8������4���F�2��w�@ƿlؒ�X�(�5=���2MB�����(�a��?T�Zdi(G|IU�Ec���.؞C��-'	l�(Χ�+n��&�h�S�~����ǍɕҰ��A��m�UEb�@Z�WGf�!T�h�X|�	C�Ơ�bĘ�*���hyj�V�iT�	��ZM��A�J�`��e��ٲ7��Ef=S�[u��ٗ�N��
G�<�о�h_$s���5����3C~����N��|Gy��+�v��*���˘�>��]�ru��%�	�@6mV�Ϛu_�5��CEj���c�l��	���?+}*J������7U������G8��D���љ�1҈��:2�Ǐ���T���%�'I��x�	Z�} ����.1��hD2�!ZU�wZ8�n�o���S٠��R�Έyq�2�8����}@�w��7Y�m�i �����R�%:8ǵ�|�5����u���e��ծo'���;)T��j�r�?��]����G0B����C����n�N�Ո�l�#���&@��#U!t��0PǁL6$�2c@`��`KC���1|R���c�
����E�7�hG��#��/7&��BR�����p�f,N�ï��T��O�����7cdK��'��bД���7~я��~�����\��*$&�@�g�lc#����m��l2sʅ��^(�zQ�06��=ch�t���37�~��Z�Y��⸇��U���S��w�J���h�53���Z�~�RњD�O=����`G�9Y�{SB�R�W��qڹE�T8D�����v�w�i<46�kd��}'v-��b�/��R���9*�v����h�6r�)ੵ�O`��O�~�	8��e��:�Y'���ʕ�U�s��m#�
�-x���{N���w����y��?zg�sr��:̃�(��R 9ᥕ�_A�U�0�M8d0����,��/�%�L�6�DQ�
�[�� �7��w�S��+��HI�@U^|�_xͶ����G����D~Oc����^���P��'��RC�%��L�(�Z�c	�n�x:ݵm���J�$��z��=���ic�P�N=�}u
��#��oӑ���T�#N����՞t�2m;��l&��q�c:cX*�\�ǰw�n��:$$�J�K��o���m"Ԑa�	U�#��э:��l�/n����5��
��)�� ,�-"}O����xЛP$�]��ք����Z��o� ѩǰE�x�r*	G������a
k����Jj�6bd�ibq���4'ȶ���wǈ!`��<�]N��o��CFO�Π�_��)�=G�x��")	�<9�@[���L�V�����5o�"��U�+�V-��l�J���9Az�O�ױ`���h[P������G�[���	[�?�Uջg�
�n�5jΉ��<0�n:��T��B8X��|ʤ[np�b���J����s�	�s{��.k<c���es�:��
�-J�����R�����9���u���?�c��QL�-�,�ù=�� N[W{�x���t�:r �_���2���qV�~��rJ��p1]�iK�¹�~|����ZX��5�:@��/Odn#�}�Z�P��
��?po?����p��)t�R.V|`\4���F��3}��m�+�bj�E'=�V���̀����w�ި�����r����q9�{{(���_d��M��XN��w�ݜ�
o�a�Z��q2аq����^���mp�����oK��q4�X�QM<g���I��`3��L�!	/��2
���JGjv1�aV���վc�@��+�V��F��R҄ѝ*(_r�h�Y�31�O� ދ�_堊Z���QP��k���A_��TO_��ּu՛n9����r,����NQ(�����w�V�w��F��H�Tj�N/� ���TAj����-�W��i�:T�V�P8��nŕCH��� �n��I Ş[��D+?�0��v&��>2��E?є���d�"9�����KyBs��ճ~���ײ�y�����%��.�ysN�ͥ÷�3|����o;*�m��V�^"����ha�*s@0�1@i^B�(���#C�3��TlHz�պt�3�I���L2�=�S����0�,����U����5�-��$�n܋0�vZƢ�����v8ؽs�g���}-��žԁ�������Q��ȸ�4��b<G��G>@��^��}�A3.9�z�Ѐ�R~0�(c�F����qR��7���L�lT|q�C�_^�]@#C��]��b	!�R�F4�n�M�����w��+EV�X�B�bܟC�_��N�`�u{D�sX\mT�=�x2���Vj��	�%��L�,7�!v*��Y��07�،)ݰge� �	�w�NX����<n	K���?3����;�Ys{Y\	c��t����ڴ ت.�x0�_��^�Y�� �)��8UWe�L���NPC�t9ɦ`Q�xtT|Rj;|z��*q �Za@f�<m�fO��'�+���E��js@k�Y��f���OH��i1d֣Gr0�,֤���S:�;���>��n&�P�[U(0l�� \�P�F�Z��֔��xw�=^�Rq{���Skj|�������XPy���v�;�qGH�%���&��t�m�l�v��N� 	گR	k�1s�,ˏ�)�^|` Ǘ������MB�&d��hȾ�0�ؾc؀�+���J�wAYv��X�ӳ�e���5f�C�T�{a�$�:d�ۈ���_�Q
���V�w"��:F{��KՃ�Z-�:�ȑ�0�}�pϑ�A_�YB����}�,e6�Q�T^�5��Ȣ�����)rZq>�s��866��y��`�!b�~nUZS������/�v��y�0���N���{!Ic�z�=t�"��4����b��r�NQsQ)S�?�6x���.�p/��*�둬���3��yI�cە��6� �����#��(�nD]���Qe���ej�#�wE(�Lb]޻OJt���[�KV���=�G�W�j�wV�B��6_�O�w��X� ��X�o[ך���8�R��5����ؤ\�|�؉7S�S/;�4���5���1��+R
��7�:\?�|�Y
����Dϻ�?��0�3�Xv���L�v��b�|��2�T�-����&7E�1�*�iد��4$z��ފ�vݜ���ս����H���.�1�Nj������<����#�:�t)���z��76�	���W�W���vx�rq���Zc��,{���qi�y�bLsy�������(�&��oc�ko���@x"ʕ���{1g&3��+aeA�!��|�S�#O��� ��]�Ք�PpJr�ەlq�/��scq�^.j�BY��z!��E�燫�;���叁t�gp��M6@�OM��x���K�ec�u0�mὓq&�DyL�`����e����9�Sd�������;������0ϐ[+/��鐾�6_�k1���H��X�Џ|sd�MDݞ��Gr�Z��*�o����=�ԝ�Q�o�|@�2`���ޡBŖ�g�8TaZ0�1�]���H֡�����1
,a�꽆C:!�hkޜ���/L���k����qA�AS�U�Ʈ=����@`�V�B0}�|�N�BtY�ӏ����j|<�ITE${�Q.eȚ���<xO���fP��O���o�EsV����y㓠ߑ3IF��j�ɾ�B3i���R����I���)���h����1F�_15K�X<Ht�ݒ�O����Q6��M���u�:/&��:0�3�OO��⡾�Zt¥!���0��`�T�>�%\~}��v�|��;e vJ{1�y��爋,潟�B�����^D�ƙT��J�AK��LV�GYŊ��ρ�$��q'��<��$�B��Gſ��l���$�C8EO&\�Ƒq́���;u�^IY��ۄ��b��X. ����F�ݾ�w�m�E)F�Ä
XY^��j{ܢ�J�����aOLuM��Vm�.�m
�{Dܧ��|�PK|�6 �%0�����m�����'�����>����:#E�|�s۳G�?P�]����-�����tF|�֨5LՑ���|���Qi>�t���N�����W)�O��~SU�
�S[8~�⌮�_�a��_f�܊����!L(�pħ���(9\�`ś�?t�q5���,���1�=0r����n�5�=@ϭdO#���[�~�uQ�F�e=D1�|�h�&=�����2Z��J�R߹*<�t�{U���t�o!�0_r�"��X�s��U�8$��#�*�ꇘ�I�ݨp��wڱ2Q4�=����:*����%�bD�zb�b���������)���w��S9�<�-� �����#�\!m���\�Ӿ1��@��G(�ǄB��}rlx<7�8,�4�/[?��N&�}������*{��%}b%y�Ś���џ�\�^7�%9~���8B��@QF��|!����2�=D��� �U�Gڧ�w��a��M� 3>6�����s«����E:/�����<�\U����nZ6�{)��b#X���������_�&}2(�
�lUK��O)$	@U�1�~{�����{}�鉟V�\~:��o����Ƀ8�����cs�l�=�tǯ��2Y���_���!�\0�VG�9~41$TBn2�a	�7�4Ͳ8�H�[=����D=@u}G�5�5�ۍ��Ύ�I��� 4dqo��Z`L�*{�b9;�~U�8=�>4��OȈ�5J��T�Nz�P���}�G�V���Dr�eE+�!~"Y����/��'dc�OOEqb����˞�����w˹�Qթ�=�w%�|�LF%�]@�.����H����]�VX�Q������Žj�Zj�6SX��dJɳ�ͪ�A$7�^r�A��"�_�X�ۇ?|7gM��J
�*lWS��q�K.w?ƅܴ�
�<�[Rw�n����C�Gg��\BYv��sjvͤ 3v�e#�l5�eE���{��ڊ�M
�ui�s���?�0d3�� tD��̂yLg��9�ٟ5N&ܩ���J�@�,j�d�dA��R��� �v�y��� aKQ��{��X,�.o�Z[Ѓ�
��u�\��kr�е5�:���#�����F��Ʊ�Du`�����G���	KVBg#����l�;Ƞ�:�=�h��:��Se��GH=���ʕ��*�P�-)d��h�% ��em���0]h�;�7��\oF��'|�
~��YQ:���sI����E?�I(/��""r0�4S��05�����\��EZ�������?�"�Yƒ"���U�bK}lʲ�U��ȶ����
��hF���I�^0h���ekMas��{��XKV|�<a��H��b�)��O]�5�g'��� �$�!NTg��g�m�w��3�3Q ��:(���W�I�Wp+�gk���L﬎��W��n1f0閄���\q���HC�Se#+�&��?�� �����Lty��i�b��5����2�l�y܊F:�
���9Q� ����1�M���9L,��n͊��b@��9�K����r%��Bװ��zE����O;	q��IH(8�FAW����ݗKP���R1ZK�g
c��A:�/�}F��U$8m�J�U:\��[1q^w��/{�7���~f�V�8�F�g�)!��͊��wT��-ʢ[H���,�7I���V+@>O�XA�V��E0׿_�5� If�4��I2�
�~L�����u������U(vGW�[Q/�.Q k{e]Є�M^�7́l�&��o	�k��X+S� �H�����r��y%�ҹ��|L�������Jː'���J�m���7kVL���x�Т8ɛ$��'�v%�X�}�U�����]8�J�f�P�݊p]]�6�9��bz�c2����?tr�r
��c:����Ƙ:��w�rp�ӕ��)���0E��
�yЄ�%��3���9�7 
<Z�/6��r�o�X��g4(~�P��c���)�״��k�H��x��^�Z�k#�?��*�hf'���f$S��	�Ȫ7NH�<�Ӏ������a�?E�i>i**���e�EuG�iq��r|4�LD��)�����:7��ځ� U�ZWs'�JYˌ��!���ȥ�L�F�������g��EkF��#��Њ��r��.jNs�`͈�+\C�V��0�;�h(�M���U5�	x��ɯ���3���m�c�^���Q�́3LٽFE����q�fa����3���u�<$/t����b[,1/�$9�Ӡ;��	����4�?63y�/�ݵ֫��[�	��F����&�O.��j��������v9��Nd��/	SǱ�D	����~�*�j���-h��Ѐ�`� �ӆ��
>:��X@�=g][s�}-W���gגs�JD��'�6��,�S�7�Bh��r��K��T7
�[i7�t�r��2���Vi-v$�zQ|��W���:M�YE�@]�M ���U�N�e[�/IPa}m�LW�;pJ{a)a�
:	^�C�q``<w�H���\j�r�-��C��j֑��h���୛�^��s �)n��B&�A=�eլ��ɞ�I�}'��uV��"6��Z��N"��v�J�\�L���U2����a��|�iB�hT��3V��ݺ|�x��`��J)��5���J��dO��йzg�y8����Y�o��a�F�1K'���|���x!��MT2��(����n?`d�J����u�N��ބq�SaE�{�؂"F��>f��ȗ���u����;�L��XG4^��a�*J=�'��{'��;�|�!�](УS�L��J܄���Aϣf�b����BX�C=�t[i�L���ڡY��	�k��U���PGqR�n����"��^���[��+�U�9Xf3�18���azx|Zu�t�ey�A�z\�F/G^mn�Y�������)�,�N�!���p�L�&��׵���-���س��F���l��]��j�:��^�y�M��^�6�C�^��!���/�#��l���*������� ���]�R󄿬����/:����7|�R��݋
�u}7]B�"	K�!��^�;TBWK`؈�X0ǥ,��G�C�p�3��:w@H��[�Gh��������� u#')��7�F9E:;� ��L�U���6�!Ē"i$��4�Lc��Jd֛��44Cs-��P�e�E#��qo�/$A �����m������l����av�[Q��Q_$/��ժ�i��71��	]?�õ-6����:>�QkjG��r;o���%�)1	]��%����ƞ�o�7F�G�#U1�}�R���.7�'�S�}}����-��������"�L���}�Ρ�n0���Z2�ILSH���A�=A���?t��D�9���N��9���+�@��L����h7�?s^6������}$>��|�\��iq��,��㨀����d_i��3!��CJ���?�<Ne�sT�g/���|�Y,��!�c��f���ۜT@U���hTCC�+��f�h��~٢���9� v�X�k�,OVL�v#ά�=��vҔ��O�§x9l��N�&l�^���)�Y.㩂r���#n;��bs���69�$����V����4��G+��Hש��y0��tb����0�Q�u�䝤|���ݚ/� R®�&N��� 1�~�P���yC�7���������?�<�a&�Y�.M�4�Af���Zt�����}���܄��)���+�~��M�!���As�^�^p�*���ڄ�\!�c1��`�bM�v��xWv�V�Y$�y|�H
U�#�g��<�9MQ����B����x�)���9��ֶ�S��KG�o �x;�ӻB^�qS�e�;��1S�O$w7��C[`8�*��%��8�	"��#�Ϸ�D_��i������7���U�8~$p�\�\��K ��b)+9/ԁ�1Ig����o�@V������]yy�������E���E����o��=�ɯ�O���}۰�4nL��)`ʙ'^��J`�dG�CC�:��>-�fT�L��������*�.�H|S���ᇞ+SȄo�nE{�4ۏxed�u�aƺw����\��jA��{V�o�XCX�<m[�EC�:��[��+�>,w:t<gK��"��\@`Q�5q�̳��Ɂ�B*Ns�b��,�q�Znb8���@�O������u.g��@䙰Gެ�(��B|Qլ���wG`_͵
��!��ͅlL�����3w��e�v��)�O{��5 �*tM�� �y�w`��%���Fk4�!���L�~�jLa���'�ʻMz5������SjI�^��[���̚Na���b���vײ�@DA���
c3'�����˽ �ub뱞��@BcQ���D���oD������uqF��)G�o�n��cy�yq�h��������%'��ۀ����E,�~�Yᖑ����h^[^��{ҥ� �~�y�8$����x��1��An�h֪,3�Ð�j�	A��<�o���iJ�	yrXg���G$�����٦O�}�t��;���B�1�YK<�<�z36�b�=E06Kn���
�8�[B�]H�X��.*�=�t�WZJSƲ�����p�|�M��:F2�\�i�d���y�Eζ�(��)j���w�Vt;��Yxc������������_6���R屟�����L?�C�0n��	�ªU�u������v,5��lە�ق����$�(��KP8�G�$�h�^��+_�)[|df/嘅�e�|3벰��+Pw
"��d8]���t��*['U%���(�����8��"4J�v��H%�z�c0� t�}�>P훰,����vM��j����ʸ�N�Z'.ߟ~�8��t��ob,���̏��4@H��G�� ��~w�B�b���\1����$W�G����0Xp���@�m�ۮímͯ�z�=e�I�H����>>k���-�����t K�|<Q9ɟ��W�b�JjR��
j��͏��V�B�w��U��=q�� �,����+�Nj�X\�����Ѳ� �ڵ��o�f��Ji%�����4�v�I���%i�S�O;�O9߆q7�LX�������@�r��;�����n���������';������P���/uɧ��Q�^���Z�-j�l+�8���?�/�v#99�>���(AztԄ��t�Ow�Kg�E��<�L�GT���Fh��n���QS�@.����*J`����N~JFv�j��$(k7'Pt4��J�E�4����Ԭ�( Oa[���wk��?=�s�'_�S��cR�K�-�����T��(BC�p+���N�]�^� 1����L�+�r�d;�y�>��eU�� fZ�tB5��yb�Z��w�^F�)�{f��s�;���$�O���(�B���=�'g9�B�߬2]��JQ���X�_.cVrӺ�B���E��K���?�匥�4�|�W���y�"�ߗ��E5x'�T�`R�HC�X�좖�ް~M��x����g2��ɥ��t�@.}�� ��H�0� G}4�i冉��W������`�U��|�X��iD��J|K���@H��i���υ����q�ăumXM��J�|�:����:�%e�S{q����N��Xs��[�m�,y��F1��GLsDX�P�٧d��d><���w&+�k�����w0H�F-���H΋�>Ixs���i�+����<���f�dtYb<�K�6وZO�k��z�1������d�D��>h�_e�(E��)�QjKj1�/���|��)�8mk�[|G�8��鐨d�uy���b���MJ�1a#).*�����6��U'��u���Ș?�e���([�+�i6�Z<�Nj��k�2��;�>��5������c{�.a��ݾN�{��VZ&.렔0�Wj���ΐ������Hhŷwǔ��䩷�iQh��7uB�\*{N��% b�td@i@78��J�T��B�E���]�^�x2Q֏�����l�K��l�0�UAV�y2�oP�i�J��Ƶ�q������?ğ��l�rX�/� �R+�u9��plk��nɴN���� �cg����}ݼ=��T!Q.�eO��R�v��		�~�4ô��7���F
���҈(��̟�/֜��U���v�Lk��;��"�f��y��`�J���$�e#�U�G-*u��$����8o���|�I��� Mʍ�-n��_7�az�)���^(���p�)_�3T��?B��Ǻ������,��z2b�a�B~�{�x5(���1��㤫�bR�@]~w�+�ī�nH���Z���[ȷ/� Y2ci�� h�p�?�������f�׼X��!���v�����JV��˫!�JL#����
��3o����yO�'�5��Mf��R��
�"R�l,+���m�u)�M*�(\��u6�?r��!��'�I�J���E���A��I�I)������(���utx�X�n�U�s��(�R�����	^�a}�� ��jDRm�X��_a-</��A̚u�#u	���n�Zy1L�؃5�ԙ"@�#�r��d�}���$ȷNS���	O������l�h�'�����G|��(�̭������%T��ވ�@ �Fy �w 5{�>e�Q`�����7�&�s�������ۏ��᝹WXZ?3�(�p=��;�M�!��#ߧ����VuH��.Np#���YRm���B����HB�0��6��$�IW^K��n\�������D:v�9�y&�H��l���W{Gj��S%h�v�S?GC�����]��Հނ��j's��c��*�֢�պ�w���kL�;�������^�&o�I�P��h��)Ӑ���d"*�m�6�x������?��p���8�oq���a_�6�bp�t��t��6qL8�VI�����Ė&Z�قi�}�t3;��i�Y��ŀ2�
���_���/礓�s�~�q�e�5��"+h�$|�N�Io�b���ƴ��־��?	�!���ngH�xj�r�h^Y}�� �Q���d�A�5e}���Om'��}2�8�cj�rQ(��Q2���*�H��Wv�3�����\�}��uL"�Z���Lb�l�G`>������M�Kg�gcP!�[����_��y��Poe����{��;�۵b�	��B왱�+�O/����k�=/P�"��CFG�4�ĥF�綃Ŗգ���InU�*(8r�8����W���M4���,9���n�X?�c>�ޝ����<H���@vd�k��piR�~WUb� #����qb��˫��aO���w�P��F���/� ?"[p%�	��!�2s���n<7�i��l���K)���ZV@��ۼ��߻�	���[�(a<Y�q�_hI�<�Ξ`7�C(U��J���B�F<�F��Y�2���y$��:F�����OtԎ��	�ɬ�o��h��M���u8�7�"m�@��"ye�o�_�[�Ź�{[�$��*^�	��F�Ϻ���8/���s�I!�4QW^ST�D�.tt�3/�SQ�U���S�+�!�`��B�r��:�_D^���/�ݮ��q��c)�J�F���]'#xn$#�t�S��پ�X������l?Q,!O�iilJs�u��(~3N�!.%a�d���nR��pA�rB6)�!��H2����^݆տZN�%��/�wW�-�*��\����,	�z��>��h��(������*")S^�|���0��T�E�6&��<��L��3h����`���1P�,����q�����2AN�0���Ҧe��)����yM	��@*^�#ڱ�׏��8_x��j�oAx"^<�����q�w�]%�*L�� &��,A�q'Q\¤����G��6�W])@Z>�~�!0m� ���GU 0������\�e�m[�q 8��W�8P��w�>�^2����w��3!19L9��Dă6��Q*ye9����e�m5G^��Ls���̵��1�Dy�F95���j�r�p��-�u�z�i���\���zt��`H�ӂ�x����f��i2\-�c����q���%��F�YS`)^���E4󎱽$�ak��C����[+D�<(xDn�SiҎkH�i�Δ�F7��nhRW͐p�Hڏ��E�[䴢�}(�c��V��g�!H��ɖOS��D�����d�C������ڼb��Xݛ2pYC����E"���
]2<���Q�˳7l���B1�(�\_�L��'���½T���tH$�з��]���9Scn��Q)�N`�]9��UgX(Ċ�v�x'���]�huCe
�]2�>�i�����B"�`��% �8��ݵp*R[��x:��\��?/�Ma����^�eU4oο�M��!�@��Vi�����l{���g�*i���):��1.G�����]�L�R	��{!r�U��Fn�Up��(j	��-�Y�%ǀ*�򠌀�"T!|f�&��\Z|��-4������i����Z�un ��ճ� ��Q�㖟��$	i_��r��KRm�L59y�W�GB�U㚕���5�P[������c�4t y�72��.{�Wkt'5#]v0z����N��d<�M�7������
<,�~�[�D|ط	�nv�mI�E��)͕��lNi�%5"1���A��,�@3ޖ|�s-�R6�������B���@�`t�#�
�ml�%\��4W�nl�����ۡw�8~a �]��#.������E�s�Gߵ$6P�h0�lQ ;nr�Aj���{a�O���6_�n�7��2���9������_���~�Z����4h� ��� ��`����jy>�$�A$Q�?���$O~���|�X�
%� �M0�u�ۺ���� z[0Q���s��'2{�h���n���=�A\}!ܫ`�wy����`�}r"rL��.��;8`��Q�v�>D���+U�U�[i��3���N�yuYx�DKG�v����P��C����+���ܲv���~��`�oevnh��Jӄ	ܙ9Xf�Vi3�}n'�����4
=J��;�奴�t�e�{���
����9��?�fb)��
����g��os��BY
{�y+�5������#�7(�ά��%Nk�'�v�D_^I��h#z��V/����_j�4��eX�,��-F�KBe�%���vT�&9^�舺i,���XӪ��d��LId��-�Rk��B]�: �E�9����6b�T��g"Hh6_�g�fu�4xe!���)����i[s�C�6�����k�G;\0�޺�AX#Ux�\E;'�U�>a��J�@�@��`��k!Ho~�~�LY�E��̛T�����Ok��T���(/=I#��3������	�(��H������+T�$Rf�F�2��7=*�Rp3؏�
�j�$�,[Q_�h�@� p�b�6��iOM�p���j��+Q��d��e:+�8�k��$�'+Z��S��t'O��j���hO�ڎ�vY��j�������v�V��{v�+-^kGPxjR�ǝ�2�(�yH�r������F�?'>��X�bڰ��kzK�6@�T����1I)Le��ه�N���s�ؾ�����K�	�Tx\��^͓"/.��Jj��5G5Qʿg\8Z[���Z��S|ͩ��VǶZ��H{���p�`346�3]y7��U���WB����}�7��:G:p	u��5- P���R�1jU�i�9��;%D�,�U��1�d������V���(rCףR����E'N�E��(\U�p&$����$�
}S��Gæq��nMF�q��p<�+�)H$��`�N�F��-ߥ����B���F����&�&��=&#�֓Ѡ�nY\��+�BsVbAJ�j�f���U�C7Q��x��4�\��K��l��s��� %p^�)�S"O��ſ����A�3Ωg�%��+bAz�-�h��v�����2�o!����Hq�	D�p����B�>��ѝ"�J�Ja#$b����C
�5ۻ���ĳ���{�2P��a��������!� �E*�^n��C�<�Hdh��>E\*�ȇaz0�v�=x�@����D�����=1A��#m�'�H���m���q�zo�8]��H�Tt����K+36�f�����ƘT�7��ؕ
!�=/�7;/��3�2ڮ���k̈�ٞ�:t�5|��xl:C�	P�#�)]S�i[2$�=�vð-��n� ݧ	X��D�
��ׅ9���GǞ�]`8��ܣs0��	�k�����|�\7^
�����7L��ݦ��ߺ��4r������wk�\m�<�jat�\q��MW�9����0�N��,��9�!6��D?2��I���?��t�|��;�2Zc~��?�T�;u)t��L���K��7aʿQUY����ۆDc�{SB925��4�u�ly�n�Ʌ�)���x�{-�2��ٷt��+����y{o}��x���>~���E�gd2ɴ�t��_�Q����J�|U��կ0A�p�0Hڥ��7��%�ó�
�����$���l��P�\�O�C�3��-AsCi&56M��zL��y�{ d���d�����2)���F,-�I�1c!N��L 'o�΄L瀋�pY7���|B$o<*ؙjs����UF�骬���˵�\�aa!3�y�lx���z_�e)��)=l��#:��R���#�y��xU��#�^��ς(���i0K���췷B�Q����=��X)z�M�@(�����NZ�2$)�x����ls�.�P��T;�.x?Y�l]N7�,Nv����(�Yn󌪅�d��t�a�ˬ���kF��N��EB�toA�U*�=[����Vm��^�1�r�sO[n���V��d�;���}��a d.�U�����t7�s�h��N�8�)6o%�d+���A����#vaa%@���:"n�+C*�B>����.�~�̂�O<��z�#Hzh�IS�.���I��)�:WQ�%��3o�[^��9���Q�V��]�0I��#�z�AY=˦>��<�
8�i�V}�e��ʡ5��V�8��=��wo��-֊��5��:�25I��n8Z�E�4��X;ßFv�[ �v�6�{����B�#D��w�u4�w{���01��� Ǘ $����+���֎�
�x��ʣƹ���!4 �e>�����K"����?�w���q1�9Ӌ��s����u�rdm�$�
�ZĜ�R$ t*u������ǁ3,�Yޱ���]�-q��ϋC��*\/|, �j��@c�=ū��8�B��O���![�1k���	?��K[h�;&��7�#�ϋN�"�!s-�������$�ɪs/E+od��݄g僨֕�~[�K� �t��+NZHxn=I�ig�.�
���
p���zw����%�\i���+�&[�p�ͥAjc m^�$x�,#��h�	o�T�$�"{�@��o�T��䆗�a������4�D,��2��N� D8���<.^�1F�6f�O̬�bd��{���qRG�?|�{u����0"=���Ŀ灲[�����*�[�
9S%�@D����؂��م�茓����UV�@�ƣ�p�8�8h?1��O+cYid{��1��>��o��\�ą�Īԋ����T����7)� �l�Iii==|p��>����?$3k��ժ�^-�Bf�8m�X�����Jr�����:\00��VqP/q�BS^~t�0���J�7^�C�,�8,x����B��a��������XP3�mW|��&��]�M|��~�Hw�c̮�	]U
�a�(����u��F��7l��Y;$W��x�'�C�SA�����[d���g�:�|���ĸ!�WKi��60��}EF��[,�Z�D�L�����Kd�A���~w�E�G�DR����&��$%\�B2�W��'���l��ꁌ r�ͱ?ǰ|�2�Z_jl3!.,�����~y���/q9 vnF�fC4⻚t&��Lݿ��8H�G��nZ��/�b�v�\Ľ�O�
�[܏���J���6�ܨ�T�}��(P�@��~��?����Ι��ǂ��<�XX��J�6A���i�N�2&�¯<��x
�GY�!�p�/��2N�S*-�_�l�T1zk�$�K����x�KM(��F[
E���X�h1/�ʲ���_bx˪.�C�����Z��
c�Ac5�U�b�\H>^�̎�\�Kt�?z:UtF�a�4�3?���h����T�s�(~�u��&'��խ�/���Z��R�y�T�
�?���
�
���eMƗ>��6���2cAk�1�a�eQ��B�Ʌ6��c�րc��kM��6��PL��t�]�K5�8H�,%��]!����i�2c�奅hO/�p���8��Y{_d�����p��$������\wSK��]R훙��J��lk�3�"�CA
H@R�#yK�}��8�lܧXGx��-I����f�]��]'r"l69�c��{�~PA�|�@�������Hߢ:t���f��>P��T��P�<4)���] ��KCd�̿�!:�2�l�c�#D���e��I�L�Y��7��K���<��))�<�^ۑ�Ԥ�Cz����Qt?j��=Dc"�诖O�ޡMtB�fɈ�������u��A�*�׷����)b�t�rA�$LGZ�������^!�o����0�}��|�h�0�;�qڞ8���=3T��x.k�'��xL��R*7�9q6F� ��v����0�����:��u<����"����-/\Ao	���
0��Q�EW|��R�>�� ?4�M�mm�.��B�\����7�)ӏ�nf[��<H��g�HwX�t']<�M�����������Q*$GHl�M�w�Wu��_;�z	��H����`�������ċe��GB��ߒ%�Ï|i�� �bo�E�{~|5�J
�<[��/Lc��=.����n��DP[d�<�$hFt�#z�̛O"=�7�.Z�~��d�����4.$#�̧��^�����j��0�"��UGz�y�]k�J&n��p�,�Q&�SK��U[��v5�nlb��;�[Q�/���օ�2��]�V�H�N���'�~��e�֟�/��	x-p�Q�1U��
���Vg=�S��c�J��ʌ� ��֡���i!�o�n�k}�p�M���Kk��&$����'��3��*ɮ�@��/�͛��������n��������m;��c�&���f����H�$wQ1q7��(�p��3�ZA}p�@+��neAf�l(�c���z����,�,�U����Z���G)}�R�%AT����ޤd�_�����򔚣�$���Ϻ��_w���D�'|j��Q�IR��UO�4SK/#EoAO�&����W�g��xN����mi�R�^����s�(!��J�����$ w"u4�݃�VO�N{����'���](h�O4b_�hL��Dэ�'��7�s��]����e̜r�=!G'A��.3ƪ����pV?�a�u����G�3�`�N%c7B�Fe����?(�f�{��+Jv8!�}dѨ�9w�Y�RLqL���L��U�.���-�ĖW3�#�\G$�"Zؿ`,�� ���Ň��5�����Aq������L����Fz�r����;˙9{� �ÃjU���7��[I�ZL��w�s�G��-2� h�O�O}������A�,�3�FU��?vg�+�B(��?���EI�j�d��d��}���H�8�ʂ��>��aXNu���I�|x&v������S֥���\ܒ�����<�{B[N�1oٓ�?�E[���_�˓�3}@�o\�j_;�SI[�DE�U�Y 0%(&o=yAI���� �S�&O3oIr�&D��c�XCƇ����Z�����:��Z�1*� &��/E��<=���L{K�5�s��Ҙ��ᮣ�=y�y20��K�43JL>A�^����ge�|>�����aHH_�rI(�V�#�xyv1���!3?�B������F����.Sӎ-�n�C��.�1X������*�����%�$6�+:w%J�,,�� ǯ�9��{�Q�f_�&�^�Pr%|�Y~jy#L�b�����Sg��r~N]�7D�y�>�zy���}������z�R����_H�(~�^+�{���@���Os-B�JY��`������,�	è5����l3�;�%����"ż��Bh�Q�&S	�RE� zk���#Jk�!Y�~��{	
�@<(������m}�>�$C���oR0�OC�b 0����������-���w�����ZtF\
E- �P��q��S̢��V�W��I��@v���PUٺ�m~^ٲ�2��ݬg&-l�J�|�3 +"z�%>�_��!��m-�=F���|H/�}t���!��i�bF�% ��!'P�����x�1�&��o_���|�UE/��d�ET���=0C�p���#ڑ���ٝA����4����v����I�G�e������7uA�ޫW���r�!�kU�J�>�۔/�'2@��~K�/����/�v����v���.{��j�V��Ƅ�'�>9l�3�6�a����	*nF܃jT��.�`f�����6���|���"�L�i��0���ɉ����lh2st<���b���=J�k-�E�Yķ+��t,F[e�"h�أ$�	�w3F��V]X:&�g�X��"s���$0j�A&\h���"M�,n��AԺ���G5aTƔ�~�`~��U$R��
�`�U��\�F�֋6�/��W�Us�M@�����-��Ƚ�|Mp84����4�=��uyH_RF-��%�0�[�	6��4^���#K.�/I�D&w�V�kƱ�z��#�$�	TU��ɣR�1gRR��A
E>��<e�cB)p{@����_�ܥ����vO�� N��zHu!���y����5zg��gSH��z�Bփ�c�
 �,�˼I+�BP�5ކ.>�uuCd�%��m�8���Fr2���5�����F:�JZ������[tDƽu O�ӄ`J�_x��攭�p'-�R:X�+�\�}�P����+Z���	�3���J�����,8��{\̈́#��#(����^5�J.h/`�fs�S'E��b" D�I|F��D�vE'B�W��UuI�A�a=�Yoδd+wss�Wg��5�+6�|r/�n)!	����˦�6.�,�L=�R6
�%�4��0�m8�l�+��!�U(T�AXx��E1 ���1ݱ���~H��MciD��<���uo�s����=�k������L"���k�$�%P�
�G��}�=`JtL���Z����2�����$$(π#����i�0�ʜ���A��_���MV�{�<��T�ǖ�g{��@�n~t���*�,��t	�|��<���"i(	
r�g)���؏c:�3��y�4:��z�Q����Ȩ,���\��xx^��~�b^���R{&�����1�Fy8��bU����eL3����l����O�j��v�Ybp	�#��n@�:��RP��<��M #�u?[l���y�j�c�2���̜�ݪ�*��%��8K7�NU���)�1���q{�u��,�������7�)���O�D�S� ���F��'�Jg?�Q�n������*[�����K#�?NQ�lpH7��&n�f[�%:�3գK�qlG���"��Bh�ϦY���r�d��Ĥ�ᙰ)3�W�F�����3��95��Wf�iN��ߑ�x�V��13q�.���hٽ(�s	��ʎ78g��Bu������#��O^��a S�� ��qIc���ݧ������#p��jլ݈�/��cd)�������.A��R���-�����>(?��Jud�郐�!��2(��/�Y�)��-MLW3��489����ےv�������Fw���^sv*dfGM����&{ժ�)� �0�}H�u�Ȟ� �]ZC,�>Q?g�M����
^;ф\&vdv)�k�^c�3�k�ۃ\�;�6S�>�дH$�Ȯ�-�'��� �T����V~_��0�n�lK��������<^��H�y��bQ�*��B�g�7#U���r�m���o	�Ē��x�>+���wl��A��GA��dMi��v���d!/)O��2r�*�����0? ����nbϏy�%ȑP�l���-6������	��bx'h�b��b>�����0�@$�f�5՘Ԩv�
o��U@�, j��}�_�z����/v4�Ӳr��:Ey�FM�B��|���$�2J=���G1~hنp<��-:�~Q���hAC� lX���S%�,��k��SL�७9��G���_�DY�0輔�OmHSR.�AW>�Lw֯�C���[ ���SȻ�4�>_�<���}v��n��uf�^�W
v��w'X�'�(�EQ>�wN"6m<_��q��ϊ�����K�8Z�_6��]����=f:K�Ҋ�S�ṌoF��@��U��	m��oS����l	�b5���?��If�s��&�t��>��(1J�XE
�;<���wN��~���28e9����!��Ue1'wg��7�ts�0C�|)}����Q؜^��`feJ6�-
����ZcW�@�B�<p��[�NکOK�k�����<�~�<_��s�UW?����l�V��M���S@�>O��H�}�e��^d�������_��{/c��qm�-E��,�ņ�\�;ȸ��s�G��)<I�m�i�s\30"D޵L񅪇�~�`ɐM]t`�o�m+K�W&r@<�u��{�O�;�M�z�mwR���������oe��Ǣ��½����ע�U�h�gf�$z����G�]S5�I�B�҃]KEM4�tP|�vx�T�1y@�Q� �I���K��~�M�e��v8g��s*���sS#}K ��P��,V�I�(n��#EXNk-R�bU�%�dL��́��\@��=[ !k8a�����I�}��o��#Đ6�p2�}ӂ�찊`��_0wO#{qf|��Z���p�4)��u}4"�$��A�%�EӥN�c���=ƭ�����.)�p�~!���ϡ����l�`�U��@��<�-<�R���l��vD�)県#���[�������|����/��,�-dQ=*N���f��lg	��m�����'�OqI^�=�k���;�6�ˀm�" �z�d�[�s|����3�LswL'�O���EUD�~Qɲ��|�=�����łq&ƚ�G��%�p?���^]�3x��}����n.-"��[�����{�J�����ľ[�����Γ�l�M�5��ʒ2>��h����Cn}�Jc#��w�Y#��3~�
<�� ƿyq~��%���� ��,��	���泝���yDO�J��-���<#�ȣ�Hl�\�T���dh����} �{;���d闑�0��p��x@�'/J|0{�Tn�����-��Oe��=Q�kɦ6 𾒥X��%�5e���,�2�/�߇���Ub�O�rxp�C�̯S����=�0�橚��}pa)�M����(<|��G2.���4�~��фJ{<����Z�#/��݅]ݲ��\�5i��T[��07�0�,��7Mf@*�?Q8����z3_${F�:(�
�����g��"���NΥ�.	@o"ᵓ�<=�.�"���_�����%A-
b�jM��GJXh�kiy���_�^b6��	�H�����Z�p��k#�� �<�^�z1��l-O��Ҙ�Y� �'iR���Xe<#^q�ct"��|�^B�=x�Y��������<���κ��c�F!������ �����wz���Z��ϖo?���o=�ђ�;�5����U���0t��r���K���ny����J��"uI�����b]�ڞ�#��gNgu]�9&�ɜ8���/�����k�֨c��"�.�J?�y:�a΢�ГC���}S��� J,̈b򉃐[�pS���#��x���&t��"2|_R�����J�u��Z%hǯL�*]����U��$ �> ASǃ$�%��wq�mP����o���=���c�H�scrD�5K���DȽ���{��x9�M����#�@� +iQ4��U��N�EǞ�����+i(8�����ƿk��wx"`�ON A:
@��18�w��x)��F���t^MV���!զ�Dn���f�|'������bD弅���#��m�*��^ڐr����N�3A;��/�&Q�VPl�65~�;ޣ������ۃ4%yG�����B����*]�u��wŵ.V��4�;y��x.-�J0�#F��,i����x�{kaG���n�<JoZ��8K`�W���;�{����^RVP'.Y��@�R��d1=�r��8��q_���j��T�a-*�_2M�?F�0̿l�;�1���s�1U+q2�uD����P��߫�y��\��T� ���+�qP���F�k����8�c�)z�&ō�,/�/��R�_%�d6��Ϸ��@��5��H�u�S8V��Z��&�H`1������Z�;x�D�����*��\��}�i�#J0Z7���a�T�"�D	h9�8��Ni�s����3$�|��N�,����(-A�{���^b�Ku���§p��[�9.H��A�kֿ\���J���a�$G���Σ��o�������D`�)M��7/7��;��"P��F�)5A�}ƅ`�\���� Z|U��� %ƌ���;]%vp1���Cj��i*@'�t��Y���;/y�^��vО� ����ݴ����J�S����C(�aKf�ӣ�X91�4.Cnn���u���`�J��w#�C�?���'�VѺ�;
�Ѩ��S���C9�܍����Е%-3e�
Q�E�z��*aP����'�'�C|o���i�g�A@v%�!2aL[�n�P��ś�
�P��=��WRrc���0���H#��{, ������,S����Wզ:�V���:f?�ak[*�"�6)��|�}���e������$6�#��`F9d/+QD��ՐʦZP�	,���,��(�/��������W���ɦ^~P6���r������ӎ�c3��5�?mj�H�g�T�w~n5�?ci�����D�=�����tIxH�{ �?��w7�!6T�D�$#�F<�w��?ͱ�hL��M��.W�����7R Aw`�k�ْ1A�C8x�z�w��s����ͽ���~�p�#?/�0������X&��6r�h�(*~�0�U;��՜pE_`,����&(x�1M���#"�-6\jсdU�l�]ܭ�Q�D����>��d���ׇ�Ls�γ3���d�QJX\�O��������#*�������"jՓ:wy�N��cGjbu�E���:��L�WXs�ۛ���`��쾽 INL���%E��D��G����B��g�tF�X��@o	�eIQ]�����R���l�5�y�����%��ȷgQ�����b:w�M�K�%4�耫��b�8�z
�X{r!�]��E���i�^��g�# ԥN�k���L�<��p�O���]�%n�2�]g�8�Y˦���P��Ecr�tha*l��=��ot`8>_�M߆�491�(��,9U%}�@������S'(�iٿ�P\�V��ތP��*r,Xr��./���P�]c����ްK�C�B��_�_�.vF��v��B��@�W�dDq\3�#��UY5~{C΃�kZ�h�]��aTR'�������Y�x����peY��s������qZ����ymB���&��T�6���Ƅ�N�]?n��Q��Ϻ�ccH$#eP�q�M�d�XC�ؾ��?�y�[W2��;?&���ĎQ�9��U�UM*�k(+�C5rя�~�.U1���J����7�9mi��9U�?S��}�M��|�2��ay`X��y�#���֤���zkT�9Q�ZZ�My��=��(��#�d�@M�Oׂ)�?��r쟱�jn�$��� �t0[�.��}�31"?�V�@�Ѭx�q��R�44��3���#.����@���ܖ����$�(~���e�����#~:RAqgZ�)M�/14�MҭU���w|���Aj�� ~�s&z�D�q���];^�7��3~�ℱ���%R:�tT���5����O��8�2����J�tm��S�?D[�|�\Y�'�����˟20>j�m*�&ۇ�F�<)�"Ux�W[�bK��pg��{W�Hj���q�@M���z7b�������r��HY�H詒Ȃ�6]��qNJ�us餦7�
S��
�o����L�Z&�M|���%�0T��Ñ���y �����x���\<N�o���b�w$��{Y������q���4�H��ځ�J���hٖ67K|^Oؾ�����p����l��w�W���mm�5����3>��ĊVo?�lM^�R/���M @'a$�1��o�.����.}��������Oo��OT}��������l��>F5�r�v��?���0)T�=7P�!�֍x���H��K��� 0��il��D}����u��캙:ӓ��U�N����=�|Yv���.�f�n���D�ܖ�9<�$���8i���?�� �-x�� �BrK���� 1:�ʢ����BƢ�B��&�umF2�X�K0�Ƣ�\��7����l�6+�%ao�s-��!�j�-�!��(�1S���Z=9�f�/�]����1pgz��ߛ'�G`[uh9p�ȧ�Ѥ�/&����Ԕ'H�N!%��ʰϙ!�qG�EF��K �M��s2��o�5���uv�R���F�5���**eS��;�W��$��[�{���=#$�BcZ���ڰ�߄Q��Y�	B��������6�k�9h��� �bZ� �9%���®����P��x��w�~>�v������Լ�H7����E����z5�ۋ^�	|��4$�j3�Ă�<[����G�]�@m.�9���(h/N�w�/��T>Wq	����~�}H �����x�	�L�㹌�����Ъ떤�xx��2���c�x���Yr��w0���^%�/ѝ3����eUȡ��,����jn8���L�Ws흕���E?4ț�ټ���s�=�;�������FQ��}��1���YD,�r��y��ǿ:'�D&nh�Zz���	�14��Dl
��@Vٽu$C;�hx'����9��wWG�
둔�T��S��&�Xu4��g���Ex�۟X���@9ןkB�:��26��ȴVS���>�ﰓ�0�2���m7 �� �gA^h ��s�z���f�\K�d�5���A�s��Y�T�E�B�l�H��#(�%�G]�u��Q�LF���v�Y�F7���H�zT��@�����+<� q�s�TBO�kk��?w��u7̽��W,��=�o-�#n�('���H���Y�H�"�O-٠Єz	<W��e�R�!��^i��� Mt0��oi��}	��Ԛ��x��;�7F	ƶAU�E������)	�Q�j�1X���%�|Hx�`��V7����h�B���Tbf�5v�2[D�P��Nb��t4kO��3Y���$Mz<� 7/7(fW%��'�L0A��&��l�?�'+�^o�C���ݏ��~J:�Q?�l�ћ��p!x����fy����������B�9L�����X�Q��^R��+e�0�׵D]\@��͕9��؄[d« �wcH((��bW�uv�	�����h���Ʊ��}{�XN���%1�PEy��R.~M�^b�F�w�z_	������*1����FQS��dx�C���9_,
U?@�A>Qf�2��o>;ͦb�3M�wu��g������eS ��2{���PkW�Ġ_��
n��B�~��_ƓA�ڑ=Yl�R�z�tU1��%�(��Y�dj��-Q��ș�$\�isHz`���U��я�;X	w���$����qjҳR?��r�MR"H��\oq�쵍�m8Q��%×ï��-E��RӠ��oTX���J�+���Kq�5�OW�П�x�2�RG����G�	��:>�Eim���Ө�E��6(Py�4�_@�v�5"I�XA��g4���Dg�tIW�JY�65�����=C�mP��(n�������#��ɶ:GC���i�g���Q3Q���IrfiY��V������b0n� ��:D ��ks��߰h��=~gx�4֏�\ų&��������Ŋ�rWّ���:Ա�aO�~������>����r�YMC�7R�?`�G����Qc{�u�V�@��6��=\-p(2�-{�d�@��c�=��T�5��ej-y\�p����9�So�zrt�K��J:2вJ��{�.cթ%�����;\`A�|�6%g|o%��]�!��*3�8�/_�?�А��6�o_
��
	���>��V�O�䏈�H�<���wNw[U��� Ə'F2�o��Y�R$�n�X|c��Ŏ�7"�����D�H�=�l�0�@�?	�y8-
x$<'��~��b51��yv�~v&�	"i�sl�0���
s�L��x�,t�j�;k��,��ȭ;�&Y|㑭`�Vad4�FZM�^Ms��c�*��(����+�	O�%)���Q�v������%�\�STh������:L�h-��"Ǹ�����j۵^]��������V�݆�U��l{հv�,>�$�0UAvk���`~}+s�o���?ų���M�j|Y�C�hf[k����{W�/�W�)ƿ�(i�k���D����$�b,���sIL~t51n�}������ɀ��+#�U�gU�V������raq]`�e�m�:�Fm�/�@k��7�c b +I��0��=wOE�e-r���Ch^����u��qH�r�p�Bɝ 5�����v��b$q��>���ܔ��������n�a����:xXQ�Z3����C�E�{<ٔ;�T)طt�6T^Y�<j���r��&���7"2(�¯CT�����i
�чv�������1E[�x�.ش`=�]+L=�M����&[TF��|�Ռ�M~�k���k*�����q��y|����$���U8{k�l���E�[23��6�����p� ������U�Ǥ9\��C��oŸ7+�˼�t���o����2яyR}'gzQRf6���	)@�чQ3K7�9z�V�;�AR�G��o��X��;Զ���&��?d�� }p_:������O1�Q�������㑾�J*�a�F��M���i���͡��l�{E_��2��e�/���G�Z�ȖS��eD�a�㤰���9�AF=k���AF��p"��m�9dν&,�2��%2�a��p�0�4'�W���q�A�h����ȝ��^�Ye����cM�V���kE�}��v��	e���h:D�!�T�#�7�Ηӳ�b��	2��v��Sx�YS�U}̿���-� >bK.V-�	�'�Ǟ�=�o�p�c0��8"�H���xɯ�S�Mx��z���5"�V�_���Գ�X��'�W`�c`�Kw_�5�o�)61+9ӹ�c��7�J3󏁬�a����qU#��{<�ڧ�heq&���I�ι/�ʻ�}<6)=9&l����g�WaO:q4]b�U%����`���D��?�7��~��y���7��S��$}�~��v����)�PƑF��j>����!����~3J'��"��f���Z��6m���-*ĥŀJ�d��9J��㴒v�et^�C�9f��x'9!�"�8�����S�����e����0�����j	�#2����lh�aw	Q2����;K��t��Gp�O_���S��~fƗ#�Y5��;^��U���W�~��j���-���S_x�B&k볗�kPS�*#t`\�����S�|ى��*�}��3�O��̈́���_5�����ăy�Y�Ϲ�=������"q�v��o��j��acR�_~N�N2G8�b�j���EZ��$ɸ�oz�C<7�_�1�059��i�V�C�^�{���W�h,y�G����x����Ư�Vy�.x�VDkkTUk� �8�_`|�X׌���OMa��I">��f )w~�َ=?�'ɉu�F��n�A��:�>{���q:
f�CU��$Zo;>��c�-��Q۹�ɻ��i�r��]������e��4�$.FWĎ��8���5܈�v�P"�"� �m����୨z�?Fp=q%�»H9C��t,�겟h�>���E�ϖauD!����Q���������'�4��k+1T�a����Y\9ǀ��L`-^�
y܏�Z���C~P�}���h3��Yaڂ�g�c�5�ʥ�E���!.V�0rAQ���t/�oR��}���L���l�Op�Jgs��խ�QjH��f�A�踑鷦x�F�PBR���ñs|�-UF,Q�W�m	��CpRE����+�����Ƃ e �-\����O����=����쓚��?_j�����T��.j�{1���jh�upC��C��N"�Yw�u�=��� �MjN0\,�{=1}�q��{�J�~��i>���ƌe�~6Lc�Shh��Yu*r������Y	��'ސ�4O#�	#Qf]x1��H�7I��I��@ݤ����ks�5KxX�NSL�+a5p�=�[xI����	����I��eryӲ�49d�T�tu�$O�i,Ose���)��)y,����`Ȟ�r�P��d,b���������<)%$n -d�j�3�=A8����9UTa�R�
�޺�G��ޮۋ�ߛ�
,��G�S�f	;[\,mTߒU���`p_����U�Wfa�/vÎ�/����S����2z<d?*&J9$�+����-�9��7�l)����WP2�vvs~�D��\��#�Vݙ�9�ih���Sk�;��#���������ı�W��>���N��O' b@��m2����?��u�=��z�q�������� �+0�Q��#�����X��G��kS�T[I���Sy�i3�C{Odm�Zh�T�j�^��j�ċ�`c�j�҄0�K���kGe�5���Y�W՘p��4t���8�8�S�����vxqLw�Kw2�t���M��9?'E����Q��cd��g�rO^P"ا�8�>�H�":�X)�r6f��U�}hg��0���E&_
S؍-[6�Kɖ+��&�[M�2_9Y	;
U�B�G;J�n�g^�Z�����=*�XK�������)`���=������<��;� �Җ��C[)�K�V�}��'g67��$���P�˹��_bƧ��8`Cj(����&dz}5��Ƙ�L6�D\��c$�?��]�W�Os�.HEh�9H���Z��P�Y<!9�%���^v&>f;�j��y#�*�ݧ�3�.������q��o?�ɨ?�hZ�0)&S�,���E���4,��W�2>ku���M��v��3�Uw*��6( ��1�����x��Pa��\;�+a�>�Ũ4�����j�nf�!v�*#+��i��]g7�ۀ�{y�~.�EC�ћ��������!�/U�̷��r��$iތH������+�e���J,��7�z�Na�{TȥǨ��a,}��#��.����(��X��K#GN�����BV�f$F��.K���,��gMoP���tl��|Ax�,�s'!`tn��ʠ���ǫ�=9h4��r� :�u~R�Y)tU>�:V�M�ϣ�pHJ��>ΰ��'����N��IO`����4�K��{a�7��@_�1i5e�@�.[P��F��q���A�;on���
�j���3YK���Y��(R5��Kdۍ]n�f9���[�_���k@[�:���:�:��M^6����}�}��\d�`
���	#;�	��3^�/�1������D�����A2Z�9;c��{Q.>V���N����4r�M#�Ow�oW//*j��g�|k�S�׃��o?3S��ol����W��}�ݷH���ya���d٩υ���b�����5F�wڦ���4����,��8GY�T��<m�xzɍщw�q &�r�{Hw��T*�P�S��c�������l�O��&�Ρ�9[MGКd�KOu����u���k�A���[��+�j�K$��2S�!���	���&BT�����G\%D)l��i�EŰ���BZ�Mɻ:��A{NH|,? Ǻ��- g��m�թ��1�>��6#����i�K��������ȉzy��Bͮ��(����[�k� `�:�qvЕ�Z���@F�ڪN��SG�D�ryX�uM�D�N�qr��SWH�#��,�6zd�r��:)�S�� �A^���lg3�p$Y���ۥ�s�8z��8&��sH VSe�P0�WI8&����1��ٺG�����H��Ŷ4N������O��O�s"կ[;�xO�����K���)�%=z���`��rZHkP_Q:��l��߭�;�L�c�2�/��Z���R��K�`�N~`�W?/�2,NE���5����)�5���
.5!��C�ZQ����"�'��G3�yN2�
B+Y��a��p���t-C�e!�4�+���st�rKF,�S�rá�<Y}b���ѷ8���V��	6.�k�UT՛2�k����*R���l7�k)R3f'���e�^��t�1
�sL��������0��VL��T�x?���Й�3^�H�^�|g�T&&���{�T�z�\�'bƸtuA�o<��]��#G��	��؂������cV ��mM��s�Y��0f<��O�GP�k*#�cbDR�K�ėV���&�5e|��iWJ �
ef��j���ė��|�#&��O��b��	"=�z��/��1qeX���@6ʦ��~F�sK��9aD���d��R�-:�A� R!�3���>.H��jdo�����:|c.حCv���}��U�C�V��Sw�+1A�*��N�vE�&}�nF���}T�?�ٵh@� "�j1+3�j��"OHo��盒A-��}�z�{FS&��8垈��ǀi�I��I淁2ko�� ���� ��&T���i<EL`��}�W�E�ݠ�
?e(<��F)d/���Ϥ����:����f��6M�?�<|mc��^�b����^�?г���T���ag�O�o�qb6��]��TPdq���)�"��%�~h�ƃ���2I��+����J��Aez�-�C��oV�{����Q�r��
!V5���@v
��L�ܳQ�4yX���fpÐ��C�����e+��v�� 
��a��]z�(��.,l�	�m��u�Ë%�����] ��$�'����5�U�����کC{��1Kα&U��>�B���}qɠU�V�i���WV�+B*�`�4�}��X���� �x+|�8�ҋ��1%�&��HS���ψ&[�mu,���:"k�3� li��b��[�L����{A4؎Hd��'�e��.���2x��8X�욒J�]NH^�{=�j�)��3���L){t��y:�j6�L!T��O	��Z�,���rV��\�MN�'�<�2�u�B������7]�5� ;+Eo���s�ȓ� $�
��ĬN9�! ���Je׊���c|��絻0�(�`���
�}뮮G;C�,"�<���vǹ	8Rf/#��)bL��}3����@%�Yxh�Y�a�uݠ���l]&�y�l��Ñ4���U7ݓ��>��7J�\��g��p��9+��M��JbҤ�~�0�ُȺ�-J�$�YH1b.��5��nSY�񘾈)om��s�H�t�Tۑ�'4�������g�� D��c1:�s�3ɖS�%U a��Ԡ�%�Ϡ�����u�=t_�;����)��^�[�g9^[>��߮��W�6��V�P����jńj�7�c�"\AG͜1@@`�M,�ǅ�s�����'f�j�O l��P$�����"�S��I��v��a�3������յ���m��&"e=���_���|�m���CK;��3ke�Mg�`3�W�*�TG^	F��g�I�B]a��ƀW�nmן���w��J��(���E�uX�=��Q�{�rL�wFm��!m*��Uę�b3������S�� �ѹ�?|��X���l�����7=Y�Ƙ��5��x{��wx�n��쪑c��:GX6��3Ъ�.x�5�u�f����=���X��7$u)2a#8���4���g�e�`t�e�Ξ��y�N�wS��h�E��i����po�|�/��(g�	�gOW��S�Aʒ�3���$6p��YM�-��
5=zK֤���OKW�Q��R���QTM�#)$+��^7�SV�ɝ-ќ�y�z�*˙�]�^">�~��3*���h;�V��WE��#����ء@;&њ��]A�ĳ\֩�e��z�S�,J����<˸^H�"�n���΋(�*�0�`Pփ>��z0�w����h��*.c2����Ƃ�%�?&.������X�rO9m'
O��"(�<.�銨Ea�`���e�r�d���Cc��_
g2��FC�#t��X�����Ud*��_ށ��=D��C���9�O��MN�PCOha*P�òZ����qm�~�J�*�R���]lj��i�ɴ�z�YI�f �ad9:���biմe�r�t��H_.-D�����|?���	�p��7~��D�.ys�\��>�~P�F����I���-Y���g`�"�T�یH��g�erZ�H+I�I��=���J>��#t��jGBz̵=<��f٤������v��#��ډÅh�ߒ\#K9�0�kv��]v��gC�	e�b�Xg�U����9���pj*��V�Q� =�Q��Y�@Q�bUs����։�6uc���-��$=���s�?��_֥u�]�%�q����R�Gt�Ҩ�v�p5�@_����7M�4��i5&&Z�)�nQ�7\)0;y3�<������Gy���ޘ{O���!��=�0��`"��im�D�Po�ާ}�ܳ���e�,��Ux���/	{+ہ��G�
0B���އ��|���������=^�z������4�D�l"8��!�W/�,�bw��Ω
��^��8�J�]D���O;y��b������l.Ї�����J�E�4��'^�A�1šG=:q�L����T�+������7��9+]�����_�{��9a��lR�����eJ[�ڥ�"~Ci��sP5����(x�j.�E�y��d��oH�ؘ��y��O"���#�I�����W0O�7��	��^�.4�ֈ����3��΍���A6h�j��@9����E 'O�2\�	0�����J�M�z�K�1��7F��q4�2q��R���p����#D�>�'�8
VzeC�:���q#Y�0�I��[ꛠ#�B�le#@H3���z%LْE죥x# D���H��T�J��H�#����	�Zg�&X��2���4閿�)��ƮJjL�Z��\Sr%oTjsSxJ�^ �x<~p��b�� ƕB%�x	�!-������|k�W7�$b٠��1ʖXh^*:�%��{Ǯ�Hr�+Y����1�@��T�Ubj����xEv���=^��%�L������l�0�b�=���MZH�n�jI�s9*����B��C��Gi�@����J7�:pJ/bF��Q��p I�X�[��5�`Ϩ�}տ�ZV���HQ���҆�Gŉ9�- :DGʶh���m6��&6oO��^�e�ϫ�h���"	��EB�6�N�;p��c	�D�t�J�����eF~��d��#���#o��n:",f[�W��n�Z� ޤ'��� �!P�����t���CC��ސ��xx���$�k��>vy��1�u�-:�o�� ��P+�Sp<sUk�`��E~{n�~�\7�b�ː,���qH���.�i�+��J��.4R30�>���9�b��h*j��9H�p�m�uP��h<2u�����{� EªE��ZD��vҾ�)�Z���O��X	�����nuwY����gl}�ȯ(j#���&�X��-��⑌7�ӜB_��}�͒VL����Y�lC<}5芮ԵI�+f��M�J�h��%L���hU57_Fc19���yx���VR�k��)˴�P�����]m��#�(uV��/}A,�q�	���{X�Z;��R�Z��Q�q�vf����K}*�_�,.'؊b�Ȧ���p�s����%��f~%2?3���
p���
'�C���4pc�O����3��.#ŧ=��̢kmJD�i�I�~������6�I����r첁]���P��}���uzPxN�p�r�L�]��-�	�r�f��8����#�t7�߂-rh�,!�~�����%��1ЅsO	y����7��F���`+�|��:Ҽ6�B�j�+)���#������m^���L���><FV4Ȗ����<^�-�����Z��G_��X�F]j��Yu
�?������aV>�B�kv�6F�[$jP\ ���^�1����wV���C�����\��`*��,�M�+~��R6��r�s���Y%����E�g��6��T�r��J�$f��Et�ޅlu�v)��=��e�2_�뛧^�mu����B�VN��B��ݎ��j�T�3�l�a�
��q^�M4�y��m�ŲC�6�O�O���8<�r��r��A��V����&��0�:�Pk�f��r2��!m>�Hql_IcD@���m�����ޑdD�(����]o�� _�Q�G�:��;*pH�ȼp�3ר�;`oJ�^�l�|���v�:�D.E��JYI(���ʩz���sR��aIj+v�!�Gp�{��9j)=N0���ʲG{��J����uD�'E���Q�5t��6��|F���@�g"�W˴h$W�R5[K��쾵�Q"vt�Z��������Y�%�Z�*���G��xN�\:�_�{��E�����ł�N�b���pϲ@qQ��M9;��P�����I�9F�)��XYG�FVvE�,e���<b�(\�ZA�'U6L�q�7�U�Ό���yo0G#E=��s������蠌??r_�q{�C��,�}���B|�mlzz�B��r�@��^�s/BX���DF�Ȋ���A-�n�"��U�o��C�?�g@Mt�q�,jK��[�[�o,�oJˇ�5���BR��qݯ>~m!�D>�V��CT�P��oE$����W0#���Y^v�湁�YUr���p9W++r�l����`�Ͻ���:�4P�Y:��\;]s��zຜE�"���;,���J�?���@��Z�{���?�3XA��V�=ώ�<��m/!�[�~�Sl��I^\���ڷJ@��3��+Dl���;cE:C��=��Q�mNj����dņy�㔼)�k�W�ؚ�B6cS�Uȁ�_������&3��`wM�S��{X�/���ߙ�*�_���p鄘�f�i�:�s9��U$�<���r��͕n�LCO�Lk�K?
�?�[e�b�u�	|g��Aa������OR����LF�h]®ڜ�*���;� |Mn욠ڞ�Ê�g�-�S�vH@��1�g���!�e� �Nۦ�m��C9�nm^jLKN��ѵHR��avU�!5��z�4$�U�i�MO`J� -z;
F��E������������ƦM���_i��]��QC�+�B�c��	C�_Isu�-T���5o����$�$/>�G�Q{��H�[��:|��k�u޼8 ��o�����_�h$�����qh�G+۳�W�0�y��1����o�)���v���{c9�����p�  �<p��d�\��[y�A�W�g;|�zV��5�l�,V�N�֪�?ٰ�ݺ�^tE͗�8��b��0�����"�j�"� -����)�')�9���\M��͖��^Qupd	q��Fz�I(jeQ2�Wovq2s�x	����F�s�)�e�ܐ��c4��u�����~mKރ7Q j�=��e�����Ư��h��O`byڍ�J-��98)�@�8�Cc����[7��B��j�`���/��yw��.�[��i��ZOs@O{�Q�?ߘ��h/�1.&��V`͑�eE-�V��X��gT�K�LP���I��qǢ�į�&�(o]�[���`�� ��lH����5�U�2��MR��8���(s`s�Vip1]�o�9�;��cɲ\�hY%09��݇�fR����t��BY�IG$�=��@��D�:���$Y�=;z]b����G� �6ҋ݊��6����}f��(�l:��d����A���Z����&硨��� ���1y���l��nt_0���H~E������l�!�r;i`%X\_���DC� 6�Z>ӏ1���N��0H��#�*�^��e�����Ĳ�8�5�h�ec�����I����\v�$�D;�t!Q�If�W8��2&�:C*RdTZ�W�,-f��'��h��@^ᩚ�r�#m+�&�߁��Q5x�;�)��{C!fi�7[\Mts�[�W�~n���u�<^G���b�h�͘�3f='?[]�m��W��L�]1��tIR�J|�.tQ�G�VBHY��Y�pR&0�?v��M�k$g���WHSoHz�ꍋ��H��xT�P�~���R]	�6��͜�DX�� ($�A�XC���<�
g3Л��H���?/�1$����P�_U(I��Ҋ��,rxlb���<����kF�������M�{z��!�J8�~/�{o�b�D���ܹ��K�̮�-��r=$��{�|m0�{p�P�}�E� ��^
��ʾ��3Uަ���W !�_Q��i�7ݑ�=d*��l[����W'�ݽq�ků��o�<"u=�bK�n�2�$Q������(�?��&�f��M7̅��ˢ�����y�i^NN'T嶌%33e$ۻ��ş���u}J��ѝ� O���)�/!�>,t*�G���K�+��l�3�(��@��TH�Qħ�	A*�~�bۑC�_�2C�[�;����N+�%��Nғ`9�{�~bY���%C��{��9�@bƑZ���������?�����1%1<�II �����y�p���~�Y���U����z�ŨC���$?RRyӐ���=�V �eS4Y��cW�lWnpDb(��R^��IS
<,��}�OA����:��5�i���ԯ�����4��j��Ǒ=p�d�����}�d����i��aTS�:��g>E�U���+�r��*�m�����P�b����y�<u
���֪�����q1��o0!�
�jGvp�_ (����\G	�L�u?��1?%���B�8qH����S�@�бX���dk�]>��p��o�D��9Q1�y�F<��MVF�������zpҚ�D�P��f֌e�-�$Tjn�� �{����p��[Ӱ�B��h9���j.W�I�����ւ�`#��{nH��e���.�j�!8$���+^.^v� ���4�(�V�1��J�0���"?�I�� <UwPk(~�5La)&����A����m:�b�z�oN|�2��'�N
8h�U�6�2��
�G�,�x�MdxW{Onir����.�dԩ��s*y �LEg`�648-��^SY�����i�pLwC��f�q�	�;�F�0E�*0;�N�*�Ml} �<���˩K��D���ʬ�_V�K>p�0��J[P5��]9�REI@6�ho1�ϛ&'�L(��[������S�^��A�.�	䲵�����M���'�}�%ŧQc?q��#��^y���- �|G+��+ԗ]�~������8��or}�(�^�M���<�?2�d�OR;��/׼�S���������vN��rYf�BBd7���pO|J�:�Fs�(����9��y�Rvq@o��K+i�1��qb����);�@�Xel޷yf>~�Qn���hE�� =�n�dl�% �˭C�K���z"�5�C�!Ф���Ţ?���bn��L l��b��q�����o�7v�1e&?�J<�jwt���� |��4@���
��S%(jL1����YAћ�8�o^�o�o��ai�?;G��҈D�%J$�i0��>&:&I��L[�:��Rk�f!&�DԷ�ƽuz�.n���_*��\��_�W���:���yJ��f�p��;�/��jCn��^#?��Z��JA� �Ac���g6��VP��h��P��^�n�4M&��5��z�3��?��u��N��<[�
@�����b��V�auɱ�� ��#7S<�֩ؐP �ESz4l�u�z�[�=��F
m��4�fц?�iE�e:�F�)_��D�(�j�D|��X��o�7)t�5WT�\�*cF�i�������G��X�r�pa�?zn��O�4�C�؄\)� N�ҝ&� �
�XL�.�J0B�:K�tW�T䉅G;5\���*�_���PYN��_���y������.Q�4�Ǆ*}l/�A���^ {8���!4�	��:�r#jE��5\�	��3_ ;aG���1�ք �����[~Zhm00��$�0fI�^̑�=�����K/;D��J�=����1:�3�� P�
��޽Q�_�?;n���0�Xv�;�R�i�ͷ��
�K-�������ն���V��6�u���]��?��/��?�T����|��jM���s�޾6�Y���G��}8�5!<��+"]k�3�Z/W�~�a|^ò�]ĭ&��k�]gD��CT�Jf�ZLPy�vy�)�f�5���Pu�EnP����^�V��.�3�/��Dz%1��Zڈ�x���`9��ȡn�2���&� 0A��l�kîZM�{b��fn8(�H߮5eR���g��:KNt���d�/�xSd��,Zv�=.��}�r���pվ%U ��6�k�3��ߕp�z�s�4
|3��,W��ݍ�|�l�����ԏg4<*�?zqg&�ƓJ3na�A�uT�~sΠ����<F���(׏�Ii�nY%f����h��=x�eAB�=�M��$y��M�۹�������R&���{q!6�J��u�m�,Xŉ���JX._/f�	���޴�c�L�H-[�^�%���C�	�fE����=#�do<�L��P���E.�������a��0.ne�f�QW#��,�'S�	��3;���ih���cD�i��z�`)^yǷ�0��`�@�|6�#�޻z�,]>�+(O������܂i7����4')�̔{��IN���w+�d����C�v<�U���w�5�v��^Χ����(̎�b����HL�+)B��ZL�p���zH��>�	�1�הBl�[�a��W���m�@��1I{�A�G!���_ �=2����H��lP�t�������n@Y��fw�Rk��ԅ�~�0���$�ɑA��*j�qE�k�v8>����d�����̏v�����[�H�tz�n����������*.�̑`	�гr	��ژ����.����~>d	�mNL�}C\���%��f6������(��v@s�^��!\N�{�}n�5ik$?ղ�~��u����6CݷZɝ�P�^4#�8�������2�׀�2m�<>�̧��Y�d����`�T��.	�ۼ��t3m��ٱ^rr��ۜ�AM���m	t�Df�A�v"O�}�g�-?����S��3�9fa�媍��D+��i%.�:Y�F^䬹�>a���)�>z��[U5╀��\ɪ�C�j	�0�z,i;m�`#�9ν��X��E�6��,k)�b�`�q���k�lE��,>��!	MfN��|1eg:�S��UOa&��N�KT��zcv����T3,�tq�z\�ZЌ�lk�B���^X[�|}t����{�[��@U��t,Qz2����Kw�Zܐ���&'0���Ƣ�<����|(��=A��nk-�nc��]�]���l �m"G|�ɣ��ۅ���]0�ֈmY{��� ��� `3U�nb��UEɅm�1�؃j_]��ɷs� �t�_���>F�Fg�@0�]a�ϟI@�ֱl y���ސ���0�=��,�ú��DdO#���Y���?e�`�a�z�ŭ�-��3z��ۜ��N�l�kq�bp�3��Xe�J��<~o��������k�@��@\��G�ؚ�RS���$jYv���E�\5�Ψ����z�x��z�Ŋ5I�
�ǆ�����c�k?�iտ�$彋� �a���xm�<���nwթ���򄣋�����4`5M�X��h�CH������<���cv�V�9-8t��A�t����4��V���Km�Zת��r�Q1qOצv�2�Ԁ�nTflLJ�a3Z���.F��%��N���$���i���c�X�N�r+pn"�*x=���� QMN�P���ɔu9��-oִ&*����׫�;K�H�o$T���b1-��)�]��EԤ0	+���� �d�~�tv: �(�D�^E���Rys���K/���Z@���H\;!{;ߣ��M;@��C��1���L�so�ʺv�1qc���K�n� 4?uJ>�G���PVk�����OxtU��C�Z_��1SX=��IE�(b8 �� K6^ ������Sx���j»�Oیc���o���L�������[��S�#��Tg��c$�=�iI���/3i
�����O@��$��uV
�����W���pOu�E�n2:f.
��q�f�p ���v��$�@|����O�ƥ�/�>�0�n�\��<��r-m��T"QY!���X�o<� �C=���n
��=�y�Rm�E��4�ǅ�1O�5����I�#|��#��:ȅ� �J:"?�T�Yb��>�n�{�R���!@�aZ��ǻכ�PD/n�w���C���QA~��p*)�}D��Y��C��H.�e�<�l�,@�BY2��3,�ڣ�"�q�9�&%�&��Lh��o�ϫHp��v]"�A������bU)yk�# ��$F�`�1�
�}z��O��ݡP%�)f���|��Grz��2Ӑ�3��a��"Cv2�y��'�)�
"�:ϒ\�e��m�e�$��Z���>px~
ʃm�#&�4U�{�+�&1q��!d^&�X0��,$��R#��/�$��N�qM~�T[8��('��Y&�߄ҩ������Ԑ�=E��5!TS*��A�4��X+�2
�'������'
O��X%	���~�30���~F%��Hb(�z�:TYs��p�Q���)��J5[Y73��(=VC��<����-P���W��ń0�=fBP�Ԋ���WC�� /4�n�1�����zt�,)g���Ј���ލ��������/���q3k�\XYZ-ߌ����s]�IS��DԿ
�C\`y�v>��m�w�I�&��m?5���a��j�ڙ�:����ǜYG�'v��V�vj�B��xd#�5>/�l���&��=�]��gC.
�)4<_`�E�fY�BX^]�:���B�x���c-d��H�kb�=�a��w���l]�B�a��R����P{���z�;��D���J�?U4�f�trvJ= �ZO�.����/����lд�Xu����#`8Q�~oqr�.4�Rl4�;�%��t�^+J)G�S-�^�T�GN�{�y��7�o`R�Oob0�n�܌~�7���#�y
�Нu�',��x�Y� 
ғ>�=Tb�l���y�o���Q$����p���6����zxF.a���T���a�C�E��;� %2�Q�5n8���M`?PzeϹ��s��,}�0f��� �/;����2��r�e(��f�3/���\,�@т_�Q75�Rl;Yѡ�:=P������ʚj�T�fqٲy�� Vf1@�;1�1!c���[ ΡC�1u+y[���ls*v[�)N�^�Þ��Kیp��\,Y������o���A�o
�c�i	��KA�i�5��v����ȝ�c��"�P��@\���,@n�SV4���%����p�oqh��D��[�-+*����w'��������͙:�E��ڙ�Q_¢S�z��ױ���b��w>D1v�;�($�$FxdA!�W9j)�!/�N���9�k�)����u��N�?�σ���I�����%�R��A�F����qJ����'¤�C��D�h?d�>qs�%�(Z��H||.�ؖ�h�,w�̖�gt��SK�
U-���ܗֱyv�1�cpP	9�=4HFc�S���_R* �_9��I����˞o��$��jP"B#uk����\���KoC���<~�ɉ�C��+�  ǹ�oj�kJ��5	#om��_A�� xAC_W胐E��7z���JV~���VXSX���i/W��A[iz>A�LRm����D�T�(�Y�R㢋����� ��F�VF��Y���}U��z�Ze6���b#%�[=)q�v�}�Bu��;�X��3����4�}esc������T
7����q����2/;T4�i� n���J����?WH�Jg��N�8a�����TD�h�>��0�:�"��{�0�E��t*X${�歲N(��Ȟҧ�3oTbO�B���m��p�"'-,�22to�6'�1�3G�\��l���$X]�����t�d.���yY�j�u�V��~+"�U�A�]�bY�*K�l��@�n�/�j��/�`G{0u�"܅��.��Ě̤�6i|�3N���r}Ұ
�!���~x��kAXA�	�* ,�cG�1�f��t����|>�̑Fu�O���U65�yZ/��	-�9�b<��ǁq��o����K{�[y��>(od���
v�͏��6T�\��VɊu`�'ӱzS�FŴ\���C��T�y�0Q�f�U��콮Xl7�t��a�Fv�m?d	�EQ.��4�<d��Pe�s���u0A��}�!"Y� a�;�J�sd�Įx�����3����$�=�k�J���	�f��A0�޻g��A-���ٹ:0���Ϫ��/��ↂ��L���¨*/ބ�b���Eh�z�< 5�F�O��*��o��a~&�O�Q�b ��^�gF���R��j�8�-��ρ�Nuq���b���V�%4t�/=(�*h���-��0��P��fP+!����HQ�iK�]u�,�ˇ{��yՇ�9:a���l֝m��X��H����U�*;Ӥ�|�q$�1w4`$��K}yo�?˯�6��E$�_s��BK�~�m�eJ$O1�YbdQ��\��Z|���f�[K�=�a��%����~L?pj��%%���������3K�1���߃!h1�w��ҌwsЗ禨]�-��-D����'�l�Q-Ji{1#���,�(��!oA�]i�[�;e_r_�b	��/�d�@O�y�{?3�Z� ��p=�F2Ͳ1�?MHt���[��i`��A���2����}�9����!-�TJ�27�s;JIK���0�F��� �K�����A��y����BW�	� ����}�b��:ȁ(V:��B��3`)��DZ�oWjvi�~��"�0t��e9hF����WQ|k<^�>�.�H�Lut'�eH��5�_��6s/j$�$�>}Ԓ+��<"�wR�}���6����I�_/�Հ�<����W1pl�JO�lߙ�&�쮴]�T���~n�5�RF����h�qD�	ĉ��4b5z� ;���))����("ڢ�� ߸�x�My�V}�=�2���.G�2*��B���k��Y���ΛO�ԗYdHq%uŴzҦy�<�wkf*ε�|��؁�\�FR%��j�G%�ZE�-x���^/K�n�����Edbσ�)���*�; �J੐���:1��w|\������n�M=�� ���E�W����伃�֢b&"���S�J� .�?���)#`�jY�MU�&̜�;��S/�@��f��7>�8�z�H�>^X����}��<z<I�\�.�N(�;�G�w���d�������n��U��܋�J���_W�Ž�֢A�y���i���J�.u���M|[�.ǲQ4�t��v����l�����O~_���R�l�Ӱm�t�Jط���Ѧ�����R�!��Z�=EM�[�m&�3h�a��>�0:9D�8���Qŋ��?K�</H�,誽/�1p�O���_�졝cZzd�]���������:O�ʌ^迚]�"Jz/�p9���Z�\����h��'F��![��篝�����&-b����X��{I{-/C�BdK ї4_�S�Xk	"����?�W���?:�������oT��i� �� �T��{R&i���W#mƃ�
5F���{����������g���~�7z�5���%�/<bqj:4�0���LLCb�&�ӊB+�]�~0�c�ph|�'�uD������`P$8��}�#	=���_��@'(8��T��X@�P��<�"�t����_�弨��:��$mDZ���r�R` ���� ��w���F!_%�0%�/	!��8�X{�v��B�"L�PR��_��%k���8��P�`�7򢂻0�Z�m��r[t��y�ŋ�!vm��Om\0���mp����v��Q0j���Ӈ6��֌I���z�|�l8`$�Lt'�:M�U�o�+^��m]#eIY�`�'MBu%~���: J��K�in1���P�;�7�LWe9!��9O��~�Uԛq&����ަ��"��Lr�f�>xKr&����ͱ� \���l|EB�H��w�3䕺nn���-y���I9�D�Ƕ�Y&�g���$�y-��=Fs��{�߄�l�/2~YP����8Lr|(�.���m+@'�9{lr�V1�cx�3�)F��>�U_��Ԫ��������	8Zs�,};�����1�8����9gh��iv=>5oW��Խ�J�T�u�2�l3J�mn)�+O�U�_5�#��?(�)��z*���RXd<]�.��ɯ1�H��޸E���4����c���;�,��~ȕ��/����/)���K?1������f�_�M���,\���vA�jiQ
�,������j�;~u	k|lD�"J�*�W�r[S�)U�RDh�hƬ_�|r��%z��|t��i�!��ڀ�T�m%}��Ə��gL��+��r}�����n����C�g�о�1۴Њîʵ�a)K�yg*D'��Hz�?��GO������V�~��'F�1n�Ӓ���GKx�S
���ӗ�Fvp�����ŗ|��L�g��Go��Tz*=��P�����橨B1dO�P�z%����]�F08�z�V��b�zQ6��̝@V�U�Il�N�/j����/6���j׆���ءg��j՗ǝ��s���G���mA��+Y[*�Y��B�G$�Qrz)�����r���	^ٍk0���V�&�g��Ë@����?F����ܐ��>�E�����A�Si�n?V�cF�$�e)�`�G��˙D}� y���5��z������֖�\M<yvA���7�}�)B�{���n���>� u�"�<"l���&���EU����-C�G�)� �&c7�W���z,��7-�QgOV��$��ĩQ6B�QW�J�mú�4�6P�7%��Iz��(�.����S�{��E�ߛ��M�"�����}�@KK���uw2�����yzF����L`�k�>���F
	
ͩ��9�4��'�94�Ҋj���
C����R���8�O'��	���w���W7���bW�w��;��3l.,��%@�Y�fx&p��C�U��� �d
������D(w"q��N�(%�-�M�`h+}V���������Bȹ�k�����Z�O[���Ȝ�}ZDr��)��V���k�hZ��n���Q�1qQ'��ֶt�+B��F�/��M6{�����U�c�_��&d��m��aa�=9}h�6�7��t#\�G:����=�D�A]l���L�h�.�[���7�Lȏ��\��5k��e��S�E��}�C����ľ��囪�H "�<h���������8'�T�2����{����X�Y�j�*�u�ۀI���e�B�X�8l���G�,�"���z���S �Έ%�4�����s�AE�x�%+eT����s\�����8����Icd�A�օy�����h����[i�����y����i��^���%�쓿,@@��4�}���x�Z��!N�Q�m�bTr�a�4��r��o�~`Ѹ����E�N(P$�78���Vy�ġ<���VP U��-f`��	��� ����!��L����m6�iK~����~#R�]k;�>!Z�MQ����OaQ�1]5�ǕC+9�?�w�f�d���Κ9��m��b*^�|DW�+��Q��* ?�����P;lO$r+*�C��������� &ܦ���Ssi�� �HǲB%X�G��<��ΰ�������yHӄ��J����i��c��{�YS%1��Q�*��.lx�2@򤃎�H�e�r��a���i����T��3-A�趈c���f=�Ge�W����>[���ȉjw�vJ�na��Q��3$WF�|��(g:�V�=7D�-��VCSH��B�|+�L2�F����d���LH��",���ew���v֣���)k�ʟ�����A�L�l��
.}��u,�
��'��&&*��N4���V;"z`�׬�UҶۼ��S8�H)�@��44�@`�W���_��� �{gӞ��K&Z���Q�>R%86�d�_�/֎�O!�%��8�%�0�b����ԥo�h�3)��1�?p�,��y5��9�Z�=,�h!�C�}P��XD�i��f#BG���W�qc\O)�P���:���6�0caIH�m�[���W����T,1��_W9�_�^�&�՞aa
�у��;S�E����+O��y��b��j#P+t�:��=�ra�T,��$; ��G8�YK9��K������1_g�ja)�nۜ��B�]m��4���4(�1OL=H�/�)�Y�h�+��qI�c�7��/&<+�VϨ��`��Iw����?��sZ��5�� Nk���t�(r�"�2��˳O�P��!B��JHQȰWڲ��j<�},����ٝ16�	��b9P���c�%�+:����p����e���Y)q��[��H���_nN�l��צ��Yd_d��F�|�l�C�E��2�ۡ��Ѹ���,�*�W^�y�����.H8<jQݖ���A%�X��rZ���r��[��[
l3�r�Yrڗ��E�$AQ�y/�'j�R����[(P��ՈSz1��u�Q3
����(,�otOM����6I I�auM����*)Od��sr��	u2�Ԃg�K+s�L;{� &E���\ώ�>����E4��N�FG�u���u~F5��Ԡ/�#�i�r������]�y�;���h�-!dά����f�B�Gs���!���.�Η��@�>zp!��.�_yW<R5@��k�݅I��M���DZ�oF4���H���mᏆBx����8�Z��q�
$�%��,\�P�6�q�����G��,�Ã���*oi�G�٠_�y��L���c/1rg�(إ�;e��v�
1��զ���;f[4	�r�����µ�(�Q���/���a��f��Aꑕ���Qh?Y���@�*�S�?��w��b�X������9����gin|b����!�m��@�N,[^Λ�y$��9�=o��.�r����e�yJ]*���AK�!�C�}��;RmB+Z5B�6��D3�����o\��@+�}�_���d�G7��[@\_�A��}>;~u5����N�?�v���=<[}@���b?
�ˢ2{S_��Tc�h�,@ځ��|��n����%�G�`,�i�h��Ov+���N4y�����	���r�j4DILd-o	h�w�"��+B骒�<ؖ�Ӱ�K�-�����%8�ƺi���U*k�Y&�rl�PU�cZN2��!ɦ(J�0Q��r��� �[p�_�]^{�	�{ 9B)��Bl�J�J�-�O����;���4\��4W�%�F����i���G�z�����^Nx:��.}sa轊_>1�H"��:�A#�<��U�E&�pה=��Rd�����f8��?r��|�U�Z������Ƭ��#�ֺ-�:�"��0��Y�#��A&���qg�˵+�h����τ=����#�NqoV���F<��h���Ze~m��"f&��
�b0V��,�̘�x^��6��J�����K宩o>Ƭ���	":�������\��4g8�;Qf<�aҧs��ݵR�YP��,�s7){��<t���7V��:A9�!6�RW&e����:ltS�v��Om3F:K���MX���Ӻ��ٟ9�������.4�\�H;� |ctx�:N��O�Q~�U� {Զ�A�^�DB�%JK�ei�
KM^�Yk�S�7�h�|�&��i�Ge�Җ_�=�-�

�)Wq����eX� sP	ab.���@A��&��W��*�~����P���8�I�>�M8�1+�o[�
7����q��Z]݆C�\ v�Y���#�HgrBR	V`3Ik#5�^�nb��l8lR��-i��9�}sɶ^��#�.�Er���\K�����K XZm~WaY�'�ǝR�����������vi���$Y���D|p���=��9��ݲs策5μ�6���u�WL�P��"`� ��dGl�
������l���Yv@vOſq`�����P5C�l���*d�Ӻ���y������D�� *��.R����c�	~!i��b�
�f���KQ� ��/�\qy-\"�8�
"��G�m�W�ye�#���衜D�+K�c|#�X�\�T�M���\�I�@L�?�70���:LgdM A�3�]Z�:{Q�7�7*T�V�g���D<Gcz?�l��k��x&.���`�F`�Wď�>D�������PR�^���m�]�`��~�R=�!A��������@�&a�1�%��)FD3��BR��*E��\
�A��L��]��p����q+�>���}��ϹgI�� yh��`��&�i/�R�{�G���7�t��_�D\8�*��W�c�]����3�}����Qɲ\t�3���Wb�Ő ���|X̵�9�q(�:��K�b"0,��W�Gfᅔj�E�~g����)�3<0ƳjZe}��^��^�ǡ�i�I} ��擄^b8����� ����Is�Ej�a�7ՃsF��ۺ
6��s�no|K�9�6��M�y'��y�5回u;[���tţ=� ���gk���"`���l�e�ּb
v�n����RF��H*���!h {�:f�2�������aq��<: 9ua�{Y�bN��Gc�Rd�l�>��S��o�~j��|�W��y ����S��[�U�s+��[�O�|�¡n��
)�`PnzÎ�X�8��>�|+��n��#K���?ڣlEԙ�R�'���2>*�ܐ'OF�GW6���0�ʦG}���8������8�)�����d/w�8}��z�)�y���	UX�>�1��X�������c2��P�Mm��dD���֩[�?r��y�����9L�'\ä��)�F�
;�o��`��)�鿒��PMs���Sy��m:����H��&�z��̈�~��q9��^Z�l{	��/�_Tb�� X�/��C<�N�`���[{`���݄�/J�tz��ug�����O�z�c#@�kܶ�^�9�G�|.�*ɂ�u4#\r�IHO�T����6�z��"������f�_�7SXm�Bs+<��P�l�L��Ü��Q�p,�&�3�A�KNk�K<7����S��E�F��a���Qʩ���� ���s�,���?=e�n۔۞�aZyh8ر�]�\���u^�!.QhZ{�M�tyE�C6tj����u�WMə?c��k�53k&|^W1>���	�V�\YZ���t�ӵ�G'G4��忳ߕqRa�:q�T,��Q1 j��c=|��{E�w'%g�d���G��5%����%VO�#;,-�qm�j��z���@�q:����p��P<�@ț�Q��/��E3,oo8���@�!�6�����Y�'?�u���k���dYx�/*�M��Ļ`¸�i8��<'ѳ���X���y��T��6\���or����+ 	:�������#�se/�{�G j�K�l��������i�g��V��lJמ��s۹���+R�>;���o��v~���/��]�I�SY���w�P�$MN�U������I�.E��5���n`0���<�-eZ�i��axp+��w�'S!�H��d�F�܌�oC��������w��𰨯3ݷ�RFw���.^�w�~�����XX/8؃Pة���ʦ��@��u2����奁�{̉ԾKǩ˺��.�V] ��������.	`��5%R�"�e4V8��,
��<�ңS��
�% Fh9���<�c����ˈ넛A	96���-��X2)��������(�5��-���Kf[�!��B������\�M$���vf�/�� �������If�;��S|]�V��Q��`AR)<j��4���p�&�OS���<h�9�q������ ģ����y8Yyl0~��x��Ƌ�~�;lYo��G\W3�B �Vk�!1��Z2���5:_@�0Im&��C:84�z����$:�g?�6��)B��<ݶMn-ht����n�FB6���P$=�0��+�;ء/�`|C��ӎ�9M���v�!@Bq1C�D��%�أ�w#0Z5�ݶ��j��9�f7�w˞��YM�>
�F=)j�+?cK0���u�C��</+6k:W� �J���.�2�'�(vR�M��uC_b���k�Jg�2]9���8L�t�>#s�͞A�.d�-bX��G��9��Q`D𽧾��g��s��u�j�p�-2SĀ+.Zm$쑗!���_e,��:~�w{'_e��h� �!>\��^B,���J���+�̧�cR���JX�3���If��,�R�����?(ԌDa�/$��U�R�  5w(OM���L�x/�8-?k���Z�"q���������8÷�O�/�	ԥ.��؆�ٚ��Vh5�kC�?\d;�;�F{	���]��^�K��қ߼w#�W���C��	�T����}�:i�Ŗ��S��O:���
6@��Y�$A��
�W�.��ۼP�[�Ex�&	�Axix	s�lV:$FJf+������QZw]1\�$� oZtdc|�$�w�,a��}��7T��{��!6���j��}Y������̴�������-:�g�e�:�Jt=Ⱥ@�L������U	=�7�4�׎7��:%�"�r���I��k�= ��ѱucC/O�N	���Fn���$��-_�C���L���IМ��+�'Ovm����K�������>�[0�T��1q�[j&Ku����#֢�+��C��ˎ�L]�{��
�8�6Sᣩ詜����|\/�e��Pt�LBH��Nv�O�is�C�<���;�谿N��y��y0'������Zp�y�to!U�&Xs�=�����9-V������;ʗ���Y�;CI��0���l�)O��05�5��>�4^��! ��h6�	���A�]T��Y�j�hTȉ�2<�/�(�&�i�H�R]�ՠ��Pg{��'D�礼pN��a"���9
{�U�L��Nb:q}v��;Qm�e�@��O���";�9 ����ͶY����M�^s򵈥)� :��άX�Z��������B?�w*�ǖ:���(�_@.\���@}�Y��{�`��m�������kN��� {��c����� ٚO�$T��\\cR� �� d[�Cn�4}�S�`���7���3z'e�kV8�F@Z�
���b��4迾��x��V�7+��u[���jõ��5�����N��"��<R�k�\��KM���t�&7��Lz#�&N��J���aUJ=|ܢ5����:��*?:h��*�)�I�A	|�Ջ�KL����F(�G=`3�@2b����'�1^8��z{.R�%&N��a@�vx)^n�{�@�N�=r������t��ەo)��;q��-?	�ώ6��e1�����������T�L0FFi�2f����KI�0q���Uta�Q������8��k�Xe$[��V6����J ]mF��iJ��D��`Ti� �NB�~Q7qQw�����:w�/o�x�Oҋ~$��,5w= A}��ր��ϋ�d�њ�-}���r�(��h�˻�ݩ�-���� k`�A�ԁi�&�^-�tþ9�?�Zi�y]�[��Zd�o�/�|e�I�Yy�U'3}���	^-]Q?�3"{U�[A[����d��ij��V-8��	y)�-�V%F|��|q��J0u��!P��C�!7��\����b�u+��O]�tC�&�3&�(��^��U�#�
�0����n2�k��f����oD�:�����ͧ;Yq1�����\g��p���lbށe*JU�U��"@��F�P��K��UIC<���$����M�g/CY\$ˉyi{��r�zSܰ~`��H��+:c Ç,��<�/Q�ˣ��N����"x�OBR���`vj��}����Ĳi���k�c���5d����ɑ<�=�G�"����\���
Y4���P�⭩8v���9�s
1���q#�U��A���Ro���
��ֶee[��@y��Օ���*���ϐB��w�x>�_��F����;Q�ls6�oQ����*fthx[���L��G��x(�/J:�fY]8zm��r(K�R���_|��@U`Lߐ
�O��Lj#TV��c�)����o�#����|(2.瞜�� 7���	G���j��>�D�uW�ߟU�0ޛi�<2���wn���^*��.z�u��C#C��z�\�%c��S���qY�j7���t��0� N��F��&������	��l(A���v��*�I��.*ͩ)@�m��;h��#5�d{|��KV���QE�o{��%��zM��[y&SGg֤��=
h�Y�G��}X��� F�p8�Ed�8{�H%d�@a�Jlt��3�ac?b�,nH!b%N�=��M����E���7� ک�c����P�^(�~^�n_&��,��WK��B<`�-&,�UH�5Z�������P3�!���/!�#��r�=�N���D��9+�� ��ԓ~��[rr�l�-� ��CL��s:D�& {�mu)�H;�J[���L�9��Nɔ1�
�ز�+��L�`���o�X�k�0H�|	��>�t:�8Os���KŻ~�)��#J<��%���P6��I��7%��Uxqƻ�)�:ً�ޥ?)��R����n�A9�����Y�O�ui�[-%´'F�zH'#CH@�u#���u�aI�_Z�K�)����5+b�
1�����3Î�,�8��o�M���<�3��߳�V��?F���'b�pj��g�T�f�X6m����ٝ��k�DW��]�L�0�w>`������{���}g˖�6.��T�O�<մei��{쓯��PM��`SOY�њ�Dϡ��v�u��],�VR_�Q.�~7Ҩ����m&�Ss>,�Z�Jtd���D�v��>cD��x�����͢[���s�4��:8�5o	���8\����l�v�G�Sb���&���Q��c$�����?>	���XFNX��Oc�QE�>#\V_��>%MB
T!j4���͛��{�����!�i��"�Z��B0F�Χ���m��a員��ʳ;� 7o��1e����Zf�r�nK��$2N������h6�N����A����ɝ��R:��.WYg��y���ߣ7� ��GpM��\�ᤂ�$S�M5�-ЬM-��U9��
5K/�<#z=i�Ӆ�4���߆E��e�ˏn;bػ���������ru	4�����G)��o���Kt�&�sB�a���we��p��R[���%c����-�8�dh�Lc���m�:c��T n�_2�R����)��i
�����<H�TՖ�Z�Cpv𸔚��}�}ݘ�u1�d�Ҝs"��6	�F��?��{Q�9�ב���i�t4�<��4�
3b�u��sdR�T��3W`�äۓ��
e���b��z��X�I,��l,jQ��T���utr��,)6�;�S����?	�X�=5�Yҿm�O�V� !��n�^/Me�=���,	Vw�(��\cr�7ɢ���'"~�^+�'3��5ؽ��5�#�H�u�SWS�����S�h���m�$���\�Z��%�/юf��3dl�)��=�sJ?_�3��r"1�]y5uL(D��h�6����߈�1 ���>�l�ord�L��;��0#0�qWm��*{K'W�1t�y`�~�nz�_�U7(� 6q���J�2^3�����6ܖw���o��r��E�=��(50oc��QÔĞ�5�rQ]sԞ �(1$k7�#�T��P>&,��9���a��C-�8�+;	���6���O��%�Xn��+]�$���'��� %+�@�|�Ո"D��'Ðշ$fA�YQ��nP������Wd��ZMݽ��E�Dd�IS�[�G����Z���-һV9�n��)�æ����1�zd��StލV�{r�h��g`���+ڄ�/&��WwF~ER���P�!� ���|�5�>��`�+����g4{-8���{;0�U.�8.�C�doۢ�̟ E���1v=�>�qҖ�
ʲf����TKc�]�+�:VT��V��Uu�)��E��~�IⲏqL��ɺ��
��cm0��.�y���ڀ��T ePrp��Z�\�I�%F���#���`�k����W����_�I4��f�83��}��~j�؃8��~�F�fS���0-!I%�W��*�.�̦���:�����v�U�W��L����0ѵ��IR}���h�������mk�%uh���D4{,��׷_��i����E�n��nY��5.�.�U��D(��~ �ky�1�Dc�M`>�qخ�ϵ�@26�(�w��G�}��o�r��XF!��ƙd%��o�0�|5���?e�g
����=��Լ�#�7	BN���VW��r_:V��P g���S������?�m��U�4��>ȔF��}�3ƪ'j	��Y�lϓ%�T��Ch�Jlbj;N:���t_�f�3g���&39��[V�i����;�z{U�Q;v撬6�t�5�i[Mu��s�	f;�;�i�:ȧ�W�<�vֻh�����w����I`���������r��1�YQ�~�Cӫv���a����do=�
aZȒ�����%���5���Z>�dx|�RQ2ϗ'�5�~����G�#�e�6��%S��g1�O(�0��v�R�Gpag�qmBv"��;E~߫ �4�tIH�|&�I#���Q%�����^׺�&Ze�-�S=�|��a��^�H�wR�УmT!I&��B�b�NJ9��E�J���O��<�K��N!�A�rֹ�b�'��6�Dk�׹�	2wB鵴;���HVu�:��dF�>�ٷ"�g�C?\�a��u�����A��?1�g2Ν�\�x@,�g&��[Z� �l�������I���+H�LN�	�H��V�D��㊅��T�[�n�y�-:j�U�;8m���N{���ӛ<��{s<������D1�č�F������!�5���H�0 ��<	YgR\E�ΨΩx����5����롖��4��Af�#)Z_Y=f/�$�������V�]H�$��nO��S�(�����UF]�������M�PH�N�	�M�t:4"�A"��<�S���K �}�@�H	�ؚ����x��Z�?Q�����+�D��3X��(ʠG�����ko[��'t_93��Go�*������H�U%(7 DPr���۵u�{?NT����v�	v��**O@z���Ñ}��i�Q��qk*��b��ƶ`N���Ԃ�D�8r�PM�1�ǯ���T��[��G�}:�\�|'l�k4n?Séd�%n
,�-b��3��ZVl��V.���8lNX��|<df�!:�f����$�>���$��`[Y�%��� �)�$�uS�q��|�4��ݜ5��i���A�ǆrڞ-#�6sG�gb �Ȧ�d� ��J2�y:A;��l<�W�J�Z/j�u�bo���f5�M�^�S /�u�O\��k_��RwM������{g�˔��p�+u �A�+4�߾z����	����!\�g=�'�r,�rSz\SP�p�Zx�Cq-W��^NO�o�V����v�������dۆЄ�z���(c�� ��_���E�Ó��	�n}[�<j۰�4ꗃ'��/��ԛ
��Æ0��C�gQٶwL�f�_>Zv_��P���]����I{l�j<k�5�!/�qp��=t)	GL����q>��j���?�-���	IGb�@w�Z��	�᭎���� �{1�V���ߗ�BkG�}�Յ^N�����(��1�*�$4���"W��[���F,��q'ы�n�?�ƈ�3��A��80Tf�?-�j�G}�K_����o��%Y3�2�F_�����nĴ.8�&���\gcΦɂnU�T�YĂ���Sg�Wu]2�Y�z��sÊ�|�WcY
�3hL�^��9O;�Z��&��̚�&�/Pb��\�0�.�-�)f�L�x-�{I[{�s��WuB)����_��=�/�bq-�	�Є�e�S�T)�H%���@1B��BKM���\d��+@�@d#�u��ᇨ� 0U�hF�/�|Db�b�k�f@S�S�m��5M"5r�%Kf��T��į���ܥ���:*��s�5�������H�^]�����@u�x� <�t���{!7]�c��T�dS��r �����,��G���ts���Z�^>Mx��/�����|	�H5�"��~�nP&p,������}�N�F��po�9�������V��ڧ.RN�͋�T�^r
��J�Z4�qŉ��P0\`.u�'���!�wAi?k�#s�����<�H0�F� a["�a��ZҜ�b�Z���Qw�Ӳ�JK�"ttv��4�!�D��hg��rF��<(�楞�(�$�4*C#����`+,U	��/�_fg��Y�t�����TW�|?>}ɝ��q=xK#�l����&�P�ѷP�V��UV���: T��2�{����s��YW		3��{�^i���rs_?]��k��;13�kҚ\{�>��vzͦ�?:�,B�s?Q��O/���+C���>�¨��h	S��5#��	 M����f��')x�r�
�S�����P�@h��dx�Z��[���_.�V����a�]F�y�y�Y�q[��m��Gv�w��� ��a/i�7���|��XЊk��6_2�n�2��Q4�d,�'�5yqy�x^�'����r��	ؑ��i�HaBg�+\�V��F�Q�l����-j��<03%����TwD;/.LT��J�U%�E��%l��zFJj��B�[�w�o��oG\�+�
���5�'�4ѻ��^������움P<�3A0���~T��'�tC2���n�C;�ᜩ%��(�S���cȹ�ʶ�X�C(|lY��2��)ݯy!����K%�����Z� ���;X��Q	���We���"F�0�z\�q��~����p��i���,���1r9lS�RY`���k���0��T����x��Z��Dd�/��?1�:B��}2��K���/��1���e3�K���QH����WHF��|�^08ћ�0��#ǎ��ʕ�9��,�~��^G�?c���5��(���8U�7 vS��Z��3{㸻Z��H�X�Ւ�.?�c;Vj���~cf����-�*�m����D�?y�����ݽ�MEiI���RH�>�'f@�f����8@����I�MS-�Q�(d��B�V�Geh���K%�~_T%B&'�v�`�}[�;�#��R�9��ű*��*�6Z�%�/�"�*�M&�#<�´�[�-[��Yg��J��ݕ�(�;�`'�[5���#��٣P=pW�~�q����	�g\7�+ԁ��,���C!6���	L�a��a����x��0]�}�TƟ7Q4q�J!��L�>W��U

��B�Wlyz�'\�)�'7����p5� �_�uA<�gc�s�}'	�4�y���R��L��u��F����!�CŒ�j�F�}�*���*_��~2;�ظ\b-2�\�~ׇ��/\7-ݶ��Q�#9[�`����\����%����[����y�M�2��RmPߞ���(C��_����_����@84�l-��=3�������81���SG��ax����$O|r�<�����<B���K�ωk��7f#�)��%����O�$��F�]J& P���%C�����l���KE��ZR�e(����)��_<(I��5do��c��Ԡ�B�����L�L�?#0`���}�7����MDXe4ϻQ���+�b���G��tCof~ݼ��N��?�$�½�G�C�����/���uB\G��~X_m����U0��!H�aLU�5*V�[{�����c�bEW�°��4'g��U0��i���DqΉ��v�vke�R�j��`���e��I?�1��%iH%o.��_k7Ώ�O����$�, 
�
���c������8�����1�a
i�pd>���+?��Z#��?���Wo�ے(��i�g*,TZ\%#dm�T źf���Z1$`��f^]���R���Ò�t+���'�s���f$z��/@��_ү�q�L�+��l��/�Se��(?$�z('�0�̪(�	�f�����ԏo��\~�����w�H�F<ݠW�/L��n9�G�ȣ��]ֻ3*(���؆s}���=��.��wX�5��3!��0=�c��(".���cZe�Ǟ �C���a�����vq3&�6�8��@b���v3��Z1.��gfl�k�$_�����*�,\��ꉱ�nog��&�ؖ��ʖ���p� �KnO�'�^�q�qy���2�Ͻ0ޥL%���&��mF ɒ��W&�
c�ĜJ#R,�I��oZo�Zs3-U�D�.�:	#a�Y)x�.?cV~���K��U�T�qr褮�m�<�L�Y�s3�#�K�y����(�l��:��౳PLUD�^�j~B�ث�x�ԤdB������-�]�ȧQ�{t��\BK#���2㷄2��#7Wˌ(�ci;��-�OWv�"zQd�&��X!4KW�C�.�����\���M����^�K��ŏ�~D)��}�r���C���6�`�U3k����7���=���XȜwt�PP�R8;�T�7q��!e���j*F���(X�	�(�SĂ����#���"��2��\��c�o�3&ݜW���=B��� r�vm)?�a���,%Iq<vE�b�)1K[	�9{�T��9M�E�|\�U�ga4�M���.[Lb��\��Y]�T6O��%,'�/��AgG�3\J5��Y!7p�E���FW���:��M/Y��WS�(*�Z��z���Kڬ���D��U*��j]��<��:1�~*3E��S��7��e�~�Hg���E,QD�#�Q�I����DB_]�k����,)6�����ByRUI�2��q^~щ�і&�*՜;�Ąi2���VT3H/P��4\)��?%�B��Y?���w�J��\�6<���������-#ԡ�5�����w�V���L{�ĝ�fZe[zZp��-�^Ų��?^Ƕ�	(�)���E�/-CK۷�H&4�UT��&���"3����%�ec/Y�1��0�����l�3_�~M�/���X~K�y�J Z�xbR�џ"@3Ӧ�OkO;�.�W�iG�a���W5�p(�|H��/6�1����������F���y�pC?�G�O�t+��6%���=sc�OP�`�z�R*`�J���\A�D��I�5n�G�X����H�����Z��9kd\ުތGm�gBg��.�
{9��(�2�0�e��f�V��P=z��%����;zQ��5�+���۟�v1U���� �$[�����x�?���@�|���3��MK��ۮ�q-U�ށx)~��p+��ʉ�47��y��*N�k>�c�,��Y�Wz��
^�y�Á�V��KZ�D>}��L�ۯ��Q/�0�$,;��4ƪ���3K!�WNb\܌������b/��SAȐ�Ń;J�r�0�໣ـ���t��PŌԆ���#�7�Aߒi���T���`B�0�!���`��Q��ga�"U����{��sW�^�#DlZ�ճ[�0�(X���	��bڒ�&9yz�&>��W����,��mEWI�`�r�,Uo�i5�H-t{�t�2�%r�c��a���?�{��,hi��S����@le2�;��������
.�Q���0����]�����WQh��\�"����l�!l/+��ΰX�m�k\R/y���DuC�?C����3�&1N*6ڝ���K�&o҆�7����z���Ϋn�~IM��nE���n� �~�	���IW�*� 9�7���{o
6�Iv�`Gf�p�P��oo���B�@����^�Q�Z����Xz�cDPB=��0|nڨ����r߿��HV��|�t��� �KRqq�*wU��&�v�o�������E\�i�.VC�'(e�O?�%��V��8S��8��l�v�/� 艋|](
j>������� 1!�M٥�`랗t�] !d�A�A?�I��P����N��Y5|��\�����2W(�nfuKa��p5N�K�ùُ��/�>Gl��� �|��T��ȶ�)ǎ?�-��d|�d�@�����B�������K�  �*4�B�[�F��P������_�	�z먼��)i=
Fb鎢B�'��#v>��捴�����.��*҈�`�?����EdAv��59�BQ�&F�J2W)Y���M�k���������G��MG�%[��\���f9�W;�����:a��Zo1�G{6vus�z�=~=�<p�;��g�����˦� II��³9JHv�+K6V����"PΘ�	y�ݵ���X����ݓ�w��ᙬ�ʿN�V�?�>qR��5'�<�7$C`���ƪ!��P��D�m`,r0��W�,yEZ71�j|�qv�ȿ��]Q0N�rZ��"���1��sh�<�5$�2���r�K�+l���W>��j�CI ����s�(]qt�iiGeO���C�M�n��^�@]�L���(!XV�c�+vep�'
��8� ��1��F�p�A���J��$�T��&�tR��r�d�PnK0@��EF;�I��{������v��'j�Pb�0���,�������Ǉ�K�5�5�X���
�C��ynek���0oc��(�2c{P	a��L���٫V��Q
"U��x�|D�9�1P�vE�����a��:.^hĥ�A��"��:j��[�[�P�'L�^J>���^P:�"	���E\zX��o��t�+*�Nf�(��hғ{VN<�h�g �9uӭIR�+z��G��w�%��dz����(�H�6�|���)-�FJ,��]]>;9. �Oa�W��۾`��u�+<��_x�s��4��ki�$Yn�6mre��&��}Y��(�s4�h���km�!헞3PvQ���B�G�2�{q�8Z��$.9�R�h
Z��o������q�t�O��25h
��44/,Z��f��M%���/g��@j>��dD<ry��?-)��n��J��:o�t��Ag;��&1�5��ܪ@���~��
FUm�����&�J O+�,(z g���J2�u7m���=��_���f����
�[��{���-�� ����YN��JA����.��o��M�w Y�9E��pگ�§�C�U���N����}/g�z-��\�%;!��!���<۸��
��'L�N�Rx���1������9X�شNO�����Q�TSP$>45��X1Ԟ�9O�6��k|���DZJ�Ӿ�22�v.u�Ҵ�nM-_`�%P���gP�ό��	2Tw�S�)*Z�j���(V����(G��	&���p��5�A�g���L��UB5U�)��F��/z��"L�?|���o�MS�2�7�����ʗ'����I�����D��>������Zgd �� g���Æ�oу,B�Jt��XO
e�
1+���ن6�$r�T�Gv;t���&���a=��H~��p���g�6���站����e�����}�]���`W;:�T)��Z@�#{iIh7�8�rr�F\�&���C�bڗ�FA|�<�1���ޠal!p���\4��}I���R���i���W ���<�k`:��`M���i��jm ^���~����}��R�{6п�zr���f'<�i������AJKս5��AڹB����ܣ�+b�D���D��Oq�x$e4�%��џ��2�������G��|!�&�ո5ԟ�L�z�o����Z���(�Y%b�e�7��d�J��^�����,�5�߷��Q��cd��qy��v��!pH�{0��ΐ�9���ͽ�����'��0�3�.8�EBa��j��i��6�d{'��$�xE�$���兖�J��>^Ayu��	Y�^�u���\�&Ɠ@Sb�O�*��u1Ӫ�@Q^QE������2�}"�C� ��5-q�:(���<)5�t��LX8�� ����kzրI�R� �E�g��k����(aΉ�e0P1��9��ai����=Y��(uKN[�,��2���U��c&���7�ij\�$]���f����W�'�2���;5T!P��pk�l���nwt����!4&*ք�ˑ& �X�g
v��Q1�U�_�#�����I,|cWƖP��[!��>�y�N>��p��dN�`mR�B������C�S��{�bZ)����� �ѫ�g���=�m�c��� ����Zл8IwJr��SPG�%�u �k�̯a�?id�G��2�\�L,U��6Ҳ�d�vo���D�֧:�n<�S].��L��-����7��WG��g{cv~���<��D ~.����O���'��'5�Z
;i��X�n��i��%��k���g�5��^��I�!�	�g�no<Ns��z;<�>S�K�����mK�����E�������
�Z)I�^�Ĩ�a�[\����ԁ-#R��3�b��`�M8�=i�͜��f�K����������:�8oY���$c�Q�\��c7L��T3T�4����78@@�63(t�	+)�RB�;@���� S��
�WGc�cM�
Y�|t�$"gI����
���s(��ruA��]�}�����=�^�K��*�g����CF�Ӵ�%1�c��R�)�S�uj*W`/c��t��:�f�z�C�9��޿N��ʚ�O�ZU�'�{,�౾\$ �e�M�	�p�R
(�B/����W�}�Rj����:�l��r���}3�d�Q����2�
����)�z�e&�AͶ+��\�m�^�~-���gv�
O����@�#�܎I���D�5V+�b�u��Op�ɨ��"ǘH��RX�Kn�p|��m�O;S&���{���DL{�RP��� �7�Ƃ�v^GI�{T���� �c�|c����g�+�M>(wPy޶�f� �90qK����W�H�B��'���s1\�K�rNg��ü��� �i���{05����n�t�##d����/>%�^�L��~5�I�0DZ��
*gyn�u�S��M���g����>��n=T���:�K$�e���Y�0A_y;7qK����1j>uT��C���+�ebi����
���������e��
S5��S��I�B5�kr�������8�2K����-��-��)WOZ��.�y~)R$}a����m���87���LNsV0_sO�ﭬs&eh��6��uP�\�{5���ͅ��٩�;�WO�����5Hcɣ����A{�	��w���B�V*.�����F��t:����Eu�>�[Rs�@�ֵ� ��4�2bD����+;��L��U#��##��NǇ5Kr8/��x���iR,��(!�B���lh�ֶ���Qԩ�X�\�����Uq"K���)[:2E�"�<ס����,���3�k�.�n���7_����Չcsv\�����͢��I���[֣���Wv*
��l��	���0��VMF%�:j���y����Ϳ��JA�b`�K�n&g�ӗ.bt���IX��9�dA۾�	w��@.�#�N����-�:��Y�����ћ��x�/�x����8a�q§��CV�XpI�)`��2b����<7ٵgh#�N!Ǡ�V�)g��b-��r/'�Y�����8=L>��2z[[�����o7�Ś��6Ǒ��xt̙9ta2fp� 9�8��lq$�o�J��X�X��޸�@,n���D"�'��vit�TM{y�Nu���~��P�DЅ?[�D%	�	 �:ew�q� B�9��v�ϊf��|���e�b m��j����Zv��Cz��c�����Ȟ��aHG���T��T�/N�b�Px�
�����;ۗ��5���ĉ;w���)chB�I%(��Ⱥ�8��w�1�C�qU��/��������3SPK� E�J�m������EV����P����Bg�u�����$�Ou�]�(70G��{�ݴ����.a~a�<��E�͍0C5�IT��f�}�d�S*-����챕�g��d�9G
����)R�
=�{=v�M�� &���_�����K׾{BY�J�	& ���×Z(��e�4�A<l�ڠ�5e���@�4���\+�߼�IH��*��y7��ãV���;Q��¹+^O���ѯ,''�M&�Cq���+���5F%^��������쓯vA�x�z�+��ߢ�����<�=ヮČ�.v5=���p�U��c1c���)�Ι]�qb;�����H�)��ؕs���4�ӱ�7U�d�|�>��3�\m�
�Թ���?�@p&�� Sw��?�\]�rF�{KnP����~��`+J��=o��4��m�r{<d��}'D<f*7��)�t��6~��"��N7{��w@9�qh���A?��K����M�Y<k��(O����c�4�aSԝ���C��
-U�o��ĺ7ˠ�:{^;�^5�bcGg�R�4�gޞC���	.r������y�=������<�m%@f�$O1��X�mvR5��V��v�qإ���y�"��B��u�E�#8՚
��O�A!�l�[�/�y�v�����،	ԭ�H����j4����S�'�v|bK� =�#�ePF���I�A+�-z��e 2�_y��ʏ���Oe>Kdw� v���VtKڊI�^� �Z����Y0�ZBb�`e�H�k������G��y��kK���^��b��B)�40����G*Q�����P<�D}�uFU��@���+���n\MZmB��,���=E��ȝG�h��
f���GK$e���|0a��^)'6S���U;�:������d���Ќ�����x1W����k+zw�5�!�)aJ�}Q|�B_v�Ciaߩ[��2+Pn�?ߵ�<�z�����*�|/��S/�W�Ic��(������2`��')��	�u�.�^�F��vs�<�T��"�շl��2e��z���N*���44�Ձ�ǩ�0+�������!&��B�������p����r�,,�0>�=@F�����}*3�"s�0/�[1��r�,�ٴ��\��T#h=W H��Y�S?J�î�]/�#�6!3�#,Qg%�Jb7����NLyh�����Mt���bC�<�km^R�"�=x,ʉ�H�Sal�C�VGfȺ��bJH��2����J�7sTB&F�$ic��Q����ݤ�����f̎�����>��.�����zW������I�Գ��T-̡�&���U.�f�W�z0/�=�F[�~����;f����m!�����؏���x�w��s��6. ~��=��4�����R�����=��//�`'@�ln��x��˷I*-�4�z\;,:W��,������v�u�]�t��@��Oq ��q#G5���{l������]W2O�~k��1�Sy�
�-
�<��vĢ,�ʆ���	n
�;��,H��&�te��������Qv�����9��դN����H�����ye��7��_��^���S�Jw�'�"�U�SȲ���9���d�_|�wN�@�i��ɣ�nM�N�+(��g|p�l�JM���e��zi�Ke��w�%R_����CPnC������TN�x�	m�Ϗ���B����iR6�)�)	��Y�u	*���D�0)(V�6[���F_"��ĉ���ļ�DC����q��eR#H# �L6��Zy��M��z��̪1�2.Yr|(��4V�Dh���J.gԼ�N�ϑ�=ψn�G�t8c�;WXE��̹P�����'T���wN��G�6�~�:i7�:�]�C�6�`�y��'����ow���g�*˘�cx����S*�����=�Sf0�},�����RI"��� ��hC3������ ����~wȽ*Q��|Ȏ	Md���D�8�����u�z�,�[�򪆇�O)�7�+:~k���h�"YYt2�|�o-Z�~��_�k�z�4�g��r�N��ʦ�;x&�NƓ�q8c(�F`��D
�P�g-�
C"�J(��
G�@�+������s	6	&�7D{�+�1]��LzQt�:k6q@�昃�F2x�x&+�9���A����1��o���WA��e�Hоa��2)PoP��~�9�Pa`����f�	0IXDIH��?���:|d����$i���l��Ǟ7<�)|��W��z�&(���쭀d�1�X��f�df.I�D�?(޸��j���FVF��A�SYb�ss }t2� �xO�]�,�:�Տ)	�j%�WN����O�| ���|t��EM4
�����-�U�&h-��ݻ�B?���;�/v��Y���ύ����R��� if�Z##���/�t2�x�ƨ9��v-��	_��A��o03�8b���9���q�,�t��\ޒ�����h��3E�h�졪7!�+��>��x�SP�%���1n�e&B't�=dz�C�z�b�؉��K��d!�%l���t��sh8��k�nF���g�|�n|D�9?>��u?S��D��ۦJ��䃵�~D����\SWp¨�1�r��	���K_��j���@����W��&и�0�=�m� 3X��]���]v�+���
��.ʃ�U֜2m�����/����vu���r{�x�����e)�8
B���%�E⃶�u���mj�̡���˰C�L��3P�Zx�����5"���rI2��k�x�%EOL����O�S�%W�&�!�غ���֋�	K|���E�,���^���ZǗ�z�|�|��������������a]m�@Q~������F��U�3\tϥX���u7eyݯ�j��c���LW\rmvS�R���~ʳ�ѓ�d?���1s�P����t�@��t�8.�3@��3�dl0��ʁNp�d��䅭��T�WG�dF/�l��:b����4���*]0*���W+����bc��M�B����h�7�_�����6
���V/�(��zammθ�2�O�'��H)�W�f="�l�[8зh��V���^��s ��w���͞c,W9�8�m���GG���n�-w���5�"}W�X�RV,�[JX���joC�J�p)�b�y�7���
7Qi�C�=B%��Z�e�|wocz�8��L����E)&l�Al��C�m�_��qo��[j��n��
w�F��N�p��8�ੋpg��'79Lv��K���R5\5�e�,��V�Ӥ�%�z����?�E�Q��!5�ĻM������-pd�͏�_;�	d* s����+���ל�P�k���7�>jtƘ�	F>�s ��e%�[�1Ҁ��Pb�@p���P�����n�>�g���g�
L^�ޜ�G.M�?xxF��S�.W���A�5��5���v{����C�؆�@c�u�.w!e�xar,M�ࢇ��g���0qe/^#p3(�f���JY2�*�R=��
�x	�e�,<�V��=�Bm%kǰ��X�E\
�ŷz|h�M�U�:�:שD26�段�S$��_<��Ò�U�g���r�v�F���d�!U_��5ݪ�(R��1�7-�����G�%��LfPSYC�iL�,���(N�x�|�=�k��3��W{?e#s+�O��.��5��5!�§]�W�!H8���,�*�Mk�];�K1ѐ����OkTa`�ݥ�ry�cp�u���
N���d d@(<���8N=���͙N�Vԃ�6<#rG�`��j�Ƥ�&b�֜�f��}�Cy�u��PB��-(��PRŽ�� Y�2�7���
��߾�sT7^X��G��(�ǂyasg�a0�n��7
�S�҂���6:�m��h�i^���ZZ��-�r��4w4�[o`v�75V�g�h|��L��@�&Hæm��e��ںh��}�a���ѵ���(����@8�bz%��;w9�[8��K0��g�B�*��=��|��yp�՝ˮ�^b�: ����2��`��r�<�/�|�Ζ,*d1�^�#��[�y�\3L�6cd�����W�̂$�/�+dk�FJ6�D\{+��B4�;(��)�W؟Ӊ��}s����*�q�;:�y����}�/�%�D ����|�	�{��N�b9�_��l�1��=��z�̮V_OܷOp��*f\��3!J}��~J�:�lo�+�ALE��B��|g�����(����=�p$/�M�.��4BЄ�م���ʳ��.��:HQF:ژC'�r��e����)���E�-�er���ۊp�L�޶V;�$��+�q��zӕ�n�'��K�\4�V�>���,��=ɐ�q?[9���v�܎��{駁�i/�������{sc�h"�������M1�NI��I
г�u#P�}�"�oF>��h��V-9ܖ.䟼��,��kX�?>
�M��7)��+9F���F�|��4��*��t�j1�o�r	ܫ�DQ�
�ڟ�]Ű�it��i�IH�o�!��xT0z�uUb6�������t��"�ƥ
��su�ҾY�g�����k�� ��"��}�<�_Zu-��D]c�nrO��N���ԴV&�ݓ���J_��:�/p���eg���;��O�)�h*-x���Du󠾅�-��e�X��;�0��o ��ר~rOz��
�t*>"S�j]su��n���J�m<7�^P�����ir<���x|�n^�aըx�Ɨ�"u��`<I`a�kEW2��d����Ò��c}�V�$��&�Hm�
���wXLM&�Y$��I��ا�r!�+"�\H��Eo)�R0Z��P?���M�Z;*�����s�[hqV��0��%%�L���?�h}lO��&��DW�Ҽ ZY�u���Z�����ַ�77rKC@#��WKJ��	0�dKe!��|��nԂM5�蔡߬Y���e据(0R��E!�_����N�[� �8���m-w-p��+	 ����+!�!��x��w�%�z��ݲ����fd��Z��ѱ���d:	\t�J�e�vU����.����т]�^��rp}�Ji�M��X�we v?O�yt&<b�`,�c��������>��(��Z��E&n�ː�U��Km:BG�5Ok1=�,9���e猑fu?�`��?a�\���$x�i!��7ҩ�9�e~�=p��l�!:C�K���1
��0����c}vR.�������e�S�.���7�Y����=�r%.��]1�����m��R�r�����܉��\�\�)b�W�EeQ�l0v�XF���$�H�>�+ݿ���Q�,�7�8#�0}�z���Ip�T�ڽ���L� ��HR�rd�u����H���*����}�#�@��?1�~�gh{'gSW�{nB��X�;|޻��A���<U~��U�w��u�C(�m�~14��Dy��M�#��0��m��I�?�ະAR;v�R��[~a���O���N��>W�>���>� ���B9{s	uQ Ͱ8�.��@,�ĉԝ�z����ګMo��Itn̕~w�ps?S6�ɲ�l;t3:�𑦙3$�Sf�[�E���E�5�}��f��j�[w���C�.rQ��9��~��z�m�[PP3��p��㊸A�^��c�	>{\���a9E��q7|��0�;id�vkj_��Y��>���11c���!�N�w�h�X-X�d��P��x��Y�lkg��f�G��-
O������p��k ��[��)�0Ԍ�7�
�a�w��ub|��z����K��
�m_}��%>�\x�y �"�(*�SOoP2��ݍU�1sp �8���0<��A�
�'����7��^Ct# �jY�6N�߂���c?5ɚj���yaO� �B�ܤ��ov�M�~!%a�a�L��b�9��n����
�ᆒB&���t�4w��N���R����Z�Ad��:؞7����ݝ�i��A�[���b[�T�[u�A���)3������b�v�l��Ut}]�^C����؝�9���R[�#ƽ��Yh��Y���{�����@�����v%`r�~@D���΢TS�l�A�A�K.t����r�� ��DrA�-Und��%)N��WO�*�0�x�7��]���]�u!���昻�/�&t�G��ҽ���a�kV_`	�n��˾�z�^ꞵ�Wc,x���/��#�mM|�xSZMZI��tt
!��/خZ�ć
���K��9��<L��v�>P�~�7y��(��:�A���z`�6���,m|$�f� U��5�%��%�Vj��É{~R��7N���^\VZ\a�1���V�u���M�$�U����-�a4�	4n�÷���h�}�ԩ8����2�����@���2HI�h��-�բL�*�Z��Y�ʝ�4�غUUG5wT�96�$���n�	�!�CF�un^����޻�p���#��ݽ��ɖe�@NZ�|i��٤�D����%&"<�d���<�y��R��sU\y��R��c�{wr��	�IQ
��_�v5� ۹����ԲF�H3��)g=�N�%�uu,����TC�u��go�A�`V�&�bZj�Yku���̪YD9�%[��8U�Ǌ��*����G������Ѱ�,�d�bďK�������C{� ���կM��O,�ًg�������|j�XͲ��|����A��8��� �[*�|��B�Ld�c��ƛ����I�Ѡ򑿋��D��=������ާq�_��W�ǃ��m8*�aآA:�0��Nѓ���G�X��ܘ\~(c���&r���Np-�hs���&�$�S}ԭ�H{�#�&C�K<��I��g��C���*.����^1�>��{��t��,�`p˺��J6&2� X��xL�Dr�K-y9~��d*G�KJ�A1\pt��"/`w/�o>Ei_���@}�"sߌ=u��!�[mA�"�����e�O�'yh��|��~��X�'�E^\ޥ�~p*9�켯P�+��=Mu��˘S��1��X?��N.H{A��a�x����!*�e7I�"�ͳY\��R
��� �-�X��� ab��>$�G<K&]����3�Ո[��,lћ��5-߄�@-�p�\L���t�Oc۽�xv�?��ӎ�Z�4��UX_t)/�a,��Ӯ�C�tH�:O�	�&+�l�Oa�(=�IWN6i�]��p1K%wB�+(�{���؊���*��7b��~\�8����i@?�29>+l݂��rn.*��h��I�b�@ۻ�+�x1���x[�Pg,�����'�|�V�a�EE�������2/�	(�B��9F$^cCE@鬂���^�{��+�4���"�����s%�ؽ�f���k7O�?o�=�B�K�o��݄�&��׷��\@%��@����WJ���-���|P�,7{h���E��	���q���@�e�m��T��bt����:�ʿ�T�u����bO�s>�6X�&lW���i�1�)�9�W8^��� ��pJ�;¥�}�pL��"��gF�mgG��&�2 <�ۚF�"��V�b�i�
����!BG��E$�6|
��Vtn =�Úuw���
������_�!0�qcZ�I���[#3���e�g�<� ƜիK���[s�n��L�4��l�����]0.{���jD��P<�j�"��(�<�I�y�(���kw3�w�X��N�ťo�
�����4g�C�l�4;�Q\<)�i}�����X�g'b���%�?l�
׾6����g��t򓜓�A�(1�I�5���g&������Hok�\;�f���-��(��
 UF�C���9<SdIy��:���He`��,l���T�S�4����h6����E?���,���w\Z:����0��ZQ�=��`H7d�"\Yb��f��Ά�y�dу��2������KA��\b+ށl����шU;C�OXG�y�i�����	�&q+����U�9PTQ��R��N,m�4��Koow�x�NEJc|���YCh��+m��2�'���%��ն�O�������-�s��,AR�{"���Zˣ���	P#k����[���g����ĉ�'<�M?��I6�����5�����1an��8�`�m��J[����\�����%a '�k�={?�}Q�o����6�����/�M��|7g�!��y{�����3	��
�!|�>������[sN"]��k�4�(��y˹ܯ�?n<�V��WS���Ԅ�MO�z�U^] �?H~��rl����[��5$��j��a���I�IVѮ٭�F��V�JG9��e#�􌵈�}���g77�R���~�g&OfE�6X���fS���?7�Ϲ�M٠��r逛\W�����&4�|�v0嚓����D̝V��{�L�C��8���3���}�$Nf��կ�{�8�'��Du̥��$���5狈S�WM��v�(��9,�{o^Y�:��ө"-���а�sn\�H�,Z���
h�2Bm#�G*��C���4����rJ� )W���K��(w�2��0�,��`�[�+�b6�x����yrt�;�(�U�ݰF�����!q��V��u�G��ņ�=_�#���_O��<��m�G�[�^�VK5Ɏߋ��˙�O�O�E�؝�L�,��~�hM�Ҍ4����fC��ڔڳR::s*F�9�c �LZe \��ȣM�E���nK ��ϓQy��X�6?�-�m��d�D��𭾬��"�y;�P�~r3�,�|�B�}�[�!Z�|�u�<�B��} ��[�Ę`~�LJB+�}8<FE������#M9:� ��J$��)�ryxR�چC>�K6%%m��{��~��b<��"�پ{|a��e��ƌ��=I��G�גP�M��AI9�]ܨ��CS�3P�*?c��b;�&"$����FuoY�&��:�L������Ơ�-��)0:��K�~���*yб�]�j��B��b�©#��������|�:������,]�߁NX�O��ΦŸ&��zz�骧����d����=ɋ[��� � 31�H�.�v3��9���#�7���^���sR��\]~e�1䆐�ŪM.,�M9 T�������������@Wk��`��ۇ�8e��"a��#CT2{`�  �A�,؅�y��НVn�`�xIw��#���#���rӿ�������љw2J�W�Ҳ�6dC۽$�?����B�-$�2�=�z	�S�(�
!������?�kg!��_I��'+�����<f-�х\��ߝB�����W�50�Q�d���6����R8"����n��ֆj�I�mb��L��{�h�,iaњo�+'f��'̏J7���jV��hsy瀓�wOX8�Y.
LmLax�Ոyܕ��#��]��ϾK���S:�EagU]�ɋ��Oѳ�XN��:E�(g�s[; ����%���*�	�M���	g	 @�}q*`�{�� �kZ�������w����KF]~|y�W�)�}������h�<X���mtn77G�F�$\KZ�Nq;`O�m�8~i�/�a�6����!�ȃ�/jb����+��-��DB���x�;�v\�N���1��A%�\�D�+G�Wa�1�sN�8���>"�؅������rE�� %�;C�ˆyb��6��Y�3�ۺ7��� ᛊ-�y�����o����n� Ԑ��ҏ*�Z�b ����Y�����fzbK�:���8���ӉF�^��?�|�ajԷ�a��ɡ�?p+gUix��l��pm3����b��u=�(f����a�qt�})��>]�c3����=��u���a��6i�!�I��~�xrkql5SG����!#3��8]�{;��t�e�L*.{�����bV��m"(��U�u����C�"k+��G�,�)ƞnf9'
0���l���ҏ������O����L�!33$�pw�Y��xhOaU��I��+ԦS�6X��/�;T<�&�'���^�~��ET<��8E��8����>����D��ĖK�eǏ��.����n�{�3�g�K��E��h���] J7@�Cm}79!^�-0�z�-�I�-�g?�e�sOX��
ZW�D�G�¡i��g�c]�3��Q�S�@nar� �f�D���l��A��9m���f�p��[}�Zw��h�G����U�E�����x�mH-����[�#��h»���CG$v�}��&����q��uR�\;���g�8�\������L����	+7�c����m]bT�	E	����Vi�	a44�����v8nE�I�$!4��72���ӊ:el,�i��(���ً`�����f�4�7���qٜտ�c�)�y��26�o��N�@�蠰~f"���ɮQÞ�FZ�����傉��Be�=p��z�k�[�G�z�+��=-��3ߙ��pI�R����1͉���p߃a����ܫX��6���|�zg
ktѝt��d/�t�m:��̈`�9��3��±���+���,��r��S���PR�VbZY����4��a���g���˦uW�c�������-�i`��k_$�=�NÉ���8!��o�]�1}�����2@r�Ȗ�qO/���\Ӌ�T�m�� -�:?�K�̃�,�T��VF�c~�C����g �
)"B�#'a�ng��{�6��]�2�YԱxCE�o��I �㴠� ���/Cv���Z/�l%=�M1�&�� Q��4�+��!��잛7�9�� �-����Y��<m+����	>7R��>��_4�`�r���������K)*a�{�1K���ѝ��^���|�qF�����TN���&�XBE��}�)=�ߠ��$�n���,���eE�^�?o_&}�ê��LhÉ���j�bs��#Ӣ��W�[J4#F�C�H/>b��X�2��
*�Fh��:3����zͅ%~�e�2��7�NO��Xݙ�k��C�E�OY�,:Ձ�lj��\�|$��	�sIN�
e��1�i�
n��-�F�ط�l�ז�yX޾ 6Wr7��W�m8cu�C�Ŭp��Q�n�Y����ԕ����=BEJ�+��Ob���JU�I�r�
U���?�7`pi�����0�H���`X�//)q�|�Jc��Q|,�9I��l
9�v'_���M�}��J���=�V��r*:̫�)�~[>��7�^?�F*��Z���);�B�a�\�x�C�k�a�|��fM���n,�����s<�����cY^/e�ry�.FX@,�?�����EvJ׍�̫��K�_�N��!i���>N�]
�$?�q���	�2;n-9>��~��\�$��Y���s�^�)m�5�����eEy��`!�H(��������G�(�^CgV��XV˸Ύm��5�n�o5s��{A@N(�dǥs�yʙND�>����Y�4��/gA1�9+anȁ�����|��h� lX�Q��ࣝ��ۂ�A����G�ͮs	��QЃ?����i�\�������I�Te����PO

4
eQX�G>��d�f敻!2�u� U�@/˨C�Pt��*Dҫ����a9<,�,hZ'�(�I�wHG��Z�q�X�������G�v��K�,N�ff���n�d�� �zp���Z�e04�Q7��$��8�c#Ѳ��IJ{σ�"W��C�43K��th�V6�g�Z9�nk�2�W��;j "#�b/�FyE��ລ�R���W��5�.=K<3G>�D��"ndT��ע �u�����⢏l-�,�k��@&�|��YC�#x����$ty`!#�������D�)�_k�L�}��m�y��_p��:В��Ȭ�<��S F}�s ��IS�s���qi�P%ȁ��w.��>z����hb��O�~��΋��N����^~O�֌�'|@)4R[���|��A��~��yi7�먒�9�E�J,=���,6K7M�g�%�7���)�T�,���+�{��&�V1�Ћ��I��Qk��{��U>.b�@F�;3����&��m�g��M��;�!�v�BX�U����P��6L��j^_CE�3]�Zy�r��ֈ"�����a�j�h����4��ZE� JY��8G!J�.OJ������X�k@}}�<7��^&�7ԞBv�;��}�m�.+�W��lc�7$2rLd�����E	C@U��aYjPͧ+��������C��oA�!���Cv�C�w��վz��r��Ҝ�W$Bȝ����2�=z���?}y��?|Cs�53��[����� �D�?ſ,xM���`�®?�8ۉ��O1e�F&>��xwM�z�����NWդ�Э�_�dB[و��e/��v�WX���K��\�#�8l��� ��iN�1���MI��=��Vg�+�ڪG�RL�E� g��΄������l�V��o�ޫ��"g���� ��"�!02Bם\�zD8t������?����j~�|'���;�?_re�$=-(��{�����\G޵%�U*i�~Ҹ1N�ߖ���Gi���UL��U�;|����oA[�:I�����A��8R�ILR{^���o�p���lM^�ܶT�x_�s���N�uZ��ȃ���7����T}�M��Z1������x���6�; ��  JU�Q�T<���L�!e-49�J���GR���>��sI�k�/�eAU����F�ykF9f���-M(|�E�,��-9
l��P26�y���v��\�q>wJ�&޺�Ȥ�f�.��c�I���O���i�!۲&W��\�Ao���.[ (��y���U~r>̢�L�Z��<t
譀�w�Y
k��8��X�>�V�z8 ����dgi�#��t���uɞ�9��ʲ!� ni��=�a�v�~E�/��ZB`ڶΙC6�B	�Nm��c
|?���VXU��w��!@@q�ݾ��ԩ�犛�W ��W��9a?���Fm�J��[$�xC�u����qe?p;�Z�<����9KC���o$�7�O&����j㞵��RT�跗<v��T;��s���!�0~7�Y���vݧ2�i*oH���%&��Ƶ��;N��eT�>��'>�؎���|Ϩ��C�r�v��<=���i����@��Ul��6Q)��Y�d�����}�T�����t̷�:�S8��Es�"e2��T��M����8c?lKy�^F]`Y,HRͽ��H��f0v�[3��EDS.�p�ģZ"B'[�:�����ܐ��@��0��6k�D���7'��{���)믎Ȯ"�.��@��t���wK�88�Z���-��[~��卟�x���8pPz����؜ww��p�;�@���<�ſ+�,����\nG���7�	��|�b
 �Y��[.�I�r�hA��f��q���e�5��л��퓎c��*�Ϲ��_�ܶ׶�Dgz=R�y�8\?ej+5Bg�P��O�I��y�a���j�&6wo�s��6|��Ո���3>j��/������ʳ�?���a����H��s�QE�� �<x�d�������6;`d��{���nZ���g(|N�-p໘���_j�<_�l5�0��T����CgX<�)
t���U��ԟ&�v#zNz:ǽI����-d3X��N��6�ڜ���o�\��;�^R��X:�ELЅ��~Dg���g
���2�|��q/�	:�ʇ�d��/z��XK�oUH����%X��ֵݑ�w��y.S*-_�l2�3>Y��:4����ޗ�~(���Y	�<<'$��E�nOm�#m���t"�h'�>�Vt�B��EQD�����9l$�j#D�&�*�c�Wy����(h�5��Y�qgƭo��#�!��ڻ�
�� sɡeN��m�S;�l�y��pTZ#�k!�4��Xm���QAܣs��KˮR3���s����vˏ�/Υ�\��Lj�p�T��Ӿޕ\Ai9��S7�=�~P\��C�s�=jT��jr{*vR��خ���n��v��ך�a8F��2�."vQu8�\G! �����I�@fJ+��'��#�Q�F�8C��3)iڹ������jy�>��񁑯�!�S���$,r~�B2+̏�=6C*x?�����M�x�(A��e�։�ͷ)�z�SE ��8�!��}F��C�����O���Q���tg���4:����yɉg�ޕ��D]"B�O[��?�Ci�ed~XDܵ۾�g�0���}��W~��3�ʟl�/��ڏ�����7�oF����Փ��� A�J�@�:�A��3m�͞��1��ߝ�[�2j��"��Iu���O�7l�̨G
Umj*(F�TbWʒ�lp6EY���lE�O�3	�-���'��u��=G>�o��K�S�(�����A�"�Ӏ�a�͚�,�-�RΓ] oxLE��m9ꤵMCMÛ��i
�^F��A� �����M���4z�h��5� ����%�~��-�˞�l��N�O"�t�6�Ǿ�D��W�K��y�~�wvm��\!T��==R�V��'�<2����r'�R��+����X��3!�?5SRܼ�>�����&~yJ��99�fɵrT&o@���� �S�D�Q��Q�*xs��E`^v�<UK�y�r3�U�Nv��,,a�+���Οּ��4�f�9%�`ɣ�L�bN�j�s �.�+��]t�������r{�x<�h2�3[X��>Y�f�L�cq��	.$}�}a:�Cq�β��1("��������n�u�ɵ`��"sM�]E4�\,���`��9Y� ��/,ݿO�����\7Z5�qN���Ŵ(��4�׊�"�������T��O�c�*�k#c$���%�ϱ��4(�2��;��P{� ���J"�=�	�{G�[������2�9�m�c�Wl��&����)>m��*�L�v|�j�2����QY���l��j,5���\mx�g)yQt�]q%�_#&���_Ȥ]���?�{��7l�i����j;[聹 M&GG���BĈ�]m� n��#�4����|]trh��ٸߡ�6B�8�>�P$�º;�+K�/O?�#��w�����-���ɟ����uX�w��TrZ�ƚ����<�������t��]z�*u�2v���qq.+�-c4�䓍(T�@��x(��[�YP�Ly��[�AW�{����I�d�����)��%W�s�*�(��W��:���Ɵ�W!�24y�:d�u�Ņak���z��9��h7k����{�R��{����dH���!g�?ٜL�8s����wz���1�4}�?���#ʮ=����lث����`���`�
t߇�+�D�{���껾�u�ȇ���*z �sS������_nY�xO[�3D;y
��%���@��� _�I2�n���lq\~L�~���<{����?G`]A�+���&
hJbcE�������8�8�4��{ux �w6/�� �c�wμ���F���+���|߁�idh��L,�����uM�(N��
��~��n���<���'#���ĹB�j����>�$����|��"+�G-Q���y�|� >�k��	��#T�=������w��s��Ф��`C˸�ӪdQt�"n��a��#XL<�0��b�ȴ/n	��G�Sin��{Q��h����Ȼ�?�z'���}/�-���v�q�YnS�>:LшhF�}6��|��K�����4����݆���ģc���%�dOS~��G�I�%�#Od�ڎ�Qp�\+?�8����)
�H��h�M��O\O:4Ay���Jʵ���ej]���	^��ȿ���c:Pދ�6�'L�����t�!{P�g7��A���i�1*/���O�5�n��4��|4P㻭ih�G)�-�+�	��G��g�3�wF�d(���J�~lX��/�Q�ߴ���h�rO)Ϝ��d�!Y���33>Swu����Ē�Ŵ�j �r�櫀7�;��4�j=I>����WQ�.6n�~�P5��I�.ԭ�\��쯟uH�!�Ӱ����(��~�̬f=�p�}��i74)[|�(�s�VȚ��xve����r! �j�kr��$"@PO���x�8\D�Li.�*���&M�u�������-QF6jܝ��H���"-�ۧ����䈓�p*�AϠ�H1�s�V :��
`F�e�'�϶�8$�1�V�C�?��L�G�[x���������4T�s�K�G�7���r�s,��U�NY_p��_B	J���K�a`z���Dc3B|�M��5I��&��6�P�R�f0�tk\	,FP���v;4Z0�DdG���)����'���
d�Й�q�c�Wۃ��>}�sP0��]=�q��<5�;*- �Θ�u^������� �EW��KO�$\o)NOd7�m����e��:�Z�G� �B��YH�W�b_g@�[�4�=/e%���tv��<'K/<s}���^�{/K���]�KC�1v��h����i-�iʌ�u��0,P�ծ���c�Ǳl�szQ�|�I��YL�!X���K�_�z*�����~�|B�)��}Q�}QV�[�"���f(i5�6g�r���{2��Y��ӓz*�8`���[�)�\�ٔw��ӥ�z�h�W� {�媐վ���������L����O�7kZiԃ&��ʭDE2�M�H7��Q�����&��n$��r�q�.�vQ�i�O��.Pj�?wz�έ���2��r��24��������� ���������	�G[�ш>&�MP���5K�)�2��Q��<�xբ4�'`ip�b�~��@c�K��r�&C�=�<�����@
�7؃�5e�ʶ\q���2��h��z���I6 ��*k\G�
,���d�'l>��y�B�0�]m�:�#U���<8x�V~�x|] �^�ԩߨ�U�9�//��`x)'z~��\ښfT�g!%�l<N��\mɢ�_���<�f rv��ҷT�1ev.�)�}�P5¡ziewG�Y�t�E˩��mb�m�%h��5� q�?�7�xr�߱*�.}f�A})�>cަ1�&,�;L���(�.�\H�m\�+H�,Om��0~v�4�m>3���۲b
:M����������	�$Y�)�Y|�
<7�����M������F����T�y��ҹ����D�����p�
�j�������|y�	����m��PE��Xȹt2�m�Q��5�@aJ~���{��d%Y�Q�g�BQ2�Z��˵ߋ��F��A�^�j��ړ6R&::��U^�9�B��]�߿�L�U&��������.�U�v�w<4+I��O���/
��]�,o�Ri���g��֣��B���o���n���m<ߜE����D�N�R�������?Ê
�G	�����GD��M.��(�ȹ�Q�]�]:{o/6ǎ�Hbi��/��:��`2�(a'u|�\�2:�׶O��A� %�d���Ғm^�4�h���>��%��:i���8ˣk���� B�"�Z5�&�0��/Uzj�A^�v�:GK�kvm��i��'��^�S	zi�=+�~��Z\����+Gt1H�a�pc�����T�éhTht�Q����T�0�J��{w�.3%J�(�����G+�� ϋ��@ԋ�/42y�z�����N �?�,�^)�����z*�����|ؠ�Cc��7vO��+��FG�t�I�yNc�����6��������)x�K�_���#��P�~ |`W��r�PӀ_�77����d�a��Bv�������[�c1&���w��1!���Q�]���:�.�ldH萤M��_�X�mK��6��e�-u��`���A	ri2�+��NA�ځ��=��Ƿ{���NuLze�@U�X�+�VQn���ʛ��T1HͶa�K�=~R�q��� ��L#��q�q��~b�iJ�jGS�=��;�U�G�ʿ��V�^��IG���kh����ٔ���Qϭ�G�H�a隤%:l~8Q�ŏ�0���}P��O��BC��G�'���� f5�`�]�V��{��qqe�� ���������ӑl���M~Ng6&�'��.ɴ�_Fh�o��M��r�@~��u�R������тD^
���ƣ﹕㍷n��oV;��h��w��ܬ1���$-g|�X����}����|Y0������N��[�l}��T�)���@D{XP-���� �n%.
�a��b����<��v�
�]�e�"���R��-�	ɟǄ������I�)�BE35T���&/]��BĆ*�Йs~Z������������s'^y$������c�h;s��O�����'�����b:�qcف���M�����^��Ȋ��ȭЅ����RT���+��>t+`��T��N	���̽���i�	�f-��ج�YvJ'(#���t f��Q�=|���_�_坂Z��8Õ:^ݞ�6����}��`5Y"{�S�h��w��1(D4�e��<#��jj!��a���sώb����k'��g,����ſ=~���ސ�P�	J$�4�#~�֯w�D)��]RC���r��5K[���Ϊ3S���Qc?�ǁze�ү���d��5Χu��ёs��i�� ���dGA$=.��Ţ���=yqض�8r	�E'�徺]�m�fx�x��IEOj�uf�L�j�P��/���_e���gC/�E��ф�CB�b�fv�<u㓂�k���W6�+�q_��]���E��MvYR��ns�0C���o�Ň���	5i��j2��ۮ�w����޷��X�4%iĵ��2��F= �����]�y肳.�����੊���G0��y���Tit�I��N,����"��Yy��"���,f\4���+u�_If�W"�I����?�������P_�L�P�rUFΣ�<{| �k���:a��Y�bK�M\�Ŕ�F�Ķ���^���{3Q�a?%��L��_誰CV���:ck,�4���o�WO8�k"b7�S�����`�AgC��"x8@��U���m�l%x�h�Z,�EU�G��Zh^���1#1�Ā5C(e���i�&�h�a����9���Ry5�[+�$ey�[�CB3�Qȝ��@�=o��->GA;s�b�MO��;UE�=٦?��ە ��#	��
;�W;3�q��������M���V��'Q�=u�Xù��'�������aXjP3���-�p�H^�bl�qܥ�M)�+�i�F����=�GSf�9�&�ɐj�5�����\t~簶����2�_�H�<cF��cLX�tB4�|�jz�%(�~��Hj)���66|"5kĕ#��A����DD��L��3M�@��J�1ܸFr!����1�yh��ԂMu�k}]�KF��+���9C$�)���t��-�'W>��qۼ��f'��kR6h���
f�G��˖��������X�e�Ғ�K�`�Q�(����x�4:9���E����#�
�X>Qi�,�҅UD�d�袥�� ED��3;N#R��[p�w�.h����UQW�Q�Z����b4g3];��cX�������{̉/��RM�I'[��S�}�=7��Lx��C���yR�6��# ��/�7� H7 ��4��(���ԕX�c�������W�u�v�E�u���c��4j.Ah�	v������{�#+3M� �u3��-ד��F8N�q9�5�Jū��a��	4?I�AyN]G� �p�_~5Z>T)9_A*wĜ�O�����W\Ó���GN��PG���ׅi�%z:���/c����&�r�����)�TO<P������^�p�
8��2Qdc�a�o_���f���t�=�
%�w���׆ɞ�*�P ��_�_�t��wc�?Q��{��o;��nx
Ḥ�Q�2=&i��0�z9&LI6%+��eCY K����w�>�D�O<X��J6dK'Me���j�E�σT˸a�-���-�ԃ�I���3T�p��oQ׋�����1Mj��"�
��c����5���0ܹR7��-k%�k<��%@�?�������´������f��>����G���_���@�b*8��e�����Òs�����,x�o�ҙ�+�pᆽ}1z��x�۽h@!�+Tx\o���Wu@���t �����_�"ղ��� �������X(v�VY� !��uX5)��|nv]���]�S�8���}���VX���R�<�� ��W,�o�4��T��H�O�#`�6�D���:�}v	��,�^m	�}i���L�_M��w�dŖ��3�_Q�Z?_-ܯ-��%�U.�K���؜8l+�NW��4ѣ�4��˩ˬ��B�H����ڞ�x:$2�Ka��6v1��42�n���Sv�=�o�7�u;�~I�SP�����#\AӒ��b�"�DDŁ�'�����EL�qI�_8)��~6?��G�y!̛�>��,��P���|���ĝ�a���|s���z�s��N���9>�}d�I�x8�[)'o$J:?��&h���{D�����S�w��\��9uyF�Ҭ�>����CX�,�p�4%�,�����xdO徿� �n�� ��� Wl�O��Ml� ���=f)(��h婹��)��Őt��!�������)��3[5�$�scR�A?>�3��lo�<�Gs%��C��k �a�8E�w<�Wu�~|gp�>���~���b�
������K�h�B��
��33�EWX���qg �X*I�X֯�(���#��T�T�KneKͼ�1�&�d�������e�2�̣#����oErԐG�
Vm<�6
4�oW")��h>O �ֽД��n�m���m�1jk������H�0���ABg�Q9�a�)`�@��w6.�2�ɒ�΍H�}&byϣx&�x�q�!��/p�}o��3�r.��%�wr��a�7m
�PSg+��[��Rvd�2��-v�]�Ҧ���w>>׌A��bu�/eT�~��KQE�Y�v`v�Q���|^�m8��f�s{|�����p&���Z�7WC��6�F�R9��e�mM)�(д	�د_~�j���o������R%������9�(%6�Ě�A����6>������HH����ޡF8h	�j>��R~'���nk�u*�m.�~ͭ%�2:� ����v��`��P.O&��WЬ�-�,F+���E Z�����W�EZ=�+!S�E��_��YϩU�Cu=��"�9��f�cO��:�Eٕ��(-b�� %������~ pv\�Z�S �N���(��3�_-�Cp��zɧ�ň��+�>qH��E�=�o�Q��?wO���T,V&Sj�J��Ra� �p�I!f+�-���NC'���)��
��RyȠ`��<�o�9��y.�#��ud��+��g��V�〤����0�ׯ@�����F}\>��yo> ��������Ly�F�Â��w���_m{8���ɜc�e<��kzìx�?k!#��b5�q\�T)2ԙ�h�����7Rv�²�~Y��}�gO>|�L_ľ�_n����>�)�T�Q/�>2J�j4������6S��L�-Թ��"������Gx�$������L�,�xo�S��@�#�w8�8�N�����ƴQ�ʛFߙ_� .< M|�N�����}��/Ǯ�r6Ю���u��*���évA.�s�W�ɵP�L�3������ۊ�,�s��~�#q�DK>��z�ʝ/�M�.@$v��M�B�8-�Sţ�#��a���o�6ο�Φ��b���$)�����P���2�`�b"l��½{���Z�C;��8aޓ���±P�˒�QW��c���^u��e�͌�\r����������f�^��4}j�S���S��6��4��w�<E�,�|s�eL;$f��!����6�*6�1�sc��	�SvĮ�k6��޿/0ƅ$���X
�5������ �f� V�H�g$CJ��� ��a	�븐���Q�'�f}ݹz`�xO�aR���7$`�3��������'2�����/y���m�O�S�%��4�%���A6�ѯ}�c��%g���� `��Tў��5��p9����J�ZiT3@���h�������l�Y�}lz�� s��^�`uj&Nr/9�1,�p��!�n�?�D`I/2$���j{�P����z�����������m��� ��*��5H����WH~ݡR6��n� l"D>?(�mg7y9��9\sT�(����+�S���V�í��ڮ�K��o!�n�"8���R�`�h�[S:b�
� ڗ��7�)��}����6M8��+>�S������p-���--н�A<����@y��;9 ]=���
Ey��O�7c3Z�ܷ�i�I��N(���6�n��*@E9B���Y�L������+l�����~e�'CU�.�`~~���`|2޳�Z��.��<c��a3I���Qm&/��Q��I����O�biG/�����4�8��+�?3q�
�2���Shnj˘��.'Œ�Ko����Jg/?�iKcˁ���.��XŇ�sإ�c�t�0�F�2T� �Џ�F��-�@P<�YBf/���Y'�抵:b�z�E�!�a��I���H��yYbzN�İ�Y����ט>I��ᚽ���Ȉ@~�J�mGv�3���I�iD84�;y�6ywG���%�R��Ii��y�
e��y�3�z��v�!
���D��	�ܮ�8;��2S�[��T0���m��<��^�U	5{)���Eͩ�������N1�]1��XN�F9���h�&4 6ι�on-��+����>���?�LfF`.��Y�f~97��l![�٨gf���@�(�}�8c�`�s��x�`�C��[ 
�"JY]�Y��%W�QMZ�{���$�U��cc�	���v��ǯ������]��mR�w��;�Q�"�@��5�>���g׳��d��c��H��<��1��J7���{��Q0�H��	���K^p3� ��N〉{Ӥ�ZhZ%�R@Q���L����	߀X�<���a�$�¡ɳv�Z������Eck��/�~J����o|�QU�U=���p3�~ӒD���e��@��SGWځ�����V3|/X�?t�Q���y%W	�a�������X�S�4q��3A���Q$C�ޅ{?ڢ��*�Be��BM����f�H�\3q�~w������e0Pч���pVƉ>�Yn�	�"�b�K�$c0SEo^.���P�.���j���ق8W����?[�o�����-<�m#��zq �=���b{��^�fqL ��~�"�?����Ѓ�d"���~����x3��4��X�����҇����
.��y-%��\h�Xw�.@�y��5:ѧ�N�K�{�nh��6 {����F�V&�C��#'}�֪�e�7Ă��g�����)�v�rB�w_*+�L1T��"  �e��N!v_4!ڊy������`�G��K���˃��=\x���Z���p��2����i����t#�iﾷ�l��D�R=fK@�CF��_�s�`1U �)������Z���ѥ|���:6��z��ub���s��~�5f����H�� ��⸛f[�7O�֓�֝��wu�%�Zh��"#� i��F;*��wq+�$�;���8IOGۋ��J��B/2S�s�y���nM�fqՏ�2T�n��"�@���-�ޜ�3r�����s��[��)��K�3n�.���lDEy���Xȫ���|r6� ,�F���(�;~��rR ��5�"�h��=�'?��E��Ti��d���|?������t�ȃ�d]��QA�Aÿ��z[��\�?��+��G,H���K#���I��Oe����^K�P�c,�u��=�O�v74\S�kx�Y�\౰	5��6�U�F�?�Y�������P�m2t�G�d�?���}tL�)�m�4L+� (�@�|L��x�8��}F	����.��� ��MM�[�}=zQ�o�l�����R�v��%JF�ׅ���|�)���d�<>��'���d}�^K�A�����q{!A��q�>L��sL*)Y� y#�̀��q[G�����s���d fU[�+~��DcM|v���ke�w~�q��Бф�/�ZJ՛<�IJU�>
1|U�\Ən}Wn䜰���ΠB�D:���Y�x03��d���j�	����Ƶ6��w��͟)ɏ��O�CNP.�7�V{,���Af9N�dp 	��ô��N?DRd�at���Y�g6,�b�������t��\A+�c���53��C,��#����)G>"�B�|5[�ҨY�("{��e�&��Y�Ā��1���8tJ��h~�_���C�d�`@�`�gm��\��I���z uȤ@�b�+(��؈�G���:��|���6��m��l%�|T���A�F1��5���
�z7����z|�ծ��m���Z7����1������S����b�J�(1�ǿ|i)OJq��,�@h��;u�p�<O�h�y9,�;,[qِ	!r&���/�k��q����p�f��� �iX�8���|��Ïѹ�8"{_����-S<d�@�9�u詿:��E|(Y�u��K��c=��[����yۯ%Ù5�҈\-4 �Kj���lv{|�
�T����յf�)8�2d���&�c�!�D�~V �6�u֖�������X���T�^i����8=�5X?L�%�W���j�Ϊd��Y���&���cLh/��n�B�z)�D��kﮭ�W�w��Y��0f|y/�1X��v,CM���=e��=�/*O��<� T�H�#�Q�R���C`V#�ۮ���fܵغz�i�W�m�[n�P8д�!�(�!�LM�����F�RT���(��ϓ#����wYC�*�4�f��� ��Ԫ`�}}*��S��?� �EO���f�}¥[cu�?4�+���嘈8aN>>�:ǯ����j��^[��
����� ,O���QB��]��Q��&:�o�e^�t�_/)�tRM��m�7ũ��$��|.�H\{�O��,������ɿ�Z������a҇�z�j�0T�܂V��Ҳ��(�,Е�/$c�;�Aa�철�Z���f��n���c��E������n�1o[㻩X��m< ��^��C����>#�m�p<���D�<�̍I9[֌_������*�T�l@����MӒI��w��X��4�6�V��[��m��@��;a���<"Aa��,�y�H5��2-�eW;xj���M:�ф�s��J��$"�5�&���<��4��L�1�8	�_�M��с�n�^��h� �}�jkΎ�i��Y��ƨ/�A/����0��ђyeU��e�v��&wv���l�|�q����[�iUUSrS�E؈/����i"\��7t�����"V�0+��V6.5s�1b��l�FM���@�w�6j�� dwl�2��T�䄛	m�5��Y0��^�Y��{�5��C��U�Ak�֪�V��0�4ǫ�r�C�؎���CIEW��Pe��l=�j�Rw��A�Ʉ��X0Ͼ�ΔA�����Z��'(��J
�å�8�@}hGL��6W��X�~[	��8�4'����CB�_���S�'!�X����k���͔�C��2�K��	�h%�Wj>��r�ɒ�s��e����#)��.��jq*��w�Xv��j�yG&|x���O�)_���HhJ��o%y��iaVd���^�$|�
j�q�w�N^�穪�����r��FN1��!Kې/w�6��J��Q�ﾺ�ii�b��F)a����Т;�d_�;�]�b���H�
v~*��b{Ɓ=+�׳�7!Ý��)���$�[Au��-0V�	�l����V�$�u�6A1&x�E�i/_1F�NN�SKD�͙s��þh��G��I���8���cw��s��X��k������7�,m{�ڡ	#i�>������#Dg��46�&k�����h~�����5Ui�Hc
�w�po�e'ּ;3�芓լ���tצ���4��s�.s"����Hk���U��������0c�|s��( �hU2��9`�F�ԄN]��ݪsz�R�#��۩E��`�����
LR%�&��cO�iݔy=�6X7�>�3�l �1-�2v�z���B,�[��[������0�]��(Mm@���=�o9��&��!�����+%����T��ղ4��yE8�߄�ٮ�"Yq�g3!�z��%C�5�4�=d�<��!��9��r�`�Wr{�'������-=K\����1���$��o�������G�=��́��%e�r��/�߈�s@k��{�VH��nXǶ{?�h�X)���������edL�=W��:��4f��~�X�n36,MW��*���9i�wd�p����иM���>K��Dn*�n�HF��nz��d�7[����Ae�.���0`k�UD�>A>&�	g�\"y\�%uvV��q������9�lph�*>��;X�A"�c"p^7tg���<p�}�	����J͉@��\c[�:�O!偯0L3d��p-Pɾ�D���"!A�K!RMy;7d�|Z,~]��`֤san�!�}������4��>�	�����������|�z0fX���ѦH�-�ǁ��:� )���q�Q���9�3�*6c�N�ק��u���<z�|l���ݿw�9�V	m��m;�Xo���m�.���ܙ���Jg���P�+�����zF����س� �jt0-�%3��3q�^ک�vCϦ��$o� O��M٠G�1�NmF�mP���Q�d��ky�DaZ[o'S:�6��(h*w���h�*�����e��Y���1De.;X�!/�6RO�h�˵�.C8x%bқAO�ci[}��m{��]v�B�j�T��.��ӆ=�K�*Vk�������A�9��x/.'Dc��l���[�f�<�ΰ�z���>6���ۚ�I�d~W��o��^®�Jg�օ-�<��aK���Q�02:CZ]� �0Ğr6��xc�)8T���N�1�!7i�0T���U��a��=T���1���NCѐDa� 514���O�~;>
�H���>J�� ���|������
���G'��4���IW�~�$��z��\��ކ��J�� U�3�/E�Ħ���77*���$ٖkX2v�O��~X�Hil��<�w��YP!�4Z蘙���NR�n^y%����Q^)�3���=�|<Lj��kh*�����*���J�r�q�3�X*��˯FA2b%7�K����x��t�D0^�� �$��������<�٢z�`πw��I@�0��i6���>վ�LL����+\,��h�##3ĞY��dL� ��-���yR~�Fx/ME�A�˷É�S�3!|�����`W��u%u7����	�$�~���w�p�ܒ��H�r�X�C\�Ah�%�k�,��j�'m��%*�J}��>��Qt�m.o����4�����jt[�K6���(���JƝl= �g��f��T�g�d��k��}�a�^=1���Wd�����9�ƅ�2_Bg��:_#c�ٮ����Iނ�1�%f]�+T�)��A���4�o�_��?[���L��5D�Cf�ϙ�e��O�L�6����?����G�(p��D^��UD���5~���Q��*�\��U{�R�P@"pf������xn#|�W�v�M|p���]�O���]���P��*�<���w�;pnb���K��w[3��,��YW31mg?g���X�����bo�L���gʧ�.x��.���^�fe���Ұ�4�?�fwS�D�Y6�.w �#m"�%l3�n���u�.n9���c��?&%�!����l��

U� �W�8��~M7�*~ge�a7��-�^�&�젨˾K8���baͼ���� JTLs8�]�_*H]�R]!c&�5)�'�;�M�F̣P0�#�-C���;��V����Ͻ"y�Y%��<��8q\�˛Y!!��m%���H�A�eE��G��r����o�Kꜙ��Zk˰N��X5�L��|����cY�ţ�ؒ�a��T3<̜�������`�x�Ѣl�����t�s�E.rA+���� ��`ٛ��H��#g�2L�rJ�.�G�?��ѐ@�������P]j�y�E{�/�ư�mf��F%�R|��D�gw?8�hY��%#����F1S4��F�T�����	v�A��	@u
�>`�1�|�����b�/�Z���:����l7wD�	<y�ؔ��O2Fu.�-��qZ&�Dƾ�a�ҽ���-����C˻����K ����,�t�Ȩ�H�Ùw��,���H�s��'3lBMd8��t)|�P=�cwr��&�QW@3�w��~zf\���_"q`���Fu��U��9M��Hl�C�l���I$nTTr�<X���K���U��{P��"�w�V���%���JA�����4�(D_ϑ�ЛM ��J���L�������u�j�U�d�ek��'�aP����,�T�Nd`���r[N�5�z8�E&[Ծ�d^g4�$ݞ��Ͱ��n��c�X�a�2�����TSL��$�T�Q�d�p��K�2���tl�� P���Ic�φ��)[,��$2gr}�Q��w��oj�����jn�i<��rVS����)�s������=�ʫ��A+/����U�����l�>���W���<��Mj��ى�3dX[ةV˟��Pe#Gf6Z�e)+�b1����o�T��q1<D\�:��'>��@��tt(�dy����J�^����T�7o^h��T�r7au��'�C�$�?(�dCI���O�F#���	��td��.�����׷L&К��D�E:�|RP+b8�v�@O��Q�]�
�#Y�2�-c�Oe��B�u��hùz����@�15�G���e�u;�E� |ƌ��PH�L��/�b]yk�M������]XB��;
G43a�g�1
�X#r81J�3��$L�ԭ�����<��u͒��~=�׏�􅬛*��4�x��C?������������@�睉}:���^oz��Oըl������<�P}�*c;R���:�9�:�]h��Q	W�H͝g�D��`V[�� kB�Q�	�S����@�Ψ���y����a�	��`ZfU�ڮ���- ~V��t�:�FSjH�ڋD95���}O`DyR���>vB�Ef�-䬲
�l����.�2a!���'�{?�)�WW]ڌ�o��b	)�vp2r.'�4)��3��l`���v�r��f5��z���������yKʑ�''m.�� ����愱���}x˼ߞ�V�H�~���� �cGW�m�
��RW�pn��<d��S���Ј}�����j��oH�������,*m�b
׿�2KWG�8+�y��`��sdM�#1��r�F��D����JN�_�ē�k�<_�@Pg_��X�G�i���0n��N��¢��"+�7�E��@���sxs]U�׋I�~6s�Q��
�`}>�m�cx�b+c ��oݱ#�JE�N���h[O�$	�N��u��B�Xa�p��{W�3�7v��O�O��0H��U3ā�4m�:�@���4(��z�������`����ӣ��hߝ;p
�������bg�f�?F��Pf�d��PJz�ME�T����J	F&�Tf�C"�6uL�I��.��0zC�,?��d'� ����
�X��l�?vCs��d�������Q�H�9�l9B��I�ފS�AT �v�E
6S��&8a(�����s\���L"Bڦ�����-"!k<�2��{q�p��8��s�>mg� �3r�ގ�k�� ��}S`<��rD���^%�c�I3�� �L��ј7��h�ˮ��s�m�B�:l��*7>�A��ĺ�X;�������`޹t��:�0>�vkN�ZR�v59;�云��B�J�)���;� <�!}����d���y�_��QG�e%�����O�>5{����yI�_��E�q����6v{>���\�_R�O�H��v)֧k����U�����$���~ �
�'�i|Lm_E<t?��P���?7x�EkJ@�Ғ9��Gm@�E�T;a?���	�nr�z�������u*���H�c�3�&EX�Ld L�i�bMfʬ�螯l%k���ⱅ�� eTpW�.�����kE�4��K��Z��A�<!�xR	A�a��P�C���2Y�z���)��r�[�u���4/١���)���4����I��J��$Դ�<��dlo�\�+-p���0��4z���Ů72���`���k������*�D�<�B��L�\�<���ݓv%t�jV7������Ȥ?��G[��� �����z��F ���;/���(}��ݝ�;�f��*��ɗn4̃==��ǘ�����yͧm��
��䞫�YB-�	�L��������tƿN8q����ej&=�A���� ڙ}"v��%��*�\�o�+bȄt��hJ&�H�Ӥ>�=�=r=OG؀��2��yS�O�̸R./�#p;�� ?���wB=�1{��Jb��{2.��'�S��%3�s�g.J�+�xBCz���u�e�8e_���W��`�,?I��]J7.2{3��������$`8����C�n��M<d� ��q*Ml~���WK�r���skA���.�����4��MZ��|�bјl���}�v8��(��D��2�ˏ�-�y�d�˶H�ϴrtZ�6i h�Y�8e(I,�>��d�a�R���1�"�X|�۾5�[�4��Eu�l��Y���"���K�9\32��~�KdGD\t�6��p9Jl����F�Ҧ�
O$S�O�
n����NWf�Ĕą����4k��h_zie�ɻ��ݨ�5�{Rm3�d�/P'íT�>PK�9��
{��%�&���H��M�����{�5�?�q^�(�ת���,HPotɈ�E9ԁ�x���͑��~v�D��!��(�`lo*'"� sL��$�vFj�V4�8�uT ǳni��_&f�L��o��DB9ҍpkI�� �	�N��M����{�_�y���x����#C6v�-&s�ܐ���w4O�������wG�Q�)�8iNo�'�9%9s����D�����w*��iI�	�SY)� ;Bz�L�j�qu�!*�ޥ'bJ��9&I�H0lR���M��%[t"#p&�[Q��vԅ]U�m⿪�Qf� ߘ�Z��5���5��/�Ѫ����ι��w����4� и�Ԟ�B����a��RK����(�9і)�d�@����:�It�甀*����GH.�F�B� ��췧���j��hɜ �+q�?�,6+B�Ve�e�<�F��o��[�f�1s�
u�4K�6���s=���d��;7?�p��S�9~:����l��Hat�\�x/�9���O���3:8W	�� �����"����j��7����Ӫ0�AEPk���q���h�RC�����������2�w�7��9�����erB�!Lx@ujN&'H�5��F�+�*\6B�y��.i[?�^k�^�P�{.�f-���"�,�#â�X�%�'���6�����snV�њ��s&�ۉR���aI7��oM��wĤ,!�~�}�9�|�>������]�]ӷt�j��fĀ���WA�#�2��a���ʋ��m�1y+�x�,D�_��r"o(=��;�$90����ctD��R^��ء�K�,0H�)�9�:5��P0CNp�l����<Hv�Ӈn t��X��un*��p!`?��W�n����c#+Y�\���f́�`��g�7"����? �Vk�	�x	B��f�/�_�+�V2�$�����4�)�b~������l���?#>�ǈr�~'}�\E^����Rl�<=^_ �Xz2�CP}43Дt��cd�#�����Ł�p�q8�0��s]��ε!U`S߈��_BI�4��`��V�4�BZ�G	�۲���(���˭W��1����Ola7�X��ݘ�p�	�����R鵛/ ��"��X�@כ����8��`���zT)f)(�>���S��c��e�#���J2�d��@5D9`}H%��3��͑��~mD}0#�{�3�J.@P��s�.QCX���ńK(=�����!��-T���4}ӯ���/������,(���pP)�s�w�I��_B5�{��QѹN#�Yg#	0��j�@K�J.�>�[�*"�*+�
pOö�4�s~��U��! <ɱ�l����g�⋌�F��u��f,Û�*;�]Si���r�B�倵t�AZ��G[<�8b�~�O��C�Qp|8(N��&�¯̹�}3��[TC��F}��t?���ݓpEQ*T���������Њ=��T_[#�%򣱮Jv�Ns7F"W<ËFJ`�CDq�tl���}W|(1�88JY?���^U}k��y����(Ͳ��6�e�"��㘐ڐ�F�Z��!ӈ.I\�9ڛe椬:�ߨ�D�7�
��\`�C� �/_F$Uo�0}�Ւ�e���T�8>�I��M�±�Av�:�c>��G������<��mK*7~~�O�P!Γr�~���I�X)�)@Uh�%�>%�_�T�F�y��N��H�ol�^>J�1��Г�_�[�;����%xbr�����Ġ(����M��G�d��U�ĩ��![�^F�E�P���f�6��C>�幃�+��q�Y��?f���5{j7v�ɂ�C���*�&��L1�c���	�����)'{�S����������Z2DUV�8�����,�w�Z����A�� �l笩�����_x̝�c3�
띃ޜx{j�c�<��Uf��qKm�Y2���BW���/E~�|�R
cI�F�̻4%�����\�i`��L �fF����j8�e���bo9�KY�I�Bp(���edI� ����yCYZU�O<ߡ.��'���W��y�p��M�Z\��5�����=��G��6���0BAs��5�_v.V��e%�����T����=�����4B�^I�g��y	��U��.�����y�8(��V�{��g6�t4�C�a&~�J�鮧-�Ǆ��.;]1`%��㮤�X1�����V�?]������A,�P�ᶿ��&gV`�u]|�J	9�vC��A!Μqs��2���)��8�\�:�PR�ai�͖�
h����*�����GL�:��¥&_�!NUB�x�,+�a��z޵��k|�1e�bR�Q���� u��N`�_A�< Bi�H��K�)��g�MK6R�y�L���^%v���PO+�w�a �F{:L�j�!8�F>L��s����$&�Ζ�;��(|z��
)7Z4h��0Gy�ݨ�t��Y�ʨ�: ���^1zHwr�$	���X��ǈO�4���M�`9+��1E�b��ߧ�u���aJO���Jj�F�0���"���r2Z:p���ޥ��yX�S��	;�9V2����Q����8���҇cʶ�Q@��t��w�p�i�]���u��_Y�z!�����1`���ߜ�w,�Tq�򕅒�P����G.���L���]��~0w_W�=��$��'��H�|1�ϻ��� /\�;j�1A�����vD%ϒ��F��`0������'^0Ѵ_�2���i>�s���5K}So�$n����W��_�-`�w:��X�z4sZ1L,a_��&-�A�{q���|
U��(b x;S�)����y��

�_�]�˰�h)�(��u6��9�翎|���V��%�E��&������l?<��u�C�<=Lb}w�J��b���٠��L"O?���-�6I���Q��	'�@À�_ى9�b���e�jᎩ����3�=�K����h~�:�ɏ~ޞ,��!�-��n#!�����tk��+�����2���KԀ����[gz{��/O����Ğ����A��$�Xº��БK2Y�z���=��4�l�����Q-�a�S%Y^�U�ܚ'��I�1�c��1)._@�E��_d�Yw2��l�`O��$������R�l��Iy���*gk�1|��n��E�$9l�0�шω���)�CfAֻ���`�P�C\����G��[%�d��ɼ�#ϑ�p��m���E¾)d��h��S�Y��Q�� V�̬g���ՇIf~e���o ���� wu��;������8긾��N0*�C؝淵�l�utx(\!m=~ٶ������ւ�91���]hA�{:��Ϲ)�&�N
ގ���կZjt�#����E����`!�o�l�頚<� +$0')�g��� ��5D�E�+=�������U���W�]��-tC��RǺA�;X7g�z��}��h+}�0�越�a��@�Y��!%}M�[ie����^�4��!�Y2Pd$DEIA�����;���'Y:�d�e����f7�%�aF��H��!�R�}*�}z��5�W+�r����ބ��<��ǭQ:�l���*O,����D�ќB!s�H��P6Q�=sRL��tǐ&
O��˟O�C�T�ů͜W���~ֶ������Y_ќ��W��O][�*<F�VߏQ����d�+���_�� ���R�hv�/}:��"i/ ��T���$y�3�:	�|/(&�u��X�A�hm�Y �R���� ����0G4�OH��Hw�Z ��D��xj"�/4��G<����]��=��T �y��q7�S���YTT�8�択B�Ty��">��� ���;��������v��^�y���]jX#(f��C�>���߻�+��ph����f��$Յ��v98�y@J\�Q��)*'��g���n][��ϰ���YzL�\��$"Xܣ�b�W�G��(�\-�|�MA=�-�Vt��w�.X)®�o(�ҭZM��o$��"ؼc�Z �����:�{��(I�R�-�w�8^׷A@�>��/����fW��&�Uocۚ��e&"�`�U�=��WMݜ@�A�����JAQ��#��V��-<f~S�4�_��v�P�rJt��F�XǢ����wC_߹&6��S.N�w�u�Yh$K���2P^rG�]��1[�������*f\�D:�ư�s�aD�/񜢯u~�(�����,L���.�凞B�����g_��Rjgu�hElѿquڨ�Ds7l~Yu�S�l>��L��X�����v�ԂI��Ѷs�F��L��i[�=����kc-����f��A9<�	�ݳ牛9���
'��QY��O�O�у�\ܾnÍ�N��� �48�9��M����C����Ğ*� S�?��j,�o�����t�x����滵��UjB(�?��3�*^�deG9Ľ��.m�3���C���fo'0:��<��Luh�o�OI�S�nǃ�i���'�����ǥ���ɝ�ᇝ���/0gc�k����M֩��D���������=�����ˣP�x���8������0�o�v��v�F����`�"�t+h�}�pT�4F&n��d�P��;�����e�D�Vz�ـF�l�a�/�D����
o͑6����vqjL���B�KX	V	Ւs5O8��37~O��� �c}�8��ڼ�P*ncT�+��AVx���Oa���ȃ��w]�V�y��s����W����<ڵ�/��o�׭H�Ť�#0��� $�(8����h��b�?(B�!�19�4mw1�x�S� Kz���9 /⑗:RpH\�B&<���5k���j��,g�z�}��a�v�)�*�f�PW^lbN�b�D��'�ŉ�X��9�;,7
^`����%�T�6�{�h*D~�DRtu���|�J6;j��#�O��]��"�x=���o�|�b��V	v��k�iRC��h�]��rQ�>�Ө�!��h�cՀ�b��v��k=��Z����l3At_A�����a�8M���04l�A����
�a����j"�lgN�
�|�w��<��S�q�Rr-�骵�Kܱ��A&D��"�le��C¥m.�[�2�+�oce���ĕs6}�Qrhچ�.5�`	^��d�i��G3o6o
� B�#A+�j��S��c�&����q�O���	YB�r�N�r$	������_�=�����K�ʃ��� �!�̌��Ⱥɱ���7���%6��3 �2�任�k�i��D  Gײ`���Zڂ�r���L��H3�ta �k2��x��1�&.g�����V�R�T��,.+�q�}�W4d-�u\Fg�sdg��X!��W��B].}�J��:.R���q&:~B%�B�<��9q��o��"{�w�A:2v�N�MN��m|L�����ct��) �������Uko&1K� e�o���b�G��al�J��(��!�c�h�HN�K�2�Mۿ��y����� �����Q�V���&ȡ^�٠*\_^�#C�Qv� G�d�>;k�9�v�#^XnB������͉3���s/�[�P�����8�ɡاS�U �e��42���L�����[��*��ue8���4G̾~��[�7���L�0���SG�Κ�b��|�iv{�2���:��,�U2�X`�ݛ	d$�Cw��~�ꞟ&=��B���;�i�NF�ǳI>�-z�N������˛ 9�,��Z- +��ֲC�O�#��������xl5n+bI�V8�-��;�\�O@1�D�;vS��HN~�"1�#8{�15�����!��(����l��=>�o2
l��p(�|u�1�l���X�UxO��o{Ğ����I��G� �+y�a�2Yp���eq
JQ�!�ko��@䎼5#�v6j��a�7P���@�9��DVË�z�9|ތ�v躏����*�0���o�1�WD�E�5	o��7?Ρ��� 5#8	���%N�ͣ�SWu������b콧��\~tU[�ÔO��2��yc8�c�#�o�O�,u�e���"ßF��>�{O8��BUo!�!�Hx�!�*�C��f<L׮�y�h����G�K���=`_�u�� ��o7�զ�����k���8�*��>�"��5Һ�������0n'=l�Ua�㼫�6�]a"�6ʲfn���9�ր(3U=��`�"���NP�j��iH����H�j;�64r�t�Skj����L�4\s7ڣ�Ay|�+ ����P3Ȩi'n�4 %K|�)����Q�ÌY�s)��^蠵�z^."��"WK.�w�x컙���Z��� ����Y۱/���'|�B,�x@�����EN>�B)xRSM�E>�*������뻪\�D���4?���I��B^ݺ�Q� ]).y�b Y\���g\�C��x|�2[?l-�8�v�Fß���X�l>?z��]���Ҷ#��3QS�2D�*�9:̞�/l�=�o��W�K�>�	��P��� N�D�3%�^�=�\4%�籪�D�PLJl��h��m�aZ����zW����ӓ0���AТ{����|��ۭMӇFBCB$�ȢP�bV�8�1&�c̈́��n�7�]�LW�$�}�b��xo#Ǯ��+[�yH�l����{����q���>��l]��\�q�����e��R���A;�"��Ӕ��1H��4a�6_�w��}t\�^&L���0���07@���ǤC�"k���4w)�����R�zd�3;��#��! :�*i:h���r>�WBq���S�X�f)�����u��~����� M�����>$�}�ߦT���	X{v��pG�?`���f�~��H���Ew�n�L�u�M�!�p*T��_I�d@�on��8����^t�R�L�E�������`���ˢ?��/J"��H�n,l*Na�����J��j_��5�]YW���O;����L�پ�����^b���+�ӻF\�� ÁW���N���\E,�^a���C>$�&/u�f6�Κxb�H�V��x���G����G�hz�VNT��O��a^Z��h
���S�q�:�@x�S�[�SH��.�}��`���z�oz��Mʢl�ADAC`�*�,Mٛܦ?�Yx���D�qpY=�3�Pq�p�J��ǔ`|�~,�3f:%��=B5�8�Ȭ���+gf�p'`[o���G�6�ޱ��h!5�p
�Gh��8	T�A��>�t��^ɺW�!;&+mL��aW�\M��暌�7Ը��%N;N�oⲺ��/B���\hs˦Y,8�����S3$��8�އb���5���6�0	���q��X�M���p���C>@��0�;���n�e]6�����4����e�P�oG��˳�	0lTInT��H�p����q���Jq�ɼ^�����5�LͶ��ƈKy��^�f�jE��˫±���/o%V�`�.�}�!x����?Ӣ}� K=�h�5	��Z�+\; 	n�W#�����m����h�����\�$�d����$O��6��X�ڼmX�|��(�ܢ�Qш�@ς cɔM9w:���KS�8��i�k�@#y!R/���8rj	��0`,چ�J���{b =����|[Ea�k���Z�>�2�m>���-{ƶm��Ri9 ���4��,�E]y��9����eB�����fL�1#Կ���7@�]�쎿^��J��AHQ�N +��f�1`M���v�x#w;�I{+A�,H������R���f�"m��S��}���G�R/��T�g�1�N��]�d�ȸw�,}Il��V�I�S���������#��B���o6m5|�6���T�%m�}`��uX��
�� ZA�1�&r�X4y�G��?�P�Ml�����=��_v��)!_�u���	��" mnh��Q��(^k'a+[@df쐄������~�|Ә�_��MF��4N!�s���`ÿ�
��ϯz�~���*@Y����}���E�rM^��NZ��CN�'�U2��_�SN*܃T=n�gq��#焊~����~�]@�/aqD�gB�&(a��+ƒ�ĜA����Q�Ϊ2�~�.������������Q�(�_nodlY���O_`UT��o��s>r��/��w�)�^p���k�
 e�r��H��0����
�V뻞@��f�#F)�e��s���D؝�K>[nyi��զ��`��������3��J�m9�nƣ����͹�1��ư4�4u��Rw�����+ׅ��\oQ�1���<f���@�&��b|��u^Χm��p���ϫ��-���L�U�W[f��nD�����ߏ����P�Nx�����O&�z�l�t���׃m�_}E`�r~<y���4���Z�����3��ʰ�%�����h\t��d���.��L&�M���/5�b���Qa��X�DTݾ*�mbN	��O��vCI	�TW��m�X%��{��!�S�O}݉�\5���Ϊ��l��F��`T��=F6��c��ziyy�?��T\�8�,�[G��Թ�áK�ӭrd������
�)���<��ؔ0}���p�K�r�zΟ�]W��{]� � ��i"	��$��&��[�L`6��:;tTŲ>�<w"A�uk>݉5u��^�����#��?#$������qE$aZ�'��VՑ7xU�Y�B�}f�?��e�<sa�ʆ��}�Q?�MB�ˢ_k[����A��s���И�i�g7V���V7����ҿV�t�U��7.Ǎ:1"t`1��|AxO s�។L�v�gc�oK�����=����k���j��!�<_W���>®6d&� �6z�	R5��[��0�/�{��uM����϶S:N"+OZ�~�,��[}���H
�$��Q�vJq}Դ"M����}MQ�# �� �U���02 �O�{��� �b;��L�!2��3>}y��tj���$��M'#�<�k�E�в������0�Cq�Ԅω�͖V��|q�ThV+G$����\Żhz�ʫ{I&�IŬa��O3GO#V׵�x`���u��'��*E).��)�og��Gf�0!<æ�����#�o�2n��y>&J&�H�{��	-�\4�, ���
�W;��2�'��{ W�W~8ޤ>$f��x�n+R��L����m�8�����fF5���*�`^b�5��ōǆ|r�O��\�$o��q����t�]$�v͠P�,t{eC����ͧ�G[��i��D��6��}[绬��8����Ѱ�� j��a�lP��zU�D�l�X���l��5D^�n" +���7�j?D>��=�?ӗ,�P���{A��P����KF]�D�Z��?�����W����E�G�8�ػ�˧��Lw�J5c��[%Ćz��ʐ����|t�5�ϫ8�J��z��l��,i�~�65�R9� �m���^��<kJ��(qځ�辠[�8��N�W�d+L[U��Y�Y�oظ}$�?��~x`�}�a�/~�.i��H��d]�R����������×�Na��&�0k����GH�\�?�s�{�/T��S}��g���_6*Wc�N�D���"�K)p��nu�Q���P�|�x{������@e�{8%-�'���;�_d�p�)�u��1AM�FD܀�vq%2�Z�\c�r�!f�k��v�#���RT+��W)���D��?���>�-�݇h����@���f��|�Z�_��o�F�~O'Ԛ�4��k.���������q'J���Y�+�4-q޹,؜+rY�)E�d��I�s�X�χY���Zs��E�8�h�,zy�,�v�����(��`�*](4#_!6u�����*`��QTTm�cH �'���J�>\v&��w\��E���dS��Q*=֗��B�W7l��b`�H�8��3rA������G��E0�S*���p���@@&&��h�[���{k�V����� ��8�=�ޓk�!:��is�:
i����I��/z7�W
)l�T41��6i0���q��QJM��� ���[�ZsˍO�p��O'��vX��M'6�Y�^x#Є�8��C�\W���A���(:�T�$���������Q�m���k�8��=b�C��Ⱥ�A�>8CA�,��6���D2��Y���dæ|�z{J��S��i*G���V���1#m���U�UϞ�5�M�@��}�H�	��OH�;r�N���>N�tϪLM�%�X�w[!�NU�, j3���]�DW~�	���}�n� �+�%�OV��u����`�.8U@\���$$��	Ϯ}�	x��+�R{�H-�.�H���o�	�ʋ@V��(�{1T�f &[�@�--��B�]�.����|�����ņ�7ʜ�a�M%Og�LX��"IF>iP[��/ �T�f#}�b���nt�?�6A���$��Cw��6e{8;NQ߼^�G�Yr��`�i1��G.!FIWќ:����s� fqca4\���ʍ��r����S6�߿-��H�QRZ����9��2�T�8����/�b�[�v^��X�3BmYe%�G���H HI�#ߌ�tB��?������rm��R�#�ir� �4p�n�4)D6G�&s��٨�ҝx������$0�ǟ��[��G~�9�� UYrx�Q��=�ì����g�E �ЕYkm}C�^-����G�6 )>������k-x`�|��h��"��	ʧgH�t��]%"�j�lS&��#�A�<�L�	��k<V�W���,D�xm��`p q��=G�Y՛J�1��z�;�^S=�V��mD�{P@�7�� zc�� �-`3��z�I���oU�I�j<E�Ѩ�*"�Rj�>���\�Z<�2?C��V�0/vh]��(Ĩ�A�����w�S0�Ǜ܁�0CHM���]�~�'��~fi1+��o.��]����=��GG,��׮"M�Q=5s�>��ow�ى�Z��Ȋ�݃����P` ª�<��ݣ��]k�Z)�SZ�l7��
�GA�S��}���Lq�J��Č�xB�>�KCn4���&�Ȏ'I<m�o@��~��GI���s�pOۇ�w�<0"�ˆ���_9�59WŰy�w��B�`�(aWDE�����D骄ź�?������c�P�SvTgZk?9����䠓�nc7�g~>�v�'����Op,����E%^T|+�~J6�О�y�713��x��[M<l�_�"iO�@�u�9LЕ�����})lY=�j�J5]?#��_����c�i�/#Ҍ��*��������	~:�3K�V�z�x�ȴ�[i���:��r:�!�G��Sv�6�BNU(8A\Pl��[2Oĉ��d�j�BC��2q0�Wk턆��{�E,;]7/mՑꕼ�΋�q8���=�{R��}�Ґ�'�5@��y�����,I�m��(.���Ƹ��
ݐ}c�f#��Lr?�5P6�NT$3��x���X�ڗ���nH<lL\�#����(�s�#�Eӄ`"��ᯓ�o%�P�^��'���M��Z�.�,�"��B�8�VJq�a��A�� �� Y^���$��M���Mw,�:݈��:CͫL���~��y�㥬W����8]m��Ӱ�eKD��L�K�j�/FM|�vC'u(Vpe˾����T� ���S��G�B�T����eW�0��G1k�G���?�	OR�Ka	���5��$Y<�����i�7
���:�����4�fb|X�*�@�;k��
�W��������g:�E�h��3��
��B�H��C~�(��pPcDװ�]�%:�kK-���A/΀�?c�2䯮���F�����=k���*rU:�m5 8����R�{��h�r��p\<�E'����@��&�ה������00T����,��}�=�����G�},c�G���bCcW�H^j��J�}�Y-�~�Cd�1DZ��l��/���<�ɦeFԠF��3bv�s���8V��k�Wb�y�L]L[f�/K)��4.�^E���g� \δA���Q�w�ƫ=���rwE�U�cI�ܝ+ʿ[/Jj�~A�Y���`0��I�����f��<ո��)���� �gU�z�a��Q���|�b��(�5�/�W��S%D�65m��Y${���:8��yQ�2��N�,N�N]J̴��N.�Q*h[��z+\��m���u�o(�_���h����}��WY���CM���W2h����a�w*���kD^��#�!�zO޽UV�
#����_�q~�(��ײ�sm��g�8
$>�W��;F�\�Js���U"��?���ϟT�����u�y���2�h�#jg��L��Ke�� ��哌D(�kP��v�>���JD�~Q����D�+�y�����?�F$L,��\XtO��gD�$�z�Ǭ�NC��"���`N&�{�̄"��C;W�
=�������^��싂m�r�N
�p� �ƹ�L�V�,��+}'M�צ�¥:�3Sh�>°����E�K��-6}�mX��}����֠��;L7m��휬��;O��P �3�ǹb>w6��ttIJH���L~�
rt`�P�C����/go_8� �!/��)Ů�Λ���R�{�� ��$�^�H�[y�u�@v�d����i����g�v�td�<���1UD8mP�{P�c'��qVfJ�Y�z�����' ^�UB��} ��v;'��N_�8���v���#c�	�i�nɚy"��[��:c��ԅ�_�+�R�#9љ#Z�f*�;s���#6L.J2�	�绽�ׁ40�~�`�ǞڻҢ��6[s���0��I�$@ပ <�j;���Q���a��!;SK���d\e�=�e���L(R:��� �1���<m������ӗ ����c4uf�	���^�G���=�s��:� �����_W�w��������&�\����6U�5� �$��ur��_�9S��JT}��؊�4�y��9��^���{Jk�9/1R�XO[�/�`F�ۖ�;��o|���^�AD�hI���e��*�D�Iݲ���?�ԶJ�&�2HL ���������_.j�e��V@K��C��9vFm����0"IF� �0n
5��H�@婃�@t\O��MK�4gcG]@������1�(�/Xr�иM-�dX����A?��k:�cm�F%���=y�I��W�޽W������oޝ]Q�YRei\���a�U)Jإ)����I�I7_�_�R��z"���T�	a�in��\�1�CC�ˁ��Z'�
�Us�1��Q �/7���b�>b�k����KC�9�;���������i�ś��+�%n{!³�Ho�awn���$�E�/�]�����S�M1�CP��D�A&Ъ�Ȥ�:�!!ο�N����s��5ʯ���Ճ.P�m"=S6��yc��+���W�,2VU�﷓<�7�t��S����ϋ��3T@�{W�hE$�#�N�:��IA�����h���$1����m���d�]u6t�߱�P�*:��E� oý	k�E�=��B�Dds$iXW,|��`�'�Uz@��&ec6��Ô=%bU6'�)p��������r�3�Ԣ$[A^4�C��9qے�El�ݮ��	���Q$0(Q�b����r�.�QT;���8�����1�{Ҭ��v�(�X�2dq�T�G��J@���u:�P�_YTi)I�E���𷅠31z>�4�B��YP=?Bz�?d�;��pĲ�nA�9��K�&O�e�����'�r�K���=��\�������q��	���D���2�!8��8��U ��gr�A��#!�|�-F����g4  ͱ����`;��ϧq�	��A��U�:�g˕`�r�XV��!�']E^���ڃL>���$���V�&'�{Y��i�W-#��'� ^!]��\��!�A|�gܝ��8�1ݓ0�EQ/Xݵ��˜x �U��?��Z�/��N)D׹���դ��\t)B��0����we�1�WZ.��������� �����D�j�/i45,�� .�1~|k]ƨ�$&��"��cz�%t�7�P�@AZ�H�-"����R*~����X��A�������}��l͜*1�۫�� j��3��<��e�g}�Vԁ趕܊R/��m	��
u�H�8hk��j3��!6�C����dĖ\���&��2(uY��������A�(el�M��Y
3�<r��j������fb����cG��Y�b$��~F�'�]���F��iGs8.&T�tML~?f�%��t��v�������1Y�� ��L��?����8����MY�6�t���Y�@Ȼ����M۫�8b���Ą�R�m��Sg��Ě��������?+yQVh@x!u��c_�^�2��{ș^-���ߛu䖻Ÿ8@��$�uY�ѹ��v!5խBB�\��xQ��߱�&���_bd��@Id��k~���yO�A��;F�"��&%O!���\7�%$�&/(�i��T�{��֟Tt3�C���A�?���ux6���16/!�7�����f�k�f�q���J|�k˂"|��o.�z�fi��̯�g�W�]J�s9ݞ����?79�C�O�Уηm鷩g�Y��t��3G%8B��$V�\�F�5t��*!���.�mAt���P,<���.ɔ�OG?�S$_�)�c\�Xf�U����O��y�&���F���>�\&��������n�=t�20zi��L �D����
���|!@�~��A�@�*�qze���I�<1X ��K�ިc!t��;�+�\�@鋎��u��S�'�X�<vb3� x�����\�89��5����'R�4
�_�rGc����ܺ�e���vk�ͲՋz���Q߃���7L$Y����U"}���u*������}�N$���׮G�0Z�2���6ÉD�F.�Ԃ��=��;ؐ$�P2T�H��͌�t��Z ϴ��nG>�s49AN�.mt�Ř-�ڥ,�X�|[P.V��Z��A��c��KOR���F*W���p���Dw	�Y�[/D��2^�S�
��:��BQ/Q(�~l��Uv���H�-`��ϣ_z�`Ό��0|[=|ð �b�[uPi��߁�kg�w����пqo��&��f�rJ�h�(/����ab��rގ�,�N�q_�!��G�&x��yҖ_��/ëe���_�[e��68�a����o&�hD[�����C�,�^��t��)L�~�<�Q����<�%j�B��xtz��gY�x�+~~�OsV�J�rU��3ɴbr9��vz�#~��7P�0��R�Q�u��� �;��FU9ds�����s����;i���	M�m�5lϜA�|��!��J�C�����U�]n�6��_�=���3l9�m��;E����k��A�V
A�xN(�=�.bng�bA����:v�q'�w�pL��s��� ���v�~������A�j&ia�?�U�m&^��jG�$�p�Bh?z�x��f,�!�є1_C]/�o`V�Wv�I/o���S��=I� �a^=��5 u@s�1�~���9[/VK$����4��C��pW�g�2/���g8����O��9�p�\�yc��$��;��^$���щ����F�"��a��/a�Ʋ�� o���6U��[�2� �i*I��&2+!���#Rʴ��ɶ'O�Q	䘩�A��x�w�)|�ӯ.i5"\�ԈI���?��֟���f��KU��U�/3��W��ye�-f�ǱƷ]YI���O��I�_�B��N���C p��N��;����e�8��b��qٌ�$I[�b���ǫF�{JC1���S���8�h\�.#}�+���\��e Hhd�xkx��?���'ɓ_�ϲ��[e���j�������S��(S���X$5��y��!<N����2�.F4��$��Y�LbH�h��9>�-�(.�C=��!۽�F���T�W�j�~��M��&��Sz�`�S��M�~�=�������8�vn�w^~L�A:���gE����8���[�%�vj�P�����2\�=ŀ�m{���Ma�[�:v�}�=�[m��b0�d�u��G���ʲ/
���g%<�=�Do �ƨxe�$�n������~c�Ekj�y�xL�-`H%���0��֩�v��SN�����J
Ǡ��"cN��d^�/��>�Q�7�%�?�x��2�]����;�)�G�xQ�o����^��B
_#�`�5h[7d�<H}��0.A\��Ro�n�P)�2+�q����1��8�gz��Q�.^�n�:��}�lۮ2��	��l
���OK�^� @'$U	�EW`�㔹�ә^��\6�e9@T��F�3Z;IГ�)���(x��;���7i�AhIu�Y�(l����wFJ#�\�?��Oo�AdS�P�[yڭˍH=��;�$��a���p6 4���C�ҜQn|�2�1�ߑop�����K�,,�pI_��}w_���P�,Ƥ�W�}(;u7���1�ђ(�5'�vl�k�"}i��IȞ ��8�|Q�\Pk`���ri@B��[D��ʲ�W�(��C	��ں��լ���n����_ն��{;������� ���V�(1����x��{���5��g/����ϴ�<�o�~4L���(�$�F�{E�N-y5��(]��p�����3S=�n�e�y��¼����KjL��?$��z�sP^ɒs}x)�6�Q�j ��jnnя���p��j[���g[�+3r�H�݊�n��ч"uc	�tG��/�B)fk�3��|�*3��H��)`�$a��0��9L8I|�S|V�p�8Ы���<!Ò�f�_+
í�_�����~C��FS�	W˷�n��$F,5l�X�r�m-W< z�֗�a�2�hp���GWp��:`XC��4z�"o��$��L(fy�2#��ʴ�鍒��N�'�p]� �X�r��q���mB��"	,���L�3�7>�Ӭy���=��V����l=�D��WAq|��u$��]�{�t�k�`���i�(�E8�j+�&��Me�!<첡���ݔ���5�ߪ4"ÒkM��t��Y�����6�Ů͘�)����+�0A7�^a	�x�i�R�J�	>�27-��*iN��-U���=8�~�fP�P�а� |��6�b7��\	��N�/���[���!�8Vlijo4]Ϯ��O��8�c�.��el��At�FI,5D�ȡ�W�Tg#�s_<�A�8��zb#cjw���0�n�&t�(�v�e>�A��`�7���e#y�9��틈�;ŽL�����S�B�!Ap{q��M�ZAn��
wv���9t�,[+Q�ޤ�)��,���q �&�E�o���w��kny��M��]�l�ѫ��ކ�D�Q�p�%E4rw�>5�,tL���MM�r/;��%]1��lN��mL!���*P�)_хwIz�䅧<�a��J�؄%��1q+���D��r;Aw�am��?-�fS�v��������X��`�+6`A`�(���:^r�z�P����V<�(d�����
��\/nl2�M؎�Jl���L_����[��}�M+��*�i'��v�/߳/�&^]����-JSEJz��6�z��U��{�gY,p�el�GM�H5������L��7�j�0��B����ʏn����w�����tu=e���,o?An�4h{��ު]�+�/,E�����K-�͵��$�p�X���j�rAoӛh��HH�`L�^?��pE��.6,c��\������5hm`wvn*�1��7�ͦϲ`�,�6�l�A=1I�E�rB4�,��Ox�X��t˷����tO�Ƕ�H\$W����'mA
%f귡����m{9G��k�>6�����q���L�`㕲��~���Jp�����_��S�5LŔg�!���}@�y�p�J�t�nc�xf|�z���;n�� �h�`��ОE���x��-P*D���M�q�(IP��j�9m���ђ�*u~ttM͹œ�ۄg��yId&���U�����s%��ϑ3V�'<w�4��9[���#o��#�$ɲ�kT��:'����?���8N��ԁV��D��t���<F� �轶T����o7��z@�u��M�>E��mL�G&V�"�,��^�b�|�w,�^� ��XQv�b�za�c��)�X��z�ENC���,�ʹ��<�Y~?��@qy(w��%�`[��P�"�8���'�<��Kk��f����Km2�����O���M������n�Z7�Z܏I$��۷>hz��s�4���*�[.��꺝G7�4��Q���)�M��r,���58w��,hl]�����FKYH��J��u`g�[��B-� �QzŒ�"�!�f�y'�"��|`�O_0�\[��G�*�RG�� �f}Lɧ�˅TMk�k����,a�^<����}���b���r�gn�Q�H&��7C�}�S�y���|�kW�q��_�veQ�h�����|�*��
�S~f3�Uu���f��>;����*I"g:��ɜ���^�18�]�d�O�W�9Xh���B�Y8�]\�l1�${�;��� @����j(��Ř0�맘"qHW�$�������C���|j[v�z/Q)ނB�j��;]�+#+���7_K���W�_��L�� �|�ã�܏ ��S,�k7����.��6x��1��^)�v���b 	�'�[���D�H��O��K���b��JX���`wg����cs���c��4�B�� x.�ˉ�&�n��_ɦ�֙�x6'5dsW�>���Q�*��i�?��w�[�e+ݽ���%��
\���ܣNm�(i]������e�D�q��f;��.�h��yXx�_�\b�؎���ׂ��>p���1�]G�=YJ�w��eV���An��(���Jj`�Q3�m/t�\���40Oc����!%f�G��_����{�YpP����zu���בD����6�0�����y�|��T!B���X8w�儞�HxRaQv���>�����4(�8|�pF�E��C�L��JeܸJ�zC���GB/���G_-W|$�1+�۫�>�.h�Gt7r3�1Of��@#T�S�؄�*����O�%�����|,��	<�{Ae͓4LyK�)�#ڇX�5�cT��"W`@n�i��1R�D��,}�/s�[\.VJ�
6�e�*:�0�K�����,�� �8�h��6��O:���rE���/�@�Ù(6��P���]o�t)GA��_X�5G,5�T�Sn��������@���y�<`@�D�	���7��<L� ֣s�2��1
���A�'[�%Y<�d�/^i}�l奭>A�v��ǛYf�U���T�f#�.�0����<� 9���jA�&�g��ώ@*���>;A\USצW��ˡ��e�t38^�g���n�ia'9r�B��V,4�;��M�Hڻ�����)²ʬ����-v�:��%��m���'Ze@��w)���tP��������p�.��[���g������B���[B2�k���Tٶ�8�a���.�_ր��K�)}:�6&�M58 Lε��fƇ6������f^���OU}/˯�j�7��9��YSZ.*�e� �r����Ar��q�-02���o8���?��Ao���
���Z�^�5���/3���09
q��ǘ䡿l�Æ�{e�R��\*Ҩ�GYZ�w �"vs����O䇍pm�I��W^�X��T.8�;�Wi�� �Ul�Cv6W40o9؍\:#�bI���1v?��8�Ȋ4Y��v�J���d�q��mmv
f%�"�Qe��f#DV��^��%Sn��6Xщ��2O��v�ע�a�e��C+$��ￜwj��#�%�L.������Lbj�^��y�����f͕���䴧��YI��(Y����a#�8gF�b�,�qX7]����%�(�������a�|1�j�v:��}���x5.�S��byT���g��/*m���j3W�����kv4l���FWwWO���2Lq&U'�y�P~pg�nz�U�K!h뚕�����ԡ���˥��ਯ[�@"�%/�J�d��ψ�
E:D������CO�4J��	y�@��ۥ���ӥ����8��d�5T����ė���@��!�nu �B�,��_�tF�w3���;�
}�쳢�J��R-��?;��DrGe�|S��ښm*��1��Uv4w���D�Eۡ�kn4�i���0\[U��!t̫�0�U��yK �|��'Ÿ��>B�m�n�٠n�����2~U�M#r��ޚr���_Z�+/~�_��_{e��]_�J1kB�і��9r ䷔e]!FLz�ԝ�Rl�'YpJ�a�ΤR�xm����똏�ܘ\ܔ�).�n7Y�uU�.�_��a`L��O�s�l�)�A����� ���U�o���k����R>�V)@6��<ge����[-�h�lߖ'ŔSm�	B�g����#�{鮨شjx��U����B�[rK{�- ���G:�U�8��S��D����J�@,R��.e�/��A�VANQ�+N{f>F�M�#��ˆ��_jEB���qcq"a��1� fF��=?����!F���_�˹V+/��N�-���~��&7��Д''�!w�yy<�1�`���$�m�������߳�liª�xij;"�q�[_{���_�����8 �~wì�0����`[LW������6��e�<ޚ;�}a����N9|bE��[{P�H�w�����Dx.ߣR���k�R�'c��]9�������6�Zc}m��]O��)A����F�1>QIRi@g65����p�jڗrP!��O}s|���ſ0�\�6#��rɇ�m�_��	�C/&0��T�!`
_�;a���Ca �n|⿽@{���у;�����l�[���P���p/ø�{F�,'6�/eeW>��!@�/;n?�hn�y��a�5��@Ah��bNɎ��k����4��u�Mg#_b߬�x�b�9/9��"�=�3�W5�xݜ��1��B��p������6�
٩¥Ã�j�.5>���8��S2H���. ~�	/�N�˯J1�`��BIhw?+�m#b�P��[W�lc{��f��gH�|�'���*����#�T�b�Ǭ;¦����{�9�F��)9+�>�{�d��J�96x�%�[����S�)^0%����Ƀ9�������ʠ�]T����>%�/q��r������m�?2iP{ԯf�y[��'|j)�6AxP����{b=�e*��3dR�����L/��aoEH;@|�N-��S6%}! �UЪf��X�w)�N!WU^�7[�6�{�ѳh�+X6��ӭ���6���TD�;�Rr��]4���*K<�: H�Yl0��^��ǔ��ye+�%�$,�.k�D�%>/���Hn���S��3���n'Gg�	��2�hѕ��� PD$����М!1����m�7�Ų�6���������{��ʴ'n�<I4��d���,,`5�T?��P��N8���o�L }0DO��p�7��{�lQ0U�y#jT�Β�}F`�d=/��q���
���W����`��������m"�7�W��R�j偱d@b��_�}U���x�{Κ@a `�ʺ���:�6�py�s�`������A�ZQ-�ڟ-<���1~�-���*/���9O�~�T���S�A�T���]9`��6��d���ݬ�\���0
��j����Pxy	�MA�N4�r)o��s3D�<sG����
��Z8��!�I�5=������[⑎��7G�]��ctB5��&}?��a��ٺ�l� ��1�R��t���'ֻ��=�&��氜���Β2G�`�Ҿ�e�h���ٽB�s�C��@��:�Mȟ�l��a=��?��#����D,�+Yl�a�
X�C�W�(���"~{>m����V�f�^\[~p%����#�ȱ)�؁�p�>�HW�m@���R�W�yeV갹��Ul�2d������d(^�6���=�jg;B�M���2��*�uzv���	�����,z���4dUO["�X|�:���� ��Q�pB�
901�� e7����1�i���C;B5Z��=�Wn�R��K'��U��8�Qf��c��W�}Csw�,5�=�àz��\t��Pױ��5M�<�)4Ch<�k���݋5No��k%w��jm���{ B���۵�� ��¶A�$���� ��ԻJ�QCElc�c���#�7�P��+�s�&�|c����hh�[~���(GoJ	�/�C���pG43E��Փ�q�VC�O]�)7���E�ժ� s(�����r��D}Bnqב�'j�(�(1�KBt�jɋ�`̵1{�xu/�h1s��;x@wp�,g�?����47\��v���끅|�Q�a��烇�����-M�u��KXQɳ�KWC�N���r/��|\Z�/�`���	(3f+���;�b���/d2 �2>H����r�.�%���":YAS�UK��NXhx_r����5��T�*�1_�|/���:�X��@Ȁ�P����c+ǟ��t1��(��,����^Gv��@�:�*���a��FX��#!�O�Z���Yi��+q��R�蕕�z��MX��H����U�%�W��-���a���(ʃ��3�B+��V¯R�P�4��v��\p>��ߪ��eX��x��@�>`�v�b�Î�7���l�������]�={vk0	��y=Xg��}����۳�&�bj�xo��(��q�V�ܯb�{㊔�n�2k,�w����<�̖�ƈ�A��jbN��Lar��\��6��}8���U�q^�6�[�mN*؁�L�+��t�@5I}���}���M7'���]���?�7p�n��{��!�g�M��4�� �U	3�Ļ�ŏ�/3����Y�:�c��{�&�Ժ�ք㷷��1@��u\�D����bo�}�� -Ɨ��R�X{a�5*�T��\�?��.ƻ#*�S��N��{��	it�{$�T*'r3�(�7}t���Vu��dhO7�G@�e�=�>P�$ ��e����S�L4�ci�g����M�x9�1�d���ޖ�K%�b*Cj��]H��N_o�-�b�S�H����x]�Wԙ��yBJs���tG>�:ø){%�H;��;��f`�v�,t�	\��z:_DU�(�HP1�w��)�ZQ�����/�[��r�g�v&� �?m8����LA��F}������^Φ��66*�9�n��@m�1MTVY�LHbT�T�C��[nrC��Aü:?�I�sv�~��x�%X0e�h�U7��90R��Te,n�%���d���z�z���辮8�a-�z7㇣JL�ym�溃��y��̠@Q3𴀲0��������kb�v_�|w|�#�� �u�[�4�]�"F0A�t̷��!��3���
1�?��{%M�>��Yk��S��@����B�����[�������r��}Yv���[B���)�}>0@6v I���+s���4�wW�l(���%�V�u�@�>���0�1�ݩ�gV�}3Mzb��a=2�7�Ty���ԍ���R	t�I:�l���
z|r���!ZzK-\�WN����8��!E��e\���ܡq��K��	���I	_ŔX9���Ȫ|%FxӶ��0f�j��ɾ�&�iꩵ�Љ֯�3� ��|�I�@������n
�9�;*���z�R�/ե\X���U�90���x���IVP��=�L�Gy�\a'�J�a�/�����ݧ���O�n�J�V��d� ��߰���e��H�3�Fp+֐��uyy�]a/l��ۗ%��*+�W�I���ۢк�v��Ju��WG!�����~�mY���\`'�g�ᨁCķ��8/�U���6��7�l,��������.|��6
���O+�xe����{�n�l�G/l]���[A9ez��M%�f�
�ʝ�ކs�a�h� >fu�BV�
���#*|��$�F��KvB�o��q7v:
�?��"R��B=�\Ą��3���G`5li� w��B�؏%Tf.d�xkN͎�N]E�|.����7���!���
9w�]���s���y�������h��Md���vpL����8���?�?��Z}o����8e��hͪ���z:����1��d�NP��b�g�����VO$�
zW1��l�l�dk�5ըZrriɒ~�C[p�![�&���P�k��<�����6]6�d���ɜY�M�z��[l�E�/j�����v|�\k��4!�}:�>��RO�1&�t:t��H��}���9�K俯�����l~W����T9����}6X�fMt02D���Ix�5H��Q3ELa}if��&�4:ԑMu
)4}��]��Lݻ钩�:�����c�p\���z=J@�W�k��&!SNX��Z�(�"]J��9c+JUNN���*�r��q'3O��$IYg��!��W��C�)�m������,J�u��IZX��� ���7����z���-��k�ۙ�Ek�G'/	�8��N�����5�R#���l�-p�򍊋�3��ض��zJ�L�B%���.]DB�o3r�!���cV���A�]~,lW���V�a(շEmC�