// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
hm0VBgjr+2kfjUOMpoMwjC0QkbEfYRD61fcqV8Pny+21ywaxHSRhzV34KAcJztt7YAmisby74fv9
8fbcnRpdG9hp2TtlFPia8GvTA1MK0iXF9VHFruIjCfmj8G5o+4vkuh3mlDQiRcew+gK9gdA2meuU
MR5wrpYMsArQkZ+i2mtfz+3nMJMuYICJCuFWlEojQ5DhI1brAY6BfcrznbpnfBsCPAdfPiUCFnBK
foIn3zDTY2GPozhVe+AUk12BOKiHyxVKwLfwtCcyr++eX2f0GTBfQ5UG2Djfq48Ec/z1/y9zUcBr
Bv+uQ4BdccKPmr3Dg3wW12V9BghibIorsFS9EQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
ihb4ilVSpq1S/7yL6p7kRaOkZq1KDTA9PNYYGTEQEel8etaBX4uMyp5+ZhBl/EvhAFwiFODzjO7G
VyfNv+A8KB0F6iryBS3KZDD0oCbd3JO7mseDJ8yfTctZna7T75HjYxU4EUE/cEUGyDsFb0mRo4a2
lUyZutcMUsDUfsPZyE4kmfVpxC11mx+sthDKq5fOg/va45suZM9hazR1GH7OijW4tPxcSS7m/ilb
fvFnEyXgy5EgHqrhsX3047Y0ttmHBJm9af4t0lvDw6DRIZNXHcXqcFUYlIgubmgH//XJgjisUctE
ankqNzakNmAEB4kWwtWfcvpS7XkBdDplBtNYgPEFl0mA+nnq+Yry82aTbcatMxKM/qxH5CJPZZiJ
wvsIeZnOeIcTD2V52qP1JHGjsY/ZYtjUQWY0dy8d3aYJkOcR+sn7PaWMSji6kRhPgxtpdDpI8a0D
NZWeZp+/jzSswppa+bknNwF7+cjEzhOT5c3gAcmGay7c/V2FnEJ7M89U2cyP+5Sq0gPVTqst0fgB
8ADOsNLnYgauNXhAtBdhzIV5eloP4hQEiQl4k82y73wHVfJERxy/BehOTZCaIZn7L5zd6JXJNCtZ
VitZx70OpCV1JVJ80p6rc+Qv0LMwHDE7KO7l8+HAOQVNElp/Pomr9Ov0ZQU1x/thVMg5zQ7Ch1m2
3qDuSjRqeJ2Nw1pksbHk/z28Lhc9M6UMbyHUuWbh1bJQCIllaMTI0o2SO90RxFNwU9MmdJFiXEhv
wLfOMGd7rm62Ly/tmRmA/+AKIfPwGhj/n+YGMRkRm1TIAGvcDXXwFlq7QexMiSgAg+wwAwvUewjZ
LV3qvde+45ZpJCYYId4k3xYh1bxUQb1HS9d3KbxMZxy3tCV9FaNbKTcwDlz4uYG3wwTBBmR8GXPO
cxldRAQzXOmvBB3KR+L0EF6EIb/8dtJfu/zFF38xitRsayyrcvFWjbguBtxgArF8RlRA7HU3ioyo
xXtTtZdOLq/xvPb5egKGAN8vayZncTE4McjEUbdBkG3hSX9L8uC+kCgQWa+CNDiP/X6eXr4qxjez
g5XkQh+pk1ts/dU1g4fYbeSHlXmX/+KwnWl45AAE8ZfgOkvlvPUuOKNCFFGCebTFGzt0dKB4T9yi
Im9trw/XM8pwswaSeOtf7Gz22HjSmElc6HyiqR73/9ab7Kvc3clEuUXVA0iMJWF2rfIE3LEV9FsQ
vvqWA2jha97uy2cY2MrXVKdbAP2WPN458IdCR0CEt4R1HROIDC70CmOecbou5r7KiS6F66IMM3EZ
4eXVdmomGHQ/xehQJ28MEQh6VBxuc7wR/aFWGLpRza3OrSNMDL5UkDZ6Ys67nrs/1yiQyPEa07bG
kgemPUni49x8Fnr9S1sRWKQtwL5bNEzfvHgpqb3gIRs3Ikxvaoz/xbLiKxXfjCPn9y8Pw3p2JwQw
RqyeE0cjVDK8EKRMHOjNUd2qLMfQJs6IjampOf4KYCxaSRlNrKf1ztUY+8VsRE6FlwfZO9y78k6d
BxqrhhkmrgI1JcvPmalXBSbFyU9TXyrISPuxUUd4dlnAJcRv4vJjeoz/7WJ5StUQ8wdmEZHCmWBO
8o8mKRdkUQ2mg3MKPEQylHTcHTEL16b79NAGXcQcZKAAtbyZJhWXHkiUZRnDw2AxPFNnaVcK1CmI
efhAgnB7Aibjtgj4X1kxBUK7X7Br3YIlRrOHdcKgPzANVoJjXGYBbRiEmfWSHh1K4hE1FjgQ3VOJ
fVltwT3cNk5nIwCizTzDL1Hb///uiLx9tlGrQ4/AD+vfb4nqokdnRdWwTeISgFXfm10VVHndqvgD
g945uKir6Rl70rqSmhVPqkVYdZPP2afJrE2iHI9OTLghjFf0jXs0yopsXmMikeEOuiADYNOMqPUV
NDuUSLX+2ztLCd0fLJk5ifvTpD2QiOOoO7sQDatXFBI6LzcF/Ubw7gfSrp2+MfISaK4GE+8xAmvk
WJBHdSgdjCJ5Fc9N1cPnKbtH6qSzwg7vePhIGj92iTEXl1xinVDcLcAV8B3+m7Ek/H+d3hyznYfD
1jTrNb/Ww1qOSI6WelaOxcZE3iT/988/pBCPVaylCJg9IQHgzQdk9ecOgZ0YCEjpkaZGsDp3V9Y0
52BD6MC5orF8aWiuJpL9BNxiDRNakfdA5WDxz2ZDX8s8tEn0x/99qFpkxjcPqWHnt7RX1sq6QGNB
6sHofV0z1KxLxdg1mHjy6Izsc6yQis/LW48U2DOSrYs4PZg2Lfq1a6rB7hZbaztJLKNWkCYJjbQn
Xi57XGZBq79pkG4eW74wFuFh4Zp27UR0nXuzA5rg8IQ9VWYyJGSclcBb636nYvCj+6mcHY5s9g2x
QzywkRWDHYe+2Ng6NdKNaNAEZ3kux9pqj2Yc9un2pDHcfcEKnCMmSQIliPaWEITGcXBZ6ctPHh2y
Um8v675eav8gEcgUuvLA1TBAw8mgdR8ivk2pfFgHA/ffCAGf3Jhw4/aozTEgQep5XuoJCTPXJZ75
0EJn5EIMdLYiRA3yVL7M3kDHj1j3CF0BOJ684scJ560mWqUQQn0fZqBhfDk4uKSlAQwGw80/E5JP
HJJHtgsJxO5hIXvnB300BVcd/4+j6231oNJ0/kXgdJH4FUyWrncyKp6wIzm1GZKc+gKsr0Higyqs
I6lEWMnvD1FiRpbDISH2fND6uVKEJX/1NdEgb9AeWBGK0ovJB+N5eyhG1X1ghpRE9sN1SIDuqNSm
NtwBGXX2mMMLWHfgSkFk2rWqLCZVSSFpifFsap++yfdaPS/iL3iYcvuTZxWfuw0M76Lrbnmw04FJ
EL3O59zDZmhmAeAOsMyE+5CBBs6u+kUgGHsFi1rUBYfxFKcTbypiPduVKFiWcn9wpuFe5b1/7k/3
faEy+1jEngCbFgdJzNui48qlYFv6fx/Vs1rhR2SGAkKNm95aqvekyxiGURLXE/wmXozagi8eWE+k
TecRrWZB3Rbh3Tyfa2jAy6CpA+ENlL1Z3zK31cOugLhpgfFfgy7xpYFrC1tGZQYILIeeLyXpGa+e
S9Ax5fp+NZJg9dmClJ1/cPAK2IC4RZa9T7aUF1ZXIOCBvufqkK7t7g94idDLCvaRsHbkZYH3fca8
Iz8eR/QjjWm9hFyWljwuYhN7WGYV9LdvT+EMuevtgaKGqkl/yb8s/MThdXyrkESA3ck7pnwPcev3
KWJMGmxQtdMUVhbqXompk3+F+dRkhEZgYxPBbLABAq53BlLUh4U0fCC7dOIr6ziGvDBml9rluoqV
O3m8CBYNG9VYd9E+b4fOLabtivoWgdR5/iVIExmy7JAZIipQtDqzmvl4YLQ+g4q5DSrMN1Wy92Ij
Bjkws2B0Kyt6GHJ2VhGqMqMZHLoOvXbB9E114K+BnBf6NSIhtQCeQrpCQk9gRGFdsf+xYLB9tK0x
6cEOc3DUs/28kPLa59LTo0cmOC5neiHVdGc9lRed73C2nGBKLw+EjvzrlXybaGWa78qqtXA6x6VR
uc84LVkkVD/9RYsE1j+Na0bLKAxMM1XHjJAmlQmxHaFsGiRb4dB39PmyxafjoCqLZ+S3/lUiYhX/
abdVOtxLCRX3gN2DZMKr0z+8UfYV7opSRy/r6bEi4A43OgfRRZ8h+LBxmK3h6C67aN+q0teEImiI
OnSWy9qL3XXz3ZbkVrnV9cfpXx2Zc8XIh/RfXO7LDZfStEaA3iVwxO63yaJa7St/DZglIImVc8Vq
8DBtDtKlppA9+/mquQXFloSAk6uRVLHweHoeTR/V88095KcVdZ1YfJL2mmGtQhtLVrXqXYr3hRCH
f6yRThDqGTleqL74VrjL5IFidoD9wjTLtsowYLwQCnKZqPNGWREncwWTABzci0r+EuiS/KIbk5jZ
gYfXmtUYCAy8sbkpGdobnIoUHCaP+dPZUz17DKURDpL1nNfSzYuyHKxKINxbmRcij1Zc0BI5eWbp
D+Vn7FpUy7Jl5IJiapJPdpxUFDyTx5Eurnpb7XxoTgALwyvQAP2Rzt9GLOPK1hOWRKhXV5xau+Lr
eKJNfQ5Wuk3LTWSiAHI5ECYAMAEaHi7k87AWjiZa+VBMZWNNtz3L2R2wEw9oucmtVzlxn7kX9IK3
zqnT907pCHojtM8ishI033FLke5Nzq2VwPkpvURgQS9pP2aMemyxz19aWUY+QBj8aUDvbkllCXke
MGmkXE3Vs5iEHwRpaQkZZIYij21lULV26A+4w46fpezBD4Jx44pYI/AQ+HIK7NjCC5zwxAZHKf8Q
iVKVKW52LQNHT3wNBIBlFlaFQql2Zkn9u1PVErk/ZxMiK+CNpLRkm3ek9+19GtQicYV2aIqLIX1K
vC+bWR6gFFUiVTyenZbbRtceRPMCJSqdmrWpSk2Yo6aGpkrJqSIZY39Pr2ycafgmDOa9lUKHzg49
+Lg9jG+j1ev4E1uheXaNjq17hpTXHozoYs8XpSshRPATvU6kDEIZT/QLn4s60XsrGEJAGmQCzkwX
DBp5GsLmfh39YYEOkky+H3VfcEvi3LrzviTVyCqy7T5a4hDDCs13jmPOlIwSTGNbrt9idfjWIQR2
LwA+Fy5ndqTvlB8Xgs8+vpBVT55GhdGJ0hG/APnyQ/c+feZ935crTF796z2SzD7oHQa7jvDHdDAF
oJOaIWfkm+5eECpaqAWoOBI09g1BN5J17ko9euMMtd12uT2blnDezDG61sI9DyjzMhvM8yCI8dDV
cfYVKgJddnhBEuBP5CYb46Lwqo0k7n4UdeGeD31gMVLg8g/w7B80PUes0psdEuCST13gFIVcXfYH
n0RJnwNwfYZaGU12PX/wQ2Kn8ESb627JkHPuPnUCsVXW8AZFt1OiyyzkzArz28hp3gNEPGfqbLZo
pXjW65JI2ep0xwH/8vj0SUVn+ZAQFDNfKA8e8jvbIMN+JuenMrsaVNmC0QbR3fc1i6u8B0/+uzuD
JnzhyhHQCvfT58JskevARfzc6adD25tBujKPlULhZl/QAGfL+Jd8EihrVT1fsGKYKUqBenDNPLqT
rS95oLsUhGDD2l31tdkRuKqRa1XGLTSwgmEIrMd0Lrqjv/5ONbgxlRWw2IoMhRhN0chpUldPSxuS
sUTDt5wTCmmQSE4Y1SuNLctDJJ5zIlGb48b7/XMK1Iqlk3mbaBRwDAA514Fd5MtiSmcVfuF9+de/
llSAVNxDRU+DNOB+hpeQVCWdbU4p1D/zANRGEdwT8IciY262tNsNFl7I0b+vMuv8MQRsAsIAjjad
W/tyoAbZtr+HXRFvcnLBeqILtqbttORyhqjdYS+wIQzAeVoEPoDGe8yM9veVbuDHDcB+vWUBSZoG
rozUHQs+x7b8dmGIvbhZoDsY/1J4pGL0VTFQK8lZX3x1pUR46DK2xuqrBv5kY6Hn32ii8is+ha7f
G3da2qeL7J8oVjNoGDNHXlJD8vHpQVRk99OE4WuMmFyf05mOA0WwFKl6vN1nl2jZqRKhAzzNm8KM
az2jO3vn6Ja9xGYzkUZ7rAAUci/fgHO4IIgDdQF12are20WY6HhOO9OfTOvXlgWvaxnTojuRMQrm
T06DSVMh0ZOiVhDoMdy4grFcxoQSlc6nX94j+N90UesObk93vhkmXm7NhTEKcSpQr/c1km7LzAzC
+STHYKwUHJqAFLbiKBQl35eDh+nYU4oRJoFYOu4dNRc4TnBNa9HuNvokeoOOzP44Q2AOcNKHh7lG
c5a9F4Lzw1WVTiMGOMZ5G4NxCiEn5w2ASTrYreAAiaR1m+XfnMMX0m/zNjmxq01rfxVstiJ6G2S6
Y0Em8CY7cdWikKLSYbP01iA2vVgGjyEW3fcTHIy/937phSsZmHwCy0xEWmmpfbPIPi/+l9GkVP8m
SS3APLYEHS1Il+IPYdu65BLl7AKMNiJQumzm6Vmaxko4MtaB5Pi9IlzCSFHkAYuVecqV2cW0Fya9
sFwyHsYDAv5O7AvThj+rTr+oCcD9DLSqq/fF1XYh+xs4oLCF3WTgWud1oO9CPcfeh6U8IOJe8/Qx
34P3DJz8YhYhE1Yq48RG8MXs6nf738hbZfI1n+5va+rW74U8yPKcP2v8e8L4oCGcXeeZK41pO6E7
iguXhGgUh15L2ONBRqu7EjGsD57Fk8RJ755fEPi9xD9amwSY4umclFMFiZnG+hDITYzSF2zyAOZE
LRqEf9CN17i9O/GbeZLNF/Ke67koyMqHlMBMS1qBqBPIPhCdQ3xf/tzZPknzFMCyDkz9X13IUHJB
BkPRewzC0tYCJRiJgsU7a/Y5lFicFzehzgKpbdVLEkug/47R7Hr0X8T4r2UyfDL5LvDgX8t/mj0g
j+mZlGuYSEno4mrlLhspiJv6CaDyjk6Lp7yuzfxcdZYRHvuMckp40T3XwWc5znMQcoE26/hXOMa9
ByqVW+V0M/PhQUMejiLjnKLJzN8x9C4iKyslkPRc4GtPJBDjEgBfNW/w04oVdt5Uh6f9hFaOswaB
XkzNpkcIYql/8NtAAq3lU64sh2uWSjTJMbHXX0tn5eG3BqcBvh/iSvzmcxhVU+2gPczIQYfQoMRc
cLOrCwBW4hMav3K5+Xe//31x0bccnc+J+ZjpZDQ7iJDVPDjYrget+1yy+CfnIsksqYN5hnyuHT4E
Qww0dtWOaCmBMl07xak4W+hRu8fKT97Wqlap/fBT5lquLOU49VxvuPPzIGS9P4908hcYaXO5RE/c
1B3giv+vbmvnu2D3d2pJ95l8kqH3yGw3lKrJK4KAOa3iNOOmVPCJO83mo/pXFmhQMgk1xxhqeTlU
/TJVyvgMbOFCG8BbZpocMP7eZGUizoty/NekIIZ/Ekum0NqsT11L3LX1ITq2RaJ8+4TUqOdML5TE
mHTxPc/ET6k/J8CZLvUS/VgmqetUWGHy6XljD5AovWP/kdxRKf9nAWESac6wSWMc42iBlwJIyEYD
eHwlz9F2ah1lIRuOOj72MZz2kAi7mLR5cixyfTjkFruCiwFugRTT0rehCYFjEZqwcyKp8OtqPla/
8FoC9s1NmrI/VcLFkd7dHaFagsphwfdXPaPmdga3H8KDcJ7vmZSsjkiJaof+qFMl1oPhrHCVpPrs
CwiodAqtOnE+65kr2dhs9EGPav9EV24RqJLu+BDEwx0iZfnQ37EluT9fO5tBoVR4xd9BQO02CGQ5
oqldTW8dlnVDMlEixPylTDQQhpFPNJIGA6EORWnC6FQNSWRjvtaeYAwixiXJkZ7EwpiKKFf3fLpj
4HDmDzdLy2r6dfqVb0aa7gclCyFHfY3twic3lUc90lA+t7mJgMOv3Nubpouv94tysjmxk48OrknN
0MiRjJuTVOr/ki2bmv0qgOTvNMuk7qU1W/IcDxfMxPP1WdqiC7eWir7S4AltIIj+WY2doV41DJNc
KPU9V8par4NPswBkz0ph4XJH0AlIk7bSFy+ctNKZvKJ33J8rqEXEcScyoHkfTfFIPpbUC5IZAAz3
gTd6n5OOARRYC/qzxHxP5aJLRUU3peADgkh+qwa8V293vYS0hBpqTn+kjgXdbtwlaqmgcqT6Y5V+
cnrUtShHeMxzvXizBbvWHVP2lhCoJhiwvjJ17oAZLkRiR6ibtiLZ0nJx84Vctjnx7eLlqOI1JdPX
tZX/YQP0Sh7FRdCejt6zIqq41kmGyYs4RuV2/MShNP6ozEP4w6ie9h0Vh/zPKaE2JoTBB/IfJ0WB
MLD+Bdf+4GAHjTBfN5tPs+6gPeuWxTbzrZKvTpPKpMe+DcQ7GfbdVuU+xRw1wwAhw9IkMh2LQ9FM
YrxsSa7lvXFOLOmUe+R6d8P/sP+Hcg03zlSv1h/TQU+U+zdxYvQZtAoRgME4z83i9PysrhHKJ/Rq
5ei5Gmg5MI1CPbJ/0tn3JPttwMUYCK88kD8W6XNrrwsJ7xJqYqcLVaHnijQFpVPuVrXqWs1RvKai
6fBpb/OYFU0zymx3og/9bl7blBBWGPxtYIqH5DDHaFz3LNFgM1OJcsvJS2vQCgB4XvBbnDQJIj/e
crnHlmGD9jJxh5gYbjV0Q+95ksNzQrG7NoLLJgX3ZCS1I3IR3L4II7UGca6Gp3FEweaXbeMkoRFj
/vPLxEPm2vdTCCMlZvR0G2nsnPNKl2fDvoZNIu6P4iooh0GKbVVVlHc8awfveoizSeEc/MZYv4P6
GbSgSiwK+AaTfdbbahLNc0XbBuV8ql1QuNWPi9Lri6+QudaAqZOslOLbrleIFcXG41/yAnTm3rKG
0YmM9QwZ5dUkwLf2gLrgy9aSG8CBZQd/usXiMZMaLGSPTAlIqqGr5tJ3Yo9ozUPMJ+MHbvKg7O7M
ztcaOrL4a10uqM3UPZAVFmNRYaFeQzC6SEAk4YgWFEvklGD4BvzAl350y8YYgz4wRHregvM1fFq7
foHDVhnc1xzCfJbLFIwseC2khZeJuQy4gvvoyZ4zzYRApt9izkoSDfxL8dN1OPQg23uTvseyryK4
9rahCeIXvdBBWkpHqN6e8J8TTocRer27cwWz8hSwJyIwvlSLfxb6XeLojGicERfRVM+SV2+/njOR
Ynk5o51bWoXDh0dq29Uymf/wfwSsNf10yfOXkLcvxWQfcyR8g3zkIlrjSKh4Ku2z7/i6xczBaglN
N72vuD1vogmham51buZkN8PL1GijFrPo6gyoc1w2HJpaFX+lcdjaww/8TqOBIlWJ+GimzPA0swZ9
7Mq1dXU0VqVyCoIVq3IfMVrkX39YTU/GENpqSiM+EUNOnMk3E3gqBYwl4TK8V7iJPEjwiLJSQkp9
lsmtiTnGJGiuY3pN8REgq933aMr9/uGBSst6ba2q3oiKHFJ/5CK60hCeRlO+sS0ryf9qEsf14u6Y
JA8vP4s9OMV8DDAW5zQbUpJEOb3vrk/ZEaC0Xss1YnN/hJ7Yk3OcJkcOrPZOSkJwVOvorVWDvFCI
cbah6c6qmdfC4BlB8ktgcCFDyOEGDNU+hULa5B02pbFT7JCQmKKzijRdBtdnZZ1yB4tcFIdQSWhC
I7kxyOmoiFDkY1t4gyjJImf2fzIC+3Flkf6ZQKxeEf3aj3I563KHhPW/wAbVzB0VjqeoZ87lYs8K
0cErTIW65BJwbmVvycaPYWz5ee9rPd1TbY+uxX6Qov6G/lk/PSkG9Z+lJr1Tin5CFAHiocYEYlGc
0S+2FUDiQZmF+OWIHuziij5hNNO3jcucSUUfDY8VwxEi6nU9/eSUoEEr3/xnrwDCtI2+BboZqGbL
Ug7a35ASkfqLEHablASdzA2oSrCIRY0Hn9sVhKE3/4YCEeKDjsVBsHtTm7MbZj5YNUsi2CLt0sSc
L0jQhK9WgZLljpiPRTfVydSg1PzdWDlRk2CN2swD4yA0K/NCuHtVilve6L+Jvv/9j2inJK4ux325
sfnY+sDOuXtW+xxBKaSYEoQ567ENjaN+IE8x9yCf1LxPQrYn+YY53UcfGJjpkJ0fE0kNp5qMNTJz
1d7R10YaFzeNSif4wwXcuPpSvnTGWLp9Qw9L0WMn/23/30UbJaYqedQaDYg3EKPAHh7X7mrzkzdB
6YL6K3dp1GKVB7tlZpAkgxioWl6XB7UOAxVoFNOvwkT/5ijSNqwUF1HIp1EscOSt9vL54M+rebZ6
sb2rX737FUnfKyZyl0rp5DhB6+SJz0l0WoOo2Vl6AabS3b+it8AWyrOsm0OUCyQq6F1ZA/SNeCHM
aMhmyG7BDiqrRAnENsmmHZCNd0KpPrPBoI9d2CYccAImz3q42aNylAXFk3DUbtIU1/0AgFo51WoG
u3RrUgSI2QeY8XdwLm/pJQbrjqgDiFeGYW7tfMu4V0LcP7gfV0Iku4NzxH5mYwmE8WVvpu4ILhjT
ZsIUoaglcXWSMrhcVEJXNgQa1y0JX1/0l3TZwRFVfPr+RvHvdv/lRibi5/BUzxxRvMO2uHaO2wwN
licUzWnUCflki9mG1E8Idh/sP1+BfGgiSCvHyQawVGDiUW3ZM/D6j6KD0smJhJVxrj+lW7z/ehlg
H2BOg6UcN3Y6Wgw9O00s6smg7pJpPJWR0rPW9OY2NxYG6357tZckHXDbxpeFOgi1JG/kM1XtLLB2
s5lzoJHC3t3FmlA36mRrpquUrcAOw41dRNU03vgnBIAhZ7GLnMS1TsDrgp6xCuAYF/zy1eCuxAzV
N/g1JFfrcQDoF4RrBQnJ1/GdP8BQqXhXcgupaKkKseDR0V/gTYC1tVhX5jmILOQi0wB4vJLojrHy
8NJKUcOjl0oH/B+4SH4fisapIEK6veS7WpsG5QMMTK8buc0PKImaDw7H1d3s5dKARvlKPZbNas8a
6oV6DQVgK7yqsUtFHgYOea8w5w6dSIgjBSUFxgnA2Ahc7inmssGg0ELcFKgCxApp1V7uIomcyCpP
ctU6riuup41bSdV1ibFevSFHa/76Mh6aL3/gGUz+EMP+fVMnLJzIFbKoUB9aewzlorgpKxWfY5NF
pSMPRKsK6+rb4UesGleDdInoz0Iw1XnVfTKUQO0k2xx7Af2dVUhJ5hVC9PYKGLQpYvdowrvzT0Gx
YTmawi+4G6vCN4SnfA2VIPyV7YYeQ4SNjBXq9rqlcPQzYqhphQ2JMq3XOjpAq+YufsFYUkWieFYJ
jUdEEOvhxeDSTRAnM5AE79sZtU3vk+QlbPOKdIlASU41/WaKfKKZaE0QLovheywxeOK6PC9zGKAG
3jP2/yNuc0laOfCIFF3j3/sBJWPnfuHECKD7QGrVicnRjv0kUScO7B0zIzXgFi1GACIc4YSy3Kkw
GB+QK/Vcy4y+N98yP6L8qTquCcM0YcIuDrQSgfxdlhNqk/SG0fQ6eQyOkVv4VKQdF1x1T3Exhujk
ZJfom63PdES6eX3mOyQLVW6DqiosMCq+Uo8IVBWbXWyLPAb+tj/mK6yRhPKAfBe7eZ9cQ+jwXL02
zW9JxRPkhz2rqEHGdkLoaxOY7xJde9OnwDotayHlKNGUtXTYA9ljnTnBkEU5uyWLYtLVIEY4t5eY
jzM6I2Dhdtiki1H0CAD1qeIhCBj3R6A3bnOoifT4OIPkIwdcOcHu85zyjD7RB1tFvvyUxZVuU8K0
ofOl69rBLmDCyYUwnH9HS0ntOY8k41SSv6p2ud0Y4jq/12p9QiX5wqTqzDzdsOMfHyK/0x019Gl/
RDl/G/zv3aa5/NuBYjhFygb5CnjGtFE2to5qGz1CqaSN2pU+mcgqgaN4SIYfvygWYhxrLkLj+Ryr
FMJr3NGNJdeNK+GbWUJcL1eU3yHkJXwfndkU+gBr8IvZGVw5hd8oNfaa/nbKr6LhZLDMYL/24C/f
gJFdAiOaCFkayU6PpDnKocgfXaFGTlN0V80Df3Rb0kt4ybl7yMkbQ6Leg+DEawVJLRmfMfdgtbec
0vyymzKnRNWwt9oH3ZWkrQQjWYLM4N404x0CTnSKUQJZOmpp91C9iCzhCW0mfTEoa9/nhs+mun15
LkRI7n7sPALg/5vcHOF4VCTOmwhv4bJ8lsIPheTokNUimIXuWSVjDGY1D4hLHr2lPW1imT9w48Ue
QR4W6tPSZWHGG09a2fIjyR2nHWEpUbeHkRiTLWk/SR4KQWzgh7FDvRHROOFF48A7w08xBfx3cu1l
0nQZoGrUConJaPMqnuq0lxeT4uVCpO3elDoPKCoekba+bbF7pnecjJUzM46IslCGqXkPnzX+GaCq
Y3T/M4BYB5XIrK6VKjbfqF7OWWPRihfLLbZuHSca76w/8aiZpte6s+kWDaDwujLdl0RbbRaRhNjb
hoVSZFiX9ae6XQibCIzRSokEWOroqZjKVVDt2LeZhpx5U44I4rTgjnCWhXbIPvShT9Afhn3QAPki
8HN/YrTFHP+A4hCanllZPXK5xOeZFOanlrwkx7ylkvd1dmUTOsqDAXCVE6E4qgSPLUpeYXRTCdBo
0H+Z+lBsrUmZ44SR09U+wXEN2YvK4v6vBuqBE6I/3Njq+3bjg8XlfMcwtc6RT9Z+8QTE9KValU+7
hxnJh+TenX/c6QDUXJqejE/ZG24VFNq+IFVCFaKgKV4fL+PwXKcE26jvf1mixOwNJBaIw8uTNxPQ
JWSu3pnZwgW3r9M7vLlmqAoEYi1NfAlnO7T9QdDgwNhCrNvk98Lyqp4KRwGhGNUwZqK6PG0N08xh
A4z1y2uUGVTYdNzCxh3zpxIzRn2pgk/B0jmiT2EO29wrO/s+MDTc/MpTPkF+h/jDacPeiGaRJ6Iz
bxRZ0h4h0j5Ka87woNEEG2tdbh8nlO0rS7p3bReoKWhP8BYbx3E2XYOdBOTgwXZqEexJYdO3IuAU
PwLotctOYaUH6rwsa67ubqk9ud08+AnDwrulotINqV46CuuFT/0hl4SiPLnZDxeRlWE4j49jht26
Fmi01BkYyBMrOXDKDK5NDHIO+vPBG7Ih1G1zuHTTmzY2GARze3T2RBt20Rba726jf+GW8XkJlFEx
bEhKp9nqhENmst7L+P0xvlwtKjg9e64fpVhm1tEuKst+kxTv3BDM5uJP5cs7WhyrU/7qmyqrq97L
dDFb2UncdM4q5NWHBawRePBZcgW1sLuuYqIu+LCUbjRqlyWCRt4N/2zU1qqVaGMpQ2tMrdNFEUKA
f/ulirZRGnWUPbBIIOyNHANDxdGVq0445E/SPq4wTQfazyrOUrvG6AJ0zZ1yr2yAbhzkRna62JlY
CGYQwYAe1zGyiVV/k2JBXqeMqd6SVIywUq9KxYQEU7JiPsoEBzHPtcF0xq+Qucr4G5qcm8cf9xDa
e3bxcG1ZiOldH1Wtzy1kmKpveck7N0WYyfVnWZhKIpZ4J1NNLrhAuDbtCG1URE+1anffFDWlog/S
xZI5+ZB+hy9q1JbfconJe1PSqXr1Zoyj3iGI7h1U0teo1M038RU90bLIq5NoLkucvp+LdMbYZ6NN
isIjYARjCU++VeS9+43QsyFk7KmJOkkgM4xvOiYRK+tQDG4rQ/RsKO+ZTECLuBFHVP9GBOVlTqEr
H1TW6l218puFkUJO9fiyNrdPYidcMeKenhnMeC4Icq6LoXo4nFPxelvdHOPcdx6uuhLafR+5iKRb
pE/oTDFCNrGNfdxoNrSuf7n3dq6pzrMVLAOEiJIQ0UYnTHBYMO4NBkKZb9vpAgFaKeE35E+FV4VA
KyZxcw3m+YD1k2RQE+C7jr1WalRxfSU/CpoZfI4HepZr+8y1SqLg7zIIzJdOFA7bu925wyMJkpHW
mGlNvnTbsuu3rwmCDu/XQ9RcF7/ip3JScZDN0DmVcWYLgeFyove7XkzKIwedjbBg2moKz5bFnxPf
YcTYaFguClF07+g0+1LcSmThmNt7mwCNo9T1SYOQpXSeD0ZVMj4EXgIiHR8QvAvowQpJPU6nGZsW
LSQKorI2uyX0u3D2ZURQFVUUroHvkrAahh6KLXN8CNdzwh5AwxdjsRRxFAa8XQN4VMN0ozLQyntl
x4X/N5bF907dNWkoHhRMmGNP7t22hW2++bteh8aQ/zhkzAYmRap6R5TOJNN1pVcRa4ayIlN0B5wG
+jr6x5SVGpBT3e1ETRueLnSd53b16QzGvxy20OgNuGpI74M4NgA0jtQ14A9dAcgU5q+OyOuiL9P6
JDCpiU1cZXLQpagk9wkezTKwRB1R3LLROpQHJPnNxnGfvlyK5s2A4M36yGrMHhnxn7JUM2oqQG7C
ikVzEDyjPH3x2GQCq+ZVNJlrGbHftG8eEwWXWZkXd3Xj8bLzEaS6WiGunkVzEsldfv1KEL43Zd4V
YxpwbXxKkfevMI1j239R7VIb+f0E8RWxhWg8x3h0Xa+h7+3d0BB/rjIUZtJZ9IisrVNEe6wMeaOR
HMTbthH5xFY3HMN0SaS/UutWwiko7y8dKVIA1JXjUVCpVMwR6FuwGfEPrNxDEYhwH2CXXGARAip3
q66wA0wIXK3ohxVNhX724V636eVt4j+mSi4Q9vHC5sQ2zxzkjpkdwYRHatnpiidyX8B7iEmBePl4
q+OY624vBiB1Jdvfs3TNnjPbUwPj4MbTjdcmRksagwpJQMNEIkYlRY8B3UmlOEop1nq2aKUccfxr
65Ru2CYe6ZP3BQlGuZHABYOFA8wjZz7HrsggJNf501QWiuin69BPeg04ECCYBpF7SRvT8gfNpXML
5C0Tkh/naXsUBoZlgQXkdOotQaoq0emOpFNi4wCbj+JuM1ECjp+r2ZnPS0U2ydfm9cyMURXM4TMj
JrZqYirD7sqtj+fU/CczRHI6aZ3q6pDX00/KZLUCF77JqmCD0HgZdxjieJY8qigIE9j4yjor3o7e
wuAIjDeNkRUQZHCesLyk/u8APiFWRwuCv2Dgdpz7IETVaHUlJoBjmW8StdY2BhL3/b7zdspC74Mq
8it5x2BLWjdTIzYkKt6mYIQeEBNnGqTjJL2BsbW4QDA0N2EIKgAn6/kIckFaTeMwp6oa2JuN3C/R
ohPouuCIKC4x56ug/nfh268iVBwcVjASLiSYtMbZ08OXKKCzp+Qx53bTI6Odj2nOEaoqAdK8tG+5
2dBwDN98z6wtVC4rEAhwKJUXpvqpDuDEHkKbl1ZTydAwdiPXan0a15kOnZXhND4W3vT1216vTPGX
lzhio/mHFIhCWLZ+NNjA+tN2cOtouvyqAi6G1RVJRunUiQeXIpE1ScjgGSJXm2YrkYV1wJ51Tvq4
lfOfTe6KFtxthZoJD5VD4w==
`pragma protect end_protected
