// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
BvSKH0dzGUoQA+iRZ7NR4k1x2V5Vs9z2Oc2R+cLVR7QrENRMVuH+YWcHpMCWyR/Q6Vilz690o2zm
NMw4gK0kcW79BPwEiDZUtMWjmmgSx3OU28v5sVf3RQdgTvprRgcegl+hFGMInuijoh8di5dvCOyq
YqniorfKigw0bsokPSCo6liCL+LogUdLJE5ZGUwkeAcKCalhWwf5UKqzWfmofNg9oDK9Mw2T8ynH
oGRp0Xp3Dg+75iCbt8qg4xXIRKjHu9LGPsWqfFhhm4QPYh2+LjFTUYCGtyi/KR0sh85yaktPe+hp
3bQrAwNtNaK96P1N9NGzeDFhP8wk0xlZPN6cSA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
RlJx0ILLSULL0tQYokYPLQ0/gLI7QY4ea/hjKXLiYjMsZgTxjdUhnU2XchcBVV0tDppDCVjB/S4Q
v0oT45XDqj48N4VbQJYu+Us9GOhklkYgtQw4onsKDk/yhTu//tlmoy1vCkywulc4Zfn6X0dVbNyb
8xUTV3vbe6/mR7S8isFdkQvQVdBJbqRV6Wi5wtemw3gT5NkJnXqeeCgfHxRVWTfev//9AR75ARV9
ncoq7wQjTx4bCVYRg+nSBZ242LAzSVrfUHrgr6cfz4e+tB3Bqaua1pAZ9+ewC0LgzEx2BrByTlhN
bPVUQphM6i/3fWs7E2wz8oVM+v5YzwlIh5KB94mKgL6DYdZwt/T3XCuKug58yROFBVg8CXtfL6+0
SSqJGzaO0Xiv0qCFhSBHvy8MavLbWyqk0XtXqaR9MDnPXIxJU91UBvxvZsFYMwbjqkIKn5G04sIz
re5GE2/94O14Y7YOpYFZpbuw0OCWItTWH/MnWqbuXSXhhnRvuRLth6cJ71eVf5+OELwc5xQ7mjRB
iqQkJ5Qn5DCz9cWK0gp5813O1iQbaMfL1wvSC3+JiEuFZYUWb3UAdQ2wZFUPfUXE1RSAqUiONg6e
Sf0YYrTEvPMr3uz5E6p+gxLVeqvIduoe5Vj0ZsxWtXfJSFGpGQcYLyN4UtQiqsDdoxE0qWrj+y13
NcKNnCJnT8SKYwUmN//m6Ogpxf+ZuBuT3YwlNjzFuCJ908k+0O0p+akKueIHg10dPiCtdbi2o3Mi
u1woAWNA0JOqo8Fsq1EsNc5PBd4oO77gf2asYJ0AMYU8x7IZppgHFqVyFi4AYWn5CXnvVIrAWm5B
1wtIzcOmVt3du0nYIgRrIRzJSIObvPrUTzEROXtiXg1vruNNIGR39q7mt5BwJEHhmCGPIfTPmQ/c
T3YEY8x6/aBjKbCZgWTBkdWFGZEhylVvkTTwEFjQThN0OThC1tKGhtVKCQRxRIAJ6XiP4HQ5zrVl
ZWpMZrMZuUXafP0d+kTjz1DS9VZtIG3TcMMOOs4+1PMBb7LvJvfNc+J9EVok4/TAbGi0evV+zhgB
9/l56F+VbIlkC+Ee+BkWsk/DLWOF0CxGYFh7AI5bxvBxrxUzmCh89ouAQaj5PtAgEJE7WXNWSFo0
CROPIPK32hhsLkhjXAiItZrHxP+rj7c/IqkjHatLU8Bp9M9sCciBgPjjVVqmBvTVScZQNeihNAos
V23wr1FdOKV8SStibnldSFgHOZWNz7Tk9YDtknpao4GonLfWuxAMJcGEbJ8htUX6RsbW9Wg+wXFW
qmywgSixDe6P4Y2uzUVDqe0fVbRGbFMU5Atz/CtIFmRB4dAw9UP0Y3S+wv1wuaqLtJciem+A2sf0
bccbiA8ihjKFfnSKppky0tkQCaKG71dlGkXOIYq8osFO16OW4aMioJGbNm/r+Jjzrdypy7l39enB
8JUmzBqUijkycogYA87zmL+b6OkhXUtT0Eu3ZIUcuv3jd8jMjuI9m53pAVdWkMLIj/oPQBdF7CjZ
qYChex988IzmwCJeAiSJ1KOB3OA+xhlf09ACuV877J6fCE/GCLlcHTSbkgTWupg0fuQYG6luQIUT
UTbwsRgMQuyfmc1Sga40UxTR47vIR2njQUv3/1Sy2nRKDq0WqD7AW62Wo1yJxLR+85z+wOcMWRbK
NVLLlZ64SU+DeJigYeG4h2JZOTzeZPhViC0sc2WYi0NZVzUyb1bgqHjpvU9relTabY0U29DrhLJM
izHDXPypfdczagrRb0gR4iBRLFqthSzF90uoccCOzRFtA2fSSt6OMm31Jsh8eO1qpiR5WK/Dr/Ey
KjZLwt+2UU0/aFR383khUQbKxVO1R/7w/z/V2M0HX6oxyo5VdpZ/v045Ih1a0mTvGj3P0HfaYxd9
ymWJEGeGjxBmkiaEYzeTHgRqoAQOd0Xavz3O220pKqpMwc/oc6DEgioWoV5k1UDiuiefXz3Y8QIF
bxSIurpnJI20RgCbnqhEAnQj096KltSlXivNjuULhwIgpPo6lLTe3blDgzys0B1uuqrRkx00Ehe3
DrjNf/Z+wvxQPCp19Db6tNNDOSIJALnSi7dQAHblvOJjwa9TtOVXvTn2/qKhZKp2FmPCIOoRm16r
0Y6czIGAtMoYZ7XUkxHb706o2eIOxNs+sO8kQJqF9DrVnhYdLYlowqKPn/wYWELnsv8LpwbjKmbY
HDTEI34dRa7M/WhMB91EXH3hMdKLklBp/ox8vnVpA3ldLV+MtSZFEn9W3MJFcJhdI2pTI2PCkWy8
CHfQe/VBdxkU0g6iByGjc8EpCERDVlKb6/UKqD+fLocP3A9aqMi2J28bv731m9FjzIfYJKOW6Tat
2Vd6qDhFZ6QXUqyXZJn72Eh/EabuNEhRfMgeEv5zbaCQrsSoh/ZCq1fSPG37z1VASlrNJ9peOUI0
cFafjh1mVVYiiYeY+JJp4UyWS5JsmWTCFUQl/9OAnGEntJKOYO0rCFIQcP6Emy914muock8RDD87
JXNhm9D6F89qECXEI9xjEQAxGCJKmUMThSZmU01ytgTD5WodMVCRhkJ++Zo606nd1HX31n96mKe1
6eH7EWSYlVzMUrWe5yFI2F8AponcX3kjrZnOH4dZo0i9xWqBitOhrrEdKRHhLEAed+2kXwnuSp1t
iy0bjM7FEl9QLY7lNDEUZ+roX8z0G1gafnOiGG0Uj8lMKTQv1Dktww6TMGoCbDmRcqMymkTj0ex9
CAKk3+/mXz8iD9cLbfIOBKo//sLNGXZqg/buEReu9FyUhIBxwqVeMEtN571fzuKGHbq61slSCTFT
Q8xWj0oYWJbvlWt9nVIIZrNwmZfVRb+BThNn4diDY5YS8AnnvKDgFkyDadB6DZta1lnm7sIhRJcY
wLvKAXH/z/d/eN72mEw0Z4DOMer4x+6fmo80NlB60ff0c2kp8lg8pqkvbbPuvS7INdTSOHmbZnhq
kM88gW/icf55ISRWmaL/Ti/fHJLlgYph+lAgg7mQvVobX33pHX1VJbwkblx5oqENinnaB8xNTNrO
uiFxQ3Td/tHfc6ez8oBIHciAh/3rgIpgG4ZrgRtXDbR7DRcrbVuj7ZRGA6iqQn/QB3fP45/+5HDn
lRY+s+ZdcpXMB4QfdCSDA0vbs5YFdgFCl3TfSlpRLaC36LyJ3/3uu6QM1g7z5IPPtxl51cHEMYt3
LjR3meS3BnxlK2cZKP/L9sitwvkZZnVPto1llwIa8+qNcfWGg++FszBeKeoLMnQmt8lzQTCB+0ue
7U/HwB4lhzZ1aK0m989Ujzaex1dvRlwIMfHAdwJPcNp+O/oedU21kU7V1t37groaiqV/COncEsqN
Hldb/ZEGCgCXox34BmHG2bbEzXO9KmEkuSkmEPSXje3xQw3XkvrWAz2bkkwmlemIzh1vYiveK6NI
FgWZ/I/lJocuMJdeaUtoO6ekJA/yY5CFPnmg9f0pCUqNhCMAfEsE8Sxd/ue8A7gu6XkT8GmAJ/RQ
Dtw1W2i2dIPAWJ4ivLBymdVuSYp3+GOrOBWw1hy7f2icQlLw42nv27BZqQhK4jRwJoGiB4Xewo2j
P+ZiBGDMQ2SkgIDdY4lazNaDKu6lfzX4C+lTWfD0fMm3OvvdLhIwe3nZ2pnL9LgIaltAPBJNVkW0
tbnyD7VzaxG7QEJXMreoR2j4h03Ig8dy+kiI5PLJ5ira+04fV1qNdlYKMRE5n7ACOY8jySdFg3K5
BVJmKNfRMXUfyJuDtotAQXK3/CxwS90w57N/jyEbzZKx3bOB2SSt+XgHIsTJgu3RzpkclwK2yiBc
bVd4zo5w7qR61F4mNY2rDsnHbZ5Av0zUaKi2tiRozC5Tp11Pi/m1JOHzcrBes2NYzgHhflijlQ3D
YEjNgSOHKgJocuSNXH7OE4gSHg81CcFwrmc7NcmAC6DZLWMufqF2iHsKbAGg9owPX+2F8R9kl5Eu
EZDVT1v1HsXrXMUUjlUpOpge5aIRGQOipe6PldGXjkeBqyy34rpTk2NtCxH3EVwnnTcAUSLhjoAw
43fzV3aCScnNdlMt2tRyawsazm25ER4AkvvUfimNLm6Q68mDm+tFtaZ1irz00TxMhYjRYaE13z3B
hQIRAlSlW++kkdbe5JtMtpayoX4xs++iQVYzdpRFXLCbFhdXvNsvrayqJOnE6xZrVSuiRdAoGNgg
UZ1RmktYG8+bwYlOl3q2kj+o4j0i+2gD8rJlHL5Fy9EHFNtfgL5GbqecZ0px0DDxuGxqK4WeY1iJ
hAXqxFXuKni8rW9nEyA52ll5a/reivjeWthd5zCAMFmmbAn3tE81ADhlk9zg+Ho+S8YqJPfdmHx4
+BskEhMYitC8QZWaR+/c6NXQHguLcwwDKPd7JceHphNBuwJFYJR/+shck7kJhq9nI2rqSt1ybTSa
AHj4PmRkItH+uj96heIbWU4RSi5FSOExnzoXnFzQMP6QoY1HDVDhheE8XBp/2CPFRAK2IkYm9X+2
j7b9XHH1s/7G2Ca4zy+fv5jiHH+ie1Vyi3x7aPrzKyFkHFBNp/GIYQcT/TJXvF8SaCsRWwX5jTvJ
tqhWYyM6uBNctP/fdP2RGjLvEhOHMxJ84VNdRymtEF0U+NFycQ1lalb5PHgKma6uTjQh/cFBAcIq
P6t2hBo4SqoG0J5AYPf8PX6gmsiI0Ys6jsq/Ch5K+0VylcQG43LnZH/JauocnbJP+TkZVGt9kez0
012WNEJLf4IBWXb2mYJpli4kjuBCo6qBKJFai5tvuW56Nc/e6jSS48Mz04lmgIOQCmW4jAUf/aUO
mkzB1VZ6v0D+ET5wM7fAjoABtf7LpBAIb3+M9cZnl+FaVMlMipcKmtZrXoM9z6nalSynNVK/rUyb
n+zt7IaVvCKGJoCU05g/tR7i32PwDnKu0t1ebFd/xPodyzK5x+r+kou2UYemIAA42wHItCaKPi2b
qWSabnB0PqLsd+DgBeYvGT1p8qMpvDfA2xc3A6kUyoZqQjAyULgmAIN68NqDxXq9moxkZ3T6fbg8
4hT/iJa/H72L4jw03kLcl+XiqWeJfB/8OPybpwonerEFG1GXIrHVNTMlE568dQ2YPD/KBFqZA0al
+/Z/uNRfs1tjZG7btG9jsdaybKUO6Fh2ZOuxY07rIsCdZGZ3rye3UFbYsIrhp6+zNPLxvy9fGmbg
KAaLbayzoDtZitRGpX7R6HwiRb9IBgHMLBqVwwaZ4wcM4ffRVSl8aqUHV3rDPPR25mPKbBiAASQg
kZL0j4xb9QVzvhle00DCCIz1AWp/NMYBITMp69KeQ8zStS1lITUJGK1Ho/ZzKXh5v+DPzJVm1gWa
gqPP0Y97WpdnEszUO5orChdtKKShBwGIEcVOGdWIwnHKCfuTnSQlqynhedNsTzA1rP1yQ66nURJu
YD35QTAEK6xU3trKvUdpol410Uwwve/ykjks8YprB/ofMFqPOGdl5NLdd8KynXYDjxu9vk20gQpg
+3KmzAPaEZZSuqgLZyfTiwkG2XTHR26Y1v1MY/mhbeJKSFIPXlvFTSnAwCCI/rrh8jVHQTKBJcCg
dBjiJET7FKJVW8Io/xns28EewN8BKYKqO2wPDV7FmMlwvjLm0UEMR673VWH7Dkxeu7Y4CPtP/1Ww
oHByiU2iC8gpYHGzvlVNGGFNWj8gup5L8R4o087ppguvx6Ki6WOfsEeKwXDCTJV2LvrAidd/k6jV
XygBsg0WpVzVnBeXJ3dlFrmZQp22Zfs6A+VZDid8iP70U/OwqV3SzLtqQDLRGQfpqyq3BGIlQfLB
eSMjuXIJAW6Z0Z04kjozWIvTH818+pQfvEao+xKfGLW/GN+BaqpvsVWpDNsaQrmQ11UZ7Y2skNMH
HQaNk6sdQDBySBL9Wzi3uAkhBvdri11JUbcHwe6ioB5SqAFzzeXaBC9ud6Ni35J4ZeDcwhme4YME
Tnah8qPTCzdgwsriq3zZw+4r7gFDOq+guLS24k6ZX15KXEmPcBjs79whDZijhb6c0bU+p+Tylod7
LimrJ2LA41yxw9zULwVzbHXy1HmVChYgOGPVPlNs+W+e9Y6ci9nP9biXS7xfEQGsfjDzcRaz+wJk
EkPbvPxYy0ypw1XcxNLmgfgEGusk4Oztza3DQclG0etSOpKCwgm5Y/MznU9hnMNRRak+EsvaH4z4
mW8UnFkiX9NsItp8Eb1HX5E0ZrpwHq15tSoopAGMeFN5CA62zpPMebrJFUBXvRzPINdKowEWknax
E27265heYuoBJPwCOezIoCeWDgzwCnGW/FPg0xUhZSBnqjZDhkLg70TBWPYfaqCoDznCysyefWoC
Yj0blY9ZtZ5Qen4OJRgV31CLnnt5GvpCAF1VnjgMxv1nbI4f4sjrd9znBWYu6+JQ4RPR43PVum31
uJ7q96qpVjh/m/Yql93pHabD0p6C8iAU+gSACkR/fqumANmja9mvkXPorHvRBeqyDgongOVcpC3s
9+LyiFkNoG3wq5+5RfaKlgZAfw+/8ZAHvYyjwjp+xEZ4JfwUN6kk5/4Re2FQW/8GDr2cOUa45de8
bmzeLF2/TPP76YmyAsp2fec52LGKxk73Hu53TFrZTEvA83V0NpM3V3gGMgkHeSFbU5ekgxiO1aaR
ArSJTHA+ryAbzf9WxdYXyadQcrQQkOvE/5eReGz5NQgmILmVAuSCltk0nU5wzuuR16gX14sWbayW
hftOND0ZqQmOLPR2lZgbSrBgp6McgFG2t+zyFyyzx8UM5Dq9/pNLSNXZVmPlwJVGnhia5Yrv2W4O
jNFDwPv0zn1CqlRuFA8kox7JDPm11217Ny9emgJxz/Pxe7ZlxXUx6KnFSzY9YPMOb+BgVp6dPTXm
TEkJQWFORjCmlTg1w3wjOFJr19hM4Tf6wZGM0MjVaZJnLadxVwZYceFAcjrV/zkHG0ZDsuCoY1iZ
PIiES4UwvQS+qKg/OFe3d0707Cy4qNVHTMXivL5tojg6fy87BQCU+d7QPyvrQ2XNGCZtmBBFXfDN
qxZLKR7VH96hOFPlmZjVRcebrG3IQeifBLOOoiHeiMAUGXbR3UlJYOydbejialM4IG++QIT97LHv
WSxqCLJ8GmHlqWxqi8mA31myx/45eu3v4/KcY27h3+blnN6zxV/0/ZYdGCJ6uCo3bEy8w9sZi8t0
SIns0oM6fZBMKAPCJl1Tlzld1r9z1Nn5Zghl7omEgl6/pmpB15fF4Rj08uxEryXJXK4ZUwIaBXoi
TN6gaq3C0QjLTOqzhx5FLo/XLzn32EgATLBF7FUTc+as4t9Im9GMVG7NrF3vRlm0gc2jx2IIx0k8
iGU7FYB7JC6PIKiVaXQU6qbXyaRTRcHWzTLvHm6hISdnGeDwLO1wKAC9n9WbHLx3R1Ar1qwRUus6
qKhq1NVdY34Yrg12cTiFvQg9hu/nWEy4HjoBM4M9rTfrp4yrgrDlfJ811Gqa4WAspWUgIYpXxWn9
j/ISeN4vZQ5J7VcObgdvSyQMo8WCUp10u3ZQWn2wrA9CSNxZBsFPr/3vap8yIQ31mtt6GQVS5uhl
L/g954H3Xf63Wck/+ca+fqYpEVnsO6KqWb4FnS7H99PrIOFWXFt2hzTZHhc5BLAfBWhU5izviBNY
iKJi4P1i2Cmy7pRz01ESNVeE8Zp8KEjt8h5iW7BRJvFphPrtUi9YYN47EOsZXpyTIO22ZMiWd8Li
A0YJ/bPZ6donsjTJ2ohUWjEqCaT8u7edqizmEBTgMQC6Sf+waEtuWnbVZV2VMC4dWzUzfMG3j3iQ
ytEGC7dvLY1lgnnHKV9wsiimYFeWJb30P98JBntDyHFQxJTmOLil+w+aedTWtfmXd41+zb33AM9t
hBEHjw1M9RRFw1ZU3PT0xLlg/6pfW9FIN0Jgds6y0DqasSFB3maVZGSKDkf3skXOZFmzHb27hskx
nHo3SHpsTHAsmnh6pxl6hnAQJOpKcP2YwDk1Zh3b8+hF/qwm1Ed83XZAEBoIQFu5OyOViv2bRMn/
3/YiS5IwvIIWgRhfrBN3cfxUaCpA6gARYGJVG3uISZm//VB0JDGvHp1qctyCWIt4fxctEoLklq7p
RoAlNuuc9KUpd6kyWHy1g7oz1eLLOO9zsNVoGyET60/tKm8p+by5DW/mIiSpVmnw9Y9lsrDq049B
DTWFWdQnJnGRoQCW9fTudb799ZJQV2lKPkOpyzHt255jcYAYTUF3OWROT1hJQIkmjJK0WVFX7jmE
tZAXlS3/eyKT3bfLSC0UhkpM7iedHaGPRylhZZW3MFchnqY4wNLkbqWAXME5sAbFjEBeTySKZRQV
FJjBXBYpS3yY3/C6pO+T+aJJNTlCiEADaC6ygvYTiqUI9rbdczSdk/cgE1m2kLoNMxdevttrxTxu
lIzy1w0HUhs7o2qN8r9gGjlhhaleNqvPW1p2umAvsufBDcmeOaoFJ9hB+RC35Xgp92xUxy81FBJs
nVCnbore3obEyd8uFiRghjsCgP02VjRDv4DULDDxLbIhdYRPYY9iW38C0YubZnzCt80DoWAEXuCP
RJ3Z+gxOchOwFwcTmXj/dk3yjaF9AF2U09P2g0Oyir0ZXN2PRHes/uvL4SOC0m3cOGbjc1d1MfGX
w10D980TawFdDdsBs5txomcgonKI2JAU6u+IHSxtRfFo/JnVnAW+7jMY8F8fz29hgK6Z0kULbGET
bAU3JEyuWEUmVtH3qU0OnWQpfvXs56dEQayuiuICmOpQ2Cz9ll9DQhUWxvKCdnHSkpF0zHQwhOkY
4eb1Djuf+9CBHPRG2LLj9Mq+kDQcJlcFcUKD+fv6QipeCC1RA1pTaOdgDE/aOEgDZ4HoODSqgzuj
xw4fXZ1sF4nuQ6mxZGR/OdVwx/BbWNc8IadpGBKVMNLjfoYMYMVOcKZPf9wBrHB1So+CUE+VD+Px
YxESW2NufBmV1ydUcOyxDtB+/OoK7Q2qoQgTPLTgARv+hbVzbEYMipjBlsMqMVCblYqngbU5BZs/
9BBb4+070tOiLtSHGP/BS1ZhNm+A1DNdxcHf4UhIc7tdWt4YQ8ZBppFVDMGgVr3k0fe3IEtdaV6a
zwCbjYeE8swj13SlRoXgdg6jYAtJoV50KxXU/zord5HFqkGgC3uBLR6qSt855B2fyY+1ZiubL7tw
2MfewUTAHCwOgIDgaih/g7K+BLB2UgGU+hp6rUgvMoCltmZ38A6m3p7Koz+2NgFd3mH4+nPXye6B
diQv7+Lh05r+msHljFdL1uuvnRcogE3J233c5UezRU/TrEloX8oQz9a+NLh54R3P52Paeex7V7xE
Da2+KXfoidNkkodVO6s2h2BMVXJdsyqL4j4pKgXB7dqQbERJBcmzj2MW6Osexe3C9eUw0gRYv39Q
+cvBOF16JkNMpAnh36J1OBJmzxB+xJfV/pnMUPAplMxaTBzeshrLD96GoEt796gcRAjiPXWHxhWu
4AgZnQKdliOXexxxo2nKDsw3A/oKwSALcUD91L6jcwRyztF0wADVhsgDDt9eyke99CRvztEFdJr/
VScjLR0aY4P3obbN8BQVz1kpOOAqR7AkDnOqIeTuVYxk5TsHDQrKkk/DuDyMIXW3kJO+z3hZHjLN
fRlNPHdnBuwho6WBKNK3eYKj6t591I+ou/o6BQTI/9wAoxFfcUg7o87kMZHGb3mJ9NKCyDsebE24
uK3AIalA0Kcuzm9wKlfIutXqiYZrqwaFKYdaKdTNbvkg1MMEsLOmLh8iKqQGYNBQ3cM7ohyFEtR5
QRaqb2rjJfcWuhzSyH9rUQ2G44dLOvVzCTmi4r0QPBuypA4ycTy9k03Vv6D8b11OwOPi2icrjyA0
zMWnMyqj87bi+pVk4ZX9Cph1TVktbKHVmj3hNvL38rHjXCwZ1rkAoaJZSNn/kfjSm+wmI0a7FoPR
Gz1GIcgq7tNRBGbKKdqqVeAScX9YBbehZ07/1HZfsXz1SqHpW/a0KejiX6HfewzInjCVWWMF8R3V
TTc9wb17s/dYPAmMpfal4ii+cHp1aHATZgvnecNY7mg1DeiFThByCkw0Hf/YsQhOOu5MVFqq7fO2
MWIgHSAV1vjEpZ5Olm0jPpYpHpVnAApJJA0mMDdDyduJ54d71DskFKEm5QL6F8jJPQz8+k/xmAij
kd/y2l7W7h58DTk2N6s4Khzxuc4HvqPaeNit7RleuK3ctPS7KNq/YtMamUs0PRfw09t0ieH52qLl
CMoDhPJhVFhIOQ+XEE+8skaNvfxI0KHiCQlpaGupPiRz8DvEyrD7v6eneghsgfogufW04kMfMS2A
yl3Ptn1xTCvGd+MYDNxaoopOGAR7/qiFsfIwcc/zeF5iZ87iXMGABZ2xdDAWCWf0fmgLF4M1pXmX
WYX92FMBMKo0NzOx65Rmw9PdV+y/VNdN6CBhduP1ZJjskGWfLGwLBiUUBPkezxtYtezmzjFth28s
rg+gUgAiHsajVRWev7OuoLPLRzZkO9KqcyJ9mc/yzIvJjM4oJO7c6neJq/5+ZBSCGmr/lgv5iWkX
NTAqakiYwPCVcCl6xm5WBs2HlZCpBq7Ngt7nqNi0KDSX/RdHWwhhcAEi+s/2NJ00LSlB3OaijoLN
GeJz1DXMe5tiJ9+w+2FBFsGfcJLUCZW256Sf/MDFDlSTVCCddmt3HIzYYkpaKa3fm7E+dgOmLuHF
ED2eY4ytooAB0k7zuoCyECiaeTh+ahS+wP8GfYJMRr08Bx6KR8kD4mSNVrWXxjycUwUdOE6TpMwJ
YGb6rqlLjDKGXjBzqX8kQ/8knndaq+EwvxTpBlxF4S+LAbJxnVRgyLwkEE7kwC4exKH0cBUYRSU/
KLRUaxkl69WgrRi0yDXTUTb3zkUNCScXJFmofXC+3zgSXHl5rC0YBCAHnOJ1bSH0UoxMdKEUfSHB
lsFHR+Pe0jSlZhJqrxrts4HjS96QvRTcZ6Y3Lw8NefTD0s9xjfOCaJhtkQQLkM6Khx7gI6DNTwQg
RO7HSD0UuEmwe0GB4Y0YsApVekcCaxlHz/8SeF2YnJei8VuDju8APELgns2E9OsF0yiatITfy2HS
9z35Qqjn+aEGu6IuJW/g7J6KPuU2oFBMLsl4S5bA4Kd3WTFBektQCH78pDt8pO2TfCuL5wModxEV
BDWslmCvzQXwCJyp3n/rY0jGzKzpnO6pJIeEwhd//IfnB5uE+4VW+EK4rLkKBB9rmpdgeXml3BNt
dNuMSO/tX7FNE7NZ1K0PLwFwzzXjVf2P/iZTL7K1gSvjwUGrzSkM7QG5j2HatRfDDTYnxVQw7MaU
fXSV3+OOYyDMYr7onn7MaH4F7iKjsCG0a8NLHC+1BKGsKJv8lROxIwj00NtPsjf+oc78cizSVjFY
yKmsw52iRQ7k4NV6vFygDaQn37r9Pxvb2y4Of5Q59eF+XackJ6K0CZ1fVZy7tTCCCbwTQpSRGxYd
xxzW10zK4mQLem4frVO+pU/gj/kD9yje0OfLJk01sL3rwQVPCEo4RCpfjUp4t+/c1G+izUUfDTny
ATL5xQKrLywCrGaoo5LJqfHrFVwW1Uum9oMPCwYaXNI7dD28x0lvM6C6YNcUVzX6sczxzCK2hV3b
OMCkE6e1rlKgAwMONqZtpTeA+4uK2vMp/yg85HrDgKuDECXjb46Ni++UoEN4MLZ/YGwOeyyVllW2
kYH7519vW5nvCJ+E/0ated/N/KYHNhSHplPmVgO6eLwQ3v/lR9NcA+jOl3meYTVVlPb05op/jz5u
76UMQ/YolHeI2AhDf7CrC9klPIwwNBC0gDEd2ATOhCvsn2gxyGtm+1tS+60aN+FsYiEFDm8DaAEF
DnrQomt/tkv5jg1j3NQ323mYK5i37vS0xz2XrJ0q5DEsCC4UfSPTbKE/dpun061kN54XRry749Yz
PPYSiD3fxBkGDewqBLX4Q3FrC5uT0tYpylvUEi+2KI+zwdMoKq8lLptpcbGDFo3wHfZ0X95LaC+O
NW7B9HHpia1K+GOlekH3uxcmWunVmV6nooxkVTnrdIdEduv0cGxuts9cbCN/xXw8+ZK/bbGuX2ho
+Tu0UxG0n7cFp8PISQlZtAFqUl87DvSf2dihu9fJT+uat930qGT53BLIjsiMhvrud3DE+MR0F8AB
6qmcDXE+427iJiq3UNZC04hCoQGKpyGczp17J/VrMjmQQMgXPPPk+49I9azAB0hlhSXciniT20Vm
+sQxpqjyTOnMAantBd5Jh0BKHgHKoABzGxphI/D+enG+kL6ua0zEhVM253+0KSeP+aESQwSQ0lj5
qJuGMXkRasQAadG6SNxIG6ZObHZVP2mh1Tqnr/Ial4rfjuir/KRWox6MBCx9IXs188vYErtTSgfl
J3anTU1Mua9jjgG2djx9CCuzOdfSR5u2cQdtjYqxbAVFCF+WCjSzPxjcWoov5Gq/IfBvMv0rcTTe
HALRqyXQJ8zGK/D9YbXENsbX5uy1GLsfmrlhiqamFIF/klo4yj6SfJEsnDqm6DZXeFSz9jiHWXFG
JNn6uEJWnpA4Xnji8rJ3aqgCgbLcAw+FZdXDQnFT79jWdTcWcg8g0NqImJTJqFMYtpGUAcGKMYIt
YYismlc9UfK+cxYWOVwYZAwKNZR7DtUtcYbaCamfnhRgQ9Z+/wvN+/5POSUPIfA2xNeeEns7a2m3
25ur/jrSswLKgknEgjVoWxM4DGT0hqLgbkxtb9o3Ol2WPvx+sB4P3DumxZPy0SGuUX1UdKNCYEc3
Cuc/AokuIw6LDmFQ0b26MBwFwGTu04ov9cX/BFOZ9NDsunWaSoB/+97lfyOLBcOiA83Wy4QpHlWk
kdEz4msfOEOjiR2qdkf5nvWjkg4qusA9YLz1vdGe5swc4/DD0mACTJszVPkII7GvEt9FNxFfeMCO
Bug0CJtnfmVjBpSwY9qQ3t3rapXapzFSU9HXrZZc07msHgWlX9iv5iwQTrBR6lMKQex5yLvDQj8m
JVWkjatG7KVfB4Fmx6BY+kq2LWhJtZXUqpNhdSNibH/84+YdsF4S61bgYgdXUyFUQAAakpcsCBqo
2joZ5MLE4KrebZ3dj7WdJsgmMwHdAC3xfoN7DXGUBRUugJ3oLQrOghKyD34PIZJ3ZO0fMnhfhjoY
NvXm/onMhM/WHAiD5O47l75qHU6pPmA3R86U3UB4oLNq8iOTQ2vCSZqmOZJ+VJRUI2V+zJ02bt7o
nTjh94040oSsBDi1naE0kRm7U8OaQ3GaMaEko5/nBCCpdCjM2l2epWoSmv3xyiSG0A/suo8pGZXU
ENmCou4d+vrIysn9ypvzLpfeAIzmlW9FFVmrzlXtkaZ01kRkMjhD1VQSVugr6ElET4596H4Xahsv
MLVKazCcrhBX5mwR/crQYsa2vMoFgtyka8Jm6PBvKTJAyBG7yt+pA80nL7+77O9BA7NXK7F0wHnv
Ri0Bf30RXARh1It8YrK/n3D0+BguSH3uAtlDMD1XpBr0ME+YxzL0IS7v9xI1b/OusJkJJdBrBT8o
0zkbo+PmFO9hRPtlQDdDfw5YD+0nv5jG61RgQzakEWz80bEolo1HzStojvfz3lcUdvcyj9E/Hyjb
KzAt9PK+CTkn5278evgfaHJtGb7KERVHAKePdsdkhHoWE9bUYbIirHz7NgBBb89AAwoFnp1R0/Pq
DXIS2uI54MTPNzRcnPlvsRkxd8kMyX9UeHfLYT62QUrnwoEgrZCtZs7AzqFCr/JvzhHK9gPAHhtt
jFHNWIvRzc1wtr+OM6IdV13ny5oQ+odKjfLGk0WSmYvd0fAWV6ySHoFsks+l+GIqb68cNuwnlhQk
Win6CC5pFyn9y2rMEJFYlktWb6YfR0CbOOcGvG9J07Yte0T/CUWmyLsF4xvIV0Vn6Gp0RllP0Eiz
sK10ks9t+1+MZQEY39sQ6bT65B1ZshqUUaJ8AZ9xFYNbA/+483uxA4CSfLDgHo36x+IiryKSgKqX
ow8yqGer08FKOgUOx12E/gL+vn4oUui/a0wX2kgQ+OVlHNiQ8pqgOhe3g2mjM+369tsIwiHvfiDh
w0OBkNQGSmbpdTmd/tlGiFgt5/G//c2E7R6ewCVzStsZ7EMehxT1ENvUBwnHDlSyQpeja/pyAkW8
zqLXs3TuHxV1PLm24vdmRZsEJvPUryFMOzdSkaox48T9Bsx2dVtdmEHLus343wcTdb0db3SSBmc6
6Zc7XVUBm75s5DmAvz0RCyGz1fZ3+BviY1S/TG1ky4jc4l59+YEeph6GsPfzwyr6sDFTVLlGesd6
2qgtEiRZJTu6dcPRlsZjvyWPxJ32Rg8uUipou6TCvxjogM3kJJefcRQeiNQ1YvPjgAQz7zjXyRya
srfXxX+ZfRPOc1IuBqX725PFi3itbAkp6usqIIBJOcaUnTWp9lKTZPWdGQfWqi5Zk+d7yBxMGXGP
98nYwecUQW1KfRZE2vu5ATd2TYDVez+hM3VTaEp+FTLy/GibOcjbtx64PMF1OlXhurNHsvrMBxDi
g2q5rOnbBXNJIHx0ykaIY+9R3ELur+GLZa3K1BozE6/cEhR70s2eLk0EzR9YC3xC6GggFXAHvQkQ
pyfsIvuf+z2FWml9nkOVVDhDTG0VijTtM7VX/j/8fosix/KQhRSFTHoM1GPtY8EjL+Bch4/ky5kb
Da3qQ1amejnb80l9qA7LFquEXWdKlN4VLTTRiyhGEl9gVSsFLCVMyi495xQNmLS3p0lZ3uowcFO9
Se5SNgz2dSZK9wFN9PHtA7FUd684LS7sagYt3r7eZx1MLblgmeU4V5KTdyLdM+3wA2pyLsHRZpOk
uMtkgOcCVwi3UZhvY30X5n9OE15yaPnw7zzxx08gCZRm8KhP83s0n+ipPlBWgqN0kvb1DhAr379e
FNItVrIgk9+dJw43toWUTtJ2RnFkolRHTUT9TTZg2goSyKvYsD19xIjKqVIWZcmG8rS1/BFqqk/I
Ru/jD7ck3uztWV8i5VGBHkNADLmntNJYQZdY4TpHTf6vhnGJnvvZZo1+T0NqVJcwOLjz+AnuFwIc
evJT8hilAGZSTjz/GpX9Zcw4Q0SHV0hC5WBWUgw5Ud5xWxEVozYcYnB1vbFmNC2qPJreRajctG59
/irNQQFxpP6bRuQjYL0xywuwK9yAUKmN6GwTU5STMQmMzMgcMojn/a5ZiHTDlhffLXyqaqbnjnms
VrhomKlk6QSNPkadY9l9sSucNypZx/Ftr8jjmdrxmDCtiAm6n10Bt2KwkgKmDDMnSRtb8F46S70j
AgkB98je0vm2zOp3oL5hJgFxQer9fIgcYyhigRoX8lctu3hvyTpSIstahMChdPwkzr/GwZxCu0vO
JXMorPXGs4o0imkxWi+mKBcDzg45XOihGm4ga/UzYkFdYAxLlT1uoFEVd0MQ62aKGIRfgCVKLhof
VCkYd2vVRfd2crFY8IOmDJmbH39YGiVCaXdyFOUBedFPha8bZbk6kwi5Vnof0KTqOwRIliHe/4sz
wTiykszuIhvuBk88lGgCXJM7sJyT90POpSNIIeZPxb6W3RFpFvyHcGfvbwIPA/41Y/GqIHgs+6Mm
WnzPiPme72MkRIY8uBjdNNkgRRjVcNd7k6LSyDWwem/KwpSv+9GaANi0SV+Nc4fQRNK835tI2pwO
be8KU1o8cBHfriawap1EGBTZIgs3XQmoPv458jHVXD0YOTLs8Nf5GOywl2NL4nlHOO+8GK9DsUPq
lo9hdNRagFZlL/R8tzlEWS8kwAy19rSxCzvP49mYNVvcoGYZwxf4yA4FI9UkA1YLcn8GgCvqNCFn
r7LpE905AU4CBKp2A3jfFbc+R+IQQNpqTTa6HsHFOM7+sbIV+iupKAdJ4iWfAeOX6M3+N5q7X41V
1tvcvye4Rbrx3xf2f4R+0dBKg97/GOT61vMtLj1p0oJt9bHOiJkk39GaYy+QzUvBx3p78p/hFYQQ
+6ApVY5O7GEKFGP6dB47NVm+berWGCUCYkpF3X0YfJqcwmWtJLk2aSV4727E0QDinAxZ8yQ+NDw0
1q8X1S/BgbD+choaX/1uqPSejD/hEu4l4Er60rPdUqNcHtXDb7l0Rdu+ofDV16XFbWI8JbsO4GJ8
Smh9/FKNEejZuQQPG4H/Wv8wARwGdp6euAUzHhTCDIYCJCyh5itnbed7l70wXkXkV36q+cToZktE
NwYy/gzYt9siEYjV5/WEEJYi/hBJpzgkfOh/Kyn4cHTBcdFm/we0+gFfYSy7yYsTlowrsG51Q678
abSnCEYcAz41S3eI5KBwf8H4Kfof4EHwYJelowy3B+VS+yRWOH3DoCuzvIwYvmQ6V5Pery5Y4Dn2
Cebqb2fallto2bbXfIljwbm/ZFlGa5REmEnJicW+Fa0Lb5fjdcPK5GiU8ayqHie20lXHp7p9hC21
D56ipGyUHkwbwUeqzRS6uft3P/rHXz4UUF+PTvwNcqYCU6LQIcA+PZ+JA1C7ko3MNrwqLO4LKmoT
gPr3Mla6C4ZoImYxCt1rUmkgWDpCvA9eM4Hz4lmh8eDGNHVm/Xd4XhAvw3611Cv6T3xkebWeK07G
Ln8lH4MO8Mkwb+z13kAzXDIVbexsnQCVgrzPJw6B7EuYeNGXVJbhUPSrwDbs7Jm3x+Vndh+iqZs3
lrt7QRSgzytASZ/aMLBhWYhvKrhncipUc7BfDEaoEe8hH96KpjktMqxm8hXxVzxZ9R0gqIPMEgmu
cxmfI0aMaW8EqJ6SnAT+PQTo/RchBRi5ehVUYLs5ZMKSG9wng0s3AZxX2IVADfvKwqjD0eTVlCL4
bsxwmUQi4GV3JgX8/m5UXHGiTlyvT/2twdXy1787U26DU/7hm6CTwOLO/r3a8PFwu6orC23P8I6W
wNHv+TywCW5KJDsQDSqDTzunv0TfOKmwnuVnKxUQKXcl4OwhAMYZEcYx0TrmphjuVk7RO+mbpafX
+/LThvx//5gOXJsfIGHq7B9dDJZtLS8I1rvU1koBGNl3c8w21RxJ3wb/x6fbRMscCbd5cPGcvB/O
RJz59b8KNDdBKSHX4Mm4MNvr/SljqrPTI8JgxaZbiWXi3wul3G9k24MbqkzZnmASAZ8R6lppoleM
zc7mNVUCFhHAssXeudxerBdkmrze/lmWS1GTQylcrbxaV0RxNuXzkGWOlvnPtfrJuq6V3ISfOfBe
bSPdlIds4/J96xaab/95bcI5nBZmj61Z2VeecOZ1Iqc2BL9gx/67/BlvYGUVtemdRYxd2XRYXyYG
8pXlin3YKQbismaN1CfCABjSj/7Bx3vr76h3vntD/cbC4/NBQ1dulV+AdDC3AOm7cuRRsRPGPSjq
eh1Bm4UV76vF5Ho1peWCNgw1Z3mynBhyp1LHoWX+d1D/PJfwfxl+BSwiY//YR+D2pWxBzjHOXwsU
c2UIdAUDqJqLeqXYFDYnb8eilFSM/v0vh2eFCkmoXHyDiOpWa3kIFhGvsHiM5umqYgHEnQIMlvUj
HGm6CwpF6TAlhl6sH5MdKvXzYj7Tz3x0WsrT+z725Y2GM7gzvDzyNZkezJMbCoD4nwpX5vehEgno
n7NBc1f2mEJYjmfbV+3rbBEeTHZnEkMJXgwtaHT7WWfmRH/DH7DRKVDMpi10mJHQjClHw1dVVc6w
EzMQ+VjGjQJIa25NgpG5N/9FzobUT+oRgI/Wo3HDTItfJZYlLy9t5W/rIyukb4M69ZuNoSJA+BtU
Fd3OyQQR7Ofezj2FSAT+LSnEfl0JYInuKo2leI8zV8ERI5rwMkuJyEvz/wzdCooBZ+ROVVTjCIqT
MwTbtShW/E9NUxZrC/KMAeOBNuaYnIkshh2P/bY8ABJTHZsnhR8ZIbpk0Me4XL5iJb7CCA4q6TEU
SIdytXcenK5kyTX/W/A93ULwD53463o6yZKXXaO5kQgx/rJ9ZVibbjpwDGCUFKQtPZHRKUkxtZl3
MYZj63ysowyqs+2TClspC6kTWacmmx4whJW6iSPl6qg0XYrFzIIhwpOejKXW8aS8CGzOqYW9rj8k
+7oM5KD1kCxoEd0OnIAc3xcKtLcC8i9BEiWU1Y95lhIsg+4Gk5hp0W2mpybtIuPbSvwEc/idd1Cq
Cux+kZMDpnHHKXJHlhx8XstVr7VQYe9bVxk1yf9pVrpj9Aokl67TYmdQif9vRXXngUBUxIhCBiRd
DXzuGbXrqov+0lbbOVGP6pfZh1AiPkb7EB2A+LVRgf1b84gES76Di04WQVPN788lHKU3qu3t4OKD
PWChTRKzQVw2BXLKD1dinhyPHnMrSV5O54q4QX903THnnBLqbGdJxJPKCNa0v5WNBiR/rnHcjooR
MQqkEHEtpxayl7EGPooaj9lNcFiL1f2PgL2mdU3ZbEia4PoAWAzzZ11c1lL6H+ovHb5U+kz39tIL
JtUzrmaHmNuoDnzVQVjqbKpvRzkAvI7ZRubimMLS3Swy1YxJZ0NQhwdVMjkQ3HEeEmdbQsQnkIPO
HRoFDOWxhfYxFL3O1DUn43xWXMQlhKjkMJn75jvU11mr1+0HLW8wGvvL0gyJp6+2zFvfiBhcf15W
eP3rCx3t7BURufk/tGWv607SQ802RIzBi2JS/lmFIfvpqq4HX1g9VflSpWUuXyqROWJQkWwm5KyM
Jer7v0uOwcqAq70NaRH7aYyF2N24eNWdfsNFZh5KKvuLvZMkQgquPRbrr+xz1fGmJkwSdHQwshRJ
xI1TGSCshJMz0+W/jTwEj0IHKKkDqt9cPoICa/KwuH0peyzk0D4x7fOG5DF3HbfczZVRYm85oGUq
1NwGgIBDi9ByEGgPwRzJgBsY3NFdoM8+RhJi7h6CdYFNhkk1Vip7bMW8tvrVfGuEPhcSZVMPl5oU
sipu58grx3EV5BOOwONE0oT9UMJ1Cpg4d464VkEnfjontKGhpid6pdqmkER40D9vgXkkGShSRaHD
YdxU6Vl+iPuTKcIOeVVea9teXHl7pGLFbNtYe3dq7SBc3uC5DRYX9Bs3VTUIWAnd+eguVMLON/sx
D/q1jdwrBMG7FH3DphC8qBpi+ES9Cc2oZULHD6vwcT+8anlgrj/sxO2eQq3zsxUJnxngRavuSMfE
ce9T7jcMSM03x9XUdhiQyi6ijnn55C+0Of0+2wSs7czfzRN7aRqYsRlEX7RL7Rj8rMDK9peC7Q3Z
6oPr8sZN5UMtAdIfMe39JkMyqEDBC2hPDBM2eRXPkhSDVPhA0WGv4GGJFpppZXET/90Qyb663ucN
x9bU8Xlm/sLohVJcJozXBDfnsj2GVNw2echReh41YWR7er19YT0tZffCoBEWByPASQO6NTamLF6j
u5EB8h+TQ/xfD8vYKcCTbZXCS0hzFVj3mK4ybXMlilmJ6hTbpPg9ly6Sj4maXxQTFpIxdna61Cci
tUmBEuhH6GeEI0z6QqukweALBuBQsu7K51JIQRBp6iOWtaYs3s7ZLX1x0tBQndca3n0smrTuVcbh
pBkHNuGuoB7SjlXZeQVfNc6SQQzba4/Eeeyp0ph6CGTGdaqUbBDWFcdoTC4d55XTIQeH+4t4qXgh
frriHo76iDKRXeuftS36gPTQ9Z/9pR8UAwkDtkVCRl13EAL51fXX6MvewJ60WeA32bOcmm3YQMTl
f7dLuYUdr6wO5RKnzmKowRi7IcqbtIT0u+vr/inGQm1Q0Ip3ERVAUZryxT0rLumxyOA2tnlLZwpV
WLwm1/oJ5dTEZBIkRX+zrKQDmsQEYPveo+PhEGrWtSwMmstjdz8unY6DP7JAgaK/azQqnpvtXqnG
7oM1FujXM0wNu9lwod8oXqdcvnbmGfENEBsKA7zLjqsR3tznxaY+uv2wfDtJIz7m1owztbNHF7eT
+nyJEABmNQl1QFGtagGwkoYJsNJY/4x7ifUwnQCZ26Qe2VFtGew/BtSeWWgTqL2S3KcbKbZnW/Mx
38H4FkUQPMFGtAN0Qo3P5BTY2N/MCpmNdF3h8t95tRxOXb4aIP0Ti2IXUAA64Z0J/YxOTqwWyTUV
919M9/NJ8a3TbZH5Dm8wIVry7whZ47k2mKQ1fcYdbIKoqPqyviiQi880r8svfxCIYmpphWB1Aq4C
L1s9jy4Q2TWfO/sDb+0VLGSaXeUQailSE2xyclM4o8zPua2t2Q3HR0ZJKb3azaBhdLXenItV1dRo
v8IbtRRo0sTZAxr1j3nXu9DSCN33QxpMtouLbrgdYAW53Bs0SF1qQ+0tMeu3kKUU7+lz0/NUePF6
L9j/Bie8/Y3+uppyxvfY+5yHHd1GAZmTL64n9H8PAmVttuym6Jqi3C8ZnRuHJ2K6sTSbc8/6hdHl
SU0fbmFes/VR5NArogiRXMJo5qaeEW71LDTRCoF/cMtjof0gRIyHVKKwkG43rf0ay35OtANHOeL9
DvG5QC5Vl3pWYluZEe5laUcRiv/p8ytBGFn6CvbK0GaD+4u/1OjafajLCIbP5w3Jwq+FyvBxoniB
f1CGXwYrVaeBbXfGqi/aIBvU/ad1rg6aV6JimL9o6UdqdcCGb5wrvU+PeTG2iKjkGuwYtyOZx2Zj
LQQAEP0DJSdbUWTM+OknAjBWqWaHRBOja4+65qzLkQRmvcvgBxCF+oZTUevsAfF/vvTC10W+ucAj
dnpxK/Z3V+Jxs0YwC/Zc+RAY2E3UH34ap4ka60z7IhWXcYi8To+8BPgkrhVvQ8G9RDLFd/9BoSfj
VbaCOw2F/4AEmMcRFLTxJ3TASoTbXXkmwsYHqTJfmoaoUnk1TKkeEMxS/uK1r+d494LeKYkuhqoR
ofkCtp6iArCIbE/N1MFTGl8D6TEhZWId6BU6rxDX7oPuOEEbRRZuX9eMRqv+zy5I0IY7wxkNnQhA
HWP0CXoIcx+Pm+kp9pVUjImMPjYwMXxJZbsqkne2K8DKe3irfXTTe0j4QVkuqFToaPaTTOgZkWFn
vCQy/MgDXnEss6M/EQx/aDlvRu9fqVjJ7xza2Vn241CTOJQ1nbbp02nYoxJs5eRn/tkpSzyisoEL
VL3rQv2i3ztu5TzOzrUpDfk17/JleUiiRlwv3y80pmCrRkIg/jgVNl0zfUEA1lIXD4TXmOs1z9re
dJN878AMfkH2Gzv6DyBD4OxpDtxhaiu73Q6OYKHpszxdBOmRrqMpYIpEBnOG9JqlUJUmhoZgOMut
Eyv53S3/8hAlGEoraEDis++GR/DfteXQrd7bCml448f+TK5Px8dMDx51bOBVIpo/0qeT5kmvMXTS
79r/FVaFnfmybwlohZPbJ+mw5QkUhQk2KkN6SqDZz/QRRmEZo4amzQhOyKcugUO/H/CjQsB+zn2M
N3H63Jdj/AxXHj4lcTfYNjb2QNXMAu7KPwsrd9DgvPQxSZPbO7XH1YvpnubQmpuZjMtBh0qBSRVG
sWcpsEFJ2EjbsmwNL2b1izb9bw3RQuB1ekWpQy0hxUpOlk3gzBUuz7u1E8YLhRnx8mFKopX4k+3y
CuVLZdWb2zlDTDQ2K+dAf7ZbKaE5gRSEKJj1vnJXTNxUQatNyavDr/Y4alk/Yd/O/qkas5l3aCbN
i0wds9edFpQ6cUSIoSponhbv+s2tum46yz8M4b8/QBiqE/Y3VA0eniEhmkppAhVVJ+7iGio8wPdJ
Mhva+GVkTgpA6eGu494fceQAirozjykf+lJwUnCCXhaU4+Xqzx9vt9fh937IPzNNbyDCqXbOgzfY
itvO6Y0UmiOxCUYr331uNYWZMdAc7FqzVyg5rVLjl/4BYE4o3zm+sCa1WpKp6xYBJ8B1Jw8jyZnS
Q7yiZuGWQVeFyhBZ+X+cKO89HseY0120JPzZ29kNxup2wUQG1G561szibdpRDAT82vyvifOyoz4j
UzDb8Krt+xVoozmm0q6JcbbRbJPWUgoAx9Blk6Tt1hEuH9WsjameE4tKkVr2ATkCxT+li39ML7lr
HewwkEVDTzhkn6DBeac/bDYk6N7xi+8ysHP1exEX93AFbYT+p2TrMT4nhzFyLNqN9OenaDXD7xPW
biQiNbr/2YMXv0WrcFngtxmamQg4CxQGljj2XD5Z60D0ZHIvDbLWOlEVhldmiq1mGob7TkHcUptX
MaEyei5iaSQsPY4Zgv3Y0/XB7uAifWsRkPXhrMyVebVHmKwo0bDqCMVdc2VP4F152FW8R0ndMkc3
iXicozURU6wv943KeZdK6lb4KavHbfcANWtUF8s827DX9t9uPicpxLElqplc6uFA7sHqMvtpwQRL
n3fMlKSP6WdgG1et0nLvLaCWOVsdXGSPx9U/rMoqUJgkVVcjZner8BFebubFP7wpSbEcy1dCtQ8K
/Vsb9EB+gDKJv8IUJ6OAdsAOa38Od9NUln617QFjIMRydprpqTkZLAJ49QweMZJSndL875bQFoC+
QJxH0k1wjl4r56RbPon5/9I5nkA5wA706/c4EPfVkYve1NCRf8L5nu4saS2cLlQkVJS5Pg2fg1LH
C2S4zh93Q3cepjZ3QaiPkUzu5fTimdg6tu17iWJoEFm2n8wQysOqzsezJSC1fyyXaGxWQgEllW/d
xrmQDRuarCmewrPFCeYPJbvlSQjSh9nk9lGSRgjFf6QaNrBiLP3+w21WYxcOR0rFIDrg/KNEa+Bu
eKn70bUW4tObE6pSxO/vJQ8dwK9tYSD6Dz7RoS4Lw8sVCp1zzTUADuAWJM0P1CZFOAX5YaVj7QXO
9D3pDc+zvNMtP4gaeWLKHqh9lOUtavERpiIHMLnJdqSf28KWpP5bTWd+Bm/aIuFbF/g6PNhyOl9Q
AxLK8yEPNFu6iALEQX7vKhJEOTjZwEnTJxqkNlscnCz/5OCPexwx5LETL9DN2miHEuF8S2k6iimx
P9Mc4y3qiD2t485Be9O5uyfUpTR38PKH9XOw6PGNIRYcXP/IKcNWi7OpNwm/nq5q1hPqBEaVXor/
6nrSqWoQPHjOSEHhq+JgSQckRVe5FOg4OmmBFk7cUhp8bH3fwR/Lu3Z3J+F+3I4esW3oy3mGScwq
D6/SI2Za5tQrqNLwUmIPgeC7NMXHuWbddfszhNsbmT6KravqySG/2Le8Sqzz0k6xT/NmrGHZx9BP
2cj1vVPHEwQXxs8V+eO2d2rl2m/PKcGyyUIuN0pQf8p89TgATrSotRg7hTQ5wwxIk2E6B96nZ1iB
9rGOAT/g3n9SLver7T6Z8QBAycH6Ovb/2Sc/KuL44c8P7lUC8RG4us4h7vhbcTDwR40pjWXI/ErP
EJxXpo8/cDEg7IPSQFQ4DyFNJEcOKtvMDOcH6Ujk5n+HIe5vNzOGrMgKPuB3vXYdOcjAZzu+Tw4p
X6KZ1I0t88sCFwq3JBRPVrKa5339MKuLmTYbZreE1x44Z0W0WAJM4NZuWqeTWmQot3nOikguJSxe
Nr7ub9wkzXNmY80VQVrEsCN0uSlzhziPng2QyQtAHS8qYRhG0fGIqreEa7RSuliSvwa0Dvy4rRZ5
33TClTaj3DBqxbVfwA/pM/Efz8LnKWRmE1Z3L0eAHYhhVIS67PxwuUtpkjoLEkEuBhqo51yl0zpg
xVIlEGiuIHzZsAOk7l+syXGc8X1QL6b8GIy2V9bH1zvp2lleot1L5ISaSeJ51SrRx3fTGlxjA44n
YqalBdXFfS5mRKxcuEYC/bDGZH/O+Lwn/kqQTDei4lAgoLjnH4EzwOY8IUFU5lUJTrSZlwt1u4am
KS1GRvuwXpnX/rlG10Lh4cmx+VF3IHWu4v+sC1LEkcYBQXd4mcqfE2My5ilOSR8EcB4I4DDqmWEZ
AIRiBX3TEOmBgfxPcBF99JboJpF9UHLZxLB3kfQY5DFBU3fxESzDvxXJOzHwnx19apgPwF9pMV3n
HBgl9s4hEPKIZkOSF7JMNZDWn1Vjw2LrgtiKZITbm9inABXRLgVCFj/UEq0ymPMd/FDqQe7EoN64
qJAeFddqARj8xp5QcsTOJoy/gNj491FfS9vCFOAbVQDUtTiOTxeTzVxgQtFIgS5xYUAiUr+zJKUl
ZQLWRcVY2/Km8/+gdmk8yIhSP2Zhd04ok+8wcCofGAgL+s+FIyqdcTmyJHRgjBBqjlSrySFSp2HW
9IIcCfLrxcigIuK26pN3MEoWswqFshrPGN7/BDHWLx/+YdCHTbBWD/tt8v2cYAbPmMOvZTYVb1aY
WsN5gXUoJELVU1Ywsx49a9fUGZoYGs/aec/dchN95UqDd98Y1SxLldhMTAfQjfAAjevo66WRcMC7
jpqDH6P2V7yuWuGcZnuy14Ndy6UMFTirivLmVfnvohJtuu8uUHj78SKcgwSPoifTBG+STA6sVL8f
v9osCK0IFa5g2I5xKOoQwFV0Yldg2K4eB5HwXVjN4d7TM82qzfl8AGpa+/y/B2VPkVbVBBlx7jZx
MXftSPuohdgX/XE5odaHA5/PMqtqXSqRgj7k1OgHx2HMxoFBJ1MJs0RA8kltwiNVBx4c8r8q2yv0
pw/xxTPimphDFqWnTEEyRZWlYwiFpuOGO4qnkRTtIsBWEPj98pe3N2O8yibkhuyspZw5pnpcVbi+
9fTffHqWjESAyTqjFFtdbO2c1bX08XVUGmzrdVeTQ+JjyXUyd6zzPmEho7Nw2Xxt16xbpRLW97Qt
JBtcUN+LjEckfiT8uCfoGC1i8kSDaNFxdp++7v4WUpeOvxlT0kmwsp1b9jEbP3S7hjkbyh1NdcDt
5qrcYVfGY62RGwAVuPCItkdtkIxAu4A/zYRmA9+Uw4y3WWb2kGsXvEqWnHQVCneywVi5MKy6UdOy
7F/s2a1h9CqbdNwhsb7NdyOWXoAGK/oTpua70OhUKc1buwhRpu/KQdL82pgZWxaJigVavsLLaeO9
caf5wGT72xPfmarxU9BPTEBQ5EDVZl8c6KnG6PAEM9NxTf5iRNBQbIJaqtxL9i8KbTo3LIFPWlZs
X6e6epAgE67J78H6rjmEw1T7KpuL8d4yAPyHCwIMSJkJTBRTfv2O+4x3JIFsOWy4J0GUHom/GvnB
/+9+5GI8et82JFLvJikUsJA8GPSzSN4fs8soWkbsxiaOHHs3MT2v17WX8+cHY41q8ZJUVA1bGr65
/UGrArGZJkrCrhE2BrqmNFzOzzvZlIEN+lE2/GoIfBkaV3DPOyUTuovMHiLXchK5yxRgJ5/5ERgt
tH/Q+8q2O4IvWnD4tNDxOTlc8MlIS/5nW84y9SOz+/iEnv4C/qqQsm0F7W6WYcyUiJY6OGc65ovm
rR6HqEfAk3WHink0cdoYtTitvVV2aeZejiAcCbBvs1Hv14Vu6FSm45B4Nkr/j39t4jfPhcqoIw//
AO4oDZQ+xMiwQmmiHBjMslfuU0EpNiQAqE6OPOzQEsmgbI9ylWlQd6nRS+JY0H8bTH2YgYoI288a
ntbgr6p2rPVUA1t3d6O8FEBvsCYmUsNLr3nb44GMztkNo3NU3dDH+8Pnhm2CSP0plWmllAL+Fw+b
Nvo2shKyMUtJ+qTRZoxf5pPmtBfOeJ4ci/foc4zvCfErWYEDEkRvqLhTIrN44/ROwcDqimWfSASD
TBfko12Tt6USXAm4WD59rfmSxfnzge9yQjuPknvElxhzMqHWTK73UvdkY3y3oP2CikNpDxXMfvJk
WVDCJ1uSaEgRpoYg7bG+GjGnTEJ3BMuOtuouYBQQ6+lW0CC11Vp0YopslWvOH9hwKWXWNmoW2Z87
UFLrBJOS+gfeGGeYs4+SWM3jyiR1wVJ4WgV3aqMoLtGR69UoZ7TyW9yOg5Xpy/YQLGUZJDdHGuzV
LDAfGVIeh0k5d4wtJg7tuA04cJRfln/EwYhuobt7AbnN5gyT62GynB+Qqx1BpNMjaeAo1S01/VfU
cGdeQjwmPunnmtrNsZlQEyGCp80/JZ1tjxj2W4MQT23nvVSGlRLX2dnwsG0xEmHaBKv+T7UwQ4Ks
lapupoOsLBIdVhtJJz7eb8XvhnUoUGmM3nGFP0Z1tpOPy1dvUP8mGWOnigDxIEtPlE1L8Lu7B81f
mWEKgqJuToE2A76L+RdDUB6iM/ygXl574sUGVpcnfNfXdQJ8d/j2GRN3qMC4fuiT8XvB2zKxrRwR
8pu/OejLrFSx/YIazTkbJLvJIGTWgqGKeJAhiG30zQmjNiG/799+xzoNl8ZjQOJGbaGZfA92guRc
Kcn8A4j0rulvUCRByY2rM2jiGXrxhu19d64Pjjtv6CzhMPU11+ukmjPrkADZuO+22RKa0ToMv+IL
R/pg7sWK0EIZH/dksgudJmMFo+Qvqv62ZHOpEnklA385cEBUEAbqPChMdcTua31z5sR+fKHcSzD4
DyZIMVsNZIwwG2NH5st9qg6xztQpD+wf71leCtMc91+JpphzaTIcC7i++i5+iUR/JbdXUSIF3pvG
7TQEr/Q/MTSZWdk3CNnVwseZ4I5qP4ybpGXbmhNR8eHl8V735m6vLp57DZhSoCCqbgWJ3R+Npo96
tJfHJh29qPsoBhzUc+xGjb7aHyIeun3UQuOq7BPzN+KHrgOw0ryuAtMuokeFJaaLQNYkx//Q5J40
ezGvfWzRJAQ9VoUbMcmFX5FJdm85wtgaos/KJgXFyzuIuMyiTVHI6Bg2Q8OXgCXVEn++XAdZ5OoJ
+bdFO1OdoqdW2rXbXbOgy48fBrwJevRfnNs3nU5c27IhkVJZhji0K9v2MCtyAmpdcOs/25KKFKbz
VdDerZVYVxMVPMqTVx6q3t0bb6Mr+8vqHjkf6MulAE112IxNupo4qYJbjVaIiUyeAXK7xLOFgc2q
+0Zm6U3phnI5RrZJE+mJX1tF4dOdhW2t5dR5UNb8AEmSdjyHuUBGiclQ3FbIvUnoV2/06PuepbyP
Nz5nt1T8gy+azOtOIs9nV2MnUlY1OmUcojbdTOMZSSUuwwvR+B4FYxF3C68mkF/y6yc0jaa30dfK
a2CO1OG0j35D7Tlvgtms765Z78pg4JmRxIQCX2/ygr6KTxolKNPbpcWKZcVTuRbJYC16WWnkGrhT
OcPUQmcsRFgHTXpWKObrPo59P+b2i4TB0F9WGDxqDN0wPgxLT6B7Uo5JDMy6Szmr515iW7K12NTG
ABaoSkBNm+9uFN+ZWcf9l2d9pl8ErwH66xgS/VTQ1IgzAQ+bnWOsrci+BVP9F7AZe4O/k9iUk9KA
pNJcSzrzRbNpP99QVkh6g7ZbY6id2cIsXOvFS1kPvqIO4pdmTDPImHURLmyvaT8D1zel3FIHBESa
cJK+purnspmrGqodkIkmp/CkCLUS8JyfLDxePyezRMsZI5AoG1IUiS+e3z9a27q+ppV4Cv19a26y
1E7n+vebsQDLi3OnTTJHiY8kGGx8vopQ/FDJ007xkGhbF0ioOqBfFMqp4veLRY9/hUmP1mi0nxiu
t1d5nQAS89a2EAnbF5nK3BmHdT2ymBAyeQX4XI2PCTV+qqF5u9UE/2kbmV5o+j+Y1tc1KRvi7T6V
08qdLKnlVsUdPUt4BThV7FRAncUK3UjP0u975zuT2WMtRJme+fpQ3Mylb5+oq4kMDoeyTH4Ib9Ub
PcLBSOaGcNj8B/Pbzdv9QAdez+BmcVBpr0c8jN27UVugtiRDJJdeAMm8LczAoon7LVlK9g5ZUEiy
0/IqoJgGGmjTqbo1hiqI47TRkKYgqUusLAuwHeZRt17ngVT/v3Viqs3cco8xdFCGiqmaA0uJdGm9
yFRgN2eIbTVDx3wp1e3Z3O0BFBuHap+Wm4GUD2kjDDrQG6i3OXZcBMhADBipD9QTghAZFYkaUtss
Ed+X1J0GroadE1tHo+qhgZkOF53c+kXZBnGvio5vZaOgvqmCD4IEZQEmTM6qUwqE2/Svewk0K2Og
vDHsgD8ATuwDjD7xEjMllmwXKDMAnABgkDqif3NrRgb1ILSv1EILFOTW6kyfsZKIrVKVyUPr2POV
PlS8vp2Jax18PqZ384M9cYJjxWkM5Bu5prRGvfd7PARm0C0lEiVoYsQfvFhfrcg/LMobMm4DkA1Q
dqxnmDXeNsrhQAkzZEMhNUYGFdmHP9RLdx/4yRGfTMGT/dGbFNvdefOD5wrEsEZaDY3aHFhUp0pw
ekmkTEECZN5a8pYhiWjeqzmk2LBM+h4PJ89+R0P/ih93tqCUjJlpShFmrb1LYnfI8f0LoCel6qEB
AP5KrHeu97VJFV9MDMmI9u6mmFOmFVRr5IC5jfXD2c+hiuCONtc99FvZveiNbz9WXhTR70sRNSKl
M+5oSj/po2acB45Uz5ryzL/vJ4EGCVfQw168rlf7oND6WU34wd3LvUXFeLmu8VKbx7koIH8PjxSi
U/xG/PYQdH1kzU7/OhupeBNwqdXOJBFj91cYl4OiCUHkRbzNaZeOh906US4p5JmuV/m9TSnqnCNZ
M9HZLQiQeyN8crQDq1HAMJ6zONInDQoJFqQA2yV7E9Nn2qjclx9KOLigcmCSOAIsGsGddG2/vuXH
AN0lIAUdeZ77990ULLGdeHGv8/7BSjSZbPbrtXRScrS9Qk3yYuqezawYN4vo3XNCbRWDeIrzX7nx
VLRlk6/tBhXwXwxWBY0kDmXPn9HzZnit7dhhTl4aL3SPl7u10J63p33jZmHQp0xFD9bl8IJcYX4f
C1UhO+smSLed2Rrj7mwfGIot2lXXNjRZJHw=
`pragma protect end_protected
