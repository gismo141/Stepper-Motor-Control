// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
cCTFMwR982HlyeVhB6gCt9tb3cf1alTP2PP44k+a8coeD9nV58p9upDa2BuHizU4HmPmm65QOmsw
i7yy4fPLQGs0+xIW+lwBOUdTiBm1oAW8zM5t4nBjRwf8USIqYLM5LpeM+NSRa9cDAN5xJhghXnVU
y0h9v9sN4bObSIIR/9mqaEDW3dHxAmO92YrbBgb9OITN4WJ6uc5Vzp05fgCtfE5EIuV6o1NuU7N8
ZGUcBvy1udyViPqBGdj9nHVQPrCR4cnoT/Eoevtj3hJpESLIG667aZhvte9y9xRaosUPOICP/E2/
XEtIc+gKAqRSDULMN+3dstn7FEFkNNfuMfP0UA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
PhUo9OMRAJTcLYXCcThwxUNQXKa+FeGMPgpVrl4LvRnKv8HbC9tzvnUHxCEeQfOZ/7YNeD52jS2T
hY5/vQH1y8qlAY2GtVYfEJyZb0YpDPNFJk4ipn2LggYhZhsngyaHb5fCPFW5VllA7VkYybkcnbDZ
AcJO9ah7cJ+bhy1sASpovUwczgvkBBiMS02CGnWGDK7fk6txO/vN3TRpg53HfkH+ejk2j2rg5FXq
EhkuWcRHGeHQleTLgk497c9Gzu8wlL97pPaH1I1mCejW7LmOJWCSFXQ6RmaHhOjyEL8bS2MRxd0N
1ffR6zLIvOTz5eEnt6G7v1McnzibhRFt0bk6WomtSYAwAe3H0R5sc2T+NVazYdRrHAPbzq89MXsv
EAzvY7WK+7LpphEg7X6ojLeGNQe4KmtEe670Mi9aOU5BBBtKNPQsvnwx5ZbpqFcTejDwgyVqndFA
/6wNlfxJcA5m5lddoaDY+g92REYJ1P7KSTHPrDmh1tupJZ4N6Oqj/A6qRkgXHVbVybehtTUgyRkJ
OdrGd7tzYnnTM5vLFkB04FpOGq/2rYUSFMCHo0MTZkLXZ6JZjr51JrmFJD5imTdB+1xEGOgy7v0C
9Dv92+V/ovEA2u+7yS5RYNDy4lKr8mwt/roeNcy70vlAfzA+pE3UM/bPzJ66171cBTLbiunIeBTc
2+RGzsdKcOjQyYIi5cDuTXIlofp03P2aLKaBOmcI5Ma+8NMNzXRWGew/szyMYaHV/YsKT9ASlaew
FtZWE4g9HE9PbWIRbHRqJTdGf6TsPsxpHgimEahL/CsP9c5Txd5t67kc8L5O8V/1ym2Bl4JNVy+U
Tq7jh2Aw2aFMWLeIwcC0oiwgS/ArbHKU9bKdPzqQAcZffuay0mImda2WK6jKhw/mMZZsK1027Pn/
Q9fOoSM+zGv2RKCY81NcWw+lookyI0jY6AuV5qwNBtM4RXocaLwxEBHFh4MzIFp0UeNkxZog3ZWN
YjnMilWtYswozcJ+Oy2wZOBeWKS7VdqLaD52snnLC59wgl8blx7hd/8tdC/VhEE5GpsS2pd1iilp
mr3RmnfZE31xe7wm2f7UWoAVJd1ClTcWmie1jBfSeC1NlpAmLI8MtLzVaVgPjSCnBomQG7oWKQMK
kPZtqQ4Gqkfz//luTqLWkP1zh0aewmbSj0GKetdHvaMJBhVGRV9dN289iIeu6khVDrSQ6cKdAajA
aVXrRjL01ztkGKTFRoLneFdm9awyt4JQbxYtBA74LUTz9VF4M0oeqZtNkM5QaIIp12ewSWVamcL4
/SKw1oiacRGdkELdv8CYro+Y0efCTVzggQTRjmS9m81hZOVZ4yEJqpve3C1dANZZZdOkkkTJqin5
c0KHLZzsx04+Hm3bH5G6qQ4gYta3TZ9C3dmkPLKXpYlUnSHMmaNL9tSTMnXaXoHLtBSE1Z6vpEJJ
ttrVulghQLYSbX7GlhQWRqxIGzY5782GbkF1hCLteWqFNBWnmTPT2OfjKnUk2C1ggPK18cxcgD8J
AXx/JFEvwvgIyPDMDWB6owALeA12COlGV8zXkiJaiJxL2MVJKCF+USHuVs+4JlxUQYUl963ZZnOg
id8nx3d4yJdFt/GbqueDVficq8culc7VZJq49BHkKwHM0rwOavjGY9uoXXeGJQJvtWeW2DE6sYtm
P8romD7PaxfhaDvXH9BSYyCUo6hOGBPAMJCMzwXf20uc4WAzlpwgsAhcctmU7/N3Gzg+pBjChASy
DTWWOf1oN1bgvKd7ecT6RCAkP+Kj3xc6+DoPJ7wUfRmQL3Sp6lUEe8Kzs9iWpgJ4lKVGg3/MBb4y
2h5VxvkLcgz0RAL0ewfnyzvVrG4PvrZjsG8w7npZLgg2Uc+PER4um2q//qaJCtg701S84E6DjIBr
LUQFVriZzUF5EgBzHDgAQhsPuH+jlwA+Y9JXV3jH65rCsX9Pau8YW7+JMt1fmWFueS4sOUMgmddP
60+3OH7lK7LNJ3UMWlXJZUKDQPwZNVT6dj2qFE/7ZjqG3eIwIulN9bgY3E08QrRt1lXcGo/9BWDQ
Zb2qK7rOkkm2C9McX0gtEKVwX4aH99Y9jJ9nj9jTUltuN5EsElKaNlBVw+Zrm3gFq65zkQJWfXD5
FOsQCO+8MWUw6G3V99kzJG+sP5dr+WUuAyKg7zgF5d5wUB0StdWPCOqwm78Z9xgeEHUCoSLXBUWW
kpHjZIsAQYtjHk9xo7G7N4awg/5Bev+6G9uU8BPivW+TqNw9XhrYTeg5TBF5alL4oBUSsru4+uPk
eCutmSZk1nGob6X0JRKVd0Yb024k33YtpUvsumvo44QhZukLtHFSxCUtSD3AGxFTZjZTk15Dsutq
s+xbYupaKVOlk2Vh/kpCTofpinpxJJVspaUEi2/LFiJUc495G5vgSeSaJpSGx9BxbA6IKtGTZC1+
DdkDmL6V7cnqVxYmohLOEZewKcC4YeAhmeIN4yjGHTIPcR0gkFwTZ/Gm1IKq4mT/karYObsa9pHe
oFppgykqrWjt7UKVpxXATm6Ic+/ctX5IKoWVUqGTrxioPPsNokZoQy+Fv2iGw9w4bB40LbvZNXr7
PsCWq/FwCb/tK7bsK3DeFa06tB6uBENx5l8YbI0zg//WSzQe375aI3KuFF9LRFUUKpLL6Ef10lys
EC6ZWKc97482ZIH5HjWejOQGi8dPy3bHhq1nH4QvhyeX4LgyKdntu+5ltaUXeAdQhsbTpwmC8caJ
KItwgXPk0UGEDs1d0RiTs06BHXv+giUT+BRItUE1chHgWNQ/8ORqfHtnYheuVUC8OcrruwwJ5+kK
VCsOvEz9fNaNAgiWdTp/fZwdSwaG6N/XDiZ/BcVetUP/VydZuGqrF4+x8FIf9oEmRHLR+1coM1LD
pFXgxncj2AjSMGvlaJNJ86jKWJ/Jf6SVyAQsL7IhZuzY3KsVFLOmtEzNzVzAAFn4iUqhVc5OoMcU
QoctJSUzRxMS1ZHus9OzexEF5vzbrXbTYR+c37Uf1Pdb5CvPC5wOfoBGpgwM5yltKvTP0lDvG2e0
V4XMx8JCUwEI47CTMwclEfMjVdECLrhZuCY/XFkliJlLYlpYTluWKKfviqID2HDAIT2LOFRYW8h4
HrotC6Ruu3Na/hjMZ4nzHap2s9BwoHvz9Ruzub4f5ciiagoxvZYW5MJncgk2SwxhY5pLPBUMI/H9
a26HLlaGbYvz6sIlI15Lyj7dnIG4wwDDaKFiG56/6AoMk58M0Zsyx9rD7j+44pgoTn3WHF29yEsQ
cvYSkk4JviUxMx+hDkXwtUd0jCg6bg/Bm37zVpKxxINU+tbr6/kvVZRZIhyx2NmgUiyOUdpif1yx
rcjZOlISLLULqAPqt9D3gx6prktT9tXqWskglmSuR2+LY19jMW2dYCmScIgs2SXHC6w+uhM+rxnL
XNrFS0LAurY8USbQA03cGIt5mGURFjOq4WYpVNCL/CszCsB5bcuxT2Aa0/7OcgMy5YVybIQLpNSk
otvliaSLrKANcbPVZNJiQ+XRMTzyIQ2P+YRWUgdGb3TR3+C77ya4TPoq/Ge+Uew8kMt706vJZcuQ
mndyoAISClvoOtDzE5dF0VgRwQPF3D+4GlP6g4dfDr3iVKaYqoqd/2c1aMPtUthfBbLSus0FLzXh
FXxXBY8j8KIsJEEmk1xFihxBS0VXicnAoCCEwF268B0I1tZREdliR6ETNzkicyHUOWHrsvFznLxe
gKzn9YUdUTLTFDGJXGhnFeRhbGVCdQZLv8hiN6f73FjBfGV2oW3DB/KfaPoLmMpWq/P4cvspKV/9
C2EgwziLzBLCgTvmkO8vwYTOk6RcQ0PqhSZysny0qQoxNfxalluUFKdXxF5kX4FF6rZlRTF2Hf1a
RbmGg7LfE8nXabGSilRyu7EpjxUj8UTN//KBM5PBQJOiTLCvkI9z7DNsS63appe78T7OpSx+Kr0D
Bhy3xSaBf9xeyR4WWYHgwl2P6YQURdAuP1cRyAiHGNHQSIK5JEHWqGWG5/0R9/m7JiD4EXuqTwuY
bv5zZ3SZ1Nka4gXlkONbJbirv4xZ+SegVgOq1ErRrMRlbIZF8bf02VesG4v6eRrQRH0G/RZ++Mf8
hFC1kLHuhqD3UYcgoK7fMC4AVzrU3sQqtyWPBNkMO6rRlbMSBrC19bqwqEk5+bEKTKz1eY2FZqKb
52mgoGWZeJfTLr843qwRA29xJi0iV3sHMgrqaGxqBXcuIUQm9i3eva4c1PeLThoRuzmgltPWT3YE
Tx25umSfIul4ucfgIaWMSrMs+aJPtf88SdzhzGSHPYAact+WpKVYCLm+449H10Td339GpSLvpFB2
tBRTctznyZioPDh4NTzR7puiXqakpkTKFNPmdAI+AXU/oHTzGQWQakS3uBal3rqTY+j/uW+XDEGt
20vrVi1jvhIeBqSnaKJf+iKKhHWiLOXyY0hqOIdXa7Vysfk4W7a6J8i7hjV6zF37IZsfiMDGqIH8
ujL6guV27l11gF0RIxJ0carBnW1kpre7vIOe1CQYccsbRzgf97wFqmmKyVty6J+Tlr9VaTjUUhLl
VeU32gJSkREg7of/9OXyBgyUNiCNm7AmwQZ973orbRrOmamXayI1xa0kTKKAShxCQPzxc86mbOY2
WLA/t/Dj86Qdw5ZI73cI9DxASPTeTpAAe0FAYw1sQXyqgLk5S93uTr/XviXRz/b8M93POk0ytlQx
ImwkY11BqLMJ/lpxKY1K5VhhRuuL7pzYBVKEjKmvx8E+aiSYUaCoc44HYepGqgfX3skswjLpnkkw
EJS4Wo5d+nkaRkpG+Lyyss/GekpUWMD/qGMqmUUehviQ90kb3a/wSNNA+Ubn2VfxXMnkQxaSmEhR
kQnAc8/TcnrjtUaJTrVd8ReqOrXUO//XHmYWz83Bqlga9ntEs+yq9olAXHAsd/JRegt11kiep1IS
evdoiNLq6L8VlDiDF1Fj5WRAE1CbWbiCJFVIgOszIJ7XOx3bOKcFfIvgbVe8KhDZcJCaCJ7ckwOH
R7BRiNHc8sPsJETMBMEMj1wsUh5wx9w8TYc+8iVrWzQWG0OdJdPNbq5FRx7zRh55rcS0Iu8DryR2
ehE0uML8B90C2/jJ5QoagW/9UuOkZn5yXfe5nT7eQwDxSLE1nBpEUwOXReTPLcnBbQZZJCRhVpJD
yk2J+A4lBwkgmj6x/TTHz8zQqdzAu8Dv08HfJMWEZcUfvLNKxd4Xx7nAl2o9HweZYqcDjVszdRlc
b7MAA1C1rXN6nYUmldAimVcHiruvzNCy+4Uezuuk6Z+JIOMyuuAyNrA99MFmnPUmQZsWMb98QFGX
JMOPhZVEk1DPoeRDkF1nVaoRmwSwku1sn+dHmeXHzU7nJSqbbecVU0VDzSIUVQXAePziZSARd+TQ
Hkd1rM/Vrjs7hpIV6sktL710dWb5T0D7fl9VziLZQpYc6SRzENYxY0MAnEyppEuPtbAGY1pv3ZhW
MrXPeAy+KSr4+Zj8IrnNsX8cpJANMu0UWqopoqv+bGp6DRhd9cFQQyd9TPwHMlCC65sRF8BITEp7
UHr8UBZKZolLjyoewCMv8CVRMIWJbr6rwqhoVUaSpOtFZTzXyXjlUX2asWMDlX54W31b6PBKEK98
0FsOrDZvIYXIB38OI2NyjErJX8RK4tgyzISyhDXCvydMlvOjXzTNYzuUmjzXjODeIoGZHBAoDM+F
q91Xt5Yr1/eVqYOgk8LYniLERgQxjYnHOrC16L2frVZI7xc28+ZouayTMlj8ect6sqV2HoFpfKMq
YuZ0WhlktVQ+x0CBKzKo2KV0Srox9m2IpE/3n2EUMylQVao+JA6YrcTxiDnYLxrN4XVxVTRqxIdQ
i5LVf/5IEq8hJ/FGeOoGxCoCZxZiz9/M6QyDP6kYAFfqH8dKSbCqqVztWmLgvoDl6vX/RMAhW5SW
ySejZ1dcJyB4o+fGztGv0IraFKXfR5L+wfEU8UDdXi1edn71nqS0Y0+2X0sCJ18TJewKaKTrAPxT
/bLs/bnt7StZ2yR2Tj3TjlGhnEeNXXZl4vhCpaayeagdhA2KA6GdSgMcdBiL6SZRWijbNnRo0MDr
hCVfT8J98Lxsc5r/TTftrpyEn42QrhQi0W5kLPbGrvB+9mnybY6NDEBQ6b7GNzeYGd94PjWJMZAh
0rvJ+cWjQq7oQ6Dtk5wKK9eS4mwA/xHrAmRklNDKLO4XgBCIoricmxMD6r5lcmQZZxldU8O8ZFao
tK3sLO1qUsWsPH3cspGkqiBNRpxiHobgtyP1oHwQNNfWkc9L+QaRH/gGiXb6O1jkhgR9facS4Psr
pVYuCRKA8FWwp93G7wI8O3LIuGcQ5sepDg5TJzRSMm/iYYsh3bi44IVord5XsTtOP8PElggK/omH
9mEXZADfsSK+8Y9pMLTRG6K5hOcUbKDygx2uBh/z9Adl+8H4RNMXwKsN5budxCDj9dA0HXc+H91x
82si9btqJqvKi0fHFi1hfAooBKp8ja5QGweqnl1XYZ9KRlmvg+lpqZU6JQx9lI4sPiSiT/Tp+e3p
z8o89VDn2BXJ4iUiLWZJSqmNdZqQz4wBrJ0CuS+wlUig4TeYlnAmXgRM+6RkDdr7pkgbempt5Ug5
n1EHR7eCNNuHIcyP2sLjEdeEn3koblmS7nhdcGiEnRqwj9QWjPSHb/TW/CBGbWSjQO8ksIxNnUXf
kXz/LOjPd6I4T0vdLACdBVccCJ7xAaPi7VPyTwjtbq24QI9WTW8VWHMqhj087ueBsH3PZgEOHbOX
1eXCdaWmZLBFhP85yURE1+GyNRuzuEt9FYsYhdTlHRcyJ/ljtJL4gcV96hHNwvCRVvmWTj+YD415
NvF1sFXWvDRUXSBqEnWiI1ghS5YY6mNDwbBf4Hj1BbFtRpVhw0TaOA9MxcXWnSnwmVT7NaO8tVTR
Jg+PCK8wLRQHquY0KTcu10JGSnqgzXqykhZnROuS/zBTf526bViPFfNOP9CUCYH2gyH+6l0Q3QuY
Z/DWCOgadItqSKurUjDKcqv93S3+oCYxy0suZeJZDozvHz/a7b7CjpDv4w8oMJdGp/leQYKWH5Dz
GRwJGUESqak2HBRdJ9XhZBgAn+WLla4G7tYxmaQ+YlD9muH3k53c2h1GPMvgu8TT4rv/klDfMPPI
Z9vu0NfIIq3Fli7VbhK1rNlZRaZh15RImWc+b4ObTr7jDqo+bAykWdRif2z4E8+K+PZVkQxCA5cZ
QwCz+GHbqgbJkKTjY4ECjOdPTDlpGj2x0ODT7xnd2+6wkU9ZsiA3xy8QYckt0SUMadyt+/pC3MZ4
ToA/LGZ0ohfwk6dYRehN7K36Whj0x9LTj4ACFnkwuGf44FmvjbxsPFZtGY0gqphzDWa7sL2ape0C
e0DvuxflbGA9aZuWNeJ0mPqnvSMpBKL2+4to9VivkgmjsQV+sZyN2d/fy/+PmO6nJvWAkzGShzoo
oS+jkFRFiWC2YJOiO95yuvxiNmbiSzr8KRwuL+JEylUJSIBKONeLx9jedHGeJFsrUkUum2WxnU/T
B598WsB05wZmjFCxMBmN+eLNUViFa25kSWMn+aAlaLXipIXG+VSJWjH7owgI9VVYKoSu/8A3u6x8
QV7P9ZSrYt/T+19Q32EH6BJGkaR7H690oRCRK9NbBvCAhAqpY+xMEFG85fyNUhaVYyjA17GBhtZp
qNk6SrvXunut8CIHd64WbmQtKS8csT8695r5a16cgI9uDUKc5h5V3IwsX7aW5tBhi9bq3gVjRtXz
liyvWxvNro90fJEogEkIGmXfQ/Og3VRQ+4vx6eJ9J6k0UEor/PNg/i5EX3mp8wSxil6oWo5IeSz9
5ex6KEg3FrOZ4iwMuJBb19ErJTv2WXT31pDHSvl9gecj4eMAKoEfuSk1vxL9SeYicC9jloS5eZjL
wye1NvAq3cesLJcErluRMhKWF/5xgDVaUAJtX2E4sX1TI5SBPV1dQikfk90B340uuTogpZ+vPq0Z
KC6rUEbcxW4qO+0HrxMhZpyav+PVt0rQyeRBXOka8igvcomqKBbjqAMvapRRGyp+ti+Aaw2CB2rJ
VYWQtQWan1uI6SZdagc+72igm6Zeavd+uS26TEYlULZLLUfBMQInntDeuXdrh2ouOCvgAh0CFLmp
4737BVrO4qAmnEHQD98Kh19R0IcJFRB4BczwAHpYZT/GtW8OjCiIRrauJciq4ScoDAfwpZpjGcnu
euMgjhWS11qu3NmvLaTS71N/eFPnnKVOfwtK2cACSVHodYUgqS/Y2m+iTKOQvD8aPm1FBRSdoDpn
BqzEg0rbWufjFq7gPV7w/zAwO/Zp72v+Pj0ROH9R0/376Oz1HTvEZQJ0wqDJGbj3SrO+rjWdSbKj
6wjW7mBQ7LURD21ckKH0JTtEHz9q8aotKOUYn8ZlMHJigSCwkvKupV9cCvFjn43Bp+ZhNFLy8iVT
mWu6t5hkN2n72/mt/871am3g0wOyHg3R4sHrDtENwWog/n4XtSiaF2kHssOuaWC4q58iHUEmrUn/
LUXc5WDHjhuambEGZZT233PdKm3Z6o/zuX8Sxd5B9fzcg0JNIjiayq406OOgLKfNRSKr0Dk20HjT
1AngfAgIqLDBTNvPx6Xhl+goTEJtlzILFbnZLUiqmz6UYaDZzT5yxBKPFv/ylzlUvUVGUjIe5bjT
dl0tr/VnY/kT9hc3rk9W4vBQN9pQogDzJQQJj2G2O1NFy9MwIr5tjBu8mLVpy0jBbOcnay/XeM4Q
B070hKsq7IX5faFEHqvaL9CVH71tt8e6v/ixuFyt1tRxLuFFIEndGE90GXm9i3TiMFcvo1R/2D+8
8Wp23flC65h6E97SFSwnHQC5qMBJh4CLJtFNc+nbwq4ROW3AsNLG8jOlWStVJN/3axsWkCAYVpya
EqiYiFl+j2tagjKv0rqvgpdNP05RrVQpVUxICfy62r1ILP+k8BFDZZitEdCDsm0jAnm5N7Gaq+pv
hCXxd1iZzhlaX+ExjdKnCNadrNwK591Xq7PJW5VSZ2lZUEMmDnKYZkyJWVP9HSg2PqVXDkziOJBV
ewGlcBX2zERQWtz+6DJM8cMa2S+GZ/UDa1jdo2MrQfFyONCG9ApM00vEzH3wCflFuDW4vpfWgfBw
QULIJcy7wtNyV8g0eQ7+urV72AVTmzhTE++myxdM97m6As2ABT+PqBj62954qSXWZQJoKerJqRIT
75+PKaYkMXHeX0VpalJ2ekdNymYNZI2b3DSAxjK5Mn6IBbxYoClNq4YYASCS0HsGRq0IGVgdUf5s
iFHN0A52qejQubX0Yg4KCxaKQTRf6MtAs95vjg6XAz3c5SzG01B7Z2sqeXKcHgTTI87XNVMKbzvN
B9Hl0MeAV2jMN35nYxqMdXYJjAFJZZmrjAUO5GwiHR0M/Eedvkw5OsSDYXnllYt4cJGsQ2w18zjB
NT4oyKDkW3A/nXS/Ohcl5KYv505dOLeE7OxHCJsGfHINACRcZ2TQV3OuIV/T045u3sCebumtjpAQ
oRe4VZKttadjYn1TawcFpmJ/m6+Ue223WF5emT0BUwghckyzNiXEsbPmaZX2jpO+KnR3yME4Dx/q
aK8nAel9r+t5wsWrRsy2yNnqwUEx436tAaNhrxDLXoEILb2A2Z7WVuWGca96BiVPPCDTih/SXTQE
oVlvVpP8wEirR9wkL3p2XNbHILzpVSomwCfctwJ3zSi64HAm9ZyCM4kdiNCWxYNGDt6HOYjnxuRR
QT0bYTzt/xS0GssYpIJ2Sd0p+hOBYGAbLM0kUcoOkpcr1Ep/PUjt54Gr7wptLQoVXMR2P9xmi+43
57nsaWmbiPeJo+PSTDRxL9R81DcTR94pwi2LlgbH5l2YNN7xKy7Oe7Jphj/KkiRFE9THYBQzOhOv
AFmuM2XtCNrj4Sp6ruVe+33tB4CT2hZk04Mtu8ixlNpoENPXDQkt+O80cDW5+1xSYMHuzrvMdf7m
iex3fTslno2vqSxtmFD7RuOwBLoWL4BLXPN4+7ryIwu0Xy13dYN9nbT8BaYiB0lK256o54l+ixKp
Z0sW+j+hGjZz1nz2jmZOcqJJ7ldapi+dPPjhlnlod2SzEldFqOyPbgMcBt5Rgx19c8Mz5NBsSboF
YgyaK8EwmxGJKmcVj5LAiSBGxykXUkmke9NV9YT7lSY15Kz3CKzTlrAeHbSIPbrnPikhnXrX4Nh4
NohgUxINu/z4IQNaDX8oF97+cKUgpSor4xiwieysIb/f113YRUVhhA4X6Db/ZqFjsWjqn/CHxoY1
eu+EbO1xTksO0e74WkqaNz+82M95L6p0HtWGNaVry1G9SUWM6JHaZynTL+eb0Ul/6rnoy4ag3dVo
41TePhTnqPx3UIVsi+6XavigeKnbczabs2zNrTC63hmc55duCtBFIs4aflu/Cx5K3gxp1TDE2pIu
EvGnIFmVRsOctaIAUjGeoj4j8FBv2G8fVPunRm10cLjGCDHPjF+KXiqZWpuvtorQUEZNuuo5UUqv
lT453fIT7uw6jbfS+EqoiGQVypcBDpl3cgM8NuK3xEjXfRheu5WvqLO928iJfvfUl0H2TEhQs4pY
QXSbotQW+FGhm8jPfNBfZrw+oArTClbszVoDh/Y39AVS6Mk1dZ0RWn9J/DL+pLoHMx8bnDfNCfro
xuYcCPfiK2JPJYP9riw0PBkORaMurYShfzQ7jMkDmvmvDWBVatl5pbfL5ROLy2iqRiSKtbkDbqiu
dEkPQrZ/+vywsd2SiH10/jjMaRuU1ESZbGbeq8jDUQN5bpDWqmIKndsYqwzh0DT/gn5Ti2ICGYzK
zliqr31HFlxEBSn9lmhBgGMXNdJBJezoldM/omzF3wDUIlbej3SwvKzypBzfcs7WvQMX1BfYXoO/
ccE5Ps55aD5YeWQDOE1yh1OHYs42k4x8Yo81j+3LsB662iGTGKRKmT14XDFUuwy8J6iDCwLAgv0m
BGJ7+sFgXVSBU5VssPrRMMTu2Hd3Y6KDqpehdr6raj5iwYzrqjZJei58UAOJ6qC3/U8oFXM+0l4N
OcMdK8aqfFQIDr7Jh4Y7JWRmWXtsxS8Tx6hs6IXAKzaSmDL6aCorjBeDzot4kDP3zuNLztf395Kg
2cXsP/PHkgszGHWF3fptBC3klG4A9z2OreGuH1Z1RxTLzhvdePkFMr3e4LdBlUXRc9a63CdsYxA6
besXSD7oDbrKGcLV5nquCscJSCMZ/w3/R5+hRTmBGSsOezznVTcAQ11mY3L79LzUwgRMYfUa59qV
y4GmiTRGoZsi+/ZKR+Gt5uVPpH+cnBVXPwD5JLjfmjwLj27GFMtDAmKu0DoG/Iia0ylSZdzoCtPB
oMkPoBEfooA8YG4GvbIcdAdhM5PNjziXogAV7sHw95ACr21cVn9rRANCA0HhPDI05UngtsfjY2Cs
+6IL3QwiGYnOg61+FY8r8fSwIbv0C6rPdMqoX4c1r2NcKP7eihxPeqAxM5dvdHb2DFkk4asqn8lg
IlGCdxNSuAIVXzUbcz+y8eGXEoFwqB4c7Pe4eZLysVJrPlZJojQWf4FpKGH8+fFu1OonNFJIys6k
2tWHVUFphPwsef0+F7rcS5mTkYg2qqfn1p/eV/CMhEVF3ouA7qJYcMTdqKzA0r1c9eIA5rtC+26b
QaDXHtjbERhgRgmdAx2sWqvHVceWZTANdOcUYYgcJn6Aqdt/LBRoeRvUElqF+/DdbUdUf1uOXvvI
oKHkYqQthXfMHtLYkVQu7Chz4qChcPLMv0bQ98jtC7Fl37ga8jkW5tnfXk6X9nIaG+2ZDc9fz/L/
EZaK4R3Kk72zyU0MBJ/5nXT5lr3F+WFaAg9sqN4VqjpiCm5nVl5ZjQGp5FhP2WgiqrRQFFx6lm9u
vniG3RZ53pY6hyKIoHGIcY7OTJpPoglNbzPLa6PadffNrnHI3T3enJKUw+3gAgO/7jjzrNvJkcrD
xnwi3eWZJnES3o6K18mon2va6QqPfYd6pftUD4nvOIYAjrDdwQ188nbB1IxSEMiJRlLXdJqG7pgL
EsACIbQaqmPKYcQ4WODxPMn6i7axTXEABfvSiVLjwOaqw4G0WXQAtHMR4Sp6g/DraSQ+LUszEzRJ
6bX9MpQLishA4bcAykh0wLJcjCcD2AIDl8V7YE3pJ8aKXwrK6yWAw+rHKIioQ8PbIgoFtBKR2Lyh
1OU8PXc4BM/mp3gWkaTxaMZvnPMrnQsx/2MYtXT4AQY74nPrUvz4sXN9qEnxKVMUZl06KZ/RI7ed
XDLKEhZ84wAxQxyBJLDuZY3oPWYIDtRqEEApKWlwFeKscEyboJPAovz/bKbOaZs+19CB/apl6eOB
0i/XLJKgsplj4/CFBJylN4V/1tbscU5ym1LMkWtsNViEMLnfVXsOMuvjCD72PCXY38ad0UckGqHh
owgjM1Ugq3dFEppEuWYl6EfH5rn4W2fJ4ShpEZEQz4WOqEJeAOR0TDnymigB2TZYA0WpiSUxhWDz
6oClOPWaLVq3bNxIrosAD4nhsg2SgmZBaBangsIhBN714RhluQrDlXhXGh+XCN4Y6rrFWEpM73q+
nxYYQbrUrsebSTGZGzrQlV4pGhwlwmlluCM17B2EhyLKg9FzR0ztZ1OY23RT+5U7jmRZHXaZ1E5u
0PAeHoKrL7/UxiOMr3eJ9zBwmuG0tzLg5ZfOt27Yxgrxx6DXn7RBLtqm1QY3+iksVkc/eKg2+TdU
J3YRRl2KemIa6UtpGeQC7PMoGLmp0G+/qrGnk1U8pcTBetwi5I9MUYVJZAs9N+v7hUsZDdn/1t2M
RAqYY6+XalNpGDER2vHSKUXiTBhbMd6SGW/yD0zNSiquGgKtiwo30T2FAaJJ1XIRxXDPhxQsMo5T
yd2gjqS3TCejqjzAec+v7NeSRnJ5HBXHEOJys+nOlgr08dt6RIKzc2JuhVcIDDmUX3Shbd6zrlhq
7d4QyS7J4hrzgwsR2dmrR7lRlpRpVJgV5ThtWR376B6iNJGqDEYH69nUkBdj3oRsZURtpfUo0ice
pvq4KxLLfj5DsFqbtBD9BBmieV4ou5E9yabt7VBRtxI+LOEy3wTZX3MDMsvHWTcjJzcH2dnLsaeR
frHJOFxmpjDNwtka5AV6FVTcfNVWFGizg6BdQ/pxnbCstIEKBzAqfMAQuLkcym0QygYHRxAQsyy0
Ln5G8kd8NmQIIwpXCXLwFFbLnJ+tEZw5O36Wt3rBsJl6O40KY4QqssKccC1Ads5tLzI+6W7Mq4px
jjZTqveXxc6CKE6BJXgOZ57JN05K9ltk4FdH0/7aeq281V6yQSALLx4oLQyp7R2DH5VZDhsZpyej
x0ioqBqrfcJ3zd12CRI7T92gdER2+hHls4MnO7olbQQ0vk4m9knaPNNh87vhghizPVDYCehcT74l
aum1OPNHp1luJ2o6ZacRCD2OZs1eE0oKqXDEUVS82znxJwE+JvyQ9HCBMT/iqpAGeYNfWcnmQTYE
suwTAH/LZodrXMepvaeyZ88UG5fGsf60V822idgllaz+vl2hsKVDTYKNF/7I+Phh6bQ0wWH/OPrt
b65LUOE+Yzj/56DYilODHnwQ5/lcHn4F1nNbT3PDH3iDdZEpFiXyTHl/XO4ty/zRlIjpTYid9c3C
26v+D8YpQLWae2TN1lbqLWPFpt5wqufaQJOD/n4AX5USTOt2OrNE6jTY+LnyChz8XOuU9h69iKCL
HVhCizHV7YxmuW+eYFChwyI/pZa+Ml8f4I8wXFEsXXcGqx0GKkcBOB1YOvWhgGgIHM3SSLhZf63Y
K+n4qCDLe8s5u9jlNO99DM+orEhwTEAXDOkcIsrB6eR5hB1nLGH8gA3RE+yCZCQNeMzBI/szTJB9
BdBOw+JPa56msnfqF0bcMJD9Cee3MN9LvZfRiELkQJ3xGJYKMq/rbDNbQARR66LFmNBisyPCqdBP
GnyoYX854ArMFxzwabBbGdH4YM1ldZOLhrmlTl5SqeYMuAjrerl9cY6JW4Uw7JxqDIq7VT/hLuLM
lhiLBX+kaAaBkrMB9ri2g6qooQhT+jYHT1k66NOS6ePN1Cxuei3Os2DGO0kkfMUIwCyrISVOH6xB
wBHuu+kiOd3eDnuz29k4R++sKGUDKV0YwkwGq2+AExMDDoso94STNuHWgn6nZDgmL5U1Jmr4egJC
OAULPR2kX1YsyMgiP796mIxOjzFxoy4kovShUC/+eog8lAXypPVzxpCYIDKhj+0RGG5ReuIFcrin
zBn6yjeW6d7/qD0zGqaYlJ5+oHBzEwsFwfXPCRyHTlrwvGEULhzEKILMbqnFYtJETLBByBnGS0eD
cJSeCWkVvAQ5erJC+Qt9qPOnSztUSQDUB4MS7GmuqilrmvwS5CvxlsTpRL1F/Su66jN/kLhSB60u
/d8wW1lyncBWV1gXk2mbItqyWkkF5cb8v4G2okzKb1aYVHsFtQWay5K5pf73Kg+16A7g1CJWbgeV
Vk45bccr15GlnZ+rp6ca1zrZqAtYF7FTDV0q67JIeKXcTybz3JxDgKBeYa7yKUBPCi5WmtI7pfCT
ql4IrUkZj99DZk6RGb7TXc7MaRIjOt/aRO9AORCohHLjhiFy3uf/LgXj2pUhlCJJJ2rMwyhpX3Bd
yv4pXPSaeTKFcEWWa0LD7QrXFPDXz1hwRicg8TdUWwkKD6KFPANQkLWVoUUlLfkCUPFcRW3m6SqU
tUZYKUksllL0ikOiLzaWJgmzzFqLo/LTCwfpEVkhTiA8fb4bqIsEvBlx72he8c/kVUxQusTMLOtE
SGLnc3C3AGloBZ7go33Q2OcQEDEBo00QaRyUkBX5GwIAbx1Otrep9rr3aDpIQVPhjbKRpqxS/YLK
TCzTFQStUOr6N19KgR9OLB/DOGXjcwZS7Ima02TPl6KF4I5LLpCsFkU+Dj4dkjZUs2C4LgFGaBov
EBFV4+U3l3+1cSVj35/3CqQnoU692qAes/uvJFsX2Z19wyMfjYXznr9KWkm0J9fsAj4NeEV2xA4a
3Se+s20QDaWVoDQbwYazWKBy1EzLmN1U3kPheP8AJBKVJQvwIFvxnziXM9EaMslz2/hAs2eS5z/C
hg47Z8ipBbw25lhh0QRoG1CTkPbkzFsXjSsCNc+Aa3W1ZZNs6fSpiSiVcOr8bEPKbifcMssf9EPs
nxgqsd7D2zcUipe0+FxBWmruD/YR3yd2KwMJHbtidieQTT+2ZGIeYXOtgAGkjvHOEo5quVxcFjHu
H8/Ol+h3kUroRVuN7klvImnoANQ0bM8qhcMluwRYm7ZsgS7GcOK8fMUWLWC/VP9w4Ga6bUYZgtX4
lDX1mQmy1ZJMPa0KH0tsDcUDzksH+ebuihA45hw+rOny4C6fv8SAHg/anuP9NOvzD7dF2GnVpAZz
9SE8oIf2EVSXI70ztym3C9OEIenY7vwQN02tjcJlnLu4ZxWQaviIjMECWlyTj5kZ38FmpX24XQed
/4Sn9EYFVm6rSqHvIPQU5oI2GHZiJJEWYz7g/FO0lTqOWfJHb1FIH36zj5Zn6G7IxGutR66G5GlI
ECCQaaHK8v4Zrkb65H5R4/lzlCtwLh7LJOu3Oo3kMOwYJ+QX4/memCCKlvDrVzE9bsjCtr73WNs+
7JRsY8/pyOApRi6RiWnqvpj8o0UEAuP0RLNnUtyyYYk+q1ILq8BAinks3NCnuLb5EDCcjIhgZ1il
QXxTR+Bd46qSJxM2Quw/McW4i8yDNwHfiUchFfFlxsGqCMJKc93RvsYcBWsG9VYjy3Wmfw+tepWr
qNG4RT4Vc3QInhEmbCJfnPqutLhJiyVe9a5L1f8NvGDaxqK7WSEaAEMc24AwAMjMHfjx1f09TdvB
0N9b8XaDvO4nPLh2YgKlK+s+6HrlveGB00s87ozwqEwsjuOvvLtHIF56H1njip9/Gq0f5nrpkX/1
yeH6hXe/L5o4o7JXkPSgaWnCVeVcr2ZGeCidUbch5qVQxrhkPHLHgO6vXMqfB3ln5gj09/Kp1ydu
FKfix69w4I8QqxVd8C3TqGf5egubMtUDcBq0DjVJ8+15pmpMmLe/SfstZLwX0DklNFcB4P1HwBQ4
mYGFytrw89K3PqqIiLs3C0nKMojljndMfFBTkGE6jAgOdJxpmvwggsKuGaietRVuaCLDi1kdi8MF
xEQ7P0o9W+jnOw+AIKiXQOTsp03t7C3Lm3tgxdulVju0w8sLZ2uw5+y1U+7biwb2rUHzachHX0sX
/HApKJ3GoHY7EECq8PaoNj2EcWZsNzR9u6q+xE8wFqo4A28QkCk0T80wjwUr+FnGzTEb5ElQpwtZ
HSvhYEauwwQa4XAASz0UE5a6+95vo4gGH9QkXukv60GenHefoECfy5EM+nDAATn4Qq6WmcX9KJtd
zi+tPsz44FcRFCVdsj4mMqnAyhVtDp5zy+qJcdXGB4SD6Wwes8DDfaKogNuvLw7EriI2W+oQVlmo
WfO8c9RPR1x+6kUltqv0AGMyFLiG2XO8nC3P/R8f4YCK4umtem03OPBe9euTZ2TsVgLP9EotEQKs
g10DfX0xOGXXNDQx/tlHkE3PKRiPUSQJlDGEFTxwgc/Bpng2PH0Q88ezGc3obvYvH5r5aUcYV2jd
6Cv7J0BKP1GhPzmQb4M99DsYi16qoOIdqSEz9P+iBasMyWDrZJYoiiL6a/VIIZSiNIxi9XhIyKDY
UF/ZRUtCsHNzovIQ+FXdFyGiZR7sDNv2ChM7COu35JjmRUQcGR/Iq66ZyiIgK7gVowelUjj5jnWX
EPQd48qdK2KfLObU7s5Dzlgiw9embwpyOI16sTTpgMMI27AVnZDXrMpUQNggSqXylHjhjOfmnkmh
3PsHaq3JMmneRfneI35729qLybraN4PltIj1saAQJO6UyGuCVLGs33r1VuhtanbOjtffC3GwAC1z
t+LDun/o75H0b8V32cg7DW3GuQs3pDJtauelUkLx5eMODLLukOupR/cTJ6sHcNc9KoX3y9CD1W4N
zV6aeMzDBWMwZj/TkUK4TYvyMIEg0GVL8h02qATqZ/IDaqtn7ysGzQX+JkexQoaKPVstMBVL3Xc5
3/SH1JC2y0MrmsBaSHxpKiwCbNQAIi3f3yvgI4rH3CVyrmwVLeWRqmyoiZefH3qQs7sK9iPHful5
cAEutxOq90xahJcJV9AkAmkC25rPatEggLwlM9Knawi3z0et515sRtZByNuOal9/Zk4OgOgIuaFh
nDgL+VpTDZ7y3wPwJo2ULLNQm3eQnEaspv4zGr6uT79fyymmEhr+mKZe3OEpIcWGyr+b3preDd/M
nTQhbkR8h8le0ULpMvF4aTHDmv5rl71lFUDxJNqm7pAnRXccgxVp1rd1WQiqBfYNoHli8o9rqYxB
YhOnQiezDfq3/nPu0oZcH1oeDidu8Vc6503ayqjP/rlwrdDL10jCb7XKk5Wy+SD+BdfLiwCTwXpG
++3NxX0c2m/mxfQ3GqLd2J9TVs+UN8zSfFcmjvqGi2jx9pcVCmyNa6lGU1zohbnquuiYZdyZRQ2N
nykRWkMaRPghods7jOZLaIxI0yub9br+ZIFVzYabLYq9Z4B5MXK0Q6B4rTeGQeN5OjYR7jw1oPGP
AbooGWKhq8pH4jEmO5ka7C0jhmCGtR47CflnY2YV0rbcxxgQSXfX831954Lxd0v2+M8N0riJfABI
Tw1+1/cpPDpRIKGWMeyUH3ZJhnxQ2FzTBIuHO1oZeHWBs3c1BrvuxOKRtWQINhoMsYkpSeCjCG3T
PHtXFmYuX+rn7MjADmGTPhKc5SJRO49rucyJclC3Wt8VsdhyiwDvV4DKLBmJDb3GgzRPmSKRAWgW
e1nx9rYUkQcBE3LkByeJfPV6MkAYdUB1o93hPd7WoRLFDf/5KEUnVfG96g4ZrRjPabWoFO0/G/Or
b4VicR0Yp4x3GhaNEsq3YDnEYngAbIrqqkWLmElQX+WCDcqjXNWDCFvImFTcYuP+0BNQdNOLYcXN
NXXWmDMKnuDZQ7s0pUhHrpTpa8KwswvzCvZTlCmZ0oQ8AfuJmVDsmWRJ07V07HZMaE9s9jADJZD3
VjJEq1m0RH41AEZwM4xrSjmBizlta1o2F6AShuwYHyBO1xPorX2qukq921wfvNr+V/ippxqNySDy
MHWLn2zYojv5CoB2bnlOrIOTlcKQb2FuAyLbq1QD+eSEHmDGaYM1xkXbz4Qiw0bBUhS9DFxUf3Ji
rGiO+S1if1LARJV6BDHTJR+11OZVu1/zARiv0qOnnFtIMmocnFk3OPg9EwO3cFPX8SfAG92e6myT
ozmNuPNKwpavbdDTPRl628nH00eJ+60AhVJjOUZSFriKG4syAANMFzGjHh+uY7Yjft39Xq6Uv8Oj
gxclzFB4HW6omZESkqwqbY18AJ1uEAZoymxHjjiM33Jzg0fpCwDEGVpTg1r+dxj/jvY63MJB7PJ8
TvDdE58Fjqe4mPqnpeAR6vfRSvkfM+rAJO2D/a8HKWn4xZsS4KOPsexmWwjd1Jifte+xr79cUOeA
SyxAqzybaUcAaOHb1mkY8OFTYKibzqzbCfpoaxaYsaRtQomA3YKsl2fDbVCGN4UAUUEVDkm3ny/J
gwhTw0GBEOeFBdip7Hj8hQUsQTsyH9znTvdFn853o20RDYk85mwI6fs0KZ0QBHDNIyvhR4RmkIva
3AWQQEH3fbJEt+40h0vHg2TJrz1Q80Lq38vJkE0IOLRIdhocYebc6ZwCGg2g1Uo0thbXxPwRGh2o
E2XQMom05OwUakHgNfH0ofapWn6rP/BA9aG/0FO2hHDr+X16YNBB1jks3qNvGU7F5s7REHH/x33l
EjamLLDeU8lMWfUGyToc7F2uriQp05CpFK5m3mJCtokjr7BtLsyoh3W7Fwdv6vJ0LdZhl8MetgTF
8Q4BkHlgr6CwBkFrrQpbeHM3nSA81N9uHu1F3wk5Rv215uVr9QhTNvyAUUKGYnuYzxumZNYMoSYJ
7FiPiVnHvKcocSf2JiGYsFCEmxEWeJORiS6IkDKcWI6Aslc5wWkQJbyBFTh+MM57oUXTOpD8cWgr
JQ90kDhdfWJAMgYtlMPj1RKl4+qw5DyHCrNMg1VRIPs+kWSeRvfjmeBau0SkbiP3sEVCym8XEsqQ
7dpeB4HqwvhHbvRg9w/Pqmv5RsTIGbDfjh0v+oCz26iwmiLe/hhmxnsM9OBrQRlLC009+eDhxD96
focrO7b7REHDpVhMGubMcjVNX4/YsnydWi2I+kDRhm32B5RV3oC+fVBs2widIzbK9Kd41Lk3jNNN
CyuGSToKAtqXSEsrwvGCpvJ++9ggLE1F9kl2T0yFoIQIl9FPWPPw74QImj0HEO5OAPwCx6gmL5ox
velghFSfGduvLuOkc9/gvb97d+w7wfkFwsWSxrkF4qjytn+yc91h7g68qFQflbLesMil0MS4yL7V
fK25uH8OO/C+oYftPfsjiB5zfgCfjmuBlVZOJQodmyfNsl875pgkSvxTQirJREOvGqzfCvql9M11
dZK3jCJzsxN1aRVQp3POeRU+PvTk0kjMJbU08Co4ptXYu10VhXddEpD0ckNYyptkXDHpWeGOg0ze
XaGs7uI3EzajyHyBtZIjroqBI4vccB/lvk26tkdXsUrU/pz0XvMeDAxY9GcqES1pGU2MnLgyL2dB
Hca4cj2J3SY6hnMd0zci2hVvIuT/LWSSc6UAhykJtLNA7Q3gfa3EGLafKBKJ0XtN1JG4P2BYRtDc
JNcE42ujoDP3dvXGUrlkk2SUq2/WB/gnUw4ADCgEEJaJ9XtiIS4IpQK8Dpo3+zlcha9GYETVrZYs
9nU0llssx26dilu3+g09+bftdawc1SY8/qoY6xtxY6r8hoUNyjLm/M8uDq7WMtFnbWVsWuggxOQ/
xi/6Ikn3LXyIY+nzGenq6RN6+exaiSQbQuq/oaiLwy0sSzhEUZaRT8YlR4bsZsNSbEpNsGMemKv0
9zhJz8BomtPxl9W2Qs+ESQm8iug/2X8athE5twqaDzFTLFY9sf64KQgm34jmVhLzspHg3pLJFYs8
IJ6l/DudDne3xMHHYcrbZVatm7/YeD4O5O5InOQ7G0nI7vmN4cxuC2HFz3FMfQg86e0GswcPK8uy
67jBojcwlhBtbnXFtNAzafcKca63DByP8eynAng/nzbAdXFbXJCIAKOap93A79LaRPTr1z+BPI3i
nGb+Fi/AZTcIZybxyJF0F2JNJgyjJguMgf7NozDF7IhozIXNOW/EtItdMaC2Z365bjLnia07Sq4Z
PLdHBK6yo1iAH0ztbZ28kB72cnQQtyDzt+xhipodFgS/FwJZJ5hAi5xdVjR7CJSB6SbN8nqgv+Wq
H8dVIBMO/aZzZ9FXmbOrpqz/B0filv4T3fOolDT9UsVzghP9NiyQ2jtcW24X6xDMSs9WA67RdH5z
rp1zVbHWvT/i/npZ4hoCSZsiaoCtPlp8c/HfXnsnZB4zrYwiB+ZFxsCyolJmB6Lhnbu/y1rcCKiN
zRN4VKQsaDCef8PN1hUvhRY8ytdKLGC2XVwk9kaQ5PGzMnwiML7HhXtLg1/Clx3FBfE12KL7KGXh
9SH7gh95nL9FodvbK9HoeDZ/h1z76qvZBUSWGHMpgerd3rzKFsTywm1kOSOWWTrNPneJFeVEvNbh
fbm3iMJ8pfAH6ZJQ9eL/bftL+x1oQOO27Dh+GIQXoU+o4CJ7M041dQk/hFm/0r1Bh1YDqLHR1lup
w+OFys7ORRfDnpcULAwzssfdIS1Qzc/e89EZLIYKS+30sTUhFAaLPQ9aIO3zC/lVPhKX4f/Gdw4R
Sr0wPI7GX24gm1eI6VvrZw25VqO4f7SEfvX4r0ChrqGUskHbGcXh+GuNO6PGI8kGTvSLCN5NWnf5
biH1EaeTC9mIcYGDj1G8NMHwS8sr+TB2LEkFBFanNds6aRGi5+pyySuhKZQo+IucGvrmfXYxe5UV
JyfsNueAo5KrOeJd0+VlHoke30ifItgPlMJnA2CSJRdlAbDbpyXrDjeeWHbPIBGdI5uUOzqhpVnB
ObFr7eSyRyxcAuC5ripHFPXg1h2qp8HQMapysOR5Tm2qAO0V/zfs2eT6JM/KF2rc1sDzwwFHMyc/
icjqkOjGS11XSnQgUfGKWe/H0zsWihyB5oUaw2RKE6TsqrgriINmMvs5FDgZ6OsQdh4XaRM/NgcA
vL8uOatJcVIVSzqtysEXtozWW6BSJ2ZiGZECarDO8LBYT1rgtYWcCM7CAXsYrLTtxY46hS/+mXpi
2bjO1uOqJGTdh7ZtcX6bfHW6rgbuytQq3cOfsZ0RYI7V6CLN/mUn/g+ZZ9FmlFZ0M5OHg5fkrgKS
0b0H3zj0Qva4uwBxl3NIv16/DyGu4XZb9/GzIa/RHWbXodhYqdAtsQPMPsXod9BdSffLfKB/Bds6
Ch+r4vSwkd/JG/QHyrZYZDp7EHddOAd67uIozbjUJlJTFtJbm4ckXGT938Uw7ubv8imsyzIRmKtt
bPsewwYzowv5HWuuU9KaAQk14E9J3P2XoCBLSexQQbyKS2z9D/l7S5bg6mX6/YGRzJY83gJBppY5
X1TIV3VX3RxYR8PVSpSTlzyqADZNhYbIZ0RRGwkxtuWW1oY30P2/bEOu1Bbx/CcVZj0bADifFevV
FDEUBpVBsdeCAO1QxbVLVk9N0YKBG9d/tAb60xXVjU/nzO+UkKUqyX1v5G7xoAOWx9S7c3dJrD4j
8bgeZWYUZv734HmgaEM8Fl/EMoR295xCN5y8CVqrbm56Iq2mrmzNfL9NEczEbT7d01p+hJJOQBSq
PKEckgTJXCUXJ/Rm+wyCKfgPkIt5d1rWaTAiODjqWys4atQC43XIrtMApziNZTQr1VIHpwEnVTQ7
gJ7bbLrmsJgLWir9mTWs+wm+TtsHs42N7El+XElyTRApaHY7zo2hKxeiO23JoeE2jG4gezZn0yPq
5oOX/sKgMlucvhzTmp5ZD32tSmliaVj9i+fjSisTwjXH9A/FQqQlDs+6NMDOPLKcw6oZUyatEwpF
QbTtQCaqXExDyaig5RBrxtE23tbdcsZ8ianbPXLcbWI+mTvJ6CsK87drHvSqyTk2hFyMCS8eh9mO
arS6bkEWfpE10ZwhbtH+mp6izzWhch+9psbJKdxRO/DZO1j8TvhEGp5Yh01L07GMrKhe0/cB4Hiq
UW0eEOJZilaACehBfwvRJOlxMksS0zIyzgj10zpXCkZJGS1AcQiX0ASiBrKHzPVTOHUlbTuFQmQw
HKCR3MNNTWcQBYnG+NTWbnjLjEhLF4YsAVz7eCs0m2OQklSUg7qeGnyba6OmCWIodlm1YUp7kGgT
brJKUHjh0PQo1aUuhGv3w1w/UW04kPh1PmrP4ojo/3Su0HYR2Zn7LicYZHvIWWkUWgdzeEiIkfrs
9sIQNZbP/sP49WKx9DPVX5KK5fc0COLhPKr2O/lemaAMCI9d93idv3g3+4vmT+/WYUuC8PZp1Mub
kuUmt0DuvgQMqwHvAWCHDnVr+qESAI3RC36COXheuhL6txXc6gtP0JeW6J9u3zz0ktyQhEOK+zuh
6+FdmJAcua8Y+RnVNbD84ecz7R4RFzxQZAKI20WqKqRmtWUjvw4A6p50LbBxNrU0EdNqNtT8nIwo
iDGViohcxu0wvsfZiM8kTV2r+4Yb8+XbPkU0zbJP995+9FbWuUCyqKnCP1ZdbmDEpuEdEXyCG7v1
hHgX+lU06A/wL2UyoeKNN2dPXQP4lzqear/IKNDYhlXKL8o4Vqm8jpKA4x9iwaV/D3eQCjqbVzEx
2WRDkh9lSe6FpUI9YJ1vebsCQCB6fmSUugtpkSemINTMtE7R3l6aq9oVpHvu0U/lCBqAi761Gwmu
gGwQ4pRibAIxHWdKEbNAhEY1peQyAk2rtjBfWD8+x3T2fXf0+IYzIVzbHMNGYwtaLJNi5/SkLXfx
r+pUEoAPgQaANe125OHcDBzyfTUb7KbvfoFZeI9BjrSw56mqPQX7QwUR7YcsYJmFWOqN0bFqPjbD
Divw/pb0oQZNqeM+bgWieldOrhvOFz8GKX40OQpAfIDdmMfVrHfr7D7G7RQTCrn59r84WpVZFdRu
jkqrjTBVQDBOjNlMmxJruHCQOMfD5Ck+tx0dNOQzvftkepCR5GY6FaeQVqOM9lMJ/U7lo303+uli
LZlrL+MnM8P4spEZXrPxZkDBDKBryQTUeCMCuiN+XIq1puGOQgB5z2ErA8x1dNveVeg6aWEqV4G6
m7ZMx1/pqg8nEdVwbQ+DYwaj/jlz14GSw/Sm/DdXNdSYgV16jQwQizBAVmqFopjSMRvcpP3vxHsf
WkM87prnv+NMuYj3oN2gnsejY6Mo32OpM8dWGxiXbQh1MnOgryzjzYGpLf4Xo+3yHoPDsySNVKWB
UewTLpU9X3hHPvoiHMmGEKDJGIzhACYtjFrQuT14u1+5TPn0jDYwY6H0kjUec+pnlXrdnqlzDBBN
S7kB9bEPAWICCu4jrak0NcyhqbnwH5jMaV+8IKqNDw3Xsbf/u1zrgqRccbG2QgSK5IMhqem2AKmO
5U71OiJ6E1VM1vBoCS2qkOSaK6gpSOz0tOHLQzRRZ5phrk34t2JcXc2lH6XRn83WOlgdbBTFalLJ
pdRiH+H4jidamBUHkAib7UGfqXcx1ztzegZuz+cj4MEd9LwpL4/5DtFweJt5CtcI/GvkHNjjEqVn
DKK/0qvbKKouInRzCv1lunLfcmc/0oDZ3nll2LfbKJeocYJcCYeDjaAziZyEtK/VlN8L7x/xJvbA
Yrw1iZlgCiuAurqQh1E+dZxT1XbzS/NGBlYntm6GZu3bs8JN3s0exKkBTX9i5Om44u2bqTNu61uA
cgrYpLH35xKw/8UskPEAw15qt5Gzu15tEeOczsn2JHUmGx3+PB4oZsUx/s8xUyFfSPBv2oVGKf1v
5RrZWOUQf6RozUStGxVxwrKKBObJYnaI8ZoH+PG3jyg4QRtyudnaNxR+G7VFHG3jaJS9JsA/f3cf
Wx3CoUgqL5vqGiVWEiO1TgRpHpkQ7lxTJ4Vb5lEFGOSaqqDK5BnqPK6+GSFedxoooLdNbeLkS0Ox
mfJJjN55kj3KMSOJdE8tsZ58rThhr/pT7YBhcF9rcGxLW4DH1uvOKb9dc3mYfE9wcN/C1Btau2MQ
bO0/R9srghHKbMeFzcPLzznMaXOYGXOClc/9fB/6YTzo4r9kvq+8pS4y6/3mXJtPVf9DKcHyQYD0
+27CI9Xj2xfiuWkwlJvTb0o4LLrda8oC2BR/leYLd89TEqKDgLzWcp7J36V1lv7eshuarjJcdv06
uYln0PYp+OQ2G92nzh95SUvjHUiGxCmaHkH7HTUjVx+jRGh36RvaJE9TjmEot5Nnn8znArhzU9Dp
DEaBxJT5GS+ULRjUexI2ubPw8raAFPS29LvJMMVaScuL3CFYguY80c9BGDfooBbpNat4yP1WEB43
XCA+bY1f//NvlkSKp6gecTXjcpIsfXPOFE9lE/ip9/jtESxoOiB9IRFYikH9RYau9ffCew1bxhH1
FvJqa23dm6bTiP3ZQ7xST4wRQqUZQhOAgLxJlO5rsEwBkxS4ITCna5n50INlTicGIUeEsZUJ0nCO
5+UzvN5lmrNk0fnE2XOv7vxD4fgsWifS4F1a6l+Dx/W6UAzsiuV8lXG4JX0Tan4SCRN6JXSMWqNk
AA7QWt594AXdIR0pMDqCzojLxJKqiAUG/e/RDung9Y5uSYZ3dhBJ9qo7Vwegdyj3MeyBO5E0vaqE
wecrKGf72LnYJUXLqNFvTthWU2LbsFIOX2b/XOXY2pw5btrZIREpXU5JYTDCTQFLYYVK6aB0TVLo
QC5V76303JbNrnyFqWImnZQfrR2JXlvHmHHwJIOq3lTNLR3pVuyUXjeFX012k48FBtdWNmInab+j
PUFKpdMjGGZ7zn2CRmN9djqCv7+O3ABMfFRnrs4Z0QlIwLnqbQD5qfVqZQfRi2UUWze5fl2NtAQ4
20J/QEkWIYdGUN5MveEfD9O+Kqx2w7gmkLsFdVET6XdH6bFGsnvs7gxukHTEmkQo3Js0D7E92Zma
1gWIFn4on2dTtyPiK2Bhu4a1qKS3xMsWBPNCvceQ1cX88WZsUoqjzX1QpEsUS+H3nKSFh8lINUoE
9nYdIc4wiEoIQ7cQUWMMJIBiNO54WsGzwgLaC8lV4XlZl0aN3mdjZ1jO4p2SUU18Px57FZ1dkGmJ
nWyftFMk4+m8gX6q6BmX/FEqAyWNyG2P+dZSmKobkwv3mPcOKluEwo6d4u3fgsp2jVOu606X8Bi2
v0LpeDdm+B0deHAKaI/u3wugNBvIaaZYo97IQl8biGkzBSJ1Zh/i5E/9Tyv2xJKJaBkzpqQnbZkW
4h8QKjsT1zvj60kKiIGcjLEBaRYCGSrW8Qr2Aanhke+6L6Emws3ZZVDnqplyFp69PUh651AWqQ2Q
H4U+Q0gLJMoH5TAz0Uy+uC0qKNsJVoPd0CFPY+KgJCoXSIgBG3qeWpLiXIWGWxgk7NXfnpGCLoue
DozlN7mTWDg2Pv+IeZ6UsHXYkTf0K9so5pn6gfF5yOYtfDaxpcvKmjdk90kDAwt5G+zgwC4OT69i
sYhJhDAXAjt5bgbxpVUGksS62RJlLTvjsJg6v2pxnOJQFRlWnJ59Dth4B8TcgqcJrYsUluvK3x/V
2/S/k4wjqniTlU1yGgBWCRT4E4uQBzGLCI1eK2fyIyyoOg5skkLg1IWLPXlDj3UN92V0ZOIFFR7/
Sz23CtRryf2qjdY3/JLVgRRr6kuwO3urFwF7fOBbS6+yjSLw7JjfibdBsQ4KeCfhXwMH8PuJ+XQG
ieyMXqYt0UJFduaCwuiviA+wEqMAWE6u73vO6AmShlHDFlTHpXthrtiI9FBDrBTrQclnwSbDZ/wZ
hkiw2BGFs573D7HGAZO/vpTWImV+jLkJdKrZ1e6aON8YAbnLlz9FUldjB7YmBkTdheHJI1PZ0gUA
p5pjboBNyBkl1d6L0KK+Xd8bU9uCCoA2CXLrq0RRiEAhW7PGItrgtbTDRU2nBe3UhNUn5wR58fNG
kKJGgBXYLBR0Ok9D0rKlLDnzb2o2yg3yUmf7hGtpVBQwhmRNv307flgBeK50+hDypIfhFOBnItUr
iw7zhT93MhU4+up0h+1BC1vlZyKFlCevKAxP3mVztqWU+lBL7qqdeRlkeyMYKdhj2U3+B1qub1q1
O8cvxgqC7ESuvVMs4bZGq/3aMqn/Gpr9B6y9swymkstpoqzqH+nztcXgAB/74h5f2tMHIjNLcaw6
3/mwikL/V44J/oyvX5pb+aB7GbdIwS8PYJHD5uZ9+4fqIb04I+eJQHagr1xs2WChJ9QdEJLaz7HF
AxnVkG0whuGM5JQIAOKkrqmrjSRSyfl0SRcatuIskeCS3Qdj8oAY51Aw/J5mnzQmdv0I4n5qfaPN
FWJXw2BDr3hM2NYJDeBrXAhDNybm+6rzwS6sfHQnvtqpBeSBRAmtb6VS36mJn2oJ8BMRrlwDKLM2
6ksUP4qTyBqaY1yVCZWPnZ9MVR9q0eNFLoVVsbOQHWiu3xTUOCBFifsaIqDlI8jR4QYOfc7Vq2Mu
jiVZT82McwABMSgVxZlTwxjpYCJLqyyDiupHrFRUi8K9RuHLw8y9oBRwlrnv7gEAJW2dtM9oOsJw
5NCIeSiFZYYmH+U9M7qMmNS/iX98bKriax6a8mUpQUXzjWNVbWi2pFUlnzDVcLJ5FVIe5Av4luhF
dn8Ym1BQZKKjGmGjA1msKlItYCJGGPCzxo/Qzeb+x6jIJsaJqrURXGM+xl5gHRib4u9/i/I0eyZ8
Sp6ntlcp5BETQqaDM9knRHgOD6mxL/ng8PxgQHCTH514lQuGvzaFajm2hlzTfHZJ7BhyCwMQMFUS
PR+Bw7biEHFKyR7P/U90pS6csb6GEV90hj5kaqtSfQqgPOeYS1AbggqrWvR5boKejdd3SMbwMcQI
W1WDhkyX6+1ybgYe51fN233KUrgmGu3yT21TDUiBEltymcyTVovKivXXUi+6EZcmSkwXpNLI9a6/
NEi/4sYqFubRzQvjDp2O/XGgY3HF+ex2YyFOvHHeOg78EL9OKso9gsc5rM+w5TRRUVrh5aeu0dfS
fpeOkmAEAOnIb9rzTagsqiyqI3eEaJcaux/LyD3eY0vjKZ7U/LernW1UxGPZN9hfwpf70seNTEW0
y1C17tKE82QKkNvhUY06dz4zp1YMpvGetd6kducuvWctSw8N8TOeWq7ANT8/+2RuAXgXKHYVza2N
WIJo1U6iWESdOzI9jradcH2D8HaBU571dYQ30K0sYkLCVr/z5h5yRzqvhLrddPQg7jEr0wy+QJKu
GPke/BpjbF8mKLS6iri2C3GgRKzV9Gg22sQpLH/pdjyC2rYvRcIfx9UnnZI/ncoOmtI11fsU+hMJ
UMipvDZGFxSg+knCWYBiiF+JXlwMwGyxHbXFVH3NHOZvW/GIF5lxqOuEdcMw+C01DNB8yQ61UV0q
n7bevkxHO943aYFRNHakqvsgIND/uRtxuH7xcySD8oQIZ23FI2Eh7rZzS7SbK28yzgmm/Q1Y8Tho
aJZimeoxb47it9YQm/KnTJhfeV3YPtJiv9p2lPPgnr1XP1CFkJ0JBWWayzJyCptX4MTRofEhi5h9
BbqNnpjVVwegV42XZ1IDgL4z2wOp3+05Q3TdZZieOhM6bHpvQqyfqj+o95VBeUwTgx36SsB4MRXn
AsgQdZrFne3VMAxlSbcdfJKL545n1ZkH+BiYCQadjRJl9Yvd22nPQevllcdk2H1eZdJx03W+yA3g
OWWUVO7fn7I2rG/BEo/Z3vLysE7tE6lhRx5RJbAOSxj53UwzUkqKoPvQ/V513SqJhgwBzoXhzKO8
0tcmKg+tuUBg2fFyz48EQvH/Vjdg0FCjlrqITwMPGsRFP6ZvVvSjsq2NoFrYo2apxL4z+4DvQK2O
hc4VmITcy8cRnTHncCFDWtYOMSN0KOrlgpj9Thui0xRuzu9FNcU1naXbwbMT3LhXAAsEBTQ1DCCK
6FFjFLsNtVJaNRh3tJ4Ryy17f0Tv0QJhCf/pea2aio5kEcMciVet3AV7imsZSiafMe4e9aKOU14E
+ZfcCdXvJyIyE0NoFKgHkK6vmWWsxFG49yiKYCwJCYiXsQoXAuzREKp+mnixzJOtNfRo19dvJ4Yo
FzfN627pujZwIYuPe1Zs3warvE801y/nrga0kJmpaLQvsQkMZVSR9luXGirtOJwUBWCm2rGt7q1A
MKCC77uBQNvQtcAErva1kQ4dQSp77giDausyBpRi69VzUgA5iLFHuFdvauMal8JssHNMDJG30vEj
7XCedI+AXgSvR1q0jNSa7J1av4oaj+d+tT58heSEBzosMC2e1bwLT+ZAFYQfHDxkkd1qLgZhP7cv
N54QKP4NAAojdloQrb4uuZ7bdHg6cpCNZfhGwwuJcgDLS94SA1DDiMVqXQhbwC/Pue8X6EtBlEbn
qzW/Z8TfpBEQB+WJpDsLRcJWjXogplj49UY428tzGOhFoF/p8/2uIzluGGLXwXVIMFtYL4wwpJTT
nhFrp2E18Id5mVBjrPbU0BwXZ5m7yax9+Evy/uer+fXswgxWUN+RdEmmvqIyAlcef/tSvbrIlnS/
xBxAfr7JTMb2IjyNqIg3/10WSI7b0pBpIqM7l5qSdva8O1G2+eU733XU7NseV+8gDzHT/+2AsHsC
1SakoVHqR+8f66BkMbK1E6Os6EnYHmEZ3V8Ldezvx1hLTzyfSJxo/zowvHMYs+MbQg21JrqRNnOU
+qmgEChbrR3D1E2LJ0A95P2i1UyNABDkUWOQ4aYApxXLxLppK7wQCQDMr40LfamImtRxsbVBvpu/
8ijBK83c7DonkqRe0+GfRlSIHYtcfuCMMejnuCtS05uQyVGD1i9JBwReDJOuo7MMd64k6cIuk0Mt
URx0AvK7P6AvZUsMxcknBhoPNbkHnrTkhsZLXgnywuzFVoiWuFG5XEvEd6Ik6y3PcXxeXHgI+JIp
9wDn/uzy69UGyADjMUe0PM2wFJr0c7xyLjEFbukAjY9kJYSrIfHNjRE4mH43TNDNj9SDpArHn4+0
ReVv/t7IIW1KadOqtTb6Uetz0+OYA19rV2MbkiK0Nv3AHwHzCzzJFWmn9hMQsHGsTOMseJS3yUva
TwmcrAAlCOWkB/YocKy8mQI/IcqDXynDgbdDRSAyOk7WaMxTEV9n3Yd2UsgCuWots32MwhhYgEuT
nfPEeidl2zhCl3MhKyuoJo0NrYLQvnMpuMM2d4WnaxbKTFXndX26kZpd6k3wpYZE+FLCOmw6oMqq
ej3gq/9CGCSEDm7RVHYGUE/i55ztseRQPzTvtIaf/s9ss/o/ZqCZxaC2CpY0ELUbXX6PGfzZFEb7
r++wPcV2r9HafDyzy0opNMjpDqhv+C48q3fC8SnewM1ppea5AM+DMwIzEbJyDShX12fXHiwsNorF
DQ46ITYThxNrnU0R4zg8fG+Lx+NrK7vZEgh301LdBjx4/sJqXqbd1npnfnx/zlvaBUVjq3o34Mwk
tUqP7nAQarjwIPcjdPSovXl1H0jxqYQ44eVXu3Fp0Jc0E8SB6+oTFmnMwohpbAw/fRpkIWxdT/Zm
Stzs+fNn4DoevoLZkHPe1CZpSDkApXh+62hWN7vwsexLMV/UnS09hzuJCzfTNSfOB1z7cHxKG3xA
FblEyAD6GxL5CQImGLnNRm8QQG/wYDPupb4pTB+pomrU1t9ij4eYSzRklTz7M2q4+JX+qWoO1ZYp
sMKisMNRPyeOUm+lOoAtcUQHQgxbqAneBJxGQbi3SRugg8ZqAJnNv0hlA3Yr/ZEPc3vw0s4uEOgW
nplCPwwTyK+orFh7WQ5szbtgvCm6SA4+w4M2ZSWQCFPsSO25US7X7YhcsniMV6ESiH3ucbSZnlS5
MXFVmFKAp27crA3H+Lm4ck9i5pOzyUd8jZttq+CcX0NIN0casHS0LytAKLeCE0ptYkmfGFxC5u5z
RFvzRW2zXo4N8VUjb7UZSWPbHCAqEYeHJzONL5g6d/+mggp8Bw7NABpzdlPNV/XfsmlW0xGF+6oh
x7RM4IrsiZKc8ciUvD9gnbczNwl+K6FqWe6RebASWeOauiJHdWhQ5D0CJH+/GA37LDr69PEBPhWA
R6jDxsWEDdNigxU036XbWzWaVx6ZeMtVzNhBeDZDpDX9dgUV90ZMAGWkpFz+UUrKGPhXg6g1UQEf
2RSu/PvQfsCoY/XbV8Zna+Nngu1/+1uq868v1hDgky0hse9sFHNZsI6C51D0xWqQGkW+9zbFEIAO
t3brVMI2sRc6/toGG7REm0HKU04D2TpcxHlLNKlMDx7bUhGZhjOl7gmoZhD42mMEBVOAA2H6ZUvz
AjylltjVsznf4Rnv98LEACYi2sMb+XiLEkR50ryb64n5OSsoUwXC5GUWuOvhxyqZt7zgOf4Yew/N
f54m8Lz71T7zcA1BDqAufOFGKSs1oQvKibDJJCawGBKwwmT4DDt0B85RmdDxnxr+w2Gaef02xlJt
3wNuNCg43hifMOFMsp3g/BU/1jqKxr1NTplmFEDuetDpI6wG0DAKzMBclDsrN1urTIx1CzYDdyrq
061GotdNfVlJ1nnMA1W7mavWS52faGvnYu1ajZIq9h78BojLOqxvH58IR97vPzXRCEU/95c93hOh
DK51JwTb4tWuieRCA5CWt+G9xKU8JQn5t4hSPfkH61vesC2uDVQjf8I6CPLK68N2iPqVcLHHxAlZ
PMboZBWWF/sxrS9fa6KbupprWoKsZTWb7Vb3d34Khuy6uZ/AcfFLVWmSJrIrTS6WT2hjpo1HECRY
SeAS9EGoutCuhGHJLOsnY0OhbdU0IzT8KztU25Ee1MftoknRMscMNLznP6+OP0JtKz6lMrC64E9/
GjLQrpcGTdSsiew73D1XI22x9Ij09NKl5X7GCKQ8lZehUiICzpPCwYktEIaHdMSZOUKP/1A7qN0y
zSHIZVE3PD0CUSJLTbxX34WVpvnkvUcYEwfpZN4uZW647TbPW26pyYVjv3aHdxCuUb+Gj8bCgcWB
ocvnMQNxBOXNgOVqTAGjBQcXCbSvgEHfABFL1YXSppCHcJgmhha/ItoEv3Cu/Vip+RGBOWchrFQR
/WuCzs3TuJldI2qMC/r7/fRNWy6BKM6kQZrPrCW1hZrzQAzVsY0W1BFu/y3L5/5U194cNZJ61hIJ
9rjJcwyLN0VrEXRyY5bvxyloIfL52nV0QmJ6yWSWRPUW0qtVTCw7ajJ0L9d8npDhmPVN1htfWxqZ
cJXcpSUM4sFNPJo/5FOJwn0fi9alr4ScWb0XAShHjBpE6ytWCiEa8pdwNS7k4cVJU4PuXKYpO/QQ
7nxEL20l4Coj6qRN1ll2m1bBkSFd5bg7by+SHZBG+h/nDAkOxHB6ImqWroUKMzRUprxoF/Xi6/7N
7VlGuKLjF8CKsnW6CPOBNlCfPu1/rW8otwvEcRs+WjpPLMd0NbZnPjG4wiXqNI2/6oqo1KH39Vlt
HfIZIUGw7Ux9iSXekJkHozofK5ZCWXcJUeUYmaE88q0sozl5j4YXMGc0fw0sBdF9q+ogtL/+BSw6
jAGcm8pGjIaqFixdEVLfvlFvLFIcnj2Spb90vQTI1SYU2nXhhKiudaxHfbjt4bkAhveNzZapkSXQ
7YsVRltrndkoYIRLkjE7tzJXNsroH3MW2cKLDaTprHpr+p7MbgAROF1yVEShG4cxffq2aChKpYPT
ga7sBOMwiCHF9JO1k17WLgnvzWn8DQ1ig+JEmPQu9XxJtGEb7E77P13nUjUmAN6wgPm2phDMzuby
NKOdCQkY0bGFsLpYPkProvw0Aedu5LQSzrjqwZ7NTUoaZ5LyLC/7uZsYavg7mMVsNb31sc50m4MB
pcgNJPt55OIXHM2UH0wPAKmSi2kl/7jhC6Su0JH7hqnIG6loQ1nJUUNjQtKkTjv1VqfcFsLBlv7r
Sw4fUITsf1hCuJJMjMGmK4XzU1vhQPGTxodXsFv5v7Tu0W248J+hcwqBqzXSsfat3n3ipUzpDmXh
s8SO7iPyWRnTQkOEGxyz8Sbn2tjSnPTg2nsrxKclpkG3BHe94/DXH1D7eH9HcmuBmnw3/WvN+h0u
JOBPMl1Kzw/1PKLig9uUMzasF59Tw8M5mtSVk6W56+UvVS+6LhBVwtzMye/UKxGXG7Lz7Z088W+p
6veFxUK5eB7AoUzp0/nZnJS0oXxqZ/SDFRgHyOVnDEUYW9oC61Y6gSvjayzXQaH+twlTDg/NL/QZ
g2Zmqb4MYvVwTz68NXDvs+eR5zaGltVfDktQsEvpoJF0PhIdfKF4B9qgUYe/JTf1mLvMAlpaq9bg
dp6kXdKnhIQi7vzqaw/+FYHWp5NWICOslOBxgWnsuLh0IWKX6oOgjGySVmKtEQKDHFdgbDqTu4dJ
+VTs/8slaqYSL/vLesW8vIX1lQW87KlxqFnR6PjvEY6IG1/FQqWRUEBklaN+Be/mowOz3SyiD/v9
uZl4I5PLKYZ9jN9wX0OZx/FFIYfzVaQgfysP4Tbjj6nSd55t3B+que9JoBiZEsYLTP5ClafUZfHq
7/ppPO4gPc2g3E2PZJqA7E97Jbta7NjEoJ3YTcMNPmGlOPgL2V+IbF0SKQW2DjBcyajGV2aLwdcc
nuB1Wi29tY/F/nTc9F/fOpZf9PekjhNyxto6OSYLx1GnSurb71Xfbt6Z6oLRRcX7x+M2l0XnJvI8
c4B/ezqvwMxIGZqbkd94dGDcJ6oG/Lp9IZu8rAYScKjyCvvHtvxdSllrIbVdbi1DE/bkziO/MS8t
8GBcQTyiv1HzSrDpGE9683eSf3Zvlaw5VmDHvtw70UE17AIKjcZrGEB/MTRpMSB1HlIiSk0+Wf1H
uHrqOsnZvlAQEqoQOj/CDnJW6D7yWYHzn2v49MeK6jLZLNZMCylab7euOcgdQimI5puwAKlx2L8j
a+8EPXNWkfEaDj2c9caS6H69RZ04KauOME29N/6Mm2zzPBj5y0bT5p+HqRgQQpXkWdHP3rBfD0Nd
rmzspHYj39/OqeOIh1Lgm8ueP+/o4czDm58ErVEpbu3hNqA6vn8JGfMYphQfQWPCf8VZMPPsqvY+
ysI3+aJOM7uTLtIgAspT3rEIQqNbtKe3LyjjgiVK06EpvpRrF58u1+gLnjXl7hN2s/uhAW46B+kz
cHaWC3uuhOIQwb4HNG1pmMPUuBjaJuK0zkpYynpTrOKh2XxGCkg4igrSiMD6+Z5g8BmxOEXYdlMn
A1yRSLSdpNr9Lt8ifesVNWtpFWkzBVLdcM6ArCMG/6KZv05QNkZVAcFJz8PaiWPLZ5y/JxF4askz
G3v3DsVZ6oKcEoQVagl8WpeLp4zq7/ymB518HhO2CzlTqdnUB7eTIptJv1Pf5kHIru6t1iYl3ZUG
2me6B8duqYIXUCd7xV9ig3C+t6knGpriREJu7G0Xp1ONbueys3Te81O/cV9bJ9tls2kgbnLmvMNy
KQ5MgvQubAImU4NVaAIYRy18O9FbG171geCqbosMtvAbBiPLFWe4LIMgaRBrdP+GGVeVCXQ4ZQmt
niwTGUk7L1eFJRPciyQaVE8wfNx+Hrz03Or1VDBA0pzZMcAqITQ1lAJoteRB9RNRVxfbN7E04M1N
xx+2wrUn0Yy+TSUYGOp4A4WaItlCIvy11C0KrGc6prqKqSuPHrkw+tfGoWkD7X2lLcfUWCpqit9M
ccl4J75XyU4uDy3uxRiO2iGa37wogZDFs3eV71DGTNwYrPuDjlpyrZIWi3W6q1nzChhpMWWIfEpE
Gb1VxcRKUllhrzAhE9hxFOTMNF4VXI5CO9KjIjURGt6GIvZkgq5NNgAUG2oc0mfxCXP35LycDVZ7
Su1aZBEc2MP8RSib9fwzFJKRbGfC43mV41ghuBvwpJ3NBp75isN2bocdEXqAQIY+t5dDMIQ49FWR
EW+4Blnr3ks1lXUhhOnUpsaKgvJBfClO/6yeN1UEEYpL6+oX8X+teKDLyVrYZcAf45E9GguWsdXk
nc45Jlpat1QrAfa50GhmPCM434xyhHqK1Av9XEFFfDRNl69m+miPv1oZPNHEzjZVn2hUiTCjvkm3
rFaMTgroE782AbGXWKwbXET1WebkexdQE2ch0TYAwdRJSx4Lrfbylhj4pXTLrF2GoVv05qwRPCvX
G+DDdft9FNaQebqTgayw4ynmtLbk97solEwu7H2I6Z7anclPolA7AR98WMXs/4iL016zzSoZUwHq
Kk2SF+gaN2hYrkWfAtE5JPZ/zLSh+JKO/OklVA3WGFq0ffqAI/fT7OP8O1ncr2pE9wXRhACiwBno
+qWGjK5ROnsV4sveDXHLIPFYEaUhxH3+H0XRC8APJv/z7H1zRTH6j6dXkBJkgKw304lK7qq52Nnw
QvMGCyKlQdUnNqOU1z8NuL1AKwPdJTx3jqz7F/pCpY8p4nEZW0lehwjA2WUjCRHWqXX65AZiqoRS
lM6CSRR+5T3C9S+PaxtAmOt5uNH2hN4y1kXhckBVf0VGebSexSRsYVTQMXJddTTIJDQpr5raO6VX
QhUn81mf0X+RI+sm6aWraEx3nPII9Bu7OIyY0G3XWtLVZrBPg4eDvmYQFtgoOthqRvIzFhO8TOmr
YWfVfLzBA93lQOYSNxqxRm2ZzxvNhTZ9SBVcZssaNkWaWfcx/pM1VwP2yaie5m9zxC3kh1aFW2E8
vlv4WXmyAkFSP5JErYD/meyUQ+tPLhtP9rvJkDg/vYmEf++Sw37hxWH6QawA/WHxPkBHKyRk9v/c
L12Ee+0CeJcjv3MctsD4HaZX1AwoBcpvaneI+fM+iZJ11aIwq933In5EtgaIP8jA3zkP334QK/Eb
RmvwCg2Dwb7KWRl5CvN3JrOdga4ZXrHjBX+jnQuAtFa1iDF0EUF0lxXZOIhIk3As7KOTvvXfFsOC
JTQ/qFjYybn8+x0oHSqPiACx/cqKPLERTdbG3MtgS3O8sohfgmv5XMc+RM2yWqVuZOQhXSle/UBa
YxV+q5eWxU6Ankv7e9pxZ1u+0N1FDKwTYpIoWvsxcG1hpHL6DuLFHVyLIw8LqA0QDU569LQjxaRP
oqBOIjlNPiX3iehlKUT6aRxF5Lu+7HU1JRBCE997sdAzu+RhQ5AwtmNM1/1TB7ruLyAjr9vJKDvs
iauVzuX8l5ZVpcIiyCIDFLukKEKCAaVBUtFJDCwdNJM5bYTxsZoClMaOCN24NmWRQMjY0WXahjPH
zH15BrMeLnft55Tw9xrIq7elJaJtP3po33YjiRQzibLnC/IlBKC+eZqdsKhj6pEEwSpo4AnyyEiS
QIWMGOYOJgOp5wahc23chC6A0kh/eY/031pFnqAx4Sf0jiCXgX+29WoWMP9bYKDerpzL257p84ig
evBix9PSeq9bJf1I8tT0lVlrhgpqs/ifqB2VM7xz2KdrZFJ436XfDIRlJY+WawSeVP3DsxFRZB+j
qUOjfmz5s9eEFurbq+H1/XwIcwHnetzWNJLJHqnVVJ6shgkzl4mNzieoDtKPpB96hLXruEXz2TgR
x9AwHe1+Mzj46Xuvo8qa7SInnkd7EeALuwYlqByuyvwLRJht6a7wbxdOi7hnR3hW8TZR0IHAJFb+
xqr3nJxcT850FRq6uAS/zZCeL/jj1M5ppM3jCmah/ZPYfomoi98LFVdgFiAlmSo7GspCNC620393
Fj1bmiBszQ1WdCDcnn4KeqiAUZbYaKMKo5cNysEpw1WBUh+omLMu3zZUyRkTJke+yC/dRM7nSKHO
tJ7rT0FftB/z0L+Ngj6RsCaNs96TEEnYuljdjGatrT/5ClgmG4znBn6zAuO/NQQlAm7hcHIZJBpI
jXNAHdQcJjdtokiH6Fh7tNbIQz7NxSKPMv+rM9HL5nxfYudMaKm9tGh7mO6nWPmI/7Mxd4WP6DLU
jVY7aNGT3AekwUrVvynVAizvDA94OTfI6hXEUQb5xF6pkLCCx1vSqUcYI34A6tx9SxD/wJNIS1Ir
sE9dE+/JwnPvsFlEr0f6CVIbbY7kr5zCQiY03WtgM89hs2FuO98FoKk7sgfJaT1x5Rc1aDj1Jpqp
bMauVBvee9s8miOHBfV2xjP/bqrFJ9eRfCtu8v/Hm3A+84ltqJaxq6k600CqviEGJsJFCDZC94az
NnwQAcy/HrwfLSNjtMo4+/cfDIpmOatdwPrjiEWluynfGtJ/1iCFn4MoZaM9dmd2Oi81qh0B/fEg
soNqLwxobXvmEE3PVbvxK/guYZch3gAeh/Z+6CJd6WYSX4/aVsCvrHnID6TMV/KH2npSFh3tdrnD
Oi3mFUw8/irG2pZssjvd0hh3L0QWbydOUS7vFqW/W01Z1YskNUpGhjNzbVYZZ2rB2NPZOQBaWuze
VkLZQj2NFLWz3sjY38Js6QFbasBMpiHBbaAMcbtbic8SNL2bs1FZ49+TVR1jUDfXYnztMLVVSFU7
VASdyvwxJ6tBwdqn0k3rZIP5BL81uBFpNl3wMIWRPFCLOvwY6FKnBxrvsn0HsWxYfbQ2eSWjmdSD
Pv5BVvms5d9I9dMgp4oyrnYIwtWHDalMlbXxpdc+B+T9x79nsaSql5x5PCLOvOsJqvLZgp1/DcYt
0+dVFIt4RO1bjfGW0byL3dg4Pndicu/Ls4qag9qWn1vYR+SlWnAjY8CnrWbYxfWtGZPNqOk2tdtg
HuhGEsr6TgGgmMsnGH1NYX+0EijDL6IgL4Z7guzBwVVH3j6QpOlWkPceLJBLsb3HPMupnlvj77wa
z0Xp0SRqSx+g1PhCw7qVOQX6EQLLKf/6VQfesreF/teAO5Pdq/qIl2Vh2CsXOKv8rMV+HBuaIG01
/34jV3fqqoGZtao2tTpFhA3kowB6jUkBYDi0L4MerFINfzNQ6y4houIc3Lq9R94mwFwBtYNsQHWn
3ggwhUOyo0pSriDYEUbummo/Rgdbv326AcJQ+WtwU9MsyiRZ5Ax56g3R8FBThhq80Iw3Z1sbNVwP
9qnq2VvCJwDCYXYez1/sTiBaz4RF7FYJmQ9N/tf56ANgaJwHNAxsBFQYSGx0TFjOb2B7+W/ttWsD
43KqqQ5Ix6qbD8Hm7+f3s6qOMO3kw94eDJ5Tytm5y4db60SGZNV377iI8jEcMqrTaRbLNbCaLz5p
oQS8nr+t+HE3tyZuAdDyMp4bgg/1zFAPrmGLkHw0S1QW1cxD16JIXhywC3GH6uHDPSK8ULciDDzZ
6uHZJUC12HFau4ymGPJG0nUX/uQlJyVJkyaA7Fs9oZPw1uHb6XZ49YE5v92Gzx6yNZyZRFrXtUcn
0+J0M8aaP70dNImeiuyVESxAOhGzjD1CXuViNp+tll+ilePCl4Bb9XuOGJV3EiBsXVyebezHIUwX
1ATmxMcvJQrUgTiN3lncr9GUCVlUfq6m5ji/mondpk9tlThkflesuXyM9t2LrMHHhes59A3DXIHh
o4mHbOgW1EalQiR5FYy6tE2EUYi0KjFg0Tp3EZVdYxgG1ocCPOIfC9wrD8HjPQxxsFfHa7sNrKK6
hnekS/HPPqnel5WG1RC+p6AS3m7bvJFM+DnTkuJ+I9f4KS0/YQkKA/HmAo8m7a6y18socjEXVkZq
i4+XQbFtIQ0VHldfw2GatcJbvCCONPbTLkQTQhE9WQZtivlehl9ecXoQQXrA4HjQikfcDcJU1c7L
0/TYwFfIfE/G1SKofqKZ1Vy5HOeW1VCU2UhtrbWK2xrEugaeSP3n8yFETte7Oo3ASRAgUpqIaZL3
H9wFc8mB/GAvzrKv6ez0vTKtxcpnu4m3ZeC0aXA69dAYQuYJBmtLZdrQlaTxnpqhY6edtZgGQ432
ZHid+wUpTOaPWdrNK424B3+vBrdjEbyogAZ16Fy2ICwYNyJLskmqMLWvHdAKpqSk7HyCyhk2JnFQ
775xHvLdnMsfZSnKKq8FWXwJD3ob9BjVaId6fFGECEFsyv+iD8EaK7sRq+O6H47BqsLVigmnOwsc
x7yzioiP8Al/SNGLMWHs1XQCIrKhEzuOZiziEvuFpMnLou3qwfmdcEbAnhel8c9l/uYx8Z0T1A58
tsPgBrRhizb15rL9bwW/jS4XjVHGOap45/5sLFGYZFohZ4tkRsjCa1fCNM0042PkMX2uZy5t2VgG
cwmLtjGdTboOJxWt6I/TSc4q2Gw3Ok4D3PR27PLX/e+YLK+xqXwAq5GiW6XwkDbKRsoKxThDRdfw
A7oL3DCnYrI9pJzA+XL/FesXXsiKcD6c3xPC8SSyj+8ffCeYUs/LgUfIy+y1ttJ2Xy07iSQXDodP
hXLlebJl2viM944K07JO6za40OiZx0tPxP6UO0OTULU5npnBg8FlQbnXDjsG+NuQRopDcw+QeXB0
hMd9dG162jlIHfCCFw9x9wBSXHbtxScljpxNpdLG66xjTcm16T/vmF0KIh1u5hg8UMkK45yh97aL
gih8CiWYsBmuSRTAQrFSkVVIISh+F2yaLNDxjhMp+vIXlSUTwecmwPgeSeN0yqEobjbEptxkHqEW
/w95hj1behIjWso7UYpJgR7G243EFIoRtgpps7By3q0VoWiwSh7F7Cxbj/8wjtp4tOwd4Vutnkxf
GusHE4IeCmQy9YoBPnFPVhwM09Me8HEampdiqhIuRmfhwXJ0fZyfyxe3vVI90daIMeHwpCv6aErM
oefeRCl7KhAS1mF35pC2QH2XGQscc1uj5YxSDg7US4PV5KNKOhqqYyOnkLqz9/syNV2Q63HWtyGG
7JD8EdtnDPZQXe8a36RF/jyvg0+PX0utV4MNk2kGpGAN5AUWi1RmvOyrBRhqJiAjlvyxXLEftk6B
fvHylP93LflGq4jzx2PjFmsFnP2awjpAUC96ifPCNRsZcP4ugLwdm8UFrLlDGryzLf4iMCNEqsas
K3gqHnFR1t765XvyIvkRWpmcLH4U3Wrm1Eixwjauxtd1H3Bpi9hX7RF/VsoNKYL8uDekQm7dt0Ue
DtNIzrsLehih5uOVeZGcvMGmX3LULs+1DYRMWn/VFXk2KMiJwl6jSPdeZ+GJIRw8z5f8KLZqaHZG
9jnrMF112dysiB7MY8rNhHMMfc6D4+GDGwmTyDz6Dq4s1vCk/BrHUeGG7IhCcjD9pTI5+rV7RvpI
gej1uuPoYryoPTmOckA9wPCV8NPqByOWmVMrDDwKJZRAMCx77DoJSTBAOYaoQRPJ8FuPWLOgZ7xO
xPwcwgnYGDZCu2EnbtB7zTEoFD66gi7aI4CtLRIXzpTqXW/yg6REDhaVixHjD6O0j/7Vr/3RVykc
j06XJlJhz1KmJBj78K2Tk5B0K3MJmwo/fzJjYAtpa6J19iH9XqXfILiVMQM8jVlcAJy9a9KpJvzR
dwf/EV4BiZbEQYtJD1aRgxMWOvM/YXjuYKHquMlTRbk7GaKec4MaAWHmTKEc9PQWmQZxRftXgvCt
my0KBVLhCPMl3LD5Swr27uY09sJ5pCHECb1rcekKDnJ9eXW2AGFzirAWcgRik3cdOHpu7m3cJWPm
he1SI/vRNz/L2zOnpSOu7rFVe18SqqWRXVPKNgls++tGGVDOzQ3VjZEL1E6die1n2Ankwj1QYoNG
jrK5DhjA1171NlEo4Yj2sz/43iY7yTQZU2dJfmIFSvE+Kndh9dgbjrBRAIMiN2NShKd0l+gXpsGs
S6O5YcsxNG1CXW/yVPILByUfwWYTJqni0Ni4HmJ5sB2E+XZqfo//EWVEvPsfFmuEvvJQGZ4ciIkb
3dBpWvPnqFgn5ifgi+yoAP6EqjF8e9ygNGIBCjziJzrLT3lJ0za3jLyWLWJ6r8Fid9oDHYd2bFKE
Ac1u+3Dki9mddmMhy8Lqks4M32SvxEKXfUu/q79GUwalQNywfvDA5Tnaf0uyf5nVjUdj8wH+fp4E
nAVEVgM43xJkTGMHtlBKyxSxjng65rFzXJbM7p2boa5pD8006kYJZu82Pm1YF33O9AKgcvp0l6VN
0eGEK9/lcTBcBZwq2Me+g7PUUlIJ+lgF/O030YNwU/PDG+MgXdU8Zf3drD1rgniXN0RqNttGagvD
do5XsF3gu0UHuWhJq+x9HyKkWAk3zWl7haNZITfkv05FXqKVwDKTyS9XIqqbk73lwJWvHzydHOOm
WUu8xgEIZ4pyp6ImTyIwNSdLzTjFp1qXj/4cTwKDbJcDuDmN7zMLAe2+ATryCO+qNFVNzIpx3/vf
l1LEpLC+CyY5nOB1zh4eSh7jM8dWfU4G8xNb1PNGYRTel+qhoXSaLftzCa6L2+GaAzbGdFYmrank
rdScMfrvy9PZp9LBnUVWEv/+bFTImAZLvPWcqCe4Mo5W0p6N3lWWJeFdjfGFtnEESrwgeWa0OUe/
BunNh27dVsPkXdbRbUk1sfgExnjAs5gQ5Q6MCNCOO8gMQ4gCncXQ/y9H5QaFYaiQ2zsaxNuR9rg0
SWC81sEocChPgJf7LCK8pzlrWq/85ajkT74v7VX+lY9cDlv92BIxqDmmsRXSzAmySVD7SqxrKfwc
lq9WuRlFLYEOXaHsAxuG+Wr3TWsReCXpnMi00OCuTKs9fmA2w5SRag0OmdPP6+v9Gh/Hf8XgRhSU
kjuW91P2l5Ihr8LP3ZoocVu9N8HOV0QPVHyheJZ8Db+gLtFx1Uz8QhQ9yJ7qjRLaUI8/wYG+3dT0
GhOabu9U4re7fCn8RUkKclMdecPO+Kg5QC/iO7dSQIIt3R5/GhW31VbFrio+2FNHPLefqV436yAj
QCDDX0ziGPlWvMZx3RqzFCVAu4pMxxVMHGH12JQlMKRy/O9/tuZw/SMQHENObp5Rool9mcDiOuOe
YhWSvSPQusi29/EaDbgG737JPx8euhmR3YQ7fMK9P8nGMcxZB6JuNtTIE9QCbCq0EMaJM/YqEffe
WV/aJAtla85IipX/cO8JDZdP2F2Ol+x5imhq5j5p3clqLW746TH4/OH7omB4+V+i4kG38/A3IlH0
ERgDvmqrZS99+63uDZMPSyMjIJNaot/ebAw9QL3Lzh4LS44uQX6IRwfv/9agChHyqjyhePsWxsAw
w7tqb7jc9A72oKxxUMkcbk1KksdFsER8QjEKDfZmMeBX2fjoN2hzwmYLudlcGxjorK2GZtJtFB4d
DsqPIwV04E2GpRAImnOFgTOHhkvV2PiGAeX7ZjbnUgFSw6FUhMASYUxWwkQmY8dXMvvevAOjoegL
EpwyyJWZt7ua912d1Qm0xRju5Oe3HEemeUS/S68/hPbVik6/AHpJmY4NvTUhReUPU877dnrAl5LX
BcxfPXc8c1nnxPYrkyOdpwRk2PWQkQTm9o5QRVcflBE7zo1RB6RjY0cWpQ5QZZ1P5ryCjT/A6dPr
uwv0AQ7gPJus9OHbJfsQxd+s7t9lqw2m0yAafo3NPmrVI+6e4G4pPmcEoJHHgQer9EIv0IwapNEA
rQ0UZLS4MG6ozw5vjVi9ioIkB6kUY7OHSMj5dHsfxl9n3yYA1mhYwMsf3+PPJ5EbLaW1Et4H5Tha
z7REvQAODo5w8Rdhgbh8ASTQyGobGE5D77b0Tct9fz1tnENLb1cUYTtWqPuXO3GRujhb3ribVPTV
s53bQxffqQjy/tctxJwytFoDgHRKw8BNjsNT0FsIrGbvsrzrBNWu//V8pUuqOanuCvsOx9RTwTdR
cXiKRAEC4APkHlOt9qUJv9ay7aFS+W0CK6/tPp4NWXHR808l2RvT99e2SXK5mNmULQjRx8jWuvZ+
HswicT/P8Xd1D7jfPYrr78NX9rsy4wwNlr5MMHEQYsHnpPGwdPWIsTfyMrtZs5Vrip8ckHR4zffy
kCxF3EXCFIwLlhGI8bvxUSGm7OHuvhL1/juPS/aDamUwTdG7lxMsmQhjpmu0zwywKjhlA4WacguS
wSuDj/0zVqzgWeDRJ5zQuiMY7EajDiLllwLwi5P+AjiSuRaJ/0Io30P0ldXLgYtufDt8a0opccgY
+TC0vgDVLqNrkAXyszxvcfOFPKBhQvzie7798ZIN0fCCASqBZ6wldWliHQeW79rr/P6zO0ZWdrsT
7i3ZpPtMbAmChvuqLsxw6g2nXqbcqSvklM2G1rjl1K/S/Zjmi4+O2ClGpj2jm0wDBX5dGBnJyI/w
6WXZx0uu3eV7C+qDqy6fFTAPoTmZxgJbdML/tangbsseNOrPlpjg8KrMATe+kqpawrTyWUgiT6/t
uEbMI3PObHsmag9vKLgWM3F1kuvH4YWILG6wvH+OgvbL9WB5u46zCpHQ6r78I9Y9hbKgTnp0OBti
vZ1tOPMvB87OiGjb8Zh/0U73FJ2CheXdkMbZZ66JNIgG0u5uKBE+Va0CXSQxltzPQ6BhmXB2rESG
gO0qa6q6QhoTW1wkqgXD3yVXrou29YdoQQ4J2Pj5VMUpK5pFHQfH520dc0io2vieYrqWv7WefL+U
V6hha1Wm11wGwLc/RucGvq7o81roSRc5DPTK0W3lflBgkmL+A26UNjihPJAGo9/taYmPIQjnU37g
otYTh+k9CV9NQ7Ypq9FsKoa9U3oDwTgsOctziKes4UGfTNCAymoNlzv6XW/OjJEezX+mnH7/b0Bi
50tUyhVCiR0s35nCLDoZ6u9vPVUAuoNcz0ImdwtLCPOceRk7G/8IdqDzmhBOLkzkGBytLuA9ZJbF
9pl6PW3shIAbYNwZuohbzbkLHDt0RtSlFXRwgyEkbETfC5Ib7h6IoTg3gk4PYhfLB9kUhxuuflpW
37hIt8W8fGOmSf2c+ok+OBSHmiNUqO8PHbsc3XNb489laYchWNyebzDh18P/B9/jL4f/wJqxtEWl
wlIiolIxCB4bRus17LNLs+5nyDw1riGjcRDBdYZbClT76Fve//cx9kjJ3NxtTW/S6g3iAMsMaTRe
FfospHEI6cK16iNyoDFyu7/HhpVaJ6OhgEgj5Qr5Cj+utU+LhJOVx4H0dPvvJQbB5hffJtgz0KLO
U6+PooAmPnYuZ4Y0fbnIn37clT0l+0LE+H6hjlWJcksx+YKoCXuRiFm3O5Nu52WhChLt5EKG89xf
g3LwzSSBa0epuzm+af4QQaj8zWIwMDf6XXIfOtlhLwpaojq8wa80M6IycqzU7eVQPT49SlEZKPMu
1Xd/bfhS9KidZ9gaaOaq3fKq0nyA0rLZR2YQMkjntCJuOxDuspONbDmHj/xEzjOexqBROl3gXEvO
zC0rkxYJ47Xg5YVVEErkKtfHoFzzr772ykWBcFjbBMmJHXHX6VkU2zLMrfdaZQ6LD5cRkpQYoMir
KzRzhrb9vI+TVUDsOuCTig48yIWpNmOF2BIZ75BGoyAQWaQWYl2CnQJSXhKKUKiitGwrZ5UmRPIL
L9dVX2rXV0rcVseXTE0JvTB6UFbDWg5M89l1+FIQSgA1tx/wcAHcx8qQkO1R5FelqxRA25/xKctn
p16SNuJzeGTWJcchc3omtC0hs0uawWhe1xQHUUgBnJ54OqcFSnEX6LsxASiKA+VCaJbwGundi3oS
f+X8AuVU8sig/epdg5mqH/Przk235PeLCSrM1BMOp5lvgRp7IHXjZnGefIB2NsCwsOvg65/Bxaec
rdbmzXx7/3ZF4Ieem3m5vNQW+iPSwOGfD6U9KYvw6twt+vA/HN60bOnCcAPik/Z5loCeKm/IHfD5
Z8KDuWTGARd9iiPlHxnmqvs3FCOLVq1b/xHKFxrSEO7RuwAiMp1I2kFJExlN2D4e35mzj/Fh8PD3
hUzQKiwOfYwLPNrw6aRArsaCk68sNMaT/iUus1S3D0/Xod4Ho8BZcBOQ+d3hi1WHRrvvGk7S+VAg
hIndGcN+toqmi5oAZpv84sFsBwVto2j0uNOR8GSvs6b2vaBcx20PBc3xc/twUirq1sn/5bPRLCIc
GklXNoOJsfhYPVB3ZwgCkWlc7vVPTs8dXz0/dI/b9Dh4SrL+JJkOyeZraQ4+ylkVb5pVn6SsXdzU
TMt0BRr5Fw8XQeCkDqOKZrUvRKw7cw0rOQWF0i+1267OTibZyTo2KVRsBn5FmVmA2lPDIP+x1bmE
WQNN2HMMAqDsn6iORc+L9W1PI4E6bdURAOxPfJ6z+CWmzQJolSjqaPIFlSPMFy2vCcXDnhXd1Pgr
Kpfxh6EMINduknBeeLnYKXLhUxxpmlrb13axTS02etkMkmlqNlw5A/6jS0ZtgiuRsJ7PB9YIk67t
3jYNgEL0EDHQRFCmeEYlGFHYW+CM9sZVoARDmaGKhFg7zmpd3y3X9FZZP2HM9dwPTmmECpbhZg6W
CCc7yo3ka8yn/CLhNsmRSH61K8G+hxmnr4Qqm7TzQzim23eDWEIjIVjhR8r2ljCwA66wxIpg6BGy
hhMBxz8yjDgiMwRzDeE85VtaEa3O9O1fDojGh8TXq426VKKx+31wU9vv2MiXnUMr1a125ePXGu/v
zjaHQxjye/y38Qj+xXp3RRYiAhh71brc+lhJlZ6uSmyRijP2GLQ/XQ+RbWMGR/fttuZ6jRadrb6T
OkJfSRavw/g2lghpAqhmMOZJjhdyWbtLWbIZVO4KRJI5SwvDgA4KHVOivuX4hXrQk4IMD00utqV2
cOXXsicUyhetIiNNDvpyXSVVBjUrlBMH5sHerMNkelq7JQXhtPLqKMwVlWVJXIb7wBRU+y/NdIf8
MpbwlR8hXETuZ7XC7UAns59eaiJh7E64h5+naXo94Bj1W28bZzE6mffkvP4JQjeJtWQlCit/vB4h
e+nTU6Vuc6eu/3xdpoEexbojlbrmAxGfgkyqwSDXqJBJYxt0CAUiV+mxVCessA2FpGytwtfvcB11
sktnnx1pSfhfgCQBHQQJHQAKW1HbNQq9ENuqZtOCEegDuTMU2dsDmT6PxYd+FEV1xmyZFRM70ivZ
Vk71y9S8Q9KYVj2D3VroHOmO0Q0kOU36yGczg3e23u9/JM02y3LN3WG2HV2uKqSidPhrD4LeYI5E
OBLvwoFLacgZB6eocO8Bts56O+DTAxELGSxZqM0D8VoC9a0Uc1x6JAEpJLVcVw5oUwyG36SgTuCq
Vr88oK/CvHp89BctaXCKsPL0IvAqHucCZYHYpRXgkY4HZh2ju5hWf3p3Pv35wYFwuvI5wM0fR5Oc
LSYxvDyQqlzuGttNqFlCgY5/A7RnEh34DTbr7bB6o//XWVGr1iDTHs+Lt++/BdF1uq6lA7Mc5cOu
sXv5FQK6bNlDG9SXSrFnctvw0FNja2GCzhAtKm5M7gRPLBZGMXhhjNZsvcwmst+z3LVHzJk7G9Gm
+7tI8o0/vRmwfMG1WfMPe2cc7zxYjPB+YEBiVMjdjuyrV9+P+HCbK4f6awVgMuiiuDNKTK6OWsjz
xw2CcKbt22v8TodexLzBVaypi/hvofeAjcuqTtsVeCDMNrUj4F476vKOmkysHA8EJGRuqe3XfF6v
XSSP7CljfRoLkNX6UR0ZKLJn+9MJjpjk5Jb46MppCVEwVzhdTmjPI2PKz+cj6wpr/cO/fvgMCB2y
3FQSq9dbgHIgZFYyLscImOnzwqSVH+RhLBuNNZhrgx6y5Hop2veaR+pYoMTl3hu4nnjoNbuOjI71
DSMxhQjWsRHETzBkmus9VNGzEwHvKQdx0LdzJyzsSEqbPGhLc11GpRsRasaaHiZ0ugxE4ORb7+Rx
8CuP/ZKByU+/unxk4+QDIjALne0RFt5IUbR7jI67Zy7npBEHEz09OLreP6/2YXTrnXEEo216+Oka
lrxMY7GCVEDC+yedGyOb+eULU7zFxs3HLfJXyOmFnESJ0/n493QhKxrpgRBoo+P3Oh1o4bbEgYVR
bjE1jzEUaVaVBkufWt0C1+X/d9kNMbQ8BD0wq0xaGnE2NyE0f1KqUVx0sDWWCICco0i7vRS/7jj0
8+/nPyTOwyp/KPC3cPPswGXKvJmtZwHGlvrXs0TXYvhWff3NiHVR7B9+9LQZnwEofxh7WJosXxVN
eczcj1sVY04ul1R/Smubd32Re314AKt2qp5gLZc06yEJy6cDMiNFA2UH++Sn+RfDtQlBvn5R1SBN
yJiZIUIxHZzjO+QmSScX6p2g7wyDPq+jwEU2VRT3JHMDkLdU6nTY1ttf0sf+U71eiCNgHGQXsOq7
Go+moXg4n6NeGRjB4wwyJw9EwnFhA93Vn2rP+YvWDvX9hhrxRJlNOttXg7ceE/w9t/0/kb9Jn5Jk
JgQM6aLFSD19rpn/jj+6R/EFLAnHJiQk6ULFskPj2qTV70uLoLDbFxQoBd9ezoBLmdgdAa+JGauq
yj7vIgn5Kd34ZeTqwkaXViPmVsk5LEQpUKZANJiaZ2L0TZFVsQ00IUrZoquLrHm77I4FjfDB8MXl
YTlxbFTIYOdsS7ksADAqBsT5eW0WX0D9Swr1fsngncqhZdhRUz06gdzKKiEmZUdF/05I66ICjSVS
e45cs/+Q+4aSePjgDvn9yOEFVgHUiUgspkKeVUbTgCTqYlMHMT4ZvnwbNdb+Ik/wfvXa4to7A9g9
MR4UJq4iYfnoyRtzFO4lV8ID61Ej0+ErKzjpmtvUFncuHVkcKDCssD9f1V4P1P76oxuTVaLNzWP+
39ReU4ku+emPf4eUyx62gWODe6Z9htHXKeyi8tseNELCAuS6rhKsPJUZlIfo9mAxGvkfszsiNoeE
f7cc6+EgCMuNhNRYIFdqwmakb2XGPITkJJZCYzlI6+G543ILbZ6+FR4yhjq9fCz9yTs5cXkmo0Bc
LQAhnw3vgYw/csA9/3Z0yaGedHU6jvV6Z4YEPxMVK12UP8fgHweF49NNhjoTvj1kyo6BsvgnXPvm
NwdwM1dFPVLXjxzXYjCArGqCvgu9lYDxBLL8X/wWe0yDE3Yyi/niML2dEgHqosA9NamlqzUGYIXP
Vo5bmqvCzhnJZW2qg7FzHMYAiy8zuWja3+9KhYUNRRHOS9YUiPa/K99tlLlsX7JvuYC9zxew1Zna
sQ52R5ZxVweHHIRtJ2l+b0v2Lfek/wHqR4/p6zV2eeaUmuDLtICC/y/mwrz38CWWc90bYJOYSLOY
l6dp16t9v3MpgaEaRsY9D7RnPyr8etc7koswW50xS8uwQJvM8L6u58JQS5Lg3zGv7AxCdYGN4x9z
DV7YX1RXpPAtqOQt9vP1eXL88P7b2XrRk2Lba45LF179UBCzwDd4pfeIAjmElu+XfA00DOuR1+Qk
RjciAZDgomNSH4rP89jkP0lwzWNosY66N21cIBdEIyOQvFaXYtovsqNzlH6p+mz70p3RdFhJ/q1M
7JSwRen3jR7mC51A6KLMhq43PoCSTJtUQ67lfvRbOQfcT+z3Pyy/sEtLcUFaXD2ctAD5t4p+4ArS
CWWwK7bw3kiXPhkL8WRRzHTPvZmtKcBRpO2JfumPpCK+ZKftESy3xUsDJiKKqVRPmR04I8onwDy0
uU6y7uVROv+6Xvo63jZgjzwSW+v4xlQCfvF3oCd940r6h1dW9ESfRUHYAjoPN31Caap0RlZzHH/k
rSH8V0GHXXNvXrZg1qEbLjbZvQN/BSgY82Ddhmxuy+aBLZDKGmau1B9lMObLnwO74wuP0/WhEZdZ
+eM7dwjWncGpVDbania/lyfg+sHLtUExuP2fk4LfHYN1vGCXSl9KN+ta5X7fUFPKZ4RWIfHdyH8G
HQo7vnVX8xdF1ycf5PZkrwNdMQ1Q4ZCx8NU/OubtUT9i64aRMkVb/u+7flHK9xZP2Rhm2B5t0o3Y
Jy420f6oz5A8Cm5wLtJafZSmS4zVoL1iGicqgAhTk+fvTrF3Cl1tVGDPvn2qyeLb/Fz1FLaCVj/m
+xouuMBg5NyHBhNnD2FN33AsoIHz0Mj3r4n6Jyv6OisZGhEaxSOubRKdmBT32MA0shBx+5CiBPNZ
cnl9lql7HfO9apqTg3IBiWfH4vptPb+6O0N88tWt6jDNq2gUe5G5NFlYS93uxgvMiKak3DuCzlbN
9oGfkhsq/PTYxdB7WZJA0wO4NX1K7JzODcZGDpqgo7oNYSgRXClU4OcpzDgKGs4JaHn4+vASe/Bm
IPbBDrP8dLAZPFIQZ9gQE5TU7nAUBrhk3ZGTROgqm3JaFPlm6LhvMRCxxmY+tGS6LdA5KMQBkpAf
3YpyxEuanw5eTTG3iMFHkkAb3qzmCLSf1tsMf0keTb6gcneo8Yy7SlUmDIY9QciQ4bE1xno8dZGS
6rvEwORCuiIywFsVcTbqo/HGf1NL7oiTJ/LZ0MowfV9dtdPYOBihtesCrnogzlqG06p6i80e1Gli
sDcPaqolveOXDn9ITztEeCE1FuPWyIYiZ3y+ggWFR8TJUPaaYBsMjN+GZet8Yl2Kdres3P/QO/K1
NMkiYnSWKRc5vFZVYlQyGfMm4Mm70zdRoECfJH9AjxMqLj1ZI6gpvJtWcnuft4slFIACKHrYFHeE
RvnJUaBpAAlpXGk09epNRdihFM24sqnLyIM0FoboMkIid/jWjYCNyYoGo/HLSpBf+Nl1ha83c3GZ
CJJUYanRcMtEuq7O4gcSCh6jEdxHht2YMpgJe0LTe4x5nfDiqjLOMVfyCv/tYTORT+44RPQdt1t6
X2dnJYZi+J1Msc5US5LIuAWfJKOG0n3IrftAf62FTYwOsj3NmhkGV4e3METFA4BYxGjqGnmt4mAU
9l8D0WTy7wgUhNdWlH0mEBN4UkD+Yn2G8Qj/Ya6MVaQbZ5fZgWI40VHkEy1Q+/vjYt6SqjRTUf2H
zuDIQxsM++Jb1oInvIl7izt4D952tgog5uXLkVFao6AKOhc+y/EKiyzguAaeLKxUy7myHxaObko1
ROB2YajarNNmfARVJyxovrnjm0HRuMoRWflAaZG3udyIl4sHXE3ZZ95VVlhbgO9izx6MOQXcxynB
87PeFF6Nm3OIrHWBv6cQK2VAFYwYaRMoDqGBnT4WB2FMrpcFpSv0UEPCCiq17UJdpq6YwlrK/EUE
uBoDsuyCU/fjAxVBSKx8Bii4VK/sjg51ggo4F0fbThQDVrOpZJjI9oVF7rHxr6Hw2/sv8+448Xzy
ZjI/KLr6NHSiNY77mRVgR5LURG0yHqMleUiBKp7vQ1CalExUJcnIJ//QVtRq1D2YwUx0GqaDoVO4
s3lm0Odg9m8wWGz/0IXGc/k0kDyAiL/8ebCdibUJEUkyoByBFkE0Mr5ZyHC6ialjantToGrHWYGY
Vz+zbTXQbMyjSKSo6MTqN8JzEi+BUhurE7xm5ZBXgelox90eBmPwMH+ySGwscKfV6utyDrKUog6O
p+UIqsfQkspNh8Tu1PBQEQtVFHesmHwYZJpfde/jnZQS+tdEqmsNDvrZRvJ/9tVvhLH1NrhKa841
ytdIOirYgkPEVlzVaTLsvv0+apSYAD9FEWkrS6I/EC1lPJ0mnU0V4A7zwoMN+vqoRyDoUZBMrF/4
9DmztnzH46qT/+aQ7PjKXhRD/m9FbJ8rmLRy9AAqTn3I9zTuVWqypWUzAqVaFmvebTL2d8BEyfpG
lA6CDgAKJUN927s0RbVE6zsi5DDIF965iDWFcpon7BFhsKvfxw78L6JHN6ToX0hlEj1270fXuDow
Ut79g7rbA3ZwFAw2N+lDuShaV6IBkaLx9VBSySEXjU8V4NNSlNNWhWgRFMZU1qzNsuCSO8wTjyES
qMSr+mY6IA+jN7cC9Cq1S+DCrnP3CXJcjI7B3cMzqxV/bNQ1EQWuLom1VW1QWOIHJNkUV3QGfAil
frgPFv72xwqdmgbGmDNI/IeppuFq3MbaLmgNWwo+H59govsUt3A4VbmBRlFmrjAZHR58AJ0jlqJX
Tah/sgXF2Zz3sZCfvbH1e44beAUs6Crs+ouUkN68Kff3BljK+oJk7msCDHSfP7FNztKU2NxZ8N+/
QUKLehSs575SYh48IahTFaMvZkN5uUMSxGheN6e3FGfSoHNysqzsPp/03MDfv9JTw27F/lZBD8l+
1t+peFi4v+W74RrSA+aARWe4wiaIu9ywgMeNNQamkvTc1TuFhynHzLmHkJiucs+2WuOgbthpPnRv
kOh02rXfXD5MGdbsBYilUEQwRnlAX4gDkXi/sx1HgF961J0Qt75F5r+Az1qQ6z8CnscXv/kBF3Aj
MKhPDOy7EfKsiDgGhcxJhcmSYtWKRTeymhbN+Tciqv/Q1OPdPiXk8Qk3byWIFImsHxn3uk3zyJ+D
YU3CaYr6TuyA/nfndw9Z5/7hMK7j6cz5MeeMnKUbxbVbXErboq/BdIyFwGDnizsP2NcCWevjLm0d
NWgFRR11nMTqyoQWLcqSqEa1qygALTKGuUXejb8mDkSJzwaWFQWu8/VLbX7BBhAmD4syjCs1TKkz
WB82EAHBO2cukQ4pm541jGWak1A7p6/9ThhBqVNaj1aXE6Yo4M2aQP9nBdJOlTLLzaliBc5kWQvy
RmMrHpNw7XGqE4DDrZeTJf2dq5lHW6IOaBHz9N9lsVyrnyyCk3TiGbHhKAD+2Zf02cdPtUPsSDIk
gt+QbuA2XO3gxLzGSmZbyQpkE7kC/0j8e3hw66T7vj/NufCG3/kaLCuOSnB2BRztE1pq8uK3rCcW
AeRvjCsTEIMFeiPP8zBCgToNkP4Cjyz6fIXCVIcx00lg1uNJVv7DTf21sYeMr2/jJ5VlAkBQZZnT
y3pz0UdGkfxyZxE31hj1f8b+gcIumzjOMvbCVJ9b02d8nU9iAKhun9U3l5DN1e4icQKZMVoMEd9r
OUyr3/El4Qr85934+Jn5DuU7b8/UCtHCMNQ3wBLVI8jEjoOOnSsGGSwW7moxaHNevdyGO3f+PDKt
dfCId4wEJ1+SPr5d0OfUR1m4GEUoPlqy5i8DUvupw+3SXlXMZdAFIW+huYc2IyzxcdmIMxsP68i+
IsJa+7bDcMXGfbqEMOCQzgADM3byqCCarz13NRRs2bVDjBu73gXpid/iFHHcIcLy6eJ20eNsjnYP
pIZGYokVi18/nHwBQf54x4WU8PXkI7Ja516m9sH8pqQAfndXPORL2gv7X715K26vxUnhXr7qW4eu
qT+M6puyDsR7VhYFvNo0msiYTxzDL5Y/HVxIooIb/ywtgd7QhE2up2VQwokYKROawD6jVIvvxJHw
rPdxY4qkSOzxj+IHLkzvz1NN5E/v4vEdJwOYim1samnCRhkNoKnNtxXqIE1ULncUwl7S1JKuyNJ3
20OW+G+Z15fAmXVJCrtlAwMGQOfrqEVEdzSggXIEsVOhOgXRFRN2y4VJRA9vVi50LH4m5/kVtWk/
emKBRiB7gKTaE+6IUi6dqU5lxIcSQ4ixDZk2x+TAie9O83sLWtTWYN/iMJqpFemSEMVWw4SBpMHk
gPbvWTu158Ci+HvTkwpGhJzpSVjzD45d1mAfo3CZPL4pqbggYBI0kCtPVukRms+wWI/2Pxst9zaD
IlIXt0oRWbZSP/41uCUDvZ+hEuWPmZ7ViPSga+3UeMauKx3ilx8Dbw2Utn/bqvKD11eVbKrdK/Ks
UTQTMrtU36MmtCZEQ6wNWh+SBH8t/WcByLtLyXCzjPGMOZ5K2EvbBLRa/sWA8PIEyYp2FrzgOcBK
15lCWsNEPgOty/CPzLisNw/cNBk7UIkJNejRL1pUt2uO2rL+UCqRRsWjDwRRKQWca/uG+G3GN7/l
5Dj9ZsZOiyO/jHnbGKaud0YL9UWGFhFn9k3em4avlSoYvm+4nptYlewR3ETRgGWSfeDrj75sJwYD
HmvTF0Er+DWA5lY8qiJLSZaBuDlRfxHfJhG4soLWq7ahIH1p4B0dJRYG+jiDaGgJxz7hdpd25cYn
iKgc9dzPhVpZrn5I2QBrSFnLQD1t1cA3F/YlwQz2UJvHpkPvh3Prwnf2/4H95N4Mqy8AAe8Wk2gn
/ytJWg28rXOcFw2oVtR8rIix0HkF5TXCYKES4lM8a+sJyyIcaRSScRPwG4b0tKZ9QBaku2fizA0a
NasKJUlV04r2umzhTJEsziM417yoIP+hiMAh2fu89Iw7vAIFopSXdjT6wu5s/LL9FrfnTwzMuj0w
niEo+u8g2t3rz44hcCpqWZ5jOjDrWTiLTVpmsUTNlClSTZg3X7Nr9u8GAXIpY5goNxUhCJGT77DY
GhN8QvdhSTIz2Ju6UX/FzQ8/lrB4twttc1lO3j2d4jrOiSQbXJ6tyI0HooJrM0uG4l9mi0SYXAV6
uJn6Hb4c9v94AI+XKBvibAVftNP1xnArJ/1qG5lT4oCP/vGAiAKTZWE1BYrZiVl3dRfg5jvGbUXG
oQhpqcYjdK7KfTREYXP77Fi/pPGXb2pMg00XgVbFO/RGuZqLUYvezOd8WFPjcwra7dkQoOY0xolQ
/ahIRhNQDRlzt4gBY5ycK3VEQx5Hw9yrgragAgkF6RmhQTo7oR2w8A/CTEWQoecaA72NbAlUe/gA
EU6laxTdlEYvFlexVmOjFrGxwzN59T69kxqf/2Zaz9mbxL4x61FSSpL6fmSSRAqWIZ0c87gs92AA
ej49a3jCE2eyHFq81z9eDQVzeQXLFMLL/e4vGXXbmxXfKS1rFWtdetHWKl6M8NRJiN6UqjjZtR0Q
LbVYsGyEIsuF2rOKBR6EcAtsTo4uYDmEUIshXVmVaTmNFqK+U3wrfs7MgK0C94chTze1jfH632mV
HqKn3HCLD3yBOGZPmZJqiVqg0UFG81HZLq6ANJdUWaAIXiRj2Jayb4sXhqkuBGCnldhF3UDoFfeD
mAgXnpa701RhX+iWw14N09kZ/CbwPgWVYYmbBy+4Anc4XOmbacuSDAMBlmfzTFCi+zY6r6AbLJfd
Ok4yoxHRg/5yQgJGHIFVzYw5eqIYMSDtQIMOCEpfajH9WWmcTHmAK0A+DdD16G9qoey0Sue/FWgy
WFcOSKRdfg1ku/GqrAZAkQ+kH4jDoocPxxxYNLaXH2k/u4FOKY87GYLjnOF4pfhW4cZiAwQCWBoX
pG8Z8MnniAr/ldCZvFSTUC6iyPJ/B+Lb3O5zBFkyFGUYbEEzLmRxq+jIhVuT3p6k9mh2uhiG4ar+
ch4MfKIE8MGP1EME3tz/sglUoWHxyCHBkTC7gzOywPo8SLi96Yk0tH2cDjQLxIV+y57H6qkGUEq3
Y5uU/62hssDehDrFsYY/tGCvKk3FjNcfuEfKa0YZP+B383k1uUaol5cxXd64v4LqtHgBkC4g0p/5
FVRNqETLUVHaHoGfwoIYHn9icxNnMzyzo42rQe2EuDGY3+TOvfQu3GJISWTfD/gz6k6a07ldEcha
fiZOhA3c2o1bqXftxQkZ5B9Tqd28PE9Hyh975+LZvBGak250wVGDFA5RNEHudEvPA/GEBZHON/6y
5tm9Mb8DsvCvazD4wQl2LaswslmODk/GqIAtulW6l9kCg5wTD6KXewMjYlZteC8wKbRGHRqFJDiJ
iJrUco44Lp+QISkRM2EQxtNZ3Unnh15WnIlpdYoVHq52RmJ/750yFlh27lS+NLkAA4NoY1Xi0j7p
PIalwQsL8do60YOnpLPQk/AcRfb4tirMpcbh/af1bh44X7vYEvXuCTb5WNYn1s80SM1OHA+qFN6C
DC561KY2reeJR/d6p0zaex+SUoOq4Q0RHhy8WgygCoNo9evgoDh4EDPcQs1rttyHFwMscWFE7frL
JOLD/T3PcbPGMmvTmHSBl8xn+/IrnOk4R9y8ETwxeMUJG9SCArrRZsOmMVUsv54fhj3DnveoNEbG
AE9xxfjFU5VrZcWVyh2s1QqYA59GNrvF6vMonYim50Da27VQETIen3NJzTAZsqgTYRzPfM3ZGclZ
O3Ty2sp/DVnfAQQ8bh3ye8yGIzW4e66792spDXrIb/aw1nrnMGncWnxP4GUkMXlYXpYfi2WLLvKJ
7e5wj7tPlYzSN9Yn7BD7L+RvqerDgOt/YcOI7BNQEddHG55Y4bPF6ZfsCZGoB+eeuTFSpz334lkh
/vA1467xvjysasByLkme/ahs1J4XQzOFbD8yU4rHVndcCw49OnCACep8MeDixJqEFlJC06gr450l
2XF/BWXD182VAjGRZN/S95S9/NgtJvWUmEn1hP/F2JWBId6DT/gaGfo8PwiZpkNFUmGJ6etBaDlY
cRNY0ojmzRZBe+nKkx3yGeI/6kATfA5iWMiSTWM9oR6g8Qo8cKb/1zPT95+soA3yOHZYMpxv+XGE
Cd7p2+UrKZhTcLEEPQ5yiy2WkLvmN2QR1roi7OX24eqnIEcBg88UfPzNAbtUhvRMlCyA3iBsw4G6
Py+Geu6BMyQJMz/CkRGF+hhSDqdKv0DafidmSkwIANVfkBGOQEcGl0iw3x7Q+wNmJSn5UKOw5eLG
m4+pO5xhSzfG2tSyeGasYKqlJ+Ne0gFOIK4FVDGcsRB29SQxNgJBGJCaqECtbL5xhiJryDR6tZ0R
S00RTgfxX4yTUGflTAWAH7NI7N68cXajoRCe98tICfSemiKnURs7niiNjs8kZPTTg9jicOYs210Q
Yhn6PdP6C1M3gmHnuUieUGUXX6SRC1IpwiOf7HaBF4yln4qYkBREDcVkn9D0+b0CS4RhxkhxxJYN
deLX/rNKThalfmAItArt+BIfJyx4NYK4uoiR9WqNSCf3A47awb0aLubGsVu71KC+sDaEWIxQDCF5
ydkfOqRqKxNPdCEkWY54Und+UmRIWYKAtlTPWZIuwai6SVuQ8RK7e3G7kXZ0fayZu8dzNQEJJ1PD
6Xrg3R9PEy4LKwD+bRz1IesGnKvrhHhNHsC+0ddKTmO5yu3zFmoTyC+UKZ+5NwpNT7k9b0W3C7Kh
8INHmxl3UOrSwvabPC0aCicbY13RofaeoDSiauFcNk+lXOhzs1Tuik7a/K1dvZ+TKXdg8R2B6sZ0
xNIYtQGVb+zKSnA49jKz8vx8zd25UbMfpe4/tgMXLLmizTEaQe3TZPPjsU5ubjHkzuGx2p0pSQ2a
dO0eOR6h4sso1eH4hVq5StXbrOgkM1zZT8R7K2XDIQdV6pjjCC3Vd+QvxNtGkJKBIdilfDpEWeiY
lcPlOLCt452O0Cnr7qH/9lofD1uBE+WZpSV/2hZpCy+xZtsuY2C4mX0D8tHAbZBNASJXDLopXHyn
1HIjTh3EMOekB61TRo7NG8/JgKvHQCX+lNSy5WdGNQNcxAdK4o96dHTJXuLlp9BZNW6sFeQZ5BGK
rnRthzWjFKSm+WvbUnooB/bAi2ZQcWXArVTcshe7lKzTpttCCRCOXkORv75d+qr3OQxPsQxsEH9D
xnJDVft8KGfYi8/zQEVMP5plso5FaPpc7Gk4fswFBOssE8jCjAM1ONP8A4oCE2aMhyaAEE9s6rPN
Q1B3OT8MGITGFX0pS2VR+a9Zx7ts3UBw27wx6/+tknrdWLVY+E/4bRC8OlT5zvQWwZI2hYfofV3d
FMauQTtwoF9CBCK6T9ikRfLf4cC+PsLUk2EBnrC1fnmVufN+c5bMswBSSNLaWP/I8EwSz9Bz3y+G
7BFmOtLsNrCKrV6l+JjnpUFGOe8nn+EhnX+BJ1MJ7RlTxAcayBSZbAHwNCoB6n5swRmUqaWdWGsQ
0CIjSsabjZbQbnc4+ow690cyIBmNVReldWbkVhRPNJOblxOpK1iUqaMfRVGkpOsdGKFOILVc68Ta
bD3snZGlgKPQbcDFjAf/nk1D8DgVeYsOzz9XiHybDd04gy29Be7FqOB0t38H6OZvGUDgv2sJzbrb
kDSNL8z8cHQtzmJt4yUguYKfnaamUXFxxEaQHLntxbFbBmlOuA1riccTwk//R+mis1Swh/ZWjUsk
4VyWDcxDmqy34d1/E9fk87o9UtjGGkuUcwOrp8uf6uiFivFeImuvoWz4XdauQY3nomp5AP4RkK1j
C34Cr52ykojU3KR1i+1iZBJ1ICbsYDVD+uZ3IyykW0tUErtxx7gRwkt4dderVQxd5R0ymvrkEnOQ
8JSZnXmaycToHnnlf1duow2O5+fz8cgqaUP5Z315juSYoc/+EVj6DE803uMhqViw4iR8ZvBkR41C
RumjEIHKYCRHL2/cpSHJ55d6SFZTdqZhHDrLlADYBgVUhdsRM2+YvFSYZJAtUxS7nJW4/oK9/fbr
TLeqak/LNkTCeTB5vxOkwOJzXmhf5/2glGFieiLh2PJcaEb65vOM1HsXJtNpl97hpeGt377+xU2s
v136vkrC3KxThbc49GEdLhTWYAPQnKfn5M261t2WG5UGO3cNB3baTtTSqDEJSiemPCQmi2HrFdYL
oIQpbR0dt9hYHhZZHHOXPmwMGG6qvFH4jNiC7syrxJpU+ZOGswktyz3odiGPHa801d/z0v3YSTkk
S5CpgCetGz6Dz1Ux1Eu86LvDuBPnhpnvVAWqOvQu8FmGW/aBdRRxyP55OyfuyBwYI+k1KBQ139hu
BCOrkCLA9iOX+RoYUPCXUfNcTZv8wgbHop1dFVGReh9eG55VTFdzy+uD7/uBRFfYqW7G6EUCqm9C
sweSHtZZf4pe7wWf2MXC3yiGKEdB9OukWr9t3zgXQFa9nrvTnRBLtgMzZ/ua78mcH0JFKGR6E1aT
n5cX07a+2JDIgCJQCdr2T3rAVbc/iR2ANVjYAIWQDVWV+jKl0nljCl+KAe7T4vYgTg94opvxFIot
0KTxPDK90dSOlNt4B7Ll+DyhJsDeOyu+dM6h5nMS9OGWw2jk3ob8TRFXrbpv0le1Wz6r6s80IJzu
VthSs9nFvtE5WDCGt63muxVOTFeozdzn96euslJX9wxhii9L9BKeLEivGyi8tK0TrCeqBGtzzu/x
IB/1zvfAJsxDRSRgfxpkrXNfmjOJuW7UTpKGFN9kzaVzkgwqFlooMcPyO6SE8+dF5ctm5r+4OxO+
+7oymitncKZC0bXL5HFTiS80pcpE07bF/E+5w+fiLYJJWpCLCFPcPecHAymQA0IqGkuyJesgOAR1
K1BzBudKIFh1awe7GfPNu1nsB5tVPl2m+lDFz6U4oM0woXsX0fdE8itvx8KHp2PIC2bKgL1uGtVY
Luc7sfUGE/ZyAdD08+UfdRanRf9yKg3wOWC0YCqBJ7sdgrSSoAjl1OnrJRlSt1hdyODKHMxg3+1h
c8AVZaNOGrD42Pakf9xoid9KC9fWAPfAjGGhyx8tEgx1D8yzCJnsFMFVuXg1XRWes0jbDeyQBqrq
0xJAmR3sCHH55C+IPqsxTLS5NY0sF96sGzU1MMnt6bqUA2jDSCEdTEU6k1O1wb1aX8IZOkFukBdq
2dS3uLaH2V1jw7tNj3nrAyzHFUCI69lZsJYrdbuxB4KcThZEK2XhYETynTPPhtD+muict9jya5aa
+pbVaSSHX+wZqcxqtGs/8htvndjJNMYEk4xf0fzGEe4EGx1gN6QVThPDkx1ukg/5kCdXSY8CbgnN
GhnYPwi5xgo6pBNr4dzEuPP8Bsto6wxeh0uK5uom3yv/vdfarNmYN2pX+uXkzjX1KEJRkikiq0R3
y1myI69qqWqorjSatNuZFaNdnsjNkmSuKuOneyLR4bJSvV44RoeLYEsf3ZsPGD8SndbaXCg6vhZe
pEEbIdUAiz8pm3upIXtwruqHsXqE5dFOVd4sGwbdJKBkzvoVjSplXS1X40ZDtdc3ci4j6y0y3GB8
bedhGsQcbZbVrlHUzFS2Qo33JZNZPD6mlBSW0zjl+54H6LLvOyoe7haI113iHYt1ZjgyU+4ISZAZ
Gcdl68X+ZoyY3lxQ+fUdDiZ4cXIG5Sim/TfAJ6nSMUtf+M/drKZDD8vSHKe5xbnHLXZk/mMtnw3+
psvB9SbsGx71PAPqgUmBU+9cCJ40ZSytiaBeDUHJ6uRb8smWS0hbxEQh+y0GKEOteQJYhlnrk60Q
to7akys7L8/mNG1AlVNm4aiYvGRtp+XMMSvKXSNERCxFl0TMzD879pPVV8F4v8aADqFoRIQhegu9
Q6oylTetyBpAqu+1QCZ4XAH/DEaNDTZY2iSVyZlnKPm9myg++dMOGhROTwBWKJ/5AuX97gnW8+V7
OFHDS949wd5t1+AhVAUGV6Jm1i2SWqBfwWeAcSQyfsXo4ZciAPvk1jXmoCNAauaLjgQHLV8pw7n7
u81QI/m9fM3n/4SCIESl7/AzfH6Z6ncJzLQTfcKkXg+qGvxDS+f3ZMbZSqDe2CIIygPuIScrcfvz
CSOhZNGIQ1KDOR1DrFAEoW0VnF1vQPihZQ/nj3fpWm/FZSW05pAz+QCDfLlKqAnZ9HoxjgNlVNMD
PA244Ledl9mvwnfN7CK/jn/UJsnownsct5bLLrf6KR5VeBTscIew/6jznVzdbpO4kM3WmTvpkeck
YcUSv346gT4WZxR25KehK5lyfvXYUrYxz1L1t5PVWqkmA0Caa+M3qKZNGqJ1jQpPxDwe1jthVcfr
78k/TeeANQIdSkMoxmbobg9xrSQ554ByrVnbPa+RgME6b8+4XTvojATzQCHIqpvn8nnVAcqvsZiv
rWhZ0a7T+GCNTeSmC4+C2U141+q55fJAdTLhl5iWo94yXIb9e26wh78/nii26dGtvTwfMdrkpglU
ZVUXT689pYA7WXmxmnY0lqwev6ljbkCPl5DcJasK/DdGDC0rZQYRMQZ6MVaHjBa2pUZsTVkLJ7+D
zSqTa4RI3ZsmabBhHK2daV7exYy3bzjE/G7C8YQ4UZuwnIgyfgDYr5hOJzrTGxBU0LL7BLpvbIYJ
PLP2ES78z5fDauH+xnsjA4gCenY6ka/MRnzMTuC7khNZfixeJbKv8u8JlB27PDPU3EJjlDBsvicu
FaIOl2VYewAXPRje+kryGi18fP/sv2+9aubzeYXm4EV6+WfAhVnTruMg9iyPA4CnimF3Bswo7MzW
RRnIMm8FfrFzMPHOAZfuX4Qjsdt+OYgJMsQsjrXbh4Azstap5kr/o1yCo+8R55su6UZPYsvljr4d
QZiD+1Ok3G1nsakna6USeU9I+EgMtzf3s7o583WbdtPS3C+jQ+6v/XyATF1MnA3pUHbtqWDI1+9V
Y8ld6/q/1az088Pmm57zVa/bJ6SgAIxe0Tkz05MoYP6n1H/FTIvjQF+d9biPapkwUli0fCtSFD+s
ibiUETyuXprzwxWgPXe4S1ZHWSSDxqav24EWN73qN64IrcU6rPUlsuXyHGfLXUhQPYO/6IbFsyI9
XJtN2/Th5ovdAH0Uervbz4qVdHpKa9I8w9kkI9XRVKFNCkh2hCIWv/YRr8FQF92rwXyYZAbY+ra3
GF22pCHVniu2lDhgKrLvSp0PkC6J53tZ5pbplEPIyZ7wErYFhQyTiNrUuwWjzbQkdEIWiW4dt1r0
Qsk2isyFvqNcraIt1pR+oWq/vU74FfYi1+Xtqmzpg3ltn7bo8+8SFr5PKASFz6rMf5crdjLCP8+N
ZRICFJGtMAjsOvVdJyqY3MEUfamGrfS/2bxuAPjCKUfTZhWYucddiZfd/iLxizzzRkabuoyl50gh
CPsBpNneMO80mkS8xeyX/YqrZCc/T34utmnIKQcKrWzmh+SK7XiDmUmyroC4toEqalP+Z/Da/07P
XAK3mp2/cJZH0RMuL2udDNGIFdYsJdqCOlZYyhH7ZvnDiTJYjon6GoWkfg1n+8RPmNUl2Z8EqZPA
9y2i+l3gzDBrFE9Ot3Xui7d9sNIsTJgbGdxoh4VxyjJxUpJ02CtCCCLNEFy3mM0u2AwVbjosQsYe
MWvPI+jQ5DSpvfedXjZizLQ6mSnWSTuWLYxDEUEtiwpN6xvTsN5HrcBygcwyqbf2tp1Z6YvyTPYg
k4i/+QDBUkSgEpCXxdg3mDxITsBtbzCJcUzyiPtsBce5UhniIpi1JSNRsU1P6DzeNIijcPWnXpJk
xP/4URq6yZmyBUtgGat37bGWI5cWbbCPV+vh5VNzypRjNt5UurBuq0Useb4xRkyVYEvnZjLN3ImQ
oDDFzGC9h7XjxrhJsKso7gAf23+xrP3kD52VbdkFjvtcCPcGGtgmSRR0WT9kqSarOEJLGLJfn9mt
ti08Dmntt9OZ8RjJDlP8Fp4Nk3tCyN0X0+vIrlC1vb+LLaBN0Y9an2wwqEaDN9X3HjL5f0Qclbsi
GXaux1nj4Ko/AsVeow+6GhtwciHdR3qTGv9lfhTSQrphlDW7QRYLz044VJ/AKweZhWshAiGqHNlO
5mfsTT82lzOIY4Iv6Q4+1O6Ez+V3E0WOp2a4rPe1kZbYeHr/5KC9wKR0UmFWUKOo7fjTqh2ms1D0
J8zIZWbSdGFgOkWoSGJbM/vcDGH+IpR5P6gA1JJDBSIkExnME2/6fctiGTFbgoIJF1LN4jGYL0er
pof2ZCyp8ai5wi+qwczPUwni5OEC0XG4nJOiRTdh9UBP/RqYtjHgCIsIcXiFoteBOeFCIFQbrVHJ
DXeVofFRa/aMl4v5qhASJ0VrjB3yTf+nlDVr5M3C3Kb3VaS08VYlQCBS54Ydw7rSyo9PELSP9jV5
JEu8ry1Tg69xb9UQXaHbnrPQb3xBHlAG0Eg0P96QIUg4GQ5m7ZMzd1WLLQ5fTigBo2NMsmbtOS1G
LhWBjlLGlibcgqXp5kKl+N7Afwu+ZOVUHLSRY2ZIDjQGVpgW3qYVwKaHrUSOvWJDOMz7JRoiMWRs
wlxGAMhcIQztSt730uHUnTHTfTnw78E8x/rOLIbkLaKBKpbW1tt2i2ot9eN3nhtR59BQytnq658r
Ups3JuD0h4wSiSrAG+KskFJNChWtN4mRAj3ZwDYLP/+Oc5w9V4SqQfjRR2TLvrd8QacVXLfspHcI
ma+lhy8SjPGLwnvMqZm9aBn742/hhjDxw595DJqQ9ve00DfM/fLAace7xNLE/txvrSVB3PxHyzjz
Py0m41FYw35VR43gVLf4v15+UZeVfDnlWcGc2gyN4y7P9k6Gz9jhvdUF9mIWL1jK5fM1u4ty0MS/
9DVj4WVvWNFaCDq8ADcixXPme7Clkkm3EdzyPQB6jiOmPdDQpSfyMKplSAPq8ApXIadVtvGSdL3J
YNFdxzwmY7Ej2AbS/0zszlc+klXNwVdQ6rLsCwHumRAf22D4eGthxjm587noGL4Majrx4XzH9CQb
tpPdwsO4XV5IVjeTxeGjB52okaQHKrF8KvUktXicdsTVIyVbwr0Vq9FO+NkH6FVKRqfpytz++JUJ
jGwetyCwLLYdEefl2fyGIJ6Zzd3oGJdALjFppmOqFPhX5ZZDcz+s88gjv3IZm+ohHK4GCbsMDYYM
OSQPR9fjm1w2FUyg07nUjMDR3ubyewq+bbq3pAZnJupHBa/HhVuvAqSxHV53yMeh68UmGSnbvF6v
YvTSWH9l9WU0mlMWlNplGX/9I57USv+YPYMhLqHUxGH54cEIWzIaBEX/EYtHuM7XLqyTMkc9aezK
jclTHmwd6Avw+sw7mz1HfstFRkMVuGJAK4NGvUQA8ZjXbazVh2hfQuT0bMMEkb+T1g0snosik6c7
6M11vvU9edpti0/wT2cFq/dei538rt9GDeLe0Yoi3A/7cXk/SerTszHJATfQ0+lZKZM4dxZLSt2R
t8ef/P+MDpYsVSfRwXX7+dcre/X2IQw1VowtxyHb40OXDoO76BYTsGN0hbBlO+lh54ZRQAYia2/a
VMRvOamcfavMaPvrm8ml1mTAi+gOVcEKWRpB0CDLmV5DS3F5Msm5NPbIegbm1sDbv0tsi6TxKoQD
3l+f8xu49753jrZ68TYKIijI2r1C9+ucUsW8/6HtsPrLUc/36zIm4n+985b1+Z90OubQnukFvBll
WUH84ZjRbN5SN74bnG+vkuBStIWCwudInVAn8Uv/Z3q4AkrPJfSSLMf55vBzEwwZpTdedeuQC+xp
AtJ8kbixk33KYl3rrOxpobDdUPIeN7DN4zK9mJpVCJg/q+ARZvyM+WULscRJWg/R4Oa4nwWv7YB3
H0f/4Zf4TYjXa67QYGnxTPYlcjt/7dlr1nptoQZyjYTXz1tLI1jbdGZWmgk69DeR1eDSfrB1Rwzr
mAVnhnCdhPgT1Sy2sAe0ZWWYFad4QRi76nIie01Ei71/o7Rd83yMds+40EjJ5W2NH6Wxto+wKz61
V2vVZauSZCaPVaW0i/+5ufnyd+hMc03aM4KbuTaXWXv1gEzvbQWMiNHmdzj7UbwYcgx7ERp2QHA9
OgRWJCGo24LqbZJX3whc6hPvN5UJK8mINTLddf6cEBx+NKqR9xIHZd+Km8I0pkhfGoMkqMXHOBYT
MZUQLaTn1w80PI28I42ii97heH0qzKfL/wm+UmTZqF5PpUVGap4T0IudNFRyHmVUTh2RFomoNn6y
01GH1O/pSBv+JvacoLYlOtvfzaDeavFKL1ZUwL+angoqZftemZAFOWYwDypZsFOUBUn/dHBYMp3P
bDBfyDYhLIsJXb8p15HblurEZFoojBOQ+9e3qLPAjRZ3pZruKLnguW/UomDSWAMk4wpePkCMPv8u
dxGjtYX7NjSyrB4w6kmcXPxlST3funRWcEgUIF62OGpC/dAPmoqiBmkCPMfgQMN38P/q+Gh3y9gd
LMnZN02cMINhPPoX/uB1L4JnXvruUVdiZR2s5ofYbxMrpEqPmp1fi3Sj/sy38rGyEPviOsqj0XPl
TTq7F0VjqDfG3vt4WyaR9SbmgL31JfCE7t8IpDrQxK47n6z42NcGSPeRsrIJtFaYaVwfSrvEVFaW
z8b9JrZM11xdZ6ceQy1gi+gnZLH4vm7k81fRAyoz3+1D7WssvFPRQjWWih2/ahZr0ZQw2NNa+NPJ
fQWIhlTyh/t+VFjeiV5F9CZ9ATfUz0AaOPjpIh9OK9i0RdTPAwCuKGU8blUq3XiNbu0+UkFBFmSi
ooGRXzlms/10nYiPFLEjCQQ/cirShw+CvjhsQm3omxoEqi3ky2rwoqnloRlwypYxY4YlqDsIThbw
sQlOaNL+CjT0tB4L3i05T5HLbnz/8Bsw0KO+ztXyLQl51qCeN46ntmLjQBgldbYtZhjRSEWhRuJu
g0xFWVuMvdt8DIX6W2PVD6iBOB4GzRcl20G5xsvBxDc7V5ZJ5W0YoxmknwH9Pw/zBJzgFxzS3fdK
Vl2USqkUUhTfT/l0VBWdYEidKeF4aztmZQqHLOrnorTmaDp4meEJE2xEZFBRg20X4LMQFAnKvOSt
F5OMyREKP8CfgBx8tv+8DUlQx/n4TtwfD34sEitrdqP/w9aAMOiaenVf/QuAlAmdyYdvi0XsCdhz
D5HPZDz2FDSMl/RYE3+A6UHUUdvBMY/5XqX08LkmpezrNv1c/D6xTbEBQq0Ezj2Q80suJuYLQ4S9
E26x4P7poFr7SIdMaPiV62PMB+4l9bBi4Mb95fSJhab7uG8sxu5JCtOyQ8nOSvZf/yX+DWA8UeFK
4hJTRyPH8hgse9vgBFRftKx0Twmz4NZwPZwxCgCV5KdTlAWbJb8OXZTJfq0+02P48p1qCXCWbubO
pQiwWHG3MUyc/urvMLUzmnjercsBcnK5KnTPLdP/BbM+ezTOGZOZ1qakfa1EnZL97WnQ6jnqTllb
PmIXpTmsuog6TI37AZ8a8W1b8cC7f/atGmjyMjQ539tJTFaUQKCVP9sged/1V6i7c8gUlWwmcEdW
LFTUJVVL9T1ZNeuYW49QrOrVGu6OGKoOgKre4CC+pM7YB+ntR/hMVdDwkeI+cukUNct0gbZl/X1/
2PMkyubJtbvPtbd4NeXlwjPoqxFGXVJDQdhgbfSBe0R/8QjAtRRBU2dJAJONdAXE70478kIxlClP
W545UeF4lncQgn+bW6jTSdnktfGq2T7rf2b4+FeMjIlx3ftLQ2LbyvmqrWz1Ea6C+70AZuRUqQA3
D0KY7REvrF98pKnAAxF7jYXH6rw3jXw7HRAr+ptB22cFkoqM0H2RnMndtx/ZqbGTXAwBzliPssh+
3l3+NwS9kqPdg/yfB05JqTPjDQ0bAOcISDiv7JZ3mouY1gmQivDo2FTh59rn3Skl0zibWb2UoaP0
widu3W3pdCxVh/kHuE6edr6Scn9k3HWD7bEe47Pxdq3tOhvrjXveoePCLN5NS8bDBoSlIQgHAwab
ofmVwJC2P5vRSfCons4MdJoCPZEcn9KtfmPWeLzCmNYKTRMSf2iNUAAB1Sfg/ghNaItqJZVGxeST
6U5qQq7lyEK/737v6gsMpzrP1FtMTyr+y1JyVGfGfGS9HcmXFGYIDDM050o/0P/aNioiTpwjwsx9
GDuZ2I8B8xE6uHEUy+F+vHuBpHD6TqbiolQS6/k4h3qwLuJHtcHQJoHZ/tCNJ2G02XwfwHuutbcb
6QpWhmm67DNX/5T3pZFZVwaT3dkulKH0dYWdQaqNy6GQKWlXUg8g9ZfVUEa10Yr65xKzXzt6II74
88wCRQMs2mtnfPBhIL5WLq24OQCn378qvhZNevne73Sa6NtpqboUMjno5xvndOtP6GUt70vxCH4R
765c7Kwzvhm2XztRNm7ZrqRGuXpQlVC5vJ5LZAI3rLxAsi/TNu/nqJsLwe2v+/VCio4t/nNrsWtz
I5J82eXvOMqc9rJ/ggqRSV4sSWw3xkW4lIVZGYyIHlPufkJ9dxgpKyU9f0H7wZ451ZCtruEasvml
IrkF10Tl4TK++anJ444QqlMc9m2AMiIonSIQnTDsyariog2+5GRvo0ZiX7ieXAjAXnevZxjzNyQQ
JQM1QwJW7MLEtpWyFERg1hMB8zzNFK2uwwA1Aq8l3Co4rHcQPzuUXH2tUT4AMFapKdQgOYYRk4bH
0AuLE83csRptIJ6ry2pguRYJ/WBskFwLpxnNOp1aAA0cR/3DK+IaChpx4pZiLNvXbbk2ObgNCqkO
GPn0fgpre60/E4rMuMKrxO4ODZZlsiY07a5hfb847ygHNTt2vKJ01frS196saQ9eAl59IqfXJK83
qpwoPz21hk6VSC6SaAxNyxMAoIDhRqCNZPqvzVlHwYpmhjAvy3H7fS2p6FPFKk8+laUwJ49RWj4g
n3wkYik5zFRSYBGkSOzxKtJCBykAwFAnP101RlQFYnTCvFuyfnWBXwF4Qxyv+C7Q8kv/XTtqED8i
E+6mPuQ0eCEb8162zIwmC1Gf6Xpurnr2XubL/Ln7cUa4sUiLgtPQ5OGltCxvAMX2SzGO6Yw9FeW4
61dRucEriYtUwZ9kPjPXGATbG+2A1H9kxgmtQ4qRWj6g7p7ZhklvDKLa1slcfnH/HnNZoUsbk/SB
Ozy34GqhpMr2ihOTUQtnYo8VCoyI9CKq+pVXWNAs3+r75rQMoPb/7vT6dr7M0/6Ea6YeDHCL/VUU
y6PAXcXQqtUpnJmFr78U2LO+1qQNUp3mPDCdQdtnbG8vHIougsK2sXXXx9wH2X8MetjNIa1cxzGK
/PTp/VoVvW6regGuY/uaMX//8Ecm1MVAk+jlTMZ2dvykRyYy7MQmtM8f+HcBbn+g/tjRNEoXkey9
23wr/VHubswuqOkVUERfanwsE5GzLCdYGOvuJA54BnvyaiY9tQJTFt5T7Nt0QXinnmocIszS2TZS
KzidOyX0zXmpzut/AOiEUneapGjRWJx62v0mVzFZG5NCSjfrm/zhjYd8eOcgat1dTkfP2v5Imprq
mGi0haUcbJEi807MXScQxTCdC0LgGuEwU/UBVtLWJRAanasqMWRGjakaMxBqW+J5ZVqTpjXEr7l0
4FQxJl5BA9yLKPI5pcZvcDmfhowgnseftQDUiHthE4VO4LNnywtzxI/xMAwSzCqKpeJ2/AIMF/cK
ZoMcCxMZHu6zyqYLCixwIv+67yhAYOKGUOHuL3EKnMa+GlBJ5x/+KTl5DDu/OBYNrQJb3nglPKjn
LrqOXusO9jK+IxSDzynb2KBmrU6PlIpANglTt1PHAmgX3TDDLVJUzASQpaBKNUXalo2XMU/HCBH+
E/9Rh07DK6iBW8qBXoL3KHRan62TubhHoyueRtHqHJf2l3riADhuxIMKTwl0Q+1grmJg97QjSSh/
Jzwqm9PbHQDJ3e7b9W9c7Rjwb1/4PhVY7Hy10vmLGktNH4jdkfbPoXfY4/G5VdN3VxXKm6YcPB6v
B0vRoOMMga6TMHN1M+D5m58ztfrqh6S3OwWWDnUu+bNY63b7PTe1cQJr/Fp97SKta8tOhBSzYdN+
TAuL2ofvWz5ZjZS/V6KWWmrpaYg099BlZpMw6C9s6Gxezt06ragRDPZsL+truH7ezalm0r8UwfTp
rLupUc0Xua83nUOFFSKEJ3JYTw4P0jBH4m/fYOXVFHdRg0K3LlC+rmYj2j4Zw4LRYvciEiiTHc8X
4JOlWDG8PI1Jb0alHICckA/cnTRggo8tc2NFUAnxDOPLjjTRR3x7Yaox0M3eok4bFKC6cHtnSwaP
YIIgDrkV94Lz5Xi9rSGZIDeCHoV2NbbhThy6YnPnikzvVYPCBiWClz9I7Ocew+1mLno07S339g3k
pEYexY+M9C/tUe50mLXOZJYF7ahGadr/bR86D88FsFF0sZxsvKq4otNsmv59dwRkrgYfbDIU8De6
+PsaSzsyuAGVwwICU0Zqnqrx2f9jmmdsraI55dkwJcFLgSdo3C8tR8oEzA9FA9zIkaFNMt+NUrZJ
s7gXH9/fH86363SdN5IHeSVHJEopT6AgFvksNJ+QukqWDtlvT/ljiggDd67yNLKi5saPkb1aAE+g
SVFu+E+WtwM7X5Oa3BdP4B+w5z/hy6htOWw9GmsW5nlIDWy+K8PA64MOcHnPFFYsaPwBE8arDeJ0
Vrl9pjcA04qg3bTQHi94ejCGGaYTFXCwhQgIjQo0eWcM06NBtb7TiyL4RAI6Jd3R1hHw64ymQhzY
59SaX3ny6xhD9mYV6M97vq0WS3rNKRGlL5Fu2xxLJzTlqjH/zYX3otNX5kDafGbJQv1J78swjzKR
uy3J4a7d3oIlOLOhYvIv+DBCZ5ZW7HoqlUKmIommoO53v++7em4ZPgl0/NhbR7zsprMcnsX+f5PP
nuUhZWWIJ3AL4abG6PMwaXvcDQvo9NDywP+YU7uFrsltcgGuJ4j9d1pKeXWMNgAPdUri5mN+J388
CoIksv5pxlCnxnGb+ibTck63/ACPzGc0fnrhAsFU9wKSSafsMNRGincO9kAgtmw+NUBil0D3gBUG
hFTje/mI1Bevz6BclG6drdoZtg+M6ap5/VKvnGbxTU2LQ6NMUJ7C5zKJqbJMtv+d9bQ2zsGPkE3T
jVwRXjoShij6xjA6UPb/lzq42iyzQRLN8dRqvmNDoA3JXgzy89E9e0hGbD0Gv2fBURxaJqFSxH/x
jvHyIWSgTANWme+XIRDYEUo5oZNq/zP9z1qne/tMbwPUZB+Mhq0cbmJ+kPsOAcFVL6XYxdJmjJSW
56rTx7pIzI3+Ku6OnkPWvxNJcO68cq7df3n3O15a2g/s+Yklgr9DqB39VjLaL5YjDwteI19POUd1
7pwhmBOXCHpPCDsk9EDV67fOyVWa7SQhbw3b0b67eZjkH6x+H+noynLve4g0e2jEUkogj4meM/qU
FuVyOT7fFIcfS4DzlsP8XnYfZtPgT1HbvQgAz16mZkUePLT7NCah/31QxkTaQ54KoAARoklBK63g
+vvCIFR5aZ9dlLN1+B9e/tNnNbYYQp+DpwFNcW8cPNCSikj/WnbC7W61la/GiS+qYLEpkfX3Ls6g
9OD6XYUc6FV97fu+dlxPMO5Os3BiSviexkjwyJBKNQyAqbcmdOlKJvhKF/3HN6sPi5opLgYpaZ+a
aBoEmnOcyJlYyXCvWFGAk/1u8r0TmUBQjNT/QhETWxClZs74ef1BJLqHaZoAbSLiBdHDhzddWxE5
12PT+gZMQtcH/ajtJHtw9Mc1mxJAFbqUJDrc78wMYT5SwM1lHnm5X3kbSKBmwO7MDT88QVQmgoJg
uLbaZPQaWWZ3llLhSOYYosggHo4WwRBVhqysWtqDzCUYB1FanoKwP/FHzlgdgEPXUSL666tKD1z7
bk74fh94/65huspPsCqctDYQLl8QvZCbpmtT0il48pPQBXnV+Ani+kuv+lKHG+jI5RGacf2sMkfV
xaepyh2SnbXWSCEBHXAVErU4SVhDqKzOMWfgbBaFhL9wsqlthAOyxQtYmSZAyageSJLohJrRGMUg
iWi0Y+pHqXOjmPeNSB0NCPmIbF+FZM7fYhif3NeVk4fTUZUe3/iL788pxvVEkOikloYFXPxLZBCJ
g/Ymeo8k7h062S1m/mqyfzQ2gvx5rE34VbB5dGZPwB/tWbJ12LB6c5aSeZUzutRSmOUYd1lZuC/C
1CJCGEY+yBhp/S+Bt/o6EfyCREsx+J5z4bTTqYj7eaz7aLrx/STg3qaG6j8hMPT3YbRGa0PiU/jQ
eTAlG9/Jwwe3nGzpyHK8eaRze2djwRMWkWaKl0CvrcwSxbBOQBq/ZzbVfGCiOiFQOHTmzXt9wxyh
baJ1f15NYI8hBm2ySDOp4S+8W68YFwqs8Krz6iIxdESD4HeHofOQJO8QgIPPTJQEQ0eDziJrt6p4
XshYXn3YFDZNs+vT+wyJzoge+AvF3RgCXpcqSD+fskmChi2dD+T+zy00qWgThUjXLf49AZb5Pyem
1i07an8ffI8GbE8MxDtgizAQnGxXwZeE73RnMdWvjRdx2cyC9eCfWgihrG8v6+BPOHur0O3obelt
aIcizBLR8usAXAc/4M159rcfQ+vmCp6rt8B1Q9kQySFNeGY4Ia1w8FCVGZLwQXNc/SbQWb56+T7e
yjwFcDP2t+fBrdNPEtjH4PEXPOke7L0GjMHfE8JCCgrhDAr/QFg97b2kv1FHVG/U+WlRIo7YTSaZ
lp5Kotd9oxF+6bv+qbgi7+Rg7zB1i6+G6p1ygDrwCxnY2K/Ma/kgAEvIjxAZz4OVRO+yRarnw7lO
sNoQfUDU0vfvhZyW93viioOuDogaB+LhEkyTp2r5wkIAzFES72ZRe1LoWHcN3Cj4upUVKFBL36BH
afo5ks7osnmAI0Nf8ZfA5Dsr36+dCNUPM0Eu1uEYNjdtKYZ4H8ESAUmzewziLbNNLM544HEU2HqG
/hOoFKsgSobMpTKvOEFIzCboJMF16xDThQMlRdH2FLWTKZyIsZ7ogUO6ZbMiJvDTyxlBMqxSXgOA
6Sca6UisbsgaIxwj60YhJ94vWsEAGPX8OMu4/legZtS1gHVgiI7GYc4ol+y15GP/to0O6l1dOZsd
iiml2Wq+mhkPZTflFfWD/lTSM2ETBquxVrlSXTusqvFLL0pNngoEL9D4m/qZDyw81/UkWzsCjLIO
dMz29mrhWigt/HCw5kjERHSgYxqEu2gFdAGgfHIWsfw8DY0IFEbtgPNh8CiHAXwcD+DhuLf3g7IN
6xaYqhwKb90M0v2jImeKT9pyD1UIgWmc/w8/kuDtvw2i+lwzQpqxCofpQWn9DA243P8DdWMvUrcg
VECY0Wd6EA6I2KLdWFFqenwa9IG0QYA2ztD0O1+phtndeONH90+IvuMK1+AJcrYIj+l4rtjLYTM/
io4DtxVKIMjVugrHkbjKvDctJQMi7lty5d8fOqml4RDJUHnP6j37//C04dnmHcV2OALlSsn61opy
GEjUpVOq7JZm9zynnLfV/QDjFLF56dV0xzjLpzbP9AKko8Tc6se/rtBCPNzTtkNc8giKSX4b12vc
CEZ7uwAJ1nrHQM6Z09wn4Kcj11mGGiOUsaEee9G8ijDcNfHCxi3fxNZnQnp3uajlSJ+gbFa2afPa
Z1ZRMizhux7eigbc4Rq3YO9HsaOHN+A0fplWnP5SDlcIw9Gy0Vqp2Yaw9CmtNhxQkplKVIiZkWbp
Sfyq87vLFzdT9BpYLZh2KPClwOlv/ooY5awK0PWKw9STFfAJmj4g+zuvVN1BmW13tO1oiBeT846f
nEeoLD9A9jY+LJ1IHfoY6rit/hztCbL3snwRAzyoGXHJ5kn//bRpzQnSYHcm1qdWtwBa8sGcvZ13
eQbQp2dWuMZ0otA/qq3Bh8a78QOeVqB0Yh2cG1xKKYusOb26Hyzv9UA2hAgurk7SVOrE5egjucSE
cqigx8fgYE8aBQJ63gvFNFGyjEJGlxAQsrCYOUzBTLWKqlzheAQe32JjyjB6cZXkYJR6Qf+q0Y3t
Xaf6W4lNNcRMpzNKHnVFZUmGDiktY50nIGmeKtfdPpT5K+vPOX5VFDdbj2N43PZ1iastdhheo12a
mAbAJxCMQmHgHvnPzMUKh6O00NGIBNgMme7poaljpByjf1WA+CRc/GsT0mh778+DvuQyut22P5Zq
Tu/cBPlfzzXfqv9MwH73VWimCwGXt53tmorV/KQTKPpoX/Iri4i94c6tunSYvY1TRWjs37i8pbBg
+kHW5xF1bfPBTvLZzHhVJObgjCY3LrHTgp9iaKXzdiI0L1drrC28lo6zvoF2E6Oz7nxGF+yWaEEk
ZoQcLBbsUBFNaks3oyMI/5WJCqxzi2rlyWgybq8siRgMISE0aClux7XS7hCx3RtTaYcQO7/pV5GH
bOVd+BBoga8f2y8ArZnhNFKUWlUoKL9Qsm17JrS461bUOiU5EA2EzpxVk+I6EGvAqquX9Vp957/u
BKqr0AgN3OKToiQfSMKPavAE0aZnUnfLJmkPtPkRt9Q3Nbfg44luXFyt631GgfSixgJRZt85Fgrk
zV5QInTAlS4wO5omHLxLpGT/3EaZQak4Jm1ip6N0ec/wUuxQQ7ZMF45IhTQRKLl1wKLNIrYVzm9N
gN2UK/hEesNs1eKWvbnzK3oKlqmLI5vd3sLcg9vVFMz95ujON28E9rh+W4bXo+JZME9nitiFIrhD
upvdWYyyF6yFEWmVfGNyLu+p8DcvgGAyv/0iN5KDhvaotj3aoawteHbn+DRVI4sXpZAJmbDrDSEc
KkZq5hl/KXHJaj03ATFL+8j8lhPcrh1NpQQwrZwM5Vvp/Rm+h7zuBRw62m3MV+fINFOdiCzrT+V6
UhlmxSpH9Ju7H4sdzJBPi4jgq11fItwRU9qFESw1I7p4EIexq/a5XjyyoW3RFSI+fI7K5Mj4M8x4
49XLZ4+6d5Zj15W2nh/f0A/xBVRxlYpCPr12x0NPwWFUy3gc6AA7SZSA2tMzhK+3dnofVdgWXyv2
wW67qQDi4cOBITpluYKTSULbbge2v2wvzPIUkTDID+jg5aTAi4XBrdW4nKbC7imuwbVyVGa0rGDy
CZfjJ8LWK38IFWEwa55vOI9xj4DNwhf+nyhbHyWeio9OYwmIqH6jlDChGbzXKXjsukqt5Mx9xOc2
oRvl8/VT5DUYG+f0i9c6WzZuV0x2iYWOGY0seFeRV5XXeaxmddGtOt/E1ADAHZjqB5nN3NHRQ2uP
F4WdXJrkOntBRunRjHYdp8XgT1qKL7TYzpL8W/sEbhFkNJjDFEOELDU++bnLns21FosBZPfaMRZZ
Q4V6B21MZiEwdDnuQL175Zpg5Twza81QPD5QTs34FucIdJXGY6veTHvHNTLkhl8WpGD3tBU7Qcc2
OP2JUIOIP7gnJ6LDhMr6IZ0fEo00ghKVjlLDGl8zCAKoL9oGgmbIFoRYOMDWuWO5VXei1FdB8nE0
XZagI/Zt1mrAn9Hm7g2FlTcKUWVTdfm5YafMJuDagonmmYlkc8DNC/bIsfUUf11IsBwdH3e4jkn6
QlMxhZah9jJVA+F8VoHWyWx5lmyhL5HUVg8gnSR9wO08MfNVK8XzC1CwldxnOlG5d4cbc0MZ5Llb
eSQikw+qKNQP4fmUmj06F2pkdXc82qzOOaVAXy0JnXcE30RAj7C1WaBo+QY5aPLPrCGjX/kpOioq
fVdt/LzqFBkmhF6wZl3FrVkTGmSoGKegeFbvLjTdp61GDol30oGMCPouYzUh75rBY9IV1HjT9L/x
TCnvOf5lpY8MV3/kmkkxq5h1Vkg0QamLeA204ONbg/Rd+LSHyBcZQXQ+IUCHa/AsJu/47tSrjjKW
FV/4tYcDP2vUvLBqKW4q2QZqkEMJcGNGFsbub9dfAlrHqXE21Aq7FilvgDCiCOGx1oLesdcc/dT4
tyYW5sTxzxogse+w4eItJvj7DO6VrcKRwYpmL3+CQX/5zn7DH/8zCOthKxwMU2NpWsA5io2wF1TB
y/3T2Atv9aKGzditVJsz4tOJvEF+EZf//3bN5cjLmZsCnAzMyvPCIXQClDrE45a+d7rXaOMC2hwt
HkSahD9UfL/ig3viBvbJXKf36WJo2aBMIgono6yFv7QMlG2sVXeJsaCLr0fBYCBGLj6kA2q8PYPH
Olm/2r3TOQmKvEuf3UGHIclbseDUzl/POuAZXiqlZVZTVN8PyyxTzKLscrGmhQ4ou0ucb4Co2zLt
Y8iTlspco/xKu5U99s9qxqv5lixiRCQE14T6Uv4Nndrt8TcKqyx77y92X/8eK4JHfwhJc52EVesW
8M71j/n7BzkYSPKH+hSyCs6TeNLTLQ2FWbKx84wF+Q8oE1nh3swV8EZmEraQNmzmWy946/crgCEw
1Zv1F6ludZct5H0vn9TDBisOEb7qHp6a6kMUbCJ3/dkGsACdO3280mZ89rOuuT1RoMZLT96oE6zp
Bb9h8caFfOYETk9E2jg5m9KScNMW7ZNnSw3qRPdfDp0ISpog7MNHdS8Ft3K8ngIOqgSGiYDd4TrK
3BlECQrDvORD69Dzs8W+oTjct5NC7m3B8sk5126egM45Gn0UuFX/30qkWR8dKWUak21UENDv/9Rd
NiM2BlPQoNThgHD2wRDiquRY5bQnwLMobhED6iuivY0roAT27fj7jgcopynBsT46u+A7NwwErut1
4Stj+PgS7SKUL5kJ34hAnFwCiRrZ67sRbKb9YdMF2pQjWcrrzcTiXM8j7U1l3n1dgWcmpJnXEeke
Bl1REjQpuFpUx3ogWLDCGGOKu6+gwyAeyz5nb0q4Mzhn2AnkHORTCdg0h3PN+fihcwDOKv9bsa/s
90U0LamImBO6l1LPZkpIecx8WTZ3AhLiETVb9RpwTZuOFT0daxY8nxcjAs6a2SFNka8bRYfaVJyn
2Xw0rHRm3WCnnI4/gtdra/7bLzdRZL74+1JAPE/pWz9J3IUlitOG37fsJXuhsU9W37MEeiYPIDtt
7xQTpbR12r9MVhYOx5PXhAmcHi6JX0sZkXW2C0RCcIHgj/8sz7q+C9SRsnBh/pqDdYE4wtAl6k9R
mGGLKcAJzFAGhuWPLSX+VUkh7bUtO7JEx9GAa0TPfiqyKlLWyQrPaVTeZL1SLfpOhIKCNKd+ibNP
3iuRAVcHZndVBoDo13wh6FmhNaoFkaJyxes4+3pCtaQDL7BUb87GpJjb4wO57AHLdgfIxT4NAJvA
2mOT0xAA7p6eFahmYaUKPLhZB8/TNrH9A6BF5h0Su7inYUd7Z91JH4U00uzAQfYBbjgPVLnKAKrv
DZ0HHq4wANrgKfuTZoq+lYiWaok0LiZ0jC7Sto2aeFCSGAvp3K/6BwmGVE+O/JG3nEaSNeta9s4l
lZjdgzIh7ceDqpJ2Jt+2/6uBGkPs9LxarFD+jjffVtjAxPBvqeiFtz3Z3tT2ovY7FmvCPPNGo3OR
k1vJ8WPAMSLtG0bHA8b6bSuuzXfLU1TdAxFcjrnZCSO+zh1jsBQ0rlohpGdEu023oxoa7KE7mZJZ
1oMzJZAj69suQ9wQk2fYa0n89DHsm5qvM5Fz2Nxymsv9WOPJbJ7SCXLEpSLszk5znVfqfhLf/NX+
RdxDZPJHui3A3ea0cogu5cGUvwJ0r42XHmyezk/Re5QWlVgsykub0TNQmL6OjKHAOCSvf5BHkFaW
pF+gmyH8AHEqIu0HBcfQppNT1Eknh5Zl6LpXcd+wrpdpDN2Or0IDvvY7yV3uROFVvdC64j7lW5rl
INnSxfnGgtpJ2iu1ZSh5UWC7Zd1HndWI3rP3R1vuIIvxSiEWO01+Dnt1uJVhipA/g1jaw27bqGrO
hX3ztoi6r8gm6paRgG3ayt3qkBm9D8h0lrXl6lSG4PRsIlQJ11hyyV142BL8007l5M8+vT/zU8lm
eqaVMSeDV3rKgESKlG4T6lZrETxoqV/tQlhZRJYNUHDDu337G3x7ECzPs23+K15TeEIM/vmZ3L4B
Xh6V/94siK6AfdRtTidwQqHAmplaIDHBnihbZLgmImNkjJRzVzJuuq+xDkgmBYycRW5bTfKbP21z
8vPgh2DdyodCGuPIbPjXezsVRYHmZ3scXzqRKOtwxaTPjlUieR46omON3829PbYWvSaGlqo3YjRf
yTai7PbmhidVpmsccVpOCRQIz+wI5h93mIZ1waX2jeMlDfdDjo0E3rVlF51U65Uxtz9ww2wBkwxW
2EskDV40RWJlAfDqQNQPDOCs00GvLGvHK8MDorGfGGW9KfcYimNoMi8sIN/Im/phtiIRzuFdq7c1
WqX+ql29BKR3Iw0+AQ/6gi4eYC9VhoeF1noHdqVbvnC1sgAtPhbp8+Pqwls3ebXIb3wRtsnlehug
YjL2dp9TFd2I83KC/3TmOvfj7KEj93+QtaS2nnCsKhlh+CUYp11pg5jX0ZriYqlWq9kXFM+tXgt9
m29zuMLGy5AsephGps8PBKzN7CWkwlewJWspX+Q4siEB8hcQ7aZmipq844ccSNS16OWuBJ6jUBFJ
C2lVMNiX4xsMYkLq9RKSrlPpynU4xd4WUCoAYm9oZC0kv5HNilJhtTHGhIua8YeSmv9lu9jvAWB5
M/JChBHaZnH5ZYBPaxa80Ki41VXbn+cuqFoty/3lWVw1S6pEzjmk6uUnKlmeUYmAM1Uo91hmSVNv
KesGG07/lUeH31UaK7ZoNcWusu2RS0wOkR/dlI6+sn2MHmHRw8FWMZeF1gRk2KxAa4YwZ4y7yG5C
2egsR66U2Su6BmwWIYl52pRpk2ZCNrgJ7kWXiNvQ0PE/S9hSOEHyfKXcRIlAH1VJrSSoTD52fEsW
xehwbBmQ8MR9i582V6htgnzq++lUCGcQyvIGEhKYhyrLtfSK42/yCY1i9tgBLkpsERv5/jrENceb
OHqG46jrp6beXoVBC3ieYbBBW5ue+y/lacT9X9+lbE1BmJYE4sqH3vrZiwFP3NWv0XIP5LpnO7Yp
Bo9haEZr8ba0KAw2dScedFin+qKl1fwpUeOTh+Z427dBEdvuj1fXu/lJpO5bLSLsPIKp00fe+1Tt
zr2v6e+Kz9/9ryo8Euz7WxJz/P1Veb1U55xoiHz4xj0b2gZBYEFpFMXMyzJClfF3aYTndBDi2f0k
yuCKWTzhfgcdY0Yz156qyGmXo/iVY3O5yiRjlyrr8Qrqljpact9pO4AqoWp5xuxhHcHlOm+1UCYu
4RK+MVtZHjEwpoIcxpWhk8uzG0q2c47adjwp5EIXcQVQw/UhggIm2zDnzZ3o63uGBmoF1SnM5Daq
60rM72eSc3IH/os/xE7Mucw4xP/59u8hPATZnIBbaj+0o0QtNblGPgPeFtj0omRDYD13MGVeOcfK
V+PAtWAooV9QDYfV0/7+t+k9v9YUPJyYDT9/TAcel9N/YOF83MVom54RUv6k3wD34F+tnvdgGj2Z
Fmg7FPmaA+M9pVHSGb1HZ/N2L92VQR+LY+JkkMIMp/MZFCx3bxqYDtPck6bG4pD4ndAA+LCXem9G
LeetDT5JU8VVKxOOXuN96jAeFE7YD2mOYtUss1MrbBd+Wp9i6sl20HqNoL4H0JEyxqTNmFH68rob
FW/R9w5d11H4BJyhaVIbmqXBHkul4YOPSO2wkVG2gYwv8Q9gPqCfSmdsN9HpcqjQt8UaouoVH2NR
uhD0o5xIcfA8agi5HQssFW1vCotTKfRnkQhzd8SKz+n1xeiIajjT1Fs5fP/WmZ+P8Bm18eWB94jN
8I2PU7NFmnxEKQwKF+F06AxF04DTW4PvJ8wznXy0Bdyh60UzcnuekbTVeVXXqCRezWdj25swVMsE
fku7BGXuIUQzPmtu9g/hhYK0FsimTbyCPO0wbxDZi0gyorNkIp+XYeDyG3UhSlqJA0VCh34Si+GL
CC5g2i+gdXy8VSxpXSUGo4xs4+6R4cVmytS+AlrNk5xk10jXk3CgRR15N5egqEmMQ/ghF1sdEcmi
LkvZ+/+kZE/XGDrp2jw/buWqbXmgra1IZdWg9SozFZDo1+AW5G2BRlxhKYA4tn15lscnN/Ubntu3
4CgYl6J2wLUGhHCOda0LFGfXJXqi69X0qv4UmDXN4zPh0RAelY1mMpfdC4B8IlNwl7vZ39VcjtSk
Si4TwrFtSQOJp0M74C4hlWjGR2XS82D4RXd7kDq+2/VJNX3S7Nj9lZQQ6NLK5+gxL9tuBOZbExqw
kFak7RBzQTLWDa+auvVxFAbbs6IWf3Vyy8sBT7L3RNOPF53nA9VZf67VqVQ2d+32ITSWlUIKy2Ft
BKau10fjdD7FkWX3mEYBiZGctDplxa8mAXY5FrYj012Lotw+DqaPRXjkQQaCJcNFzgVnLwi9pvww
9Dv0MR6NHOTrDasJHt1koG5USNiJ0uF9jUWFBxGmKUmUNFJhFGtp9umAPwZVwvg=
`pragma protect end_protected
