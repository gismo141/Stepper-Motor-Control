// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:50 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ENNRh7aWa6vdPQCKIBQmNPx7sWZOmsqf0c7eqYCNr2CcTU/7IEU6nLLdMXlS50FL
mSehtUsIHXeWFskzSHxu/SJleHCgSm7oKdpSC6+JlIBd8tu3PIRR7o/4q9Ui0T4E
0RPrw+t8EFQ4cCDwiR89o14UCbMgRxQGjC+kv5n14BI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17440)
UOVmyPto34dLvhBpIulkHh56muCG83jvRGs/ZRvaCFQ9RaiLDWCKt+VQQalQJtYl
yUPfrg0NZVJPS9R/fkG++fGHA9YHy5KkUeEQw3a/9ZreZy305i+6sROcx+iLF4cm
VdJEa2qCXDdqe+/cVQlQpCzIEWanea6kpK2WEramYzzASD5xseUqW/jhIW9ypJB3
z7esdhYpC1tP9WlFFmGhj1hAhMTpy3DxhWSJnCDB5W89W6J7ZB1hyS9tGeo/6DNI
1LVWdIHaLm9cyXCY5sZ1Kv5rrVA172p7eH5GD1CERf2HX92YiZgqNt5dp3KZ5wco
a2DcnVfo+nREgUNm3ZScz67eDAZPbzK+qy67LR20iAdaefJhbE2vEPXEt52AdZsk
B0oZMXQ+j2nTCWXzB0V87Y9dCmz6nATOakzybgL3O8f4q8pL1fZvdEMBct484rMK
c4d45vSiuKk4b/QC/uLWEfdjSTJBLVSK4LaqP3ahiTerVL6Uy+cQ1Nxp3587RX7X
azWyBApCIKcFCO8DNcOlYW5y+wwKoeDRGHzTA1HV0QnsSs2Y28gRW9f+3Cg9AfAW
fJ3mHrTdD6B3Dk41NIzyb3I2DckpOlWqjP6C5uYVwbBle/StAGXzN/WbBh33J4T5
riWrd0DuOKhP0nD2JGBHRUfJ/p/Oebr2wg7H9AvPNOCvHdFzNbuzoTAS+VSCGl1L
P4QHqW+ZkLDAHSjW3ChT2qjoJI5+WRvp7HYrAPH/sXI1NJqdOMq4ykt/ec06+6CO
5B1zl7WagO7uikerHjJCXKlYY8wYtHgIP3hTllfNoSiJi5HvV12qZDMbmfolsQcF
31TIzXH2frNntGV+553h+7asEPro8ja3M/fKH2WH9g0fvVpaFkNjOJ05bb0lRUPf
Dke9NPMeVra1hB4R3QbvWFSNnrr975R+WFDaobM6e86jbkHqFPBLmcFjSZWP7ygq
hJxs8WvBLzgdkMoAnccliB41ftKn20ScmKMgiEX0PzuQ9IUARn3RWj/YJVDA2Vfz
C9R6Njs3rOUuQoZojcbQsF2StKASdZiJ4HsKE59sm+KSltXJOlRiCgNVGL2rr5ed
+Yz0l6tSNSVWfbSgEpA+Qe27sFFV83jq/7y691yugQYm+q5VDFdzgKpPS1/yi5FQ
/QkHTeO9Xp7pCTXskfCBVLlseixvV+upjoM+c98rrT4i4NNESEOIDjfXkhvRSHtr
dX6C6E8V/EbwvQ41EnaBi1Xs68cVBOZ7ZjQh6jXiSZqpgIs/CzCV3MqgluryETTd
POBbS4Y7BnZiBiVoTc1jBzGhZ1Z5RLYiM6C0hKmwwACOGE9CUuo406uTHdg8p86m
sFet8mmY6wr0ZrpiQpDW0NNAydcPYm5Y7NKXYVlYBxMESO+z3OnB2uq7MUCvrmGI
aF4ba3mqEdULL0YEErm58pZPcD7DEAsxf1YvXV5QfW5KJkRLunwMBTt+eT/ejX3+
JnaNtU7PPpv9etD66L6ylNcSTkVoU4dV+zBtHyItuEKLoisIbcHO5hqXUEzpM3mH
H9KwW8pZcaXcR/1uAbyJt5F9Qrhe4uG7yM8QWYueim1Upw1pT5X0O/kGSVygAgJi
oCTjXmigagRdvDrjIl8Qcn/GuGZXuKNs6r/j/ZfCSG+PIH4DmoAPlrT5U/oWNXlX
XltTUM/kywfAB2ltARHixAko1Axpu5EupKCfPH4aQdJq446wv6PIScOwKl5/dB22
w+lNQcf80aq2Bsjfexl61yswsIl+AAE+5K9V+n1b3KVPgY4L1zjCW3OR78zaYTJV
7dP5OKqV335IEQ1re7Iap0Z5zTD1swpcGdjq0e/7GGu4FtpCJdhTXACmoUdEfIKU
ZhKDa/kAdDIWE6+bNtEfgJTAyrSaON9GQnK/pMzfgjucNuqo7YS571SBT2KYdiNy
LRJM1KXw+TjN4inVRqxMNiTCodk7ldLmnHmImkO96OFzqHWpSD39kwKe29ucMfHW
BAUd8Wc9NCh35WRoEQysNXYHXAny9bqmGtri3HKghTJ2ozCWPIf7qrgj1iJRDXae
hmym0dGVvAOG96czG6kviutvzU4GpdgX1fomtmp81SKyu44rSfz328UjnnfzRgp9
Dxz2f+XB+d23zLeybPhcMBb3nSfqJ/vv0j8aH1IBQl3WQfmJjYuBIOkf3nbR/Isr
To3Rb3CImXX9GF9ppLZOem9dYYnMgi2yJBq7jRXeGpcgNjnqiyWGd6SXsq/mUxRW
fAlHMXC5ytW4BZlO/ua27RugSFT4X8nkHK+RmLwOIs5/FO2sD0zL2zAXJqA59xr5
EZLSTRZn8OTU7JrYFmqdguswnibL+85sb2F+LH2LpBW4ndbNNpWNh33O93D1MUm+
2i1hmZREup9hYVbKJ06UmOt0Abnd+p2ak0LymlP74ueoazSHtstuZFYmGaBmTgum
SwtgNGKGgu+EyqihrQpUYzIJL3FWvHq20cRRL2i7wm/FXzZcFdglYwHR7AMRAiL5
nnbMcPOYUlf8T/TmaE+Kz/WEdvvqiJ8M+6CggYf93KcOUXAg7/mWMUoIfPqwcAJ+
6Euecxlx0Ubj7Sofx1lhxrlyQg4OHoVbfg8wrHhjf5VZ75ATjEsh0pMFQMRzbobq
4iC6sZarAYD913DKdaw2TFuzbdfGLaQHmm0ewDSPUK9FePBF8t+bGFUXwlI0UzLw
pfn9ZobFtRzr4gIVegJZ4RBpJJy/RC/kko15kGv/JTo2GHXxyujEoGy/nCxH9h2A
uKZaKxqd/WnlQBXa4unyWbVPdRO0XQuo/Gbi6pBiRRylSFMgtTUjSUfetXZdrsN/
jychdFYo8xvR245Z2A3gJQrLdsSqGHgcG55xQb6zrQqw/DcJe6qWv+D4jYCDjaqm
Av6sm+uW6QFNYMz/rEF2Ih4YfF9nvFtup9BTKYdRdvuGIyXgUFnJ+lLUNIJ/wEJJ
F8A4ji8N6KC6yVLBIpqb6NIrhs0cJ5CM9e32wvwMxOF+AXDEWQ733Bl7nQT3tlkZ
vk+IMl8SGmZZXGFBfyLKDNa6YtZ1NG9LsiXHbRA41g/Tvv7R8l12x1ZWZfYnBuA+
HAgrZoghEngJij69C76O0W0B5ofTcpQaNXCX1eQ3HXV4FaGgJoQzbEW3QtzIymqd
07lFhjWkDN5krfKSGww45+qVk9U6Re21ouUTs5rWrn2E5azukv8ErNlUtuPt2Yu2
WBVv9RNkX+PPJ5fhevx4xExOnxTfvr2MPS64coKqzC+/6QeLNps5jzh9lurcZJuM
yJZx8rcPIlFvCXjr9Geso1LB+6aZSec2qbL0iXU/MzYXyyldFtzPSFQWiYZfcgXp
zxpiBzJnvIe9e5k6ZEV3QQnGgdRLJCuf9YONAgKo1AKd7g6TmOXLwZ1AKdlGAVLU
a2GuwBv+uMIf5YTmXNbYSkH3ru2bC1kk2Mdoqfq02n5oW3zeq+zqvtydqullzH7v
pm+9k1OaHaB5IumepmYOPbsu7s1Rg1r1eWSMAdd0btxyXfuQzYu0a3gUXjoNSmNQ
TrB13pPnw/Tu2zzZacPvoct2NzQxADnYByIWWPSZ7a1qSWg8J6DV6gXdWVvS4u65
0kzzfAC7b++6QvJJQnZpzINykzpitfbicggzgOlq3vvq8wkdA5jzzofQwGjbo5v1
It5cdcxhnxJ1apyGbdB5NqE7ak9YKaBYiRterzptw2CeKKcMhRG74RjPC49hcA77
j/6/SGd8oNgmHsmnSQW/OX8TF2C7DJY8iCzyVuWTvwmhnLP0pnm91VqGUCrB0ix5
aNJyN5muOfB9UTuretrTDXnPzVtzchLLKOUpKQuu61xzX2eZiRWNycyLbY18qDC1
WV3IMRuy3Bn/O1FX/bLzrUFpPwxGJzRdPoG9E702+y+KM77Ww8A8tqiWT2SubnnX
ZJPFZZ/Q2fTVNLqkOBwawxeFwyMuA+B5NFnW/YSUoMZRhkTFzgNMLNdqBa/4wQ+/
lAr0eFwuLH4tLVMypemYCsoT0pPw/eTUlf1Bw6x1pieU4MO8UywgOgZdPOZFeoMC
iQF6uhI2Iv2jkJe+fQxgQX4GQxBFK/bMXauz3IFuUqPprOea+DMZkFxJ3t2V/b+0
I8mhjS74nRG3k8IB0AoOJ2lDR6l3X0liAsmcFRzK3fo4ISpCnSAqX4wwKbGQm7U4
ryL/h8+WHP4+qYflHDmdaX5GDpSzaJhHnGRvZDRfO3SZcfjrb5UQ2Op34iLL/gBD
dUMh4E86adTOJaYOoVLJoUykxu63O859KgkZvkDuT+jJNrDpJdHgnFJrHEmM1vqx
7wLqoHpPXIs61kMY0T2+0vuvwGaTWND8jeeQ+y5L2rakTboCEaGa0nXeirXLbNbp
Dgg6mDG1mHy+yEBu8Bgg8OFGDD4VVa/v48//dGvQ94hfeicDoiIeVS6EojRHtlq2
OOOXGPpsX3ECe4F0YQg7G2Y/SAba8FjxUUA4TeKEbzi6tGm85T/NglXWYGvvIlop
ycIvcbUHS3zdtvC0hIFZs/cnBD8IBuASO/ue7Mh8jwFpdbbkWbDfc8nIZl/YNo0u
HQDXq0bwpVwcVwyQQ0zOql9BL6USe91cBfiRlNoFYi8UViEUGsmwfiIjoHGpub/M
eDuJyTW6FxTDxrSRFv7cZcb8TfswMB5ueVn/0nabjZa96eaPvNEHsXgyqtLQzjOO
4bVpqC14gKS0jenU2FBRBlv6xMaqxoh7EeSkyLLU5xz+TkY/ldA2gydvgD86xKe+
FTbMOK6q8r8D+/dbYtP+lKsN+EXIZ/chw07Vztwcus/oS+smYVExI5iPIrvJPbVX
CfjWc7vVECk6/21MD2cyHkpdYNK2y6zQqbeR0p0Hg89rcbt647L4K0PXzDdpjIqg
rSGPeB1U7PmjJuxk8vVizcfw4taynSM0JTRAVLVgd3J3ypZEnCDByutSzK0qWUvt
iJEpRtwZRHxqK6ArDIlO0iq1sn9xA5lzGzbU8+u9pydIG3/xRtaj3NrlHTR+4BRv
tbD8G4c+c6xp9pA//K2yifWiUbXEIPoZA1NDQtmvoFdaLct4mR5dx8j4Bgn9hsEB
527LupKER9ey2n7rQL44zhLlQCKrFTuNRyb47cadebB32oqBMut4wx3CMm3m8v6J
k1G5p7EgEz4NQcnYjmPSwYqky+pivT0FBrltC9hDNzygUNweQUETHRAODx4ETMtH
iFEHINx6QWaGYiIIiCoUL7GR//h2JT8AeFBrXf/xxmXDL8FsW/740/hpe8Zf+H6S
ZAv7UY+MjOYCR6HtvYwEFoI/M0nmP/iPb5mwHmrR0eFIqvKSR0hhqbj1BynoNOw6
cfBcqJQfxTuosEVnNs/AfDkbF7Mw8mCDXL9vll9W5K3rb4D/VAVyDfL/zfVZEo9B
edBpKXKA/jE7Ax2/0zcB9h/VDAG/0ax4iz2R/wLyPuXbdUmKnrVYTFxJqJJ9V6oZ
PTzeWyav505UsRI9NmMD24dR+5IV9/jJM/d3PwQJkhdj/oZPiMKs4Y4M6DYNnxbA
NWeOm0CG4iBToA2LiG1b/5bYnqDczDLMVrXIdXAfQNSjrc2CiD5r5NmBkosewMwy
lATFWNolIMJgDKC8WdAQqPtC94ErM5NRx+4AYTobFrUlfHti0rnzeGvq1nCLWtja
t8ak/JZ2AW5WqO8D3+JQbGpmwRe4HiQZhKxAKcV2FXQOw9435DBC1yU6VB+G8B9z
CVDgTghemFPB+Dq0AwWlkDmS1sIbYaJr1LS7+UABsiNs6TCZWZBQpSQglGN7yW/k
CZJN4iZLF03lq3eNbMRAQuA2s5lnFqsRZBhYQm2sugZGuHOoNCHENlQACtFcySnl
VbGmpp26D4dJikBFp9fvbd9FQQwlSmRdDBdq5c23QVpCfRjtYtHouHDEYGnB7Xto
DkCGq0ucfLkLKnklShVCsbP9SR+u45QhpJUEaPHquVJTQrI3xQoB7q9v8KMAa7PW
qlkDprtBhJVDTFlGZfJRYwJR+1gPQCbbHd+TbhVeAcCvSuxQYP7z95ODJJu6lkA7
sUyg+nLm2Boci8OfUy4BWtAo/+QI03RMI3GfKW30ST31vzCeeuZSWXy/dztUdWly
w7GuCiL7QSvalED3367FXUYbYlsQruYI3qIA2ZbT492szn/PunAybpnvk1VezcpZ
Fpotc/ikjqm0vySlxLO30/A2gzbwgUjJL7QyuQIxzXn9oqKrynREYKt5yLWsB8vI
0GqXZnACJGrkd0fzmOTNtk1mTLQOwrhfWNNCHqdDTriqmonxjdJuGFCjoyf0r/07
SKbw1cvGlLW+BlJ0/jFOPzmU/yyMCKP/zNuyp27ftFS/C4m0sShgjccvSKm9s9kg
pax+DbN8gelJAI3O5xEsLxORELM7n1dcfLZ/JKBeEUfbn4koiB7il12W5XFrlaFX
JVZMiEtAt/WtNkBxvBBaJNVhr9S60YtqANhR6jYzg2Dq6LutX9IoT4/Ho1D43DOk
HUZztNFBSovkQFSEZLf2khi00ewmWfsJOZs5nGeYi1jnRfnCfPGaxsuuV+FTkimL
kjXZwUnfuYbTN2t0/WBpPaEC3762c7NrYrp3lILkK3m9RWZhi37AxSUcQ8UPlp9S
6qJy4A304u4ZRuxlP8bghB0LdbcnAZQY4Z49MocVrLt8LzYYPoghgBoILij4VIs+
B7df7xku7kLkixDm3WGWaXWGtJV1ujm1lKqCcTvMPoqlle12ZvtSdlwareCXaa2N
wNMd01jG9WqfG4W+vSx8g+onMlgRaO+bW/VtiCfApU+g+FX8d/1qbEQ+bJttSYCH
DSoGTMzWYuglrJPATwWaKIpAsWWF2X2L0YTGh2DxC8sKtRyetiSE8W0kcRBZSaVy
xOXd9dSLLF+zVy1G8/0epoJRXeTkB/DG37iGHjW+J5bp7MxuLiS4YuX2EbWDz6Oq
4xzb0973EH2I45oNuztiCRDUshqI3uc0ytJrI0xfrulUa1Lv19u5TUpl7F7Y0Pp3
s3d28DqCeaRCD1Y59dlfj3OJQgoPmpo13VRlsTjN1QWdl8o0RwZiZK2T1WNSkkGs
cPJjeLgB3KPgdtAhz55up/Bu9bnr9DvDMB/F4CiE8XPoZnyxjisIQJJFCrQMtb0i
nLIO8NkQ8iuVt+Wy2Ld0unQgvadwOm32/bjmEnmDfIKj/PVifbcdEaUwRj/7KKhc
Ky5jF3gWMigWFEjx1Ktus1bJOzJ6+wpmHrtIs4C6njLLbnc8215YhB4WHkMLcq8u
Jgor1CgrGKHW/B69zr8cJVWuyd/Sj0o0FuEz6AsVft6OtkyeY6ZfDtlOwIyHTuvW
h3CXFFABUIMLUFypi6FAEQhuGCTqsXEhHqJDLOlzeHjm7j+b510LcAoykvLaCMt5
VmqTlM7ZsDZiL+CFI2A+pYXq5+pteR/+MWw6c4dss9U5lk3aJRPxfqExWK5CIkn3
hlLGYHXVpQpJZUWjh28DSxcSgbI19VXU9wBHNV5aAt0bvvKl1pSUW5ynUqa2qHVr
oirji0x4MZivQfLBvm6WXTtDO5+kh5X18leaZSzdTUigZKZ8bAtqUubyZ9sU5l0/
+SVE+UJLKIlPY3hwgamjF6noLA4epKtXW63HPZpZPKVK4zg6r1Jro27WXpo0vx9n
QRK5wb9ou8jjYKu40SbROz3FPL6o9VK5HZQDuS+bD00QgGzJfnmEa06iEU9kTFTD
Zo4lXRQ/3QPlx9M+ip8MUvXz13Uj3rpKZbnJjYI5deqo9fMUe0LQRDmJ9w8VEExM
soT0OTqdI2ErtKipWS2dwmIfhEO8ojFMmR6ttuTzafd4SKeIAsQaB7jAqHyQ9Xwi
HvrG0yKehXTVZ1qxmp2t/f0A1vkc00yp7iekHjdl46am6vpDLr1yXJGuDGqvRuWC
VEXWj/NZszzwt/6Jex4DAa6ptznZQW2AjKqwDmJ72uy+RVKSLFJqqTn+DjdeSDPF
QN0QdPrPrGtWYTNWnl5BBh7V6v+hdCXqCeWs9gNeSzkXjcvCg5xqRy0xob6GypQC
LvQQoy1adVHe99ylslSEeBOcwtTHuM/n5Vt4nEV/lcLvffHTOQQ8HST/pDIFwXWK
JncONory6bebZ9Akug4pi1xzaiJNuauKlKLq/M/i22TTLkfyf2iAfWHlPHMx9WWa
/bU8ahuO6eGw+xcF6oODjrSfP6WDsgpVR33jsppX3BbOKkNPZdaRmC2HsTAvgyQa
5n+kWXM7cx6K0+80LghbDo6doQqw7J3o70Xjh7yRzOfNqVJxEnla1Rk+h0sD8LSP
6hjkshlIwb/m0/JE9BrJRsl3AGePm10ZTh4DBHwqCIk9Gjtcgo+DbABjo4KmJdew
XB0IJJQkHrdHcjze1NbMhur9nYLvBigmgTlEvisXq7HGXkHcyNsOw8VglI4jclZL
SKfY20O0BU2CmclKezyiI2WztqA97JoPrynfeqIrr+r+Wa1N8M4Q7CRFSvJUhWcJ
wctw7dQ1GrGJEnkMXGYJvGMr+grorDMcEYkHcKFy2+RGMbff1JHgVKTD7H38hQ5Z
+6mJawSo796H7LUc5xo6YVsftETW1MrdenOdIeiTC/SH6viM+08ZGNVDUdvQpMsd
Xbi5S5wlxRAYhqcWbrkWNeVbafxChSsVeXSUnu//XBFxO33kCYgFmcui2LR2gUOB
5+3IynT6DesWkxUbZbA67ogS4gEfMwp5n/vMQAoCfF8MLbb+LGnOID4fD/ZunncY
lI1XNLhe1Egc5nzQTI2p55AtJmhkDAS5NwpBad/+1PGQvkMKpE3BPHNB/KLTVeGB
2mrThCdCQMn6ASXANGiIheBJHDjA0phi2XE/7gr4LZ5tXQ4vnqO/dWjpKAtJkQJ+
vLqQRFboIsJRm8GzPgL3fnIFmrr2r1S8OMdFRJzunMKDfUAhtm65Uh3k3BushszW
dR61IhLu7cNZjxE4TCwUPTODFODjclGcLHcUOWRv+VlBon/VkDn463w6+giE5C+W
n1vLImK8tvFi+el9/zlqG5IFuaWInKF5hmAlx//A85NaYW2sLTzWv2krY+/OVIU4
SJ6hl2aECG5vf6Ixf4Y9koY8kkTqjfsyVd9COJ3FzLJDgu674ZGqGPtkzlY9nA4N
9IXIWEgHDbhUiJ7Svj2IWUl7SvSZophHZCPxP5YSJjfuVqZqKL03ehU73qjsNl0k
TJyX01CrJk4H0BM5TnHlIiNn7wujMSarIq57tps9lvcsPk4PLjsMS7At622gw93M
/LHlUkd5PTUFmnaaIgYKrGgQG7zmEh0OpBBMTctGCYReDTpc246e9Q9eXqQuXSOI
0dqwh2ksKncZ1nVAgJn7euMF5KAgCqBu+MRW4TL+5Y5xTFT1FKnZRMPgvKq6Ap8p
bTlBS4EJt//lAXDRR2iTF1ofwM08bstPShoPFRalIGh4eLhL5kIrj15kkTyTeIYY
wU91ovQTxYYSkfU6eLy7rHbf+jwwIcTjtTGwm3F7/ubvP/yH9eaz/QOpNAn8yQLI
BKdxgRhJaXVsGWYlFxaDTf662WzJ4ShNNZ5dkkL4yZpxuX5cTHpmECIQ2R64je3s
fSK5Q8dalyM4ro1NQilmtPwc4QCRHs8Lyu7Uqmf22ILRBWwMA0DZHjKAVfMsdXAV
mSTbEKh6gqCxDqUkasMFNzVPVqbrTf6L0/Nb1FiKi/MONeUQGw9BJQT9XlFEvW2I
gZn6rUv/38PT33O8soseF4YbZ3mp4kfTGYFTULprVYsXnLZUFWJeIrDjMtb5MlPc
aDMQjNAEzL4qq5SQDBl7X0iwfYKHWsTguxZC+CkFUBCtuly1FhvEv+mLao6T/4cH
YT0EqGKU8IRRlCagohNnoh5R7nI04PZFMjDFyZ+8uME79ClfnLMnY4WmD4ignqhO
OIDgk/o1UD6Iog60DjGM7JN6pBtTu6hh0aaYXI5J68pKeE7MBQXm/EyZt9a5JaBD
Laf3ciRSLwRCiwZ5s26KeEw6BLifbTmr9pIbej4yt7BPw7Ah82wxnvUhqQC9EWm3
JuWYJOPL/x6jaWklEZJS61eVgNjRODogyTLUis90cp2xck2lvDSbaWrVaOdfIVQc
3nFgDoNGIEvBNk2DMoYTwtR/bS9nWTUyqnQUBham73x8RM2gQa0/1Rh9gW0fXp1O
/wVDKlCEQfFMk6D7/7OpxFLCD4abqpPpczBqqKQ5xaXV4+B6bmwjmmnIPoAIkKYh
B949htxwdR5ecSmnxAMoV0+c9jSqhQ75YRVH0whhe/r7Pa5Hp5EHtASAlRqPYa0Y
2234dHuJtmLhubsCP1ft5pU2nII0dbtUCDcQQVzlFUcjD+n+XsmfKLUEux2mCR2O
z8b+VHRtm6t8YakUHDis7be79ZDcftkpseQUIYFwxaupOk0t2iV7QlovQxkXvq5M
r8t4obeKHrvwlDi3i2jnoLyHlGTZx+4RjarfwvV3MZTj685UgwWfvxWA1a5uqxTu
ouHbxGGR0XEuIV1vUfrtv82LZvMuXcNhIy7sLVdsPejR5j7SYsQ8/1CTMTh4B0H7
S+zAgL+Zk4rs6NaGmpo3UxcIrnpbTeV1GzMePaYe40/sjEl2TnIYy89gy80XqeJF
nNEdNsazMejrqXBKzps51VL1eEalV2Oa80M3TuYOMcbwKF0RQ6lDHrfmhXudMrtC
vmPxxp4p3rje/Y2Cf+9T5um67bGGGiu3EIdmLurAqS8TMshnY/OUXue9coRzi2t1
kfxmi4EespsaQ+fdazouQduAOHnZJ2a+ugoz8G3GzWHsOVjTF+vjoqAo+TpLAU0D
EgoTqHbvxQh2XOCw0nRJ4sYClNPU4fQzwVHTLWHtguI2N+w+Tz68gsE0TQgSDacS
s3ALJH6GrE4wFqESwWR3VkT3ZbzN2408oOcs3Q1kewMHAC0rqD/klviIG5BcKKIf
xaTuGsNX2gqzPBE/h4o8eHhlElTvROvM6gojWbllG2K3Yk0rgmOzC17Bg6i/lOvs
sqh6vsm/grR+Am5C0saaFvqWnVbr0rKy9Nq8NC3KZWNYi70JWyP1IBSf5O9ow4rD
y2cWwTSoCeUTDbS2aEOa5KWzmzevT0GiDe9bCHx1b26+UH0VLlPBPHfT16S2VkTL
W/UdhecsVJBTK9HtEoRSUlO1fWFfUYYultthI0Da8hdxEVEFZM0e9vJEfgXiInPZ
gWdJx+Zvj8LbFbO+krBzQZHYUZqSJOly4qmmdK8d1wKm7vSfHGtcXFGS1UCs4H0G
3MG5ICorCkzAsvMiMojdCS+UuNtUBf/jPlqdUEvlWdHyqF3t9NdyJER6jiq5hang
ye6dffXLM5KqbUKyWzcINgbuoRfXVdiR2EoSxa0dCQjB6+IraRshPZu+H2sJwMuS
vla6WzPjafF3vkE6u2iND6zPmI0fE9inkXXjrs0GzVEKHEW7c04FyheyBOpiMn6/
mM9Xh/3TuTIE/uRZ6cdsite4FxQwzH92MomE6IdgdchEL7fxlUhMqmEmSwzqjZWV
hbOudeJ5/Svk9dK9F9Fne9VhT7bkdHoWusQNh2EknegKC0FDIhoucJbnga5IA+Ba
4NmCdu8JB8vTx0e0FbfSIK/53krzrv1C4DwefiBHb4j9mHG2APx0Oz17QC+jx+qs
pqyepkAO+rmwboer8UqsG8XUKpcvyWQai5AkpvyMfxUongvktSEIuUxmKnbcN5m7
fCmQTzAs5ATJblH6TI4j7qXDawzPk0FR1edBoJpRphUsDImL22xm5Ae8YJ9M2KPH
bFAfBLZTO0Ngjx7EgrzOmUq+FuihUqbSclc219SgVBol2MxRuC6TJeKFRikHmvcB
lyZnBYNmuU9HoMTP2jbdUGNXjtYAaKV6ED1RZzqn4odBU/SX82UHdov18Wi42RxD
1jlCTjQFcY2/yzubGKz0pJ54mCJhCixwzKh6CLROokpcAlbSs2zdd+ZGU6l0Ll6n
/0st3MazErw8uAvY1KQE5UaD2PKM4LCzFq397B01ZO/ETpD8JKk0cJIMO6t23WnM
5lzoSMeBiu5w3u/QbGewfQH0CXgFPe/n9O5UvkruxnH2jDvA8wsh7RWWNFGM9Si4
q8zqhvZ327CONseKqpwzB0+klITxAxf+fb5CyamK9DRr7aP+X69aAM0Y18lGrAaK
qqUXEfrqrjFbZfbV3o0WzVVO9iXGmgWGuiziBMIWJ4kNy0s8ZWZTHBCiWyRq8Dh+
iEJcrd0g2pX/UVlxmGlsHmBiBB7yDohHeP8jVLYxSSAEqArQhbKoZ3qiqESuAGxY
qPhGgYBu+iSaCFDonwDztfqtEYUpUoW6d3bgvYilDYHzz9YURJYnwmG0jk0HYy9/
4STzALlXU5OXH7g3a+FwGqxZCGKv8Du4u0uOqc9OOzd48ERLvJBOcW2swlvZmucY
dWRlJAlZuakh2D7pynTZpNBQ6v2VGHjPnHqxcuxC42ZjHykoA6+G5QxUd+wSaWk/
j/EFe3rV5k85ARlUBXb8MXIi8Tt/zmP+PKR/hFrBXi2EyV5DlFDrqJBt/+CySVnp
wkjEigVCztN7XVruBQNzSoTifV2SywsO5nyAyC4ueL/JUmbTuTLSKJxnA5fHbm3i
JdvOop6Gw22S8nYGVNhc2Zud26zayjzaWD26W7JR5u/HSCs+SnGMqb9TTGqNAv1Y
NZ+e5/9LeD02z7AHn4ZJNdOh+tib1S0u5bZ2QltZu411fep6bELXZX15XdtSXKeq
qZZEExbmMDRTRoTfCHUUxiehFpJ/BMSJ11eBbMEGq/LcViHN3AVxf0+rkyaOXYx6
LEjTb/bVDcS3E0BQsMFCuv7B56suTBSZKD6soe1GdDrKvuimgTPChLfkXMmGwBnN
J6b8Kny9lul4JRGduZ8RYfDlDMntYO0rBtUPhj0e4XpZKN9vMH31OIaQHVbRZLbg
ATr8o6xTHlU1/Nz4XSK4UrKzo3j+27jT6kOOSTbNK5OAM38WiW49N+jQdKPE6mWR
9U+oabePvPkAAdQbGUPtQ4fTX+JF4Cdxe8P4Z48OX47uqMB7CH1GgGH0Uy1Pryio
5C+7+RoCD9XStYCqNzAnxyXSOQf5gaNA2iC2mOJDBTnowDjBCDS/1nI4flihgArv
g/4qcOq+miBN/7EnbFNEbhjDvLsOUsIzITnHLbwe4Y+QzS5FoTWnm7g49Aepo470
TfSNA5MSnMdjjarW++BqJkD/WT759o3BM+s2Q+u1Y148E0cQQqrhyfqBnQ0w2LMK
GIVL9pprbjuVrgJI1Aoh1g2CgeIBPw0GL9j+1y9hZfG/cqnPHfM6ZFkrATQfw2II
9YKhZAhikj/qLutf6l8sEXmE9IhAS1WGPjCVKtsKKtQ/ex2xg/ZmPoR1dbM5Ham0
KjA94o+TJOW6kAHPZijA6mL6HN2eESSHTGvjb3Phmox2N6hULS7SX/ha7ET93QNb
nePRE+0udYcoW7eeWJ0PLSPwxtrPndjxjXDQb+2fJ30HTFbt2Ae1Cw/i0NHZcNbK
BO98vAdCtQXcaOV09RrmsA89Cu78Zz4nUuMj9xbVd4YFbvEb2lg3dyoNrqOWii6I
E3Nbt7+fBLtIBFBVBpvPR0kkn/JuwRIV7vjmd6hKPl59jwsaT0r0YwulftS/vyVb
i8Os/zsQzgFAUkR0+6gMwPKE6FVvctvCM9AIm2uLR0OL9pTgJK3CFMrsid2u4Pmo
4pVsZ+/dT0QsEi/PAb+wynJ2SqcDNWyYRpgn12IqJKqsS1LhzWAoPIxZQlFyqqbh
S/1IrFiIsTP3+MrcIijrcAhkQsR4A48PugEbEMC9c3AErzpZUBM+NupalyjU5KC4
4UK4BVjxaMhuC/5wjfziUzZHv27pMo5V4GvAy4CQ9AN8Tos0G2xrOF6Bnf9zZg5L
ekI1Rybf5XUewKe5VLFiypOEMyCyBDg2bGaId4eovewZrW+lhpxgARpoTicUhDL8
xyQd8A0HsyU0iJ+1CMK3V8t+HzeIZWsNtIR/6F8sgNwV8+T46DA+9p9EawLybrUV
c0qXwMEma0FrQj2CgdFHwk6v3tj0Mez0mI+Umrh3UCAZ2EWf5MUQWVvKrPzQ/jYu
jfnBXi5PxyJ6zRoH7wjslJ8L0K0/mU8jEtSi6mNjnI+Ahzfg2Fi4xkFvK2toMNxs
ZpOSGFkbemre95GyT7FXF/rX5mkq5B7prj8nXiUmTCNVLS4BXbTBf54lKUtKd+mL
c8TDKAhYEQ36zEXV9DXYieHSr50HOqXMi0oMXsdF2mQ5bfqPsh2tSqhkBLOtHgd+
stwFsZTssFlc3Un37ysgLixVf4HpHC1YtHuTxAjnoFOlEBXuJtt5Ss22kKJu4KJm
c/gGBPpy1JeJHDlnpkaH8vRlYiRt/j6CYXaCbk4jZ95R0OKyiBaPj6ol/2TXAMGk
8RX7PRSWzM2Be4HZz8pW+kRZDyeQg2c905WcA2+lcGIVQlqaB8ahcMRSylU0C4vc
U9T6Di338gu0KjSQi38X2zrP2nC46JPZc55JxIkktAww2fYBa9tjLWgmsGmRYqk9
Ia94DQonW2GheE47saoYq28WotI/QfjaVpET1SJKGNpvS0SCwnd4U8h8luTjZVEC
JJJhbTZ2mSs5Y1nc9xds1IzPaHZDAdYFrxFRyMIK77BGq50yNNbgcR0C1fwj+y/k
biSf8SJn2A1+apyalupd3tl26Jf9r/h7nkMDtNsa0ChW8shHZFGB6gvgc7899er9
EZ2cLhqiN3b6j0Dsk5Y1NhyNHWovMjfivk+HMJDQNSa43IWnZAxdr5j8KvwlQ8Xd
76uuz5Dvz74JIgaixybZllvr3Fmk532YNkVXfSK18r8vt5NFiVKPEe+ND/gx9ogU
hDH7GKB3mo5FvO9goF2hLumx/83fP9ZW9xcWei1qvudwo6z0lyf4Gjuew/AOUOSZ
4hyDUhVaxfybfIbtMdBcKuEI/44mx2+uvsTR3bumIwtLYcCVMLj29bMDVh+h0Aso
DTJ6oDu/Y9BqW91q7Lx2EvzlAbaJOo/osqnPGL2tl9pBY1g+8n4LsQ1/Ntt6UNTa
wUH7q8B3FlrJQCWEq5CqSdKDaCTmxC8eRlZYwtE6KH0wdvEp+K5kTOigPEJ0RScL
6RtJCprH+O/IwmeHi99N99U+jrjBIwkKT9WdVT6eeCk0iaHIpz/ED0U1XVgpch8D
TZI4IDXKuaXeQg+d9XzMTqeJlOnf+01zl+NlKGmbSQy0NAAgWJZq/eeZr3uB/UKG
q/5vKVwepu0kU68K/6bObubfAkJ/bpJZg0JMjd8iBUGpndm2YaR/Aee4FoAgd0Xc
yZO9jfv3WnwL1XFwAaWRIYQ1ci5k7ZLmZ2Ta2EIMkn/JR14K23K85qFptQDZ1O9M
O3LRGQ8vC//3obWwLvgd6fJcCFhyChVt/aH1gumLEK9Zsj6/UpVt3o67mINe5QBC
d2CBsDbLksa8+xhEJ8I7gHIz8fd5s8TH8BHxArT2IJCEniiVzEzj/XfwehTO1teX
pIEIIL1N0Lc0EOBGsgJwqrHthTyBStl9yHx+qizDopOChwklkYPI7d1yopOfc5F4
pErYH8GC0/4NW3DEsJd4PIXmkFpnpVsseQ/64ULZA5x6x2EI4Jn47ATmY0aVR5+o
qp5MgoWfFmXUShqH0W3ByxtMj7dm9x71UYba6v7ytp3XAq+U0xX/PrAr+T63E1X3
SQraf4RGjj6zktWlKVpEuAxH0MRlm39vupeZ1XJBQwMVrQlr8UwExhp6tqJemb4G
OOLD0QW6yoQV/sSEoMCa7lXLkRibb/IBofwI3q61Y0aUhRHRGJw1DV6FvQbiBmNo
pJTmH2kwRHuj4SvOqoMnnaZIJkyuGR25s8tobXTPQgK/2OhJNRsyERs2tR39qqlV
Q9J1kGJv10/I53j9j8bG5zMOLROiGUuZ+WO4H/PyUl5irNsdNi6/7Z/ezC5PwKoK
DlyUCI5UnoIKok/TnFJU3jH97x4qAL0KowPW+Hi55jxh006YXtzSU0l+/CN6duh8
3adW4Tl8EIXszDn3sMW4LkQcQB74wciI/LU6ORmv1hg4kt2XD5a5AHfPqjh9yaoD
eCPCS9YAsHOdvVH5BVK3kkn++5TV+I7G2FNdjUVXEyRWmZw47BsbbOuifW1XdDCc
6EQc0pB0A/ss53bMLsUYDKvzPdhsVrn4vHxD+1C8Na8F8AG78AkzNgxewTQ8Yf0P
QtG79gpCQcTLw16mgXl+H0/1NoDrK5LiS+NphHMor9qpWUhy+UVVdyZTc9ChrV10
IPgQbwmNEh90fS8p1Hutto5+Ot/eNeo99MdpFbtJSP9qZbaeIktxW6c/Wx8pnwk8
pTCO8lv7hzmARIG8bmnplNiuzo41vl0OfPCHRnTEuX3Jz3hgFiSmS45zZ96zoFdS
3yKKht7b2mYXjvZU357xoNTDH6yJ+gRKLcdef0B9R9NogPN6NsD56sLPQgR5usy6
YWnWzkASF5rcKK1voh9TPvvoTezRw/uMpgcw1YpqqcoCsZgmFYtLKlLOhSZ++szC
GCGB4rR5elsbaTJ66bFDnF0Q2Xexez9Mq8xXa3uyYCHQGvPQb17hT8yt8hoGb1nQ
fzV7Pqc/L4SKD481FanyBQXEOrDFAPUTz3sFx29/Pmuu+lo4vvR3hb45HpL01R18
WCL3VSl9AL6fvgLURpBqG4kNd5AMi60SVpTu4H72sRYO/hChS1lmgjPQJ9xvzVXl
qvy/pcqid3UNOIQN7XGRHHMJ/dwio/rtiT9EtwhcAQLv8rSip9VGJJgWUcfY5vby
liFiUPBzGpO36rQmg4KGqqL0kCFUiox0gIfnkQeTBsw8CntAuOVYBQiRq/jS+bFi
0ld70hwwBWAtblLW4qBW8Ri+MW4+yKo3z/nxKXWEDUB1evolrw0lvVoTRvMlxgnz
jIX4dxDajqN69wcJsM4az3oBiEeyJdAFcgwEaua2wicu8VggItPyAnJ4RQs7qG3v
MEF0IhCV/XPMhUXms+6QKwvy1JQGSbdzj0Bi62KGsaRQCNc6rYXtb3i5hn4pGwVI
rIPrrWf1bH9zezInhe4psk1tx9697vBnbbXF9Q1IqB7WXSM+VUpj2WKpQfA7qzXC
j3PHzemXe//gHdVp7KTftSUqOfqvWcNkZ5i6av9bJShXCON0d1KnORuejCo/PdBB
JkOgkIjAaR1UPI6PxzhDmBVfH6YwCZE9884JRsnowgeDOTNg2dsjevpRe74s70s3
ecEkFyRFb+kTnyGw5CWE4N7M9MMzYJ/Y/fNiF0nCx3ve6IAJ3+1bgM5Eor0mjQFa
70gG/qIXH/c98H7mx9VwWxKo0pblKJVzxm3OFPCBVuizCd/4V0WHrIa/0OP2xDDL
T+uon8sMHCq1acqCGNYZR+2pgCC2Rz/UkOyH8TNpOJ7+C7boomuO34jvyauYfE42
+JJN4q10ez0sdQoXDUzcgPwacmJz+B7nXhbnDP6D+v0hJvFX1be26lBHCYzbBGTR
ShCqoS1e6ggyPj0yzKueXyG+P1sRHOKDCSrP5loaIT7m4t00lYZxurgxW8JcOfdG
XwNHvqLY2XNOm4YaDabae1dB4BZwhUnmpYJNvjk1pucVPFFW66VE3oFYZAXChXMr
Kac74c2FpEl9+ya5exYnnCMDUhOoHamjHZCjhCsmCghZ8ZPkpYY35GgODaHrHP4t
dh0HlZ5+NEwQig4qBuYCTk/x30MqX96Joz4y9J9qVlmO2oPczjfg4ZedQU5JD/2q
J6NSP8D25IL1M54vbD21ZBQRy3MXttRMDG+0gyAGs0ZzLVZJzhxxSq9Cyh3JlSYH
BwP672JECzPfL0PxwQKKOmpKI9KnePmE9n5HaPLroNE2ZlFZPoi12AoGfZYYpVr0
UYv8D/yJIvQuoTZhUaBF7dIr8cQss5Sxd0lk/hpg2vJt2ZYV4P4tYzptFlmXi2kQ
waRkRHTmh5uTS62JPok29ZPqqzj7GdRv0FDLVgW+qGQQX4u3xGH+GGz+sMMjMi6j
SAlTuqYOOSDA2HR/K+rPHqsPe0I9mESyMzC1K1YmpRvsDqvq9Cm6Rb42+vulVqo4
itq0izxWJ3uQQSkrlPzhCL8YNoKBZdKJuFcCcTF0SMCzDDTFODGXRbOPXTs9eVF5
RJwWCY3lzlC0/wuRzWbqGMxtILWtLBp1wYBD8utwiULVuaaQWjuHHVHhPQOS3UNY
bfX0ShJNo7v+1WXXlbq7tUMdLkCfNEJLHDLvq1Ok+Xuwvq73btLshecujyapsPlM
RHLEmT4xtT7tJW6Wq0WSB7ARhiyiFGnEW4KgUP32dwDX338+V3Zaw4xQ69Jq/xyy
v4+dFTFTVKO+zlgWTY3Eb/AlV50+Y9xeK5r/yZfNspXj1F1Dn0LD9YNUfPrEWDv4
ejzVlJGw59REBt1I0j+ZdYITgu0B56NK2DI4pqqjOn8ZywvSJeUXUhmnXaAxaSp5
TeOlgKY79C+iCiOvh+0/BwXUCLI8GpfkbCu1aR9+ZJk5w0yP8sB/AZaydi9Xl3pM
+p1/unFcdYdyDLNYstDhQHlJK+y3RRLHERxzf3tmNFY8v/E+WurUQT2GXo7WDEH8
R4vQzUhWLSJ8fbvWTth+r7c+1fB8jroi1L+d0RHqdJJUypVVlAAxEWGfi9Dx12nK
sUDPb79dp2b2SaL2/5YITLcsT8CvlQspxDYYOg9spgA+yKgJosGkGyrzZzNdm2Jd
TkoRkvCDAhSU3v3neNkGwILkeK5b8KkQkiMEUVs+XAEv/uuHFd41vA3vXr74ujSj
PElzNcgnxjljWuMeNEXZDNjTwCz9QZznPVb7IJKYLp0w65bM7XPEvFUn23SB/uni
kcGVRVrMdl/vWrLqkRyLWDBFceKtZSLo0Z6U36qFBackqtGnJMXHkzvkelKoTmHm
MAnr/D43kLQhbYVl0P3pbgw2s3/SAbK/jhqdPO+NvGA7SHmXf0uoXgoMYlpBvj7e
DtBpOht2zzpHg6tW6cAJwO9/Eyl+2Naaa+KgpLSZ4NqBvZGqZnXmdF15zCqnvfVQ
uPgAJ7xsSSbnFyabUfVJMCo59otHiQcf1eH9fvuEi8iPM6zFnx+nrSpyX7XLTGtn
dMz8+I2cy6iUl7oTbYptqlZroAN4gX8kfroTKZ04PG0mlRDbkwTtwFFwC+TmdLgC
Lr9DEEOeZS3k5HvUmptstB3Vcw6tsKr3KyVymupH5seZNY69Ao/bj4dFnjWXQ5+f
9aLBb1zRS69RWwx0bfE9Dhqmb4bCR5v4UYRnrdkohOhB5RKSjgVOemC3WX1ac4RH
gtL6oxvAj6xHI8xg8k6ET7wRC0XjcwNhRmWushq1vKq4Ph58czzB9onJwQ/EnRbT
YjmVutiBS1GfEfjcmM5ON872BgOr0AWj9Cle8NIi8pkKvt1bp7lPcv8Nq4oQt9f/
bFnFT1xv//6RRNJa9g1Dh8Qfj/85/C1ktvpgQux16EMy6U0+KpgGwnvFHxo2Wqjh
2hp6q1c21Qc7Wlx5KFnuCQ7Jocrdv0M++nh/sDsXjYuCpugrVgSBC6erlOvY3nvP
JIxgwIs3b6NlcLCmJ4hqddyq0iRr1vyP/y+Ubmmt8/YQ2tnNOaMWZCYiE+0cgAEZ
savlSbz6RmFAgWxAkcf4H7BX7EFO4+LoUDjN1DUXGSVqQt/DJcFraJ76MWNlxIsI
QPIV+r7h3g0V0G86wsxGt8ZgFw/2s/5IGYduFpoWffEmnTG7vpgMhIjIkB6sE9Xk
fof6ipjEMrrWFUUBWOL1ut7IVChKCGOgCJCMKdrwUXyHZ6krPkgKvKclyhlhB43d
feZKtejgKOAK0oIDtPhRYxC14haGHm0fUCfgZFLJzgsvRI1knsPc7pcDemUozvIX
ZlN3KCExi3j/Gw2gIYXZP4CMbG0dvVGsuRupnNLHIlm0QmLh2wnMaUaS753Yox6l
MYKSrjWglj6KH6dz/VzeUInBlKCincgoZ5dYwyR0MxZAg6ul0pedAr+VjSMvSm7L
Fs9XXLR+fZsv5GO+L6MFCzH2pjL76KL+g+MBWQ2AIDFHhc3iYp3w+iEfJjOhFmzy
nHtS2fTnfhLiljUJm1HylUv6iQQFij2wFMu4SGnyCpLwpvfcq0W8VkAn3KJ29XOx
u5Y2E9s7Viq7z0G6N7hamEPfB/P0Qdf9Xd2GAYOh8ti1kKYREpdxSyRgNlmQLevQ
tbm6yqGCwTlmTS+nmP58XlVuIGOt9F60NH1IFULPWYDz4C+yRNxM1V8lPYIF0dKz
hGRFfyfAYlAF+d9793Hp/RK/qlDwUS5HtQGBBRUl7oCPqgqlj05mwC6KsIHtHR8V
XNXq7GBwalVEaj33EP4vCLA6RQ1JNtzqu5QxwxMA1UxAgRJlHiFA6DE6049dktuv
0k6F+iP0DlTfQmmlzuaWHcmLKwvIdDYI2lywF0w4a3Ej742XSTpUC27BRbzWNQuf
QdDeV640HRWqJXpBum518V6PgZjEFiR3e6HPsv/KKKXOT6F20gFPtjmTijQjobdm
CuRTTFkgdI09W5pDl9gXhxNdJyTBSEpmq2aHraSTkzGGG/SGTtAqlQyS6kX4VXKV
kjrlU+PSv9hdWsPI8Ch+5EnLSXOeblYmv/BOSeUUihyPvOZOJIWXd5leQV67BL0w
iR8/RnCtMGeY+y+eXXVTnh8dG/u+cXqmqQkEpjVJecHmzKqbWSkJ6TVdz1uA84cN
nN4CbXU9M0JBEZDtavdFPkBuprmA9KIR6PyoiyjOHTs/Ys8CuXVW0yxnL/vs8/Ox
YUh0oGCsfZknKGaipMWonOKwxZO0oynDWztKc1a7gOHdIkyH7qoCQSRr4LQNCr2X
9h/6eLvzHrKdrdslKAKdxk+KRnyA32zy0ncEOSvpfgFDSxLuL837+n9BwasJvPQO
oWewLNLD3+xVAuRZwiAvm4g0dC+8cCgG0nYD4/WuYQJU0YHndgK1IkKnq8bZe3Sg
ZeAmpNqlT1jwXh/YBVResnWds20iEyTTvpETZzorzYsIOD5T844+ohI2TlEog7hn
t/vnIfBT8kKfjfkPs8TNQXKN1PPmWsojUywWc0hGZvr1jdI4nDz+QT2boWD7QWu7
/fsOEcbiBxZDVm3hH+qJle0owfqz+kFsvJRH86mrDxpTRp+rDpuqd8FGXD8nqrB4
cKfMrkow5XgI3OQulb1OSJ3PHXYlj5tQm11BXU7Ea8yBB81HcIBRutWCulsb1whm
lcuK1v6KfTwpJUsr5EPynDimc6fd4dzQN3by8qYwvlCu5YggYLkDjL/XnYd0PNlf
viQaVg6eAUwLYX86l7NVokRXenMCIzdid+Y6pNa7e6XJZ0wOwN9dct4JhN08/GLr
o21bJdjXVJJAezdfUQQ2qRip2d2p5FFEi3owFwq1ouhQ03w4MFoS/Zg1lPbTFNWc
MFzJE55PnlrzhT+AAMJVB0lYnhws5n9PNwtshHxYcwY00q4vAcbPPFTSqZA2PTe1
6ELBDczJJypi+0p5AYblHXpSXDTqZPbqDhplp56GETeFnhqdna5n3A11VHZVNo2F
joO10y63uMyHqQNzur4AbGEGFYHGJOg4CHKahWdS4xnlY38wgTrGFt2+4cfjw0lN
pZOby3nLYe8mW23Sduh4LxtHHdszsQGOO9I44Kr39FV49rgGMrDpKOWD9ZFZNOUU
lM6DT+/KQ94ZCfR1C0v3RAtzosuzG95IYoc2izI1bv5OrZdg4f+IdT37U5ivhRay
vmT8Sby8m7bMry8eqdQQvae1FngxdwQQI1kZBWAajAK0v0llLOO/GB3ZYqmbrfLl
qoMuByi4QQUOTmHZt7HkQnS5yhN4g1lAc/Whqz39B8l+WyF8uea9wXwVNdvP/LQF
STPcvPBpwqBC3uVjj55F/xIFzKSanQCCCglzCIIObPUHTxDVA3UdS3Qze1U/spu9
yXPnKyvBTZGR4gX9gw+Bd+N2bNG0ty7jMUUMQjuLys/B5qWTl7V4xCtuii5Ti62b
H8/OdinLSMrffDGQQuB31EzY5So7waKKUMyoLDgaTdLSWcIjvyGR3X/yQ4yfpwoT
vGuPvXMsIKYjCeeViVoyw5hXae5t7PySVYaB7WBnsQbXSW5jR429+G00l/nljNmp
wWjNuUa3GEpsOf35+VpKrmLIE8MNqfbiIo0hHVtxyzf4nu2v8fbf0h3+xDzTRvID
hpDMEydyP9hgKP0piTRar7x6AjfoS6nteA4dsjdBp7HJb9aimPA9kFNgzsBdhm9N
JqQJMMTsiAD/MNr9w61n9roXZTubcqRPb7hNZtSOH5mjPktCx5qIv3lFH/S4jOjE
7mz+jbwGowMcd4IseV0jryhaK33T7C5/5VpLmu5Xw4iEZz1ZtkL3u03hXj3KC3EF
0Wi+kF9/sl5fcjtNFAZ2zauL3dQi/E9ZVpXDfcyaWBJZ6+P9jdCpAzBVNRuU3cIA
eaAQ/eIQSI8nkXkA9qpZIAbHan/k9h68jj3KDMbJLQhFbQMDlvkYscg2lHfVLb8X
86VXB8dSBEAVCEL8vLJ+FTl23fwz8xFswjAEOpLGmJ3baKDOUgL8nJiVh/0sKMtw
Ad9Gq7OpumzX63Z5EK9hKPbeSI5x5jszbVuOnj6aAnfm/qjZxtcS0R9YZCXSJi4V
KsWJUNpwH/lKumpGdyPRVOdu88E/556htizIkMf3X5mI1/VGazK5dCIdM+uKTU5w
2RTJSpz2WcADO2ziYcUFPqoSOAuIZK3PjHFL6KARI3+cywcW34iFdkOy8NeCqYf0
6atHZKSKffTpLpoYvQgrsSDtMOqvgUMP/qLxQpxkrD2OC8+ZaXOKARAqwrVCACUv
RUb2h9d8d9ElVLG6svAunu33U9kXvw4Bxs83ZR2AXK/nfYKZjVCxTAwBbCEQ8JZN
9Sx7Y+pJ7YTLMNUoqyTsLNU6MuK7TGXAWkjlgmLpeU9Pk3HYSSWdzgH/b8J9pV7A
mYJyeviWBYxGi7zLxZ5wXjChf+tcgqeinTNts7o1S3NwqEvD2StTEy9+dW9xTM8+
pIUHQ7DRsyzLthhdt8z8oH+yN54zj0VamnGzAclFF25S4b9QP8koJqI2BI9LpFgY
uaCfsXnb89RmqC4Yjq1UA8ruTNlR4AAULGvZxwLtWfoTzoqht5ULQXv2HYgNwfTw
AJak3vI0XqclouNK6i4703Hc4t5RKDF3UCxuVsoa/Ta+NrAneSQy+CgvbuiTlKl/
me1pm0kvNlsaTkcTTT01MQ5mSkWnDPSd0zTjGg4xT/3cZSOWGYowkhK8vKg0mCKD
Wp3tilrz6158MeRqoqYUY6L5dPTLVm8/aHG6Lyul0Zf1Fwpr85M6eTWn4G0ALGzy
uxnS/zu5l1fDQJAjHvRbAQ==
`pragma protect end_protected
