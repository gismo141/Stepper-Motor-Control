// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HJWVHSHdzez1Rzr0A4uT/vpYg96KRa0GXgTaD+2WE8rXCMDdWrehYMtdCsUBAwCX
bVu7gMFhvtl57oceLOUjuqmJjllf0mEkqxSexLy4yiawR6BCZqu0f/n8/tyBO4oZ
lk4UNMRmRQNwSL7OxSNwp6py7ARf2aD3V9IaIYXZI7E=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 8224)
vKeGDoTiioxhVZXZSoNNU/1ZiypL/kYRwRBO0AFBM4pWK76/MEIuM6rgkQ5jIDFV
kq0hs1f6hFrQxeSNJUDwCiUbuJcMJGbNSC4Y/IUEFxXasTxfA+MWsdG6yw4Vk43g
RURtd6bD2GtsXDKEbBUCybTNZgH8h6ehrcYo+IjbwQJnCqGiEZPslWy0v1ibTyRV
3lsuknLcmghrZollhI77nu35yfO2nHgFQUcbaWSnFhPCQ1R98GA4FKvn/3OJBSQU
LA73BtuGfnenBiIxor7xZPkNUUjML/QevvbdHA2HeJ2xAED/pKDkhvnufUPYT2a5
q5JOpI8EIzkE4F4ttW3Fmi2+6reDROafxyk4NcG2s8SDqQKfzwOS3Dog7ix9EOxD
/7JeWopUvZ7GDuMjsCvawrykltkBA5jnuQRWJ1pebtYdOP50QF+yo44lQSU5zT88
gPas7rbVD60b3FBAWt440KwZ7x8ogtj1Xw/I7IjkfOfU419P7dwlVXJmwW8gDTfO
AglO3fXXmUOBCNJwk/sTB5JevdojyDgbf495cSEFQ7NGPwp6ZGksllQ/49OSJkb+
fsdHTNu1X/9J1249f2zdp4URud9yI7jS4ouqAAC+WZOZwcSAUJJwvjJlPtJsAwFb
Ky6y0yXcKicP9dRYeX2IztW40ZuTJ7tpyCBqhL8XuPLk8w9HIcUt2UfCaBAqLW3C
kBZUTqSRkiVpf1HRAHj+jOHoxRBZj8jMFosZ0LQyZYKeYWND0EZUxgbplndElbdr
s4hP2pdh25W0Omt0qdY90XfTvxeLhmbsg/LEv7Ce7rN5P39hS71Sjfpt2FZtSzap
2LHa2/KYSz1uXpyryhk/DBp3LyYceHKU6BM311jR/uNhCQEuA81H++EHYO8UzuFW
/kngoefVwtJpaYH3QxHVfyt+o93YGWTP5ckIrR/Z/6XQYDeTwfSpXROCrHokM2lL
RsKodjpTrcMeeZG8XdbzGJ+5So4MYss3af2Nzf0NQKCsp9+sk3WDGhLCn47k7cn3
X+dPPpTJTsXJus5vkEUnYBhSd9JEr7ZI84UowkkrCl6nNcvOI0vg10YBXg+/Y40o
XqI+uV9fAj5julUtBgto4XNPjrWEW8g1b9q5Yefh217UjRM6BBZVum0d15LxnCHR
b4DmNekFtm+3XcbR5apjcHSoY5rm7SIKJJXxRYGbK81nNj5drZcNf1ut8omp/et3
iwSIZ/KRberLTKu8iAhw8mX6DAZHywcmLiBs20t1KDVmin2ardHwm/2L3/B0V2gq
7s8IDgNoaFU8hvz0qFtOGbcBw49auL9JynRN3UmhrT/DIiOiO7jHuqQmPdoicj+l
ylTFNsyj1mu6KlaQhWiC4+Qmaiwf/Qf4wFzvtboiNjcsfXnfjNHHOSyvlEqhIXRd
WNPlwP6JdYjhMkwD9ltM3ca3RgxXByVAbXqnFP/1xT0nGL3CAzRk+X0e8CjdSzoM
k7x/xuspDggeB3B9jpT8o/Vs1g3Z9NR/7moEFFHlFcFivHsbyofZwNoykCZQPh2N
YLWcaXCcIaVgsSYQPi0NzMWDj6z6wrathSAaQsD2D8cff0SIuhu9/6VruDwyxd0k
QQwZrhcdDhhDfpdxI/HWYjTwLgn2Ld/gSAJM4fbYyk+7N6kgH53tNuANTIIPyjQh
klBlQm5v1+wwkizHF4ouJloiCPvuFVdYCZBqOrgeTr032jjrws7yK0GYxGrC2QlG
EnX2L80D2xiUp7w6r3dDnBBAPDStuagkeyMjGA0sC+FXEhJpGr8haqqxYuOcwqW4
SENLjXMu3H668kvm+LpIDCGZ96HyvED/incAkZB7+Hnitxmj7p3UJTbLnevd+HcX
gqxXswZjwwPArQ5IWAXmHmv6C4BYDaad8zsxcvWxhG2MPy2eykmfnFw4/Tk9ZcMq
beITSGp51ujSag7qaXw84vJYCKD8cysyCffBbmL6vkvcVIP9l3n9KOcfXkr9bR3v
LHouQfOsm0j5HV3K+VukDtjDsQZhpqJU2P93hYlPpX0LTAU3AK1Cj5dimgjgKnwo
BmiSiw9BFG6x/kisefvugPAQfuHQP/W9IBZh8hC7e9j8USz2LfJnxESws2Nc6yCn
1RpCmc35bLoMXniGbXKUucs11zzOpyLX/TmNJIDKD74HOr6BwLH6WYcKsAVf/49y
eXQJBIt88oEzIEIZbRt3CuJuayGBsw8grRpDbBSbwAGfZ3DjXFwU82lRgCQMMZXO
MiJZwhwawa1m+OhreTNlwyqbxCKJTOrHS0OwLuuC2XdSIQ07q1iHqpIpg1R9jYYa
Bs6Bv7njedKAld9zjnAj6hn+PxncZp+ZyPSGBpZYxFY03axsjKYIlE6vOC+fSOet
I55BklxYmmn5u81OM4RqmrlqcCI1RgYgZ2dq1l5RFf5NBKsYpt7777nSu2sdtV3e
2GdlQt9BAHRM8oi7+lrPzbOvde57HJnwbE/Wn68Te+MBgkmhSP4oHkGthXHx2fRl
DBIR/SWTxvspdDnHtf4i+LlcuToyYfKKsjpbNTSl/PU8Qm6xhN4he9fFYLiqdKR4
5osxgA55eA3oSHqBFNRZL5gNgbR2FhgXwSGYrRMd2lB2Q3zUfW4FfkyUeaVLunS3
ui4XB+iAfFJMSE6G8heg4jO5XB48vlfGxj5AmHsKi4z0Q7oXc6LJ8jLShZRwXIAj
BEVERLFEtCdBV+8+w4eSp8B7SK64ucCGN7387D7DHNGJ2krFGo/RiWWicLcwozHr
bDaXtCgO+CMVtaoXCu9AQZxH44Y/1m+kSfksgNnupTYnj61TIBK8xGgrnPCd7rSb
rhIfyWjtRVlz0kEyP2DR/DeDHXeper2OZNe+Ejvk4iOaiM37xJbggePbHlM4Ssy5
DdGie4daEFnE7KWtdY24QY/b141tVF2M0/+Q9jHEE7JaCqvV1Dg89qgKAciswIyL
8Tngr0bBUZPrbUv5wO+DF505G92ekJSmue+r+UA7bNIO2P5gsb3S85IMiLlhRHqn
us04LhQ8bHZjfto1DaxqNMGPAGMLRFd5YpUxTiOcH/pb72y55KuuPDaUFZ4XqR1B
HzbQGhM+KtYregB2mvhWnY3ybMlHqHl3hlHZQqXFasSWypqkBedXanrej23y8OaI
hj6IYAvfI4/6S9qxxPmJkjYGFlsKSjZEpLMKa5uXE3QVhdsKxwdn9IyHzUKQnPk/
pTVPWu8GXsNuB8w6erIUCxlVyormwjArtzBJUOaCLIC9JR/2n/JgBOHAgr6Glole
e65Ve/wodAKwD2E0ktWqnB/QTj3Xr7Ug4nof4jcYuas8w/xjPCJNEkPr/xPgQcIH
Ynyfq7JgEGXxKK85wgLk76/zSlsmbkpSA/NF/nuZW2NP9ujU8Mcfdi5BnkgE2BsE
oa3Xz1s6K17ewxhTiYBcsBfHf4GgvLsjbn5Mc9oEcuzHUyE8i+jhS6ifuDuhai4g
mUO+6DjgAZ3CLyHm+CvSAbkSZHelKmbbq3hYwJ+4slxgIHe5cXhzoqgI7w9EXiy/
qtFzd6rHbXkfzgfM/oDeo6eK/C6HajIHHcxilhGabWUBkTsTFPoVdx6SY4QC4R85
2rtryYygktlNWJePjR+DziotNYIU/qoUiYcG59TivZjZdW/frZ9+baKtr+MXK2P9
+wFWJk0qFHbhUZLlphl21ttRwo6NW56NDd3Xgj6iC3yRUI50CE/8CbVWGRLl5TD2
73JNvWwV5E/gjnVLV1u2Qrp5zNuQkruImNqA3bATfGgUUQgtN5rVWGNKbBSaBHAk
Ki8HvknUGM0B/ZCayaJklQCAO95fqL7KGDclfngw/TFGe9boetWevfFQOmxLZs2K
6xPj4kzZTV2v/vTaxZxgU1Tt4CciXa/y8FGWIyZ74l77Nzo7nEr/layZeBd/zET+
UU7rdITTqqXdW93WkOdmrdiJ+va/cLPhbO8GSVQ3dFLd+DFrpchQOkSt19f/ipBR
2QG+u63yrOIluGSoJgQTshm8PAaESe9UXiaum6G1EWHRouYZ+Bh0Vk+x9E0PwVlm
jX/E41I9J7md32O1+yfXqQZZeK3+nmN+t6QAcJ4KgI7LYc9uv/u/Gz5L4Nd2wYcv
NxK5R5PIn4KteCZS5UeIqS2EiiCPreDdsf/R/hs5XtXBQIeEnYf0ilTDzWYjxVzX
YiEwMSly2TKtzAoTb9vUjOJObIHIB4BkLiwx0G6tpV2KTJiC6p9TN8913nNWQCAK
AOEf+4d+wdvLBSHCYpCNh9dBlsi2RdnodEXAIsN44kVP43+to25CCfXgqQRU0NF3
D2RuF2Z5keG24+inucs+6dixNP8mnGwMfn7gUMRc1yDgkAMcLkNRrRDd77IatPfM
/D/pa0bvqVZmsNzIrYFn0yyQiwHW721yaoMqAQt5e5oPYyjN286IQ5mrCl24BHBb
B0hBSA3+YPZkriwnszEvwLLlCwR8IKRdYA9wBn0redHPvQ3jheX35/XO77BhxMdy
l2gurHpqDjsd6DZS7uF65Y1bdcbldh8Lk0PKBKmsOPdbcsbqUnK1qwYNvnMRfUTU
3UFWUS7pNmHaHhPj6jjQhW+c8iQZGQfRQuCbPC4UE9OboP5EhQwbZOVqzu6qVsmU
Kzn+1HHMje5COK/0oMgVlmWozLF1bMNlZgya3RKSiQKBluB63hlrk1cLiNkmERpZ
KPReYaur9ffzd5uv0cd6goJ2rBckLT9RtenVLeRmdJ1Z2ETD5WkQW1nH5wZMmtml
0LAxk94RuJDTbRvasYYZOsvo9H32ZEJOfTll8HQK5q5kXMvo+yOBsWWCxsxJ2lno
uHHOQxw3GQLD+xMg8M8oZx8uCK5K9I/IH+dvsrSpvYtXFbjik73CGTmhvtam1U58
XBUG7j50TYIC/5EEkQNxAnxxU5i7cmPT0beopCeP4IomXLHy1pJQq6wXNYO+TK/1
fhN+Vkzn84BZUVEoD5Ax2lWcg0k96NTx/NlmjvWEjE8yMwgA6oACcWv2X55ZPB05
4esuYIWCcH4tHoDaGCj5MB0URaTK56Z3mvGFu5TIKo14oTPUXm7EeDyZepdZob/D
JpMDtyZwW2KdawzoWHWevEAxOcskuQbYv3/cdw47ADyd9msHHAjZ1b0Xn72hnND0
OcBirUgFSH3ef4sYWmwaw8YoMZov/qSfoo+QlXiNGAf5u5vTq1d5lIO9lnN4Hh9N
0mtncmqhMLmr7kkaaefYninrA1zjsFijO6iYC5JsY0E7cPhDibemD8+FWIGL91Ud
Tpyqy5QItzpuP/VD8NfQ7dRgm8Xak0vS6X8Ab17wLjL2ijxMbv5d+oVCvEYjz9wp
fb/cuWN7+tUJtarA8KvsJ96cmM5tpibekIwaNb+2Ah6ZNreg3oQpsyQB5IoxItG8
28Rz8DOjIwLLmJYh9/hJQYnkd8RN3rbC6xvbUMpQSWgaBGYR9u+9pHPuG5WSLPHs
BB7WuKPi/1mBX0uRKWT1XrfLAzVkoIA0xZXbiAZh98LT43gHQChrE9LVmSFDVChT
T+LXYmoGRx2lWMKry9jckQ9XxXHlbELkao/L/PCUoU9SwOyx4FEMAaMQQm5mSyOo
UZl772u+2qUavs8sU0tz4z4jN7JxDh04E1oQ0Jdb33hewIyOjBSK+TUDTA0Owj5A
Tc7N5tX1svHhH20ijdROZfoEPCKfO4Gh70UgsGoBRtzus+btAkSuDIlYob+vIFT3
M2q37LQAliOeksXK0rUbfTC8Z9Pk3Z2qF82LwJ4DW1py/0pHVfakdCCTBXJFilkt
OB0uczy7Wwf4KQzw1BEaOV+/i24t3GkPtFN6axTn5NkedVbutkoEwYmD1eXOoU0J
vxd/ufMM8ATHEh4nEgBir+P0zH3DPd3dD2ydOv4qFaJ7Mq4j4v1HrdurQ5dI0p21
6xtB/qgToJTnJczf/oMwA42cD1iWrYfHNqoNOVHmFPdm4M0l2cHfIE60VCFmdiAk
FCyuKcB9QH6H7v8o+q2q/RI5gxXPI1cLP9KHAPl7rey392yUzHxoukwkbLEDR7js
EwvpwOKQQk1Ew/6o13FVpODPzNKSjyHIDq/Jdob9EYnPmtSJ0t84FZDzUuJfVK1r
txyoEc9zKvFTNoWjM89tpor7QwZMl3Bj0S5vc4YW2beO9HZKb27QdvauZu8cdSQu
zZSYMn2mUDcYXfFG0CQpEi9TgG/9TpLuxeYCNYxCZUnabGYioBB9gyT27ohXfiqO
qIhqH/hctkleCagABQJteWyDCkClYPosiDY7ZMCc+VYNCJVbqSzQRitJcFkhDpSV
YOuIQcRVllqSKAxowbiLkqRbaUJJCnPu4o6MbJP2nu96arf9bd2nqQ2fjzDvoX1z
ktAz5phlh37NuFpnkdQRYfZBhpHn+1QLuJ09HT7CHpkyhL5cJzNkpHftY8wMA96A
fn8hUMNe4QDxmyLIWXeossciXkdD5kUeUl0Qcp4+OaSeXgK9q9KSGtbyGucw0X4X
ufgk+gF3Z9GsSZBVxGjzsZG+42XbPIMpjh4MqeBMFrj0mkY/usLZGUsc7hcmaCFk
rI90CDdwM2bg3RnRIjUIDcvqoQsovmaPQAYWvw961BzWmKX/UwWG+UvlYKkPFYr+
fUmi7Wfx09Se6mzQp6QvSSjm7jRsL5qhE4wYY48ssRxO97Q0Q3xKpSpfApt80MPm
ssdK562Ce27k+5V3vD92WnUwJv4TG7Q9SGwwgXk/ODChU0K42fF7OIA6W5yoy54E
buXd6EGZhT5kRq99Heyu01wPTHEFeffA7nMoeJeHEgvivBxvR5nfjRRd+OPtPTzb
DBctwTGcsFYDBMb9p2h7gYRueyHHWe/zKCn2HBxc7YfC6NhlGizEd5KXxBoo25T6
wq3ytOp5i5tOQC/zvCKbZtbrmlRvYE1fXWQYITgsr8do99crZSNB0cE84k21iHK1
y1qwM9pI4FiHiweaRBy17GT5m0E2JrZlpiRdAme4gS4yyaXEOhGWgGmJAtRqr9Cm
oYzdsJnVWkdAYTKUH6RKK0od2NMSAOiotsFRIvnRtJj8451qExBfzG3TJ9sgSAic
Uay+i7uJMR6Sl5LIMCv9c0uRbzdz9IpNvvn1kR/uizFmPiOiAYBmKvX1gavz9cjO
fZ5iCihxdEp8wah1NaUHQAfyzq15MsUzCtEnrK+myDfgWtw+ZbPy5eFPdraeWILk
nymWRFn6LqmDX8u62BzR+nioBaF465VF/IHPP5CbiZlbpOWtmVfJBEZd9WwRjdgI
GgREhjCttz/k/F7l+WivCQxqwVatE49CM5fz0JyZU5exiYnIRnhl79B29XNYZbyI
8UbuQOtEq3rSx3TIfuhdRcSwso7vpv2L5hb2hfrl4HGXnQGBZqphfBo+QELOfrrp
15rr3Z46MCGq6M73DyqhDqrlyVSEgiyORm7wNT+EavN8PGQhIeTWDO3SfIl7y/ef
PYS2giJdBh7VQUVQnD6fsuxB35U2qF/0aeUgjtHiWm826tq6d9fWDMW6VX+E0mF1
bnhOt/y/O7BxOZ74OjMtfplr1hVJle19xzhxBECGgN0SpjIZuR//TJaZzNA5b9iZ
JLjiOgNDcyLmgQw/jyVOT2B/WNzQAzCJWT8Kns34mEggOKWT9wC6vt2RjEEy8R0L
i6lf2RG5wGxDhONv9LX2yB/3uXpP/Javd2wbPQLbaH3lOMBkBf3T1eLwdDcGZFZI
JJQXqm4gEIdgye3feF0Ni12/mevIjj3cq0w8P6lsQQ5t1O7Fhh1Wh9OphQ6gHTkc
AGOGEEahtblQi0GX+cYrrBbFl1GR/znsolp5JWonLTOA6o0+IFpINU9clma/TBeQ
9+ZrQwosNS8Nm0jzZ+NCSW272L7z8b3hty6/4I2FWdz/zUufsE6sMpF1vHzU6XHi
+ghOCc7RiushMRWynXHULnqtHQOwwP6oUoh/q2LfkXjgTDbC+ZbTDKueyvy4Z5AV
Y9ylkzC+4THrC7xRPlaKLLPvje+YYmoYPJI173yPSXWsGHNTQFyISjw733m2TZw2
cUf+fbyW4zmh9CL1dfAUeLgMxeY/BbhI87+vdfvzP/DsG9/Uzin1xM+Ju2e/23eQ
ApEDNsqdJNETzXWp/IhS9DGmkkOXHCVMfSKn6kY6FrUMOfmy6mnRqaUeVg54MOuE
tKnZt0ajgOXWZRCT5f6ro/cFVVRvkeS4OhJ+IWRdJp2s9ucp7cInV1auTKXTRowg
79Zgost1KEgZknXmML8Zfm8qnqzy0HcZ26QemHcvJW8rQWrQzdJsOiUp+tuxCaBY
P+3inuMWX9dl+uBFrZ8r6+ynh/T+eDDrwEPhdeBlkIKRY+PFQlbL4y8U/gtD3I7B
o7x6pko4ZlgfBVpMzLleHK884/DVDm/Fimhuu8lopm0Qzt69gKVUllWaRAIxa9rE
1XFwjbnxE5JkV1SbsgXwqfkJjK/hNIPJJVEb0iP8Rjs/5rm685ucmZhfyWTS5pCZ
JMbWbNA8WJnxHczCGnchriF6sE+32FwaZvyhliUT9TKErD/hde2lOl83cjx4JS42
788bgPKngwtUkee27y+gmm8WIcwB3v5Ur3lSP7gL9N4G+Xu3wqB6qAPGgNfmV56r
5TlaH+bG3NFrexlBh4wGaFTl9Acmijoux2P92WHdphvt/G7wCekxZODhtZSpDhuC
7ji14XvI3zjaSgP2aJ5YCeuzK3unGztRsU5raGdj95mDpVhQ3SHE9I/BdmCyVkrT
GGUEjwxD+/pmKCB+m+ZOzFz04UYSwH2BYW+k1MMm02lHlOOkdP4mheNSXDk4XG7F
gANZ0NCkZwmFxbAyX2VBJXLxMDseBelv5WU5lOPvOwrCE9Izyyzkh4cvR18m5maf
OxUHV2fLYJ6Nf0Xz50vyjwZUF0AevjXeHFsbOHbwF6I2Z7VeE4bMmkyDtKN0aE9m
j42s4T1AVeF3wk6hYp8tgZJ7vWmw7KwIoIbudxf8S3C4aIlyo7ZAm/U00z6GMADr
NB1JMz4ctmIidRJgfkLGqEQD8TNtgFRjX8ukU9zJY0PMcLeq2rm2bg29Mg3gi2Hx
OUIbM7jxQY+QatBEaLuQ5vmNPsbSzfuA5cFwZRxWNtXohPDCKMr+8XGCrOsTgzmT
QsPSYLdLpXTsz/EXWd1yQl/+OFUL8fV+lnfU0QC8Ru7DeRtac2K+dw8XaF6EPIgW
ETo4DTaodMxbsltxZZtlE4V41/gNlHwpRuf4ygxKfB+MXtSI5H5nhfUUXGHJFnRf
cunEk37ZqVTep4+Q1xNJ9h5jg4yzHHMGPHEPrUM5ZrBKDoKHHQVjEf/+lak+XmNb
eLe06/dMQhr5e9YHxc6t2cZqDwMaqxkhKepqpCst6KCaCQWwRL+34nmnK4ZXibvx
rk8VM4v+BvAfBcqEiiA6tVKmRZPrCYe7IbiA6FYxn9G9uWd+f6lM4O22PWlcev4H
PfNMtFH1Cdwm43GMi5Pq49r15vsZv5pZbeo+ZhFINdY9RCvff9d+neQr1dESgIQ8
Awc01MKXoojtRr7yqE+a7Tvk021DYpLQJo/AjR1WywG8mwBhsj4DcTqqgM5+qRjR
pFlGRreNp2tyegPwVkMizAWEi55SIl/HutjUUcDtYVO280Kayc4Hyep2bwnHPW1L
o7YM6TphWLYRwtnVNOULx1sB+panyI4MIseXCfCgYIy0pq91PuWYQJIbDyzTnA6D
NxvgdMiJzMREnEghNDHN572YNyDdCxG7M5Wv2DSSbRQOJTtFtRse+7xTWF34Cta5
kzcJKo1Re+pUgx/dUrGc/qNQJ1AhhjZ6oISrZX8jzQISPzaaQHi9S+T+qrFzh7ZL
asB2Ly6HbRzE25HoL05bvi7tA05ebr59OwlQP3iyu2gbTZe9yMZIKd1kEd0CKert
zKnyv1pT7Nuwj7YxPwLHtM1DyWZy/ptFnNd18t1qR2eU0LufZiNzcGg6AVBPFm9/
eNm6hVCIx0tkYIzTssv1o4kM5KVj1kuqRxJvOovRtlrW2dxSASEuE7SdA8yH74Yu
uLHHikWeIsjdCnEhsald8s/Ahh1tcc1LdidfXiIT/Wf9Jhcslt4WpGOfO7zfNebq
DS4cce9w4hxO0DG/cLFQMsYVi3YwbpyVN0FegaqZPeuY6hUtrApR9ZyFbyXcfGyr
YdaPd/S6iN0ThXOFD6juhK5HBXO2mXhKmkawgK8r9NhAdfpz5rdFsLW8Q55NIBJo
r40UgZvrgpLs4OhQAUDTf7XWY4ZXBm3eS9Tor9bymIfmtbbkpJxqISJzydr5hrY7
09Va7DlkJXRxsQmb9fe760jD2gKwhzWj27VDRM2duBZOGffg4gOtULCT5UdrFN8B
QrKePnkJZfmPG7SdADw4wdwdsMkwLyU9N+J+aPlLDqeqYflt2+AwIP16Aime3UVl
o4TWEavffrhyYWD6XkgpQfHKxH9cQa4ggUU6Mb1mnNrekQNbxKGNkblk4q+VaHWq
TdaKNSmbZR4a13tN7dZkrMaqQEK9NWhbdhXaRPRnAscEtkV78Z09KRgQXrScA+7e
IkTiscy4/msuWpK+3uBuIkFClMzp+yeKj9QigpFZa+jvi6w0sOuhDbCuaCQLj/5G
MOrYzbKiT/UOm+WtlOUElQbq96kAiXrDwfBJdyE/O6CjLDZyzpjtQHXE7fkFegAs
f/eHzMXXMlomjRAlPxL4j/1GBJlSoR5qA75p0rbtuRSqsCdzTrY4gH4wREZNes6s
APRfkeVxKsDrTVAO4UnPpskze7pLfWLtzqCzB1Lt1TNnfZkANv2mNCJ1/t5WzTUu
uFrsHRdmG0CZCiWHeWs647CENSLcYbPvIms2VXb0vP6mtP2HJr0xBPE2BCEObDZP
g4+OtSthPsi080bnRvxn+gXDp7PoKB1CT8aDF+lNZbh6c9ms9+2fz1ZjxU717Ydf
eHQx/dddW7oLTUeRQ2ockmfS+tpjKEApkYtWc50oWq75AkkvYvtTf2DQlV7kAKsi
lWQ8FEhILyj++ZcRY0eRuA==
`pragma protect end_protected
