// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:47 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nLzwHpEUy6mapWNR8lR333sO1Bk27Cs9mgMhsTnxo6ytbr05ZEiI/F1mcQ97MrmZ
sU0T/HgZAZnsHEDePBQD4Sr4YBu5e84DUwRc0CiNRQvxxC3qnr8x0BEtb2qqSv1g
v5G5GC01vZnd+RoESmr25pQ0++POMYMrtHyKW9ICSZ8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 57696)
ZB9MlikGgaSSrVuxPw2VdzsiGw6PewLzLDj17/izO8iuwY0I3yo0sLKibbb99Ma+
Y8ONTvkQga+X30ilP1NXFPTmIN2l3sRzKOwWPYuGaCIdXfmJB2X4Rcs1OPuHoKM5
BL8w0gLqNRAaGi5YfWklgGLFRGlhigKxSPoi8laNDk0lEEPlD2gXc5yvXfPmE5eY
a/G8E2H8bxz5wohYKup3eHGXqCpIGea8Mdobx17F1Vjc3DAW4GJzoSv5XdIFdukW
toFlE6tpYHXco3MevtBcihq8glf3kaBVo11rAP+/5vws6Gh0Uryz7285jGAG8MAX
+XulZt8WjXJX8ZPEl+Ew6NAM0MkqVysQNITSyL0LoCTKPPZvVOkUDyaOvhWKbxcD
IMoA6i8Y6TzwFzcVUXQeHjCZdM4pZl6R2H4W5+Cw0rt0JWLvbySx3jrg1wh9O9Ew
mUSDhQLzTsFaTz1PkyPpSj54JdiTxVfyPhqgb0/Og3skXwyPTckWmNXTLVtFJ9hm
x53mr+aOPoV6gfahfiVi/SNgqWH3nfkOJApQwO4vcCijdw9xywdq2n8LNX2gOJPg
0jgBempUcSYDnRG3Jf753vlBOm1T58maBsN2MIor/pk59RwMTaxBQh5ZPkneQ4At
AlOrtzAIzaZop18lkkQGZzIlfIofVkjCNyp6uGbHwAstAA/X8u+38hxqskYDHuI9
Wg0Eu+cZFY9lOlWqyc4gkd1Ok5jCM8uxru4A9CNqbMP/mZ6/Sa6Hijv0xUEew1XG
wKm+fXdoeGk3sKFTy8bSktGKajDNuwXwlS2JK0nHm7I1sBnXkMVLTmXokDbradoU
6oOh/RAZcPUHLuV3mqEfwirUfxSWuvv0wPEnikMdFnQOiiJ9aBX2lAmzgKH2cigu
nxGqQ+KM9Bc6ojet9Mhpqw6r1MP7GsY1tkbAhG1jMVWS+qHD2aPU9ce0uNbsmR3+
tfGzlC6yq1QIilrjpTlt/kv9Tk6WeHDQv+IM5LtxUTpC6l8R4u+7P0pmWjqHBpvp
/qkuhOERlVyi96QK6SKHe7gGEtcPzK+urtcxq1oAY870xRHjwQmQUI//xlb8kWqy
sHNpT+Uv/+WHS4I9wOYLR5ijGDg+YnBBu6JkXQS5zMV3ozqvNnS0MDdw+U3mbYzr
N1Jaefb6mVTQbeKaf83WWDFjMabI9iMi8fAi+/FIauEoYF92hiU8McCnF9+57OEm
yfCEWg+XrzMG5k0Lp+RCaS24t8ao7a1BJYV/56/j8TAo76L+/P4Mx8YifkDr+9MX
5lLtY5bdpxNjjqTcMeeCuLGw/SR3vwI+mKsLTdqQczFXQMgaeFIOV0sMmKmB/UfG
3M0l+/zqNutxokP456Xt0w11kN1lXJRWY0EdCCnN55kJNNuDEoVGdz6r3MiVQpEC
f3DXwoXP6PrXQR1GNAgBOGmSuVmzv6rQAxFvo0TRZuSypB8r9THl3CONEFcvD1jW
OCHxEsOYGSrx2/i/Jw6bTMubKNqUgcx0ghyVNsyNxeANw0o8a8bl9QExOVLs0gP1
PaZ+51Ab2w4DcMMNU9qhRNvpjoBkz18LL+Y0b31jlZH8ebdeytzxtG5rlAcf4cnW
LAQSDFwH8WAyJuhuSanbVqt/gZzdl1jFN0C12FI1zUy90RPFiVfO1RdVBhHsqyNx
9Cz26WzvnU9jAJ4s7NpudOqssuUT269R0e/bYMP2kgYwX9f3zgAkLgpF9NOgKObq
zu3mnW7Gv+JQCYD/W6Gacz9R7ZzeKE6/mo33ApAplR7WC1eWYNeZJ3m8spEBSEdC
uHsYeUwNck/G3IcHx09zdp2PAkfs98n7nshfcA27MCAVPL7WFEjwCFD8gIoSTm3L
+h/5iLAsmdgrTEgPtZ660wgE3XNZpbu+l/xA1gckuQFbFNX4jeABSw7X7MyZuKWe
CHZIGAZ3zxNA2ezUUdhegQAaviEOAnJTpOJueeLH2PQnLZ5Ekv747uTwMJrZBKEP
TjPUsmOW29Qgh+t3ceRa8bs7aX/QFahWrQyGW9dS26MXoi+WV0X3zhXYidOdXe1S
/H2UTyignaPn/hazkCTIKjyuZFcsb/c03kCBSZR1MFIf+dkzrF1Z9Ic5USWQ910I
xJ+fJYei2wTJlWlTIMX+KTYNxugYLq6eL8p1M4k4A6D1hT9exTDfkSJ280FZYXof
FKA8msRncyvTm/1zuhxgowgxBRgohFKZdkgxp7U+VkrmOM7ganeGFozBtndEIIna
MBnpIWJLFuxoEci7sft+N4ojpLMrcfbxKKTX8CHfIw7a3+hT38vQ+tw8lfabOlOH
99BiLhet3/f3c1riU36a3dxz5TRBEsB+1g/ahEPribfwhuYF4AAToFPsPgNOnYLe
gFIAWc+zXKit7PLXVl85RWbwemI+CydD2SiDaYFsKYkldtsoxt7raRVFf7nPOW/x
wJW0e1gWDcI9gNunkvDVWgfujL2oPA7X/feeXEjbqEsKkjY4+IJjzfLfkUet3PAU
RinwM3lJQfSJzKyO5KSlPvgWuotTsiwWDbcG1lpOmsz6l8ApbDHaZe73syEVCl7c
Wi8BayU8lLTQgzcS0mbbeFVDcnZHiT9fhw35H08Wxzw5DDKI9kLnawvgarQQdhR+
0OGOXRqEu7K7YY2C2oUzXhANyRRjvC65vCbz+4d0JlvrDwQLeBZbAH/dMhI758GZ
IGx4J4Spnkwg3++oQp7eBHgDRDCmGE8zBimsoq4TrdWkP4e5rhAB4zgTPvKZ/HD6
Cukbrl4pmTyUw5jNP6e/SphaFtqmCCe5wuyXXekQzGn2Bp+VONFMhvFCmddLXcVR
DBRyyigxtdUrLmb/C50RfShI9sBJZXzAcLSLmYjLMYjHvG9jBDn2yITzAqQ5fJMq
LgxbhCSnwoztJSoGwr226tTIzNqnAzPqm6KCuURC3Ben9kSkSgGWG8ANyDA+stWk
H/vwPdz3Nap46/98eonVxg2XMPunVrMCOqthbQgHQuQ8L2lg7TokuXOViBndKdD4
Q1U0xE4lCgnKi8FOaF7looo09JaGaerBvy3jeMsMTQQDWtdo2wUWkzo5mSfVIcUw
M9D9hmKdZfAe+xICb0aOsnI/ukat5Nhzc32rfu9zbkCTR7mIeL4/IqXuNwgjyiMl
xXoYTbf5tdu0jaz9kbzwbQk0aQu5A9wEHmChqRxnNSxi3U2IcXW5w02OFzCwN4uO
/eqg/Iw0+KCbLohnZC+DGbcHHzH04eQK7e96IWPWM0qbL23Cjr7LPEDsPAl/teOq
7YzPaY8haJ30l++MK4a6UEH+67+azSo0s1xh8FeD59dRo6MfqIWenNevB+JBVXDe
INzt10X/8mFMDX+tzWetTYUJ2aP1nuosFjW1rckHts49QC+viR7GmZiQM2Gu4bcO
tH7X8gubcjMbdfY8eyARwS2xcDrUwQ7PMpWjF+I3dvRWql6C3k/OSfRyaqj1Vprr
lHD3e7WrGjF/LU9qOWdOfLbs6dUWZDPj7mxQjNXoqAovT71h6y6+9dqVQHvNzKlc
2rcCLt9CCuCN3lyuE2OxAa87zpRu9k0KgXzt3JCI7sJSj/AH7hOZLXLkMNHy5Gp+
DLWbTxyAT21HOY8MascWi94grbF4Na60YpZfYN5uIEilIK7QMuqCGXvf2GKp7liR
B2QsR9gePyA5pq5maxsHxR6EPixzQ2eVs/VmdQo6m5qEUhnL83qyhyMWlWNZcGzD
N88rlYHYTEQ2SN/ZlG0YvJPQuawHNT/xJIrxC87y761y3sJw3myNCD2E+baTr2xt
URe5Pogfc6Dappe4yUWUbmN67blgVRaD3uqdhssEcFELxk72YkK+rHk/+OhaZQsb
c65LEQ3frj3vrqYGBbx9rnmpWwEGzuFpDygIiwnyklJJMtGbVVlMnpnbUz5rGlq8
xRSaLOoauyqJlj9cEAuLL+c9h+Z9RbqKc1pL31l8s+8iaWZXhAJd767AnIggQdq1
pxahzNfRvk0awGSZ3LZ2OZvW/fS4hdyUpWivJLsB0bY7Zh49qcKHTOiFmnJKNtu8
q2O1sL+jzxIRcpqIqxAxlrIE/25IS1Twtug0ANvsusL1PnaZu8VZ+I4AQoeV1W+p
MeE734lYnRzU8SHHL3IpYGVx2GrNcCrKCZn3tNW7gpEIwT2KujCCSOFn2xajhEsv
rVf+pyBs78K51Ot7lSMVn+xrjk8hm4yCohTNEYFtdmkDQizAXFTXyg0axV84HZcm
FziKrMyyaVEbvIEFbxnedpU3EjqBKro5onv77/0zYjaOGvkMykbB3kVTpDYK9kEQ
xuEMYlodXd7mqRWU432V5wHCXqK0DO32RtrkjHP04ijStOP66W2K5Z+CgjlyIAoD
gChLkfOXWPanOuiHf9rkdhIzVt+gFALgXnO88mAxJCuxViBT7A5LMbSUQ7xlBrQK
H0HBUZCUgfjfloE99xzL67kQV4x8R2UavEnv7gPVQ/n3EE83k1aGauGE8sXUEa3J
SVwxTIrho2jAN6Xjd0G9Ch24hG77lV0i+1cI/PoSj1x7goE5nfInkhtoQwtn/waO
8AjFqYL3xyAGw+aIvvM4Rukesrd5ybfwCXIdLcXflUPHOVdUQUcPSzUn9xyIUFLm
dduxXrNbEyof3YnTWifhiAv2/Ybpb/XEoGtIP2u3v9kevuZISWfqUwEjAFxwpayL
XKar/g27zo8VTcEiny/wsT8vl5SGvGjHDnqKQkEb6sfOjI9wkGy4mFtRelNSHjjq
uWZBZXCX5IMP9x9hXHVi0l7tXZ6EovREqnteKho6B22XQaF6ns2NujBkukNQZvSg
4HttiILFV4KStj0nnOYL4f4ulEK95CDjp8kAv1b3qJKS4SWdEPPQFCafs29Pq8b0
Dqp+P2dFm/enc2a40E6BGQaBacrd7aNKdWWpYwNjoRPWvPeKkCWtqLO2MLeJQKlh
mM2Dh3Cih5mqL2UX/6EBR+Fq4y4wTh0GIpEmhX5pumiEio3kWOmoovE622lbUh4k
4CqvEVvIuIDiFjPjmKo9R/HFR0uq8v1QHf8RKjDxMxG/8YrrdDfkNkXT8W7AXoOz
BDUacTQwbZ+v/qye9GwmkkdfWK95xz3dZf4HgwQ/s7wgvX1ouJCAZb4pihAhh9wX
2G7rwny4QQrUCshhocihZzkI7WXrB3F7jTaYmhNlb4PZ2tZuzmR2Gw4bqNN4w/t2
1A76JphtSCPPZ6HwEplBhNHGwEI2qZ2P3WmpSPiEB3mnfvREvRC4gzzfacvePc1D
Yf+itqmRhRT14Mo52JG5vZyPXja6Br6CvgBdPLjTfOfIDkm1eZoBGnEH5h0D2Zpc
vS88WS3p2pWNWuJsMgXZ+XxyChYpzhozKqfPorasg8lzhPXFRH/RvtLDEkIMAX7e
6ZqdtDQLYm5JP4/K0GTR1QDZBzw5OcawidVnwxEOQWcb+93S6UUUBnBO2wwBK5S4
aZBYPYLLmYJy7uqZuxn+y2TrxEDPf/WvZBfpMy90BS6OMLn6L3UGtoPtTs8PdJ1E
sma0VyIclZBwZJ5OdzhMmhrttnZG871/zny0miJeODXw8Prw94DRvdhMrU+cNf9+
yGVoPgfyNKzelrVniCGLaJTjIygsjkGBSQhZAaAWGlKsjUg05aennY/qPz76e8N6
/6G7X3B9UPEr3w36qPl1pHnBWrnNFHrtgTxVz8IqYm15ZbMZqCJyPZDAfBvQK5KF
09WSDKKPJE/6fQCqSEfptpMxvU73aLCeyfCBiwYnu5aY1OL0D5kfCsYCvkAJZGAJ
SznlD1TYWDU6CgX1h6K9aYsJQ3s1Zevq5+lmIFYjnagvBBpSxLOjKugDyhjCREBK
XlhyhuBi0NO92lpmDyQH8t7dhGnVArWsYnc0EbUrToGuG/0SSgYwY0OqW/JkJh5v
wW3lU8jBQ9hMWZXIeg1RJdSqyVAndCbh3l5JL/7wHfdHynMWn8JZOk3nBntHCTNN
HmPI7mDYsAr9+801ym0j9dPgiyebKwUAQ4e0dLQAvMV4rJD+eTjlHA39v8ohVfTD
oT1qy/+h0NjNvQUmGrbGw/sUfxK3hFzbal/5+LeoV5ed8xyeRFhwFv2mVXeQ1QIO
Z7RhKATY62jisCzA2Pe1tmJG3sHw9Hi/5gRVIi5NARcAyAb7zMYpBY/3kOh+zMK0
CTKbYfJpjeIT3RnJikeF5yg6SKZ9Q2VA5Y6dL5/VUdPBDoxRZznDorfiDaeG/0Iu
SC7rP1fzGP8oz9EZu9zU0QeS0WuXY1Olzrtpf9X17UZ/bjv3Qbyf3vFxJfVNRAtG
4JiFXz+BXKcRIutMiYEyEc2rPwGNZy03NMV/a8sk+7tKQR4zS65HtVCqwQ392GTD
f++OvWJ1WITwgx84cF6Yzq5U31KqxYsFLXWKYKGzu6TY7MmeY2YrqB1fm4p+ABAe
JBmWyUeh/6+YOKNaJgq1SZOzxTcsOaYveSjrYuhEfG2opX186eSDhOzwY6O6/HpG
RpDj+PYq6/35TZsQbyl42Zeuf/rlFZnrYsJ3Bn3bz+UymJ4Gs5fDx0Vs4ggka5sV
Vk+otIOE+rLSZh76cg8PEvzSiQLxM4UMLvV8laG3P/wbLwpNf1onVNAXlnTwLT1B
/mrykvdQo2lJpvL/r3jTBde/aRxIjDRmtalrdgV1IM14R1LbfDt/fog6YevBLhdY
Fva7UiO4a8yNJCFOVVkUOWE5oWAKZGZYnaZ0VLMMuBIZY0YY2lo8Z6NSYdetGN65
BaFbaUYOZmVEiBlvqwyDfFQaIPke4EBG0yx+RnZn79UrUmlqTSNiRXaedU+6AmvA
8tWN3Ueyb8gIAbqbb0qBGjJtKCdf/+HPG6ImnSZ7crK8mWE7nk7ai8ILFgqhW9SV
D2hSBbrFjHBOI5B4M4dVBd+nPpJ4AIei3nHyio34RRmwrIZnPp0pHIZYkiRKZ53I
ME4axAOBAm3D/+83LXqPJd870jVuQnbn9298N0Ffew4reTmlcCep8K3C7ulDY2U9
v1sPMjo3PW06RfLggbCNjA0Rh7f9KY0Gg3R4JHLrRFT5PqsVSFUU54vrwSX/M8Of
YkQ/Eo+Rbp9bZAajmo/vP82awrMCt/4FqKOeOuB3HXHKHyAiKyGKqDwSDEw7vnNZ
+wPWqIyxm4XE12pw+m8h2mvo7Op8JGvZ8tRueBsOkRVq4PXjHtD2Du9j+Wu/gFmR
uZ8tOFQVxGLHl9pRByP8iqD6ozBU163JYgWGdpzIeOBp5d7B7JRwuCSd4vX4yN4l
BCplB9CUjNvN6Bgx7HVOLtf/pCh/BPz9sYSQGtN8jtXW1yPPXaVipb+a68nL6jwj
GLG0ekDsyZU0lpr388LX6yQnkRhw8ze0WIeTeGTDExNTjOVq4oOkVH7sG9xwvkx6
AfdkV78nkP5L6FLxPiQWcg5XmQJ6cz0BM5FVEBt+DVsywVmdHz35IsM4GCiJENJ7
FCswIkxHdUg6mKUDnI4IvECkByZlLPQ2XJrh0sluAiZ7MPFDt4pzRADJQZccyS7w
FFuYvbOuBjZM4gDhRxZdkzeFePc/qyJkUCZLhUiqvfAF3dZwa7Sj6AjkXErd52qj
f0/5B/UjL0G1iT+uPcHRdgaQ+QFAzcU0u1dZVtGbGznBxCiCnng41j2A7kGvm34J
0FAy5LW0sU6jvxOLgqdZu2Yv+9weKQFVKdhV84or1EkWKELpVVjM9IxnlPEMXJVF
wHB0KiVtnEd3agTvkYM6l/luSH72RtAO0odTOQFqpVnRfpbRb3BzD1q2gAumQryg
X1zpJggsyt9cxvolMuWVTShEEJGN7iS180tEVqEpHBSUDzOHFXMpiFXU4gYQ40Iz
qcQOhKfKMHPk6PYCgsXQtTXRX79hlhhHAc0SaXLa0bDqQWDf70B5NHnrRrDZLGO1
aRNLWIxtGsTz8M/3nYfQ9AXe+rrCJUijLzqtnDm8/MYhN+Gl6E7IJqk+L4VYo5Us
1bGxwDzRn33gBOFtFLv+G9G8mprU26So62ZEjvMZ5n9HEZAKnR63LhPeqThybvEp
09IpyFO/tLhj4xrKafafrhPnUn5HNaqUwfCqzR7YskCKG7SheEixRF2OGL6r/dkq
gtsfiuz/vUVvdYa8FEm4ENZF2sxEDg1ZGtg0tdzn4KAGiwU0mHwNjGKNIJPVvVQ+
QnCUJNGsTZUI9f3oX5aBeGD+W5eobtSlKGFVy64It0bZ/5JPg3bTuYk0T8v6rx8z
WuOxBHaFPTNmec4CQAG38T6W1CWwKBV7KHxINiSZo1C8OncWRdsF6DqlJ7+5YW1V
Tth1iRdv0/eUnMORu29aJ3NR/2TN+aVUX/3h06cL1a0PPEFhic+HeER50ocIUhmf
cVCUAiyxJOnhs5BhfDq4knDRFxIcRnFNcskF/mhUE61MasxkL33R62GijaM9+/Tn
nscAaoZNDMZz2AajoV7xA6vA0udRoxVfsdxxZZRrzkroZUfJcr+McWHmLq5wNcY9
WE6YDFz8hs7vx1GqDX3rhsojK4mszwnuGwM0ZTIA4R1PiMcFS3SdqDJRpLDeN77N
DbFPulHisUnEjlX0oaSTvwCtRKN2Ngrr/sPpTZKVyPkYOViryCEY26RnAJ8PEHNa
CuWYmETriKh1PjvJv0ay/hifuddb/JbiUo5ShlPB4fpsJmaqoKu4yO4HyVIb+0vF
eD03TCxeUqtKNfehRMIBHG7s5qtk/8xHneHyvy61R1DNj3oM2qWjmm/8NuydCRRk
XsVOlKd89Gu5fxxLXHkPFexvsP1NdyI+owrk7fEeAAaIo7Ou35nJwa1bdx2RKHjR
xEHtBAeAezaqVxZ5BSEkMNN4uDw/BvIDTRmHWB6Jhhe7tUmIFiGx34C+vIkpw0N4
tnyWaPo3MsiqPMWskbybK1z5zpQYvNHpkC2JQR1VeJ2rD1Y3vfBpu+Vc1LynFrsi
8i+rLm87HP4d2p/OuOy0iBjb21WzfKc6EfZ3yAvJVollVIvoyZUp23x3pxEK65tm
U4z696Ebqdk81DbBsVUZlRFrPTZK8Wjf4EkLKYHRc/bCcBbDZoO3NbWU44WkCtOw
+sJgRqvp4gqIyYlQBFCQPU01te/3B2tQ+TGPuOUhZ28XxpplRf/rMtpTpfeh/UcB
6tC4UV68sM/yQvWF1igwNGPkKqI5aXAhyTNkoK4AyFGC3RpwCg7peGau9xS011ao
P+EuOcy8LV296wRb+tB1mEeo9GOIYveqyXQjwPaq6MhurnCpLK8RSXQ07YyUv+3Z
jy/mQyHe5wiQSJHOUpGgRfPbIwOMxqFwP/vYxSDOLNgPJNcT/m7lTLAbA5Ve0yhF
5X4cPPeOzmkesH0wuI2FXVMTZ0FMUYBwdnUGfTbBzxByWLvgd+xRfJeJ5gAs3wKd
+inGuJJIclfVSb7aQpiM3kxq8HVJ2TjcUqzVTAxaHBgF4dnWin7rz2QyAzli/iiw
9ABOu5LtSqzTMZ+jA9fW6rQNAPxFBJAOgmGXt8NWWsV6XCtf6y6bSxZJpVCbx6Bb
3fsd06bzA2J5N40tHiJrvxB7ZSSzm2Vtq70npP+6tXl34UveJT/ZfZT68ovqTnXi
7oRjsa7j8o0iMDP7w5ZZ2d0I2wV4RRL8GUD0ezFu5k2p3TUTCkBonkZLDJedbqTT
CfT2WNeP9m4ApodZ3/lkm15AGJIPTVkrXH2Gw9OzSamkzSX0QZxPMMmNLY/Kjm2h
O9sTOnHDzuUVpkz5lha5/E6ErtMOCdiCUHdm2mAxR7E9bZf4AHOSRPuwl1E5/7L4
xqgk4d1khzZVSrGxJl1qAM32oEJqSwf3j4bfMjD44JBGbK2/vXiUdEGXn0jczbZt
AEaA8KjWP1M0lcIZuVgmMvmvlzJKpSezm+vkjEVYr4NUbiB/owlJEGJvzOFJa0zr
VHENQEYSl9++qRiqy7YWy7uazl476NF1hh3DNseFFmOoDmWMavrnfempYtj9zXPN
vMkSVk/hEYMeBnqFpts2bzEXqU/FSXu6+oyXEInGmNmqTp5l5yrWf9c2VJhLpoZa
cdeXfRhULikdrrX5d9EzKSUdCw2CrndmVHynorxOREOEwPb9KvwsX4/w81/B/vw0
1JYzJ++viS6BXK8cNLj3ha/EvDSR9F6+OmDI75oCHXXkeIakKNxeN0bpiOSLU+mo
NKhUlJbmYUcBqPOeL7gKOk3RdQbuh1rVNJjC/vzNHxhklivjGGo1FRzUSoII7pEK
L8E19YH/fud4H+eOaIAkg1+pU1AeQXQCtfk0LhyNJAyEIw7AisrsG5Q6FpQd5Dn1
J3PtXuNW0cKkZM2JzKF3BVEhHLC9hfQ1GGGCuy0lStCl9tsnwAHREEq54Suy1VoS
Sx3iGJkRaeBhHk+HJ12Tw9Fdv/2L4so/C5GT5aY4c4cLo7y7PhTXEAAZ+nIqD72/
1x3G7pU+madG9zd2Yt0/xyNOwJv1917mT4cu1Wd3ch4Ll4cWVD9tnuiOYp3fP1JQ
kmN7ieCsnpViBSOLMk2rlaFrFuUAl68QOgeHrBu9THWLCXiPl8GotVHdle4nXt1Y
wAWrdaKuKq4kXxeHwzzlKycqHZMyGUXdBERtAhUcP0fqyb0puQBndcw1OS+f4ks8
/nexrcDyzlVaF6BtjSTplB5I4PNNqXB3pTaFhqHG+ZCa/AVY4R1GP+UtVg3yYe4M
YkpOAf97kJdjrJfZzzBVwAWswL1+aHMB6IY6dGwfvFUSZmp5cnzOwmdT+Dvgfhux
4iH3Wmff+FMyE30mFl+It2+7MrfSIkwoZnsEDY9QQ8sDkyV1OJoT8TFcbVRU6jF0
q7be4KbUm1meOx1jyfJibZ3uKQqiaNZr3azx7EQ+ntYKnjHiM+LPIXLHile7/T8H
3nRyr71MejZeYbL6vzG4HG0Ly81PtM02bWW80mXBYir4IT9JpOjLZgElFvxeKwIy
liQ2R2vQQJvTGJpgC+PtWLqwUEIL8cqjjasLCtOs4aJdOD+pt+NhYHw+eoiHdpuS
cfX6XAgNwOVuPRjpIkpNJ8RnoqeOuclKJ0ijfawVo2FwNJHKTf75DPMjD8Z3GDOG
HKMEwznSYnEKEP4FZW3jT4tlFjKNXBUtTDDq/zeJcer3S59LEdmuxRzz5kl8imPx
WZgL98xdieMZGTxwmMoiXJc8qoBkXF4Dmfa4JkEEzCBLZTjiKksDTrjMfISV9KU7
g1v3RD7U71+bdLdwADCq33JjYp8Hz4llFsDseWKKs4l9xkSc8nGJim2LaCLHf1jb
QDowzz//g6YZHF84RgMP3KWFxoWMJ/xVH3YYXS43Yu1vr+EpU1Sf5DABn1+ZIg5Q
spAltSNVJ1ms89vowyby8FMDTPwaJXNNmBzDcFgHzWg7SIc9DXLMDDBxxUUicSvQ
kycAIfDVEbIWHKm0NKrP8SCqDMPFDDsEAkX5U5QxmB1zkII29/9vQLdGVSvuoqn+
2sElo86CN02UYvbck9Mz8pwOwcSmoVBCtVNjR8W3l9KBrp8rIvJ4hS3z9LhVBS77
VTY+0HSRlqnOrBuCztax54NFikF/T8YhdyBEnrFpB1G7e6RY+K8ZraX/OatMwyRM
IHCz3ybYalznj4d15kEUOpmuTN3Dfzlm6NBPgQyXuf19AOhhEzurYOVuHefky2ex
PlFa6oc5SmPqeTmoj1fYMlesO9gseAmwmoLxVH6ungQ1PvlFblnvunbCefHOpN1n
h93Q4S2TEYvLC7pK6wdh99svS5vhiV2PlDkyKIvLNj2naLeCg1lM0iB3blnG+gmj
mkrIlHYzWoj/S00tuH6+RkRsemqQw/WfDRDWmkyzHkzX5/JcmxrQ4FfKm7Vn1vES
TpA1eenLFk7mLVXZbayaO3DkjPbbWSjp86VJz+q7iBhym32rWAVCPALZ1CuOFFVh
/72DVYu17bAVe1JFvPVR4i1Qz5aWucNj3XAUMps2/XQwhgF+iBKQLol9jb8shGZd
YdZlZClBVg2cA+HL1AuUgilxj/H83PGqEGbC5G4w++TCmq3LqKWNAltBEw8qY7oB
ALZLBRbcYjf3Car7888c3x/lmvvIgVKqggqXgBdijlBByFwm+s4rcW0vuncyyHTc
17Hvw1icjHirZVqBd/UoNSPZfuk7SZaM7ChXSPQyt9u791hcKmgT2XPCXqcWMsBm
zA1P9Z2kMxJZCAdBeqE8wuLgLHep4Zoh8yVzxXKtzBF2Vf6IiDmvG6ClEeoubhlY
hGEYVUybejal6/Qtl36yee0rUALkjb0YCi3xcRzFzzVIvDTYLGCNX6QdF8MCJ5dw
MUPP9krr1WA8TZrPkVTWnPk7vuXn6MlFC63J1ZpFyifVpWIPXljBgknbaDdeAugY
VMZ2dJRids7H8fRhtrDN6C9yu79tt6TGgIDcQZjVAkazkTpW2GNwmjTDAdrPhUe4
DXYcF16ZxXbyqTU7POi3Q0N+A9Gh+G5+PWUhogrPJhznDDVAwuyK3kg0g79l6N0m
fs3zfPxH5bGUEhFabkehQ1tpdjS2TRKMbhbFHlKvE6+wPQEF+h1tsXysCCC09WH7
RsCermkUA4K/gFcjS4IamYY6aJcyB6DRsutT+N7XgI7FXQeJejD6TNCoYamKO06N
doN0QQgPwzyjo/Kh8cCox2HICop+6piXbv/d2HxEgVywA2xFSWVMnwY4fo8C6dXT
g509y9Yz7zMeO1nipsFwpevHvozmgASTfP/M9e8ha4Q7TIi7nP4+C62pP0xOxeww
IORGSyyXBo/Mk8+7pzVl56RvWIccU1KLIEePLqX/YEoEtTDaIGQcyGbJuJLE3uo/
0CxHvCgXt239m68oq5oA0oMHU+vs+73tIpaLm04UoXYSpUDj79OVRyRo42zuKr/C
5A3+duo3xe8Z4gUDUlCTudzYVIJxEVXVB/E6DQMQE7/2SdKa6bhm8NqLBxKZUBUy
LYRVjT4O6la/CW4cQrLM2/0KP4uTZKar3KeIaVUpo7Aj0bWK867gbCt6hUCfGbFU
KvzOsPEyUUUs9i7Ct6U84HOnogTItaUA4yt45M4LB7rKeK29+0fdZw7sSoicSCM+
p4tbNfi2nVecLagofsiAo8vqNTXIF6/iNTr+WNgBEveGqcNVljEA3a5Bre31odVd
OIrPSVPdgtyFrc1lDKp//jKj5c4UriWA656efayjrXAOvfxGZ384zSDifrSHE72d
SmscfpWbSSzZfga4z9zRMs5VuHMzf+a0S/PG6Tj1cAZJiEFVenNJ4rRhG/Q8YMT/
WeGS8uPbvcyWOCkFsMRo7wcbOgUSUhYBOuA3F4y+iKN4Qw4pnXon2nFYAe5DIMKR
ZSTD3iYc+tRsFi1WwFrNqqXHpNvdYvhpsvZM4A4+lmaNooNj/bgVOJxGu23Pclfk
cuDLT9FhYwrVRy9vloRECPzUIsk7JXXcn/dUVJVrtDRm4iMb2jYh8ye4zsRjXxTx
i2jQRtA7O4hDGSXTWY7ddBuK1q7V8ByR6Ixg4ogSVb/muSOvn1UiJlaO6arWRmM3
nm/oquqJL+GCsWtYHmZoErjVuH52B5KTUIXUCLA0tlLwvLmixOYe0AO8wuTEaTaX
oZqDO61hkF2UsIs9jv8u/wGxOnVacMrhzzGovsigQ9PLHqTZ91j0Pi5kFGDAvazC
YP2mn4NMh/Z8pk4TjtTsvrKu98A+tKFwPhC4iH0E76QtSG9F1W3tQYgLeOJJDLVN
eJHLe9qFPIjeEDlRH8rFirrmYTp1aXces4Jp36cZee77gd/zGCHGJiXixef5PDVw
HHX4UB3vHhlBk3dVLHwdhan57bjarUy7jXedV1p3E2KJ/48xiyriZkUIa3RNN6Wv
b5Yvmz2sQMvuM48EruY22HuR/GYZe3klug3Ah5GJLZorJ0e5oP8KMjk3knvsqStu
b+CaKjL6gJe71vV2yjNBRsChEI1FtTCEGtKyoPCWAaOLhzIa/F/2Ji7Qn0fS91SO
fISrT0iUfc1ujtVBTIziudr/5MRG7TNUJk1TlIkmzMUIKV+noGm2SRVr7q493KjY
Jyk0iRfuNTPqR+A6CAaWuQ2tLLcNpcX48aZT7vd6k7ut8l/6tyC7R9tRJnNbHEeq
HdjRZ6EIAFFSMOQzeRHLg3dNsfknVYc/fjaSn2UIFAtViphKp4FSS4323Bkz96DJ
tpAQGaGV/GgbuI8Li6B6gdvbnBeNbE8gAXBjeFmuXUtLUYKdNzo7MzxoA/cDGGKU
O8kR/Ku6JQyTI0gqVC7SEngb8cTv+cjm3Ot09TK8IGakYY5nBDz+d2Md0nf3/tZD
2N32l+WkR4qWz+9Z2apliQc3sziL0tgoyeCL59fg6ZJAos6WW6pX7DJ5E1a37wkl
xv2JMd4tT1B1R2l2GA2z5zKozatlttKp9trByguZveMonih/f7l5Z+yz1PKEufmD
EIOx0B8s6g4AFiX3T47TT09GmWVcm8+a11R94sd0d+w0ANvIDZ6LDYSmtLcnX0vq
ju3SGTUW4jF94Fi9FC3f1g4fpjE4ZqngNecXIXDigJZzo1xfnbhjmBcNRKa3sWrt
+2Tl8v7NqttFBB2DsQtsSHSRDbOg03kU5dtEtgh0hKAs6PiKQT9+AIzI/Yvbd2qn
VfDTPv2HhiQENOsctNyq5FeGyxR4uK9Inj0weYza63EXhKdhH8/aBJY0/A5BSghg
2uZVcPl+gj9mIwBVmgIOMmf+UG5JwxmmEaqjB9Da+x6ULAI5p1sF8EHA4M97nuY+
n6uP6N0YrKusfr+LhjCRYxb77X/zEUGt8BoTpVq7Skj6jNa0h1VtKhwI96LOEAJd
Eacr4eQinJMw07H7RgY+nRrrGJXfmmk8ykXMW46aC77RAkPTBmmJXCVcJJ60pGrp
AfHosx93RvkA2xxRF9/TlIXUbv46ZH6e2w7Z/jR4afS6Ns45DTolrHR4eLeZb9hE
iIUUmrN/fdTFNZdk6CbwtdE+V9/ql9xx/0BjWzRkGvfGmoDWFPh9EC22F5DzHuBc
bEUOj/II5vsTh8wR3waAsvI7SOJ9J8SKcNoh+WEHEEcLXGIRgp9Vf6aNwVAlO2Cs
uqVsy71TsmNnFTVMlNX7TWVsLlNFhZ5APdVw9yxHyyIqXjeQ65Z3ULi6BGrLvyfW
JkGhpHzEB9yAs+vucT44QlK0qZpLur//EZwB3ju+oss36MsZ2cZw4Q9XJBkSI++b
fhJpGb5ZqWVjOkDxpc0whi1ivLaPNtLeDJ3onhwA2SmkQeApLD8HSOdmiYaslu9f
bMuLtgXFIzEzMqBlq+JGk4yrXcizQt2dXQQusadq2lrUPNEbIrFJIbnBlMWbh8FG
qJWONEUqo/XwYbhi64qM+M3Mwn3cflm4VdIcbGyQOyXSrFowhduANVPnjG1fe4MV
RzwPoG9XpAszNP8vDPzBpBRzNdTt1oMAP3y9d7qBm7r9R3I0sxj92N7AKZOv6pmw
MzOZMZ6VkGf5Tu7Prsa89qUcxugzNE28fuN48v7J6CWNS38ZvGnXldDX20RjBBKr
N93EnEWvfF79K72X1NQRZCOmjH8GKHTnLw+0uAGlqzAHargtnqcUbst8zzyLGGO5
6PxnUtOvqVgcK1utArBYY3ZZsccKamAmw4mrpEVS08INSz21S4Vx9/SDaQt01hjh
7SzBzvkF/7gvptLgTiNOvXlrRhSXWcyZohA5e2xykTXDg6NZGwEnjlk/AQBYI4en
Nw6nBPlmdKtM9nPAioPvkwBmRcWgBEJuSTvxVW6bGr2MxdrHduMzs0ZqUjMmqrT8
hPcdCaEqQxTGWEijplNnrKJmjQWP3FiMjT2vTVH0EspOS9lzsvPjFvEIW3hvOUFa
12l4MOmYFJ2TnKWfOpsuTU+ZHcpDu1EOfmsLu8xS32MHPdwZguO+vEGfve+9GMzW
fRhQkjvIGIRPPiJ0PhjMVq7mai+6KJlTiEEDmumq7zoYJ0cq92ZqKrpj1y6S1nC5
wRD4adKZ2Vefjk08Q6tu5PDzcyDqxX1Q3SKJwLYWoCbu9VoRy5eiHVOsHpjqc3uz
qauYG8iJmEQ2AKZRrCyeQBgKDW/cO53J/jGvuJoels1JM773a7mRUJ01kJjpnTiQ
Op+bfRf8VwXxmfrcEegOmkg+DPjxyge6d90Oyu+sL+7t+2kPz6/CID0WRrkMdLbW
bAgblmlFc3Ig2OknmV+40/N5PXevAtME3XWLp6vqn6U+NmIcqLc+Jlb7kpU5sZ/t
F4GcjR/nG29WTffDwxw5xOszaCluMLNIOCabJx9ypZ2GYf/kBrADEIiijfGfpMO3
q6y7gOeBkgbMOp+QVW3NS5ooPWDZk/FHjadezdlh1pAfpBKMcq3PZ6y/orZcGxzH
zeFtxiN94CIT5W6jMoOrdojRYl0cBwW6SNp2cpjxDivewgCYJZPHzZzQH7WHDZTz
QxENlwLY/mY6b9xsctIxWrYEdTdmb/0bxPBxxu+pZEwtPktfyFMfB3cuMLh7tk3+
IM5pblIAnjiW/wImVxOIApE7pfpDgTw1S2FIhw5MMNx6dEeneLr9h8b8T4r7t58I
8ZSLHf3VZ2KF96f0goRdxaT5+RTN2FhGk+KPLg+9fbvWjukk4EwnbGbD3V5QjP+6
ZhXeTuVPjAji9JebcTJOaM7LD1RVpPyyUMa1XfYEupA4aYUQFpTVUzDpzXZUQvOo
dvZ3IoNvts/Nm0KTCQNZL7ZinfXqBVAjWm3jr3PMYFpgVADvDKTJb0BEAl9h68r3
TmeoW98KRp1oCGU7winJNT7qXgLjxII96fkoMRMIbMPcCtZmidI8TmxiZGOwxioA
1dya2EmvVos7uxgZty9JG3LXysDZIS9/EuHNL9fvp63q4FmMIqWpPjRj2R1Ma4i6
1TBV0mVmh9JYRR9F7OXiCJJUJS9EqR1C97HGkYwpDlSQKU5Whe2pCGJCRTRgUTbN
vxUCpyBZ0DanfozHvcIMLljHTxsrqmiH3Uhz3C203glsyIZliXPpQaaOWr5rbp9k
SoG+SYsz3vGDjzJs132Mx1eKOoOSvT2ma3PVtSf2mfxY2hqCdKz6XgEJT11Gugzv
12yWkQHlu3Ga1+CgsP13lCmoPWWWjaRO4zB/RCDMSON2WLsyYGZYmfwdWQ6ZqO52
h3ZXFnfuOdct+NzDosnhgKY3DxuXIU4XzirjoYwPvZFO9Y0m+d+2mMhu0YrevTnK
D0m/cXm4tqElkSbbdMKO5qKQJGijK3MwOwGpKXd1yDwGigPRWIl8IzGVwW3XhubW
NbOc4S+ZNjjkOPNsnRMa2Li14GEJYnqvWcYbCXhEiwiTfiq8zVdMya5XxAa5z8x+
4tsa14J6Z7kR3SwiziZNXdxeA0/lvjyRO+WoL+ic16Etnh6aCiAxHpt9bjWb06RD
8UyACqNPBED5dZ5E0Vcglug/uXhgShOCEG/q9/l48dns9Cg9U6fpXGXGKORRjuXC
LwqAGEHhVB8ora/rByp33jc2N7gsPilO54hXK2ltb+FzYdOgzJ2nAtPsi+t+0vuW
QolpM53gDxwDI3/GGa5mTacPqtJTWKxjXGJy5Q9iKNEbVhAaG3VnYB7LhmS8w9ba
+1tCfOetUtdqq3lm943TiKrYBGeHyHYVV4ihgdrrY7EKr8ypa+5nTEzknw8f/BHd
yk1VSDUy4XMUUA0i+HCOfSUIuw2LaZapkrTv6AYIzZ+12YJpBEr9Sv/lpFYniBM7
lW5ybkVHlzYEblhJBM0aJPIEjASN+iXKdvcrbNyERYjBP5VSSGNZJU0AeqiSauXc
DVauxijyNPIhN9f0FnAmNaATQH280VtzKsYg6jPr9qfXaj9pYN2Tp4QJIrYBuR0G
F3Hwv9J7SNQg8gfGSF1H6yT2PEocEQMwNke0Fed7mX2XGfhfP+s+F7z9Ope3PtZ9
F5Nu0O+1t/vrbywEldjBFeLA6npACuYM0ZVA48IKVYU7iAsye2AZJR+9WRvVKLwN
S7SPudo9iS6YEnQRinkDBMGDA9+SfCEi7EtAea94O6f8wKDCsRQkIIsJefKupvup
1cayWiQp0T5mN6qvwiu3mrRKVh2ThXreYkuGlYn3Rvnxe+wHtd6Id0Jfst0xye+D
um18SBXkKFsdD5e4aDtGVPDLWpwRWHQPbElpG3Cm3MxcuNUo+6W3DRF5YgVHiCuU
kML5BHSoyB1haKKi9abhMuS30vGHln9+JHl73nfjELEqXLngGhmC+FFpIP8Rrtft
sgG3aGCxyfaItVaIypMgUZTkjKaRxmsIIba/Serk9aljCOA7EO0fnNz5BQyxX4Lb
OLa401wwI+sNdkjGHNKnK57mFVMUHtqN2HACQJBf24pwp2xP8i9euVX1GSw1KN0+
5ooZattIv3LQCLcJjMU1AGhvdRe/GgRoE/65FE4eoL1OrbRzdgLcXysi/bCkEk7u
xjBwBb55B6z1TDPq6AKmgg3w9CIuG0mQccADTdwM+pj/ie5tEU9QUzpZWYQR1ORV
Glzw6RoRBxadewFVEc68x50onKlxx6KkkG1K23LyuhaBTwDGIIRtTBKjpnTP6X1n
/7DBCrtLbs4dW+qRcYBX92VfifTTmfc4ke7s8KQ5zuEXS0dy4CkxZlizqa62rKrX
ds/yH2rQD1+8vmvw0J9oRnzZoIGEvaxqFNr133tlwPEZiB2GuNmxrX4D0xTzbn+G
Bl310pnW5t9XZ55FJxMJyixpYhEev4nQ3dKbr1dApEOF58mVn/3mSu1VexbN6MuY
fRUeFk3bqZMwAELAZD24lwlQ3BobULz7tNqJjFtafUn7QUmY0u74s4oE/KXQkn3x
l6HFkcbVxY4Pn8qt8TmoKc/x5QLMhSr6KiWRSfWJ98k6LHbvWnlg2XGJMBhpBWPc
7j2fDwTc8lyynORWvl6bkxblOvtq4jOfJx02DAK17tOK83+jrKUd9kC2blUP4Ee1
4rLdErOLn627QyvVz9kq8k8tc58TqA0VZuhgc5KW4ujuFTSZRhAKX1AOFT/ARtQD
hgZ2PEDHyndGlTv3WIcEc4Qvyxw1+KgjOKD8p8If/u7R9Bk6D/cgkg26tSiM7Dc9
IQ/OLWeMAXVD6CxE1OSiLBQc7pjwd0lSXnH/VKtsFWde8kGLWmmZelLThuu4hSqd
N9MZqkgzuQCGNbFsBtQvvmBZ7EL/99EDiIk4gnY7C7VEEtzZMZoygAo68H4geqt7
sehXwnfWqQgFlHYw1WpIli2Wxnc4AtdyxlY5DWCBBESfK15Fv+94lvkMylS2NNFw
4qJHtMUlB46Lya2FVNWo8S4/Ua9TmivOm11EJ6YLqcbswY4XK8h9EO5MN3kkwOr4
X0rA0oUZoK0NN2UIy9RIm+noy2hbbqgvNwwhl3n4HekveIHkAlpso+CzY8QP/+hv
iBUiby1dyLoz1X9NVzSBnZdsUD7wy4HxwHrOSuoh6zPtoAP/6p8zKWMh064Wr/UU
FuRtt6Cfqcw6CZp0OjOseMa24pHCjZVg55knrYeMaEzHT7cvIuckFYjKxTZKcIZ4
QUjo+Y1V92Zr5PTDyE3wTyCHfrzrIIEK65fOKJxYQcV/F1DQAWATdJJrrfy7cjid
uqUIhWFN6LBjiKPXXSHMNcrPro5JY/UoYP16tTA5nRlup8AbqFXP+/m8REmW6gug
6npGA5XIZ3MyxmTxmPnEBVL9C4f7K6fbfhqwoOs/o1rf8R+HeMK41D4V7JUgzV/b
0wqKUOlCHgb7t/XoNFKiGcX6QSJ100K8pRWj+xfkjPOucJYXduihOJ7bdX2kMx6d
WhqdTU65CXK0BVZDVdxE8Ffv/38XumLb+jEB5I8xM63R1iXNfuPGm3hWZ9hhspv0
gM7UIVeV+xBVVNjr47QqEb0Lqcu38LNBiEDEZSmriGhpPL3tjZlXpx35PMTSFDXi
IYl5uPUe1RPZYhkzFeIMGlRybnuMk0vKj3IqTTGn4oERaWVurGVFy3SHZeJOm+6o
sh88cVTonmAL7a44fOW8IhvJY86hFvGsonJxPFdBQLtQKGQOj6aZN1QbOqkpoOy7
mvlIX4EtuYJYqRMm/xY4iHuWR1kfw5441vCupJshx/hf8XOggu8FP3rc99JdKtmZ
VZ82WPmqauN2lyXNMLGVKHsnFv3D9i0teJB5HtARz7JT1Ku4kxJC94QMvxSirV3i
ubVLhb8rjqR2Gt+pb+CIFD1Xu24THc8TSUNEBEeKi4LSSkkaDPE+GfuPSL29zhgR
fHXZnzmBlt+BTEC7+fh72t2VAuKOJ0XqQNSaJgsb+Ng21n+uHdz/Y+mTsHDJG/5L
DGqa/qkZ2D6T2lUD5GgLuvWEEvBGbA0hh5DV2TWxdCioGl03OX0boIHkQEpWNRSD
vRay8pKwM5ePMz2rLK6NbdS53gml69RJCSCdeELDc7ts2LPOC5gSbm2FmBcG1ZUS
EN0pR7sijQDGdGkuncmNacIF0Ex/6QZkRitmo8M4hSCtpxI2Vj5O1S32GC09i9ZN
QDiLfWW7rGt2ZMDD8F1+6jwj/OFcTqI187DCbLe0GoQxQq7b8nKDVhCCDFBVfAuz
HxOKUgcKSUdK3J4heeLPTdlSPPx5nbmnOfm+yUd/GiCNIFLLrhb/Hlc4sxI6iiju
K6qcU47KhrQOxzqPyxFjj2+WbECe69YRE2WDsXPYknCnvVxMxLn8ZuMoaf084sbW
awpiwru8ph5OitQ/Uv4Ph0Zg8zvJi30Sv7bdNo7xnXPJ9h/bqJkFpgo4mNxBHjVp
NQNOrTDo2HreeF6ZabC+SWsTN7xYAhU7Sa9sZEa/fWZSRFYvbfFW0vqTSLgoRzYC
mXHRtWTEJTTfZJz4qwrgqmTysK+8D0lB4dY2xD5kPrjnVuJZF2OQCSj6gTQTLd33
a6T9luqdA88AvTgist+VB46yIUMj/m548oXhWqe49tZDiWAKB9g3zU75yd8SdndJ
d7xhiQgj8ThaDX9NkajQ1oOZb/F5OzaZOknx7y0YHJ98NbK0rRKNuL6dKZMGD+8O
Yxc1tUORyHtjrOuzArEhuzKgj8zU+wmJxVCz5hsK0Jcduz1wTluXtQzxbANLoDo1
c5T3xY78Po+tKTwB9/hbTcSD3oV2MjRz86sjvkjJn27Ns/vaIhQSCxJL/bZUXrHe
rACUeZtY1lwieI4sJXH53CLBHk4uEip5no8aolfTKM0nEZQEaDzNTytlAoRNrOtf
WLqDv+tI3PbbgNYMzAp6cKcSw/C1KhwCwt6Ary+xprW4t9upd8tiZIRtG5vBzed/
WpRokIxdwya7otVc0eWNFEP71qV3QS7sqmDBb27JJpShrcbjwMk03y7bu8xunw/4
zKr8MNkUOeu33iayFZuwBrapZLHOfIjolLN/cHRABxPqJoLpGWTWO548gYnQHDiy
1wbN7p48wTLKpt0dnHL9po24LyAsfGA1+IMGngWDZT+xZ0XmH8A719qf2mBqKmZd
rRMj/fON8tWmQ/qtBzmfjl9kK6d59ZFec4hB/mrq/mHe8P+yrlbX2JquOZ0tWnAF
SxG/0IC9puxPK53HASVWSU2t9ddcfAwmBedGRj87zWuOpQmIdGzKgh1ev988TRqC
TxFE0tQYkuhvXHceJh1AOv++mhZqg/6s/NkqDtGedrDb1aK26Kob+h13UxEYHCVQ
oDuKUBFc74Xd3kF9DYOoo4AbLK/DuPytluWmHtnbqRH21FeZYILUAWcboFyPPcB1
3oNz4thVyWitgfpBJ3ZqI9Tecof992UkAQPkkbd8DWyCfQWE1iYYFOtky/l/6KI4
lJEmhGaWTMiYIHGkVyFtIdm6f8WO+0L2qAeR6g7+hp52nMoqw7LTHGRAqdV6h+uk
PEYa6u3plHD6n9+3zhYH8QgWGg89M3jcx17KN/sObaItqzzhJXQwxYi5CDiwwyT2
G5Hl2QO7cLbF+2Z92bx+er+4IVY8kW1OwwCIxrtTlbcOykaupyJw7kAv0Lgk3dGE
CWzIcWaLwLtkZ62hhouK3GrmUGczp4gHEZ2RC9gk0iLjFH3X/H7RXhsXosP+q6Ri
EJi+RylKWd3p3Qryp2XxFfWrr800VH9eu5YP3ftErYGk496WlKSb8yBgCqrpIxhj
F25FIG30Bipm/ohLFOmnowo+Ru3oRdQe/Yw1SEm2xJxXpnP+NLEPHc5Jl9scD8WD
gquQ8ktipIlVIETePxXnlrRdkQZu86YkoQ/sG403Met8T9kL+TN92EiHe8KkYFk9
WZuB34LLRjA9Bt7fmHR/g1G8HK0YVb7cdRVRy4Gu44QBXtdbBw1YiP51W4WK0seN
ciws6qsRgWJwlp5dZ97Fbhx4MUN00gxSMSxVVSMtwgcYhYCqzz80agA9OhUtAPp6
K1spwLMZEI38GLZJZAIiXy0r4DqHnxxLQI4nZ530ywSb46ijpARrY5W1fv8o4kU6
d83Yjcbq8dIF6+XkAT/Zk5T+eF9kLxoG4RfCqG694H9hWBESyw9ZnpX/HFIoN4U6
fxPksMfwiiDlySlXrSGSfjFhHlCt29WcJzt2NUEsXtJdkPsuN70+6KaR/YmO75Dn
Q+6p8I+NYNyb/VQWQwqoRLm0mvRBo793kJbhu5QFRT49zJh983BNElChI1I8xw2b
g/UD/mXgU+lHdckDZOjfUI5tM9L2KDVq725m8OSE4Sgq2ENee2yzC90FGnt0BAQ4
B0grpZ8/fH0BijSFViIW1XyW1W3NOfLEbLDdXAfUyxT60N618aWs5CsQMBpRtXX1
qdFxvMJfIbT0ik60ZE4G7DQoBO1L9dJABfD15Aj4gebZT4NKHL4KQ9HYkLAhvQuv
cw6o1nlG7JViHv4erBbILAribsYFNti8nwMzdBPp2XT8SgQaTuhHNocBfzW0fiJp
uAlh9VFXR+6dG327+g/q0bvniaPmTZAKNEwGVjcEUlckjdCY8oEb6+2zYWS/NiSk
ye9LP4LxNDBGgeCbYJBPakSgBee08n/QxgJULzmtcc9cNYajn8s+TRUIbYXyHOD1
vOzxQStBUcAxaxJ9o8HBDP2EjQ1lcOa+2jgu1AHxp3f9rQUhqZ2OtYSC7/uzbGCO
hbLLfgAzUSac0Ku9dVh8Fs+8yCTjXxsTT99k1+tGzLrJZQZXZO8lgu51wkf0CkX+
gA19a9NGtXPkyu68ENDGYxcU02r9hwaVUvA+iIP4wNIdqf4YdOGrwFzEFUNp6rOT
v+wgfIpXgPNqcrT2F2pZa96hZcjeR9AWoFM5604D69WUJwV/w2xttd1BoztQiFXJ
SgsWcxDtfpdegK/Z9HRVyKPORAnxYedofDo+Eyfah9u+7keGloD2um2xnZHlQOmD
+zF8zcQwPPP/l1c3u9qPaRXu1TdhvmLRsnFfleQniyuAX+JRFmOSlMVT9Z4DIDwV
7oxV87pRj7mrsQDbqNs5gOfSwhup7142nN3tOESU7eiNnOCx9FZBNBKBsvBv6rxI
NIZdb1mkeIh4QtyabT7gkdL5zBqTJkPbCtjR98RALtlVZFvZQldthMbn3I1UMLrI
J52xqqaO/tvtB4ig/I6mCtC+10ZG9gygqQ2+nXUxw1mqAcJj14YeMLk6Y/c3x2XI
JNk/GITCTuHpisNRLutomR9XlCCz1wMu3yaCCDVUq8tcrl+4tGn0617sUl76CdNQ
RIomMafgWJacfaTrBRUtSFIYYGLxmzinNnEkXPTMot6+n+vPp75BCtUS8VgLH7vk
jne6GTyQq3t9wmR6h4/HQvyq7EtAbVwQyasTOgGA+m32PrPky6/wAOstvwxlDU6L
h7hBYgAxBngmP5RCAWW59vLzY3zcrmSrzMb97VBCdbNxe6HQJN3HtvaBtboBtw43
giAfqc1+w5ecItulyz6Py8HS6qxtjI7s+LADf1wrJmr6HpJK9FB6W9LFc1ir9Iwj
AnccqNu8VBlvzNDd2pDxCyP4kT271ds6DBgQJTgF6A8c23WeCeEq/Py0ftQNhhrA
Q4UdJsY2Ex/eEeBwmnrw8mfGNOwpWeEQ6FEYVjDlmS5yLR7xbr1lsDBPBRMXV0RF
zdVHHMAEze/i9X+oFNPN2l6OjrihDazUzS9LSKYXsoZF65FKHlsuOSPu21O1kRyA
k+CYOFz+PhqqYCMpfVR4r95HV4KIkyKLh4T2PKIWPPLAG/c9h3GGfMEE3KLIRYb/
g6iDB5oJ2urmfTbLBf0EzzV0w3dr161hIEzBio/wUhcw1zBqMe4zafPjNBJ/E/wy
suK5Qv0la/qpAv6KFf5DPbkLKSdOW0gyARyRpaGyTKHsYifKQIX8/DxtRvgnC0pV
GxdSF5QZhZmGbNPHXIVebVIL3gs5DP6O34AurvucP5WYzTMvYcI12w2+Xjp2+1Bt
vXK6eN1yjoeqveCyKCrAzdQbfxp4ArUCJHy4MF1OBiL93atemO5QG+ZWh2Oyu10e
jZb+yVwR6k2R8vddAga9B9YvF8t2TxYzAWZJH+sLJEopdAes0sH1ZEA63dmYyd+u
5UeN4dZj6zMhtl/w7jolSEmZYVyIDjFCsXerijmNSwh/UspP3hjCuhG92/4ZhnCN
jpfJEIJaYksC7rgb4dBS0qZXOsTuPEfevhRARKrwAxJit+qFqsplsrPqPbF+vP18
pindclUKWsKATJceA/JyGf7vFLGzw4bO8+OBRTNXAWrrEipYR6GotpPsXRBwDp85
08M/6f8JWU+EZBRBhh8l38POtlO8b05PMtqj2AaKzJX26VTke3cW6C/5c/Z/7Pmm
C5ijjeOS/2yewd2UbQsJcj8eMortVyN+xYNVovKBezqz8J5EvlLTcOREL0hx7JSk
vXFEDRgURMPIUj8kVffcHTGx6fuKd4ywAoU7D9+srECfuszeL/BJKuyozxEtp8kP
+uvN9qLQq2MJhEsr61vpmptfp1RNowWotfXseNABxBqwl/ILsfOpBRvah0Es8iJD
3dORDo4PEFE9Zb9CAGh/JmhudmIFJ9MK/UmH3vjhEncZ6ndvax3BMhwrY5JUkk+g
IMX2C78mHmQNOy1vLZdLxTV3dQzC/hqE5eKv62MNRiCvs9tL+40pMs7Ux4mxmL3I
1mXQORcVDHIs78jB6ApYTVUBzoq28xPAlwOyJg7Rzv3UGQgXnRTd8L1DaQJuSNJ/
Ahd5Km+q4PUSdDrv4JOGxEYo+QE0jeEjETYAbV3KT2R0S+sMDoQeVSQ9zIB7oQWa
MV259/dsDFk570uC498VgoPGS4T3xlbpDrJ/dymOJNxEYFL8RHUan8irsZ9EMpCX
WsHf3xaVUndlidHtzqEfYW4qcX6uyGc4OUsn+AJ4oQrOUb/+Uren8xDH5br7VdCS
jMiIUg0AiVUgYCyC5KUjGWapJ0qBFxRd371j6kADncyAaDuDlqLLpdU70hUP+/YF
tRoXabgi4f3gmxryBSpYiqukOXOWSiIsRA4/heJ+U1gh+1OLGcBoXpUJiD2WIu2F
I5rMoCfUzD2D8H532zV2C9HqyYmw1leIMqGRtz1gT6U4BjWSN9E3/4LxgKb5Vaqr
WrzIrsCJIVQ+peYQpbejgnRXOcKZjpyuxrPfzc0OFA7RmjEdELPWeG6hp7z2OwvV
VGPDVANOuq0QHUu8i3sWsAg7dGxibyEs/Z5BT0rlID5PysNlxxUHyZPFBSie58/1
rWNpMAmgasGatks0TEEjkd3RJBzyB9tCuhHoapAaTp44go9icPaFd8Zy8ZjqV7Fo
Tje5W0OkZL1ci4nLNHwhhYOq08EeHkqNvGWuyuuCeWV4i1UrL1uJnASX3R/pv7WH
bWPan9CwRaec7ffAQW2RdMg0hJiE0E66br66RJv1K1a+/ALbhc2j/vpJ3kcgyLLX
KEXrqq7dPPxq9tpvSBHdoJ+ICVES52+V64BCuI+ZbaAJVnHDqf/Tscr0XsLkVJl+
sx9/cPXi73ZSueAx3kTf+VEwolgM9aqPQPDqv5BcsTMwkbKZc1xlVjIVkE19479r
AP0uc4zimK6+P+yQY9PpyS/1mFm3fkD/hgUtaoTmhl/4CCMe7Zmj6O8YID19YSzr
jzaDC5gp8zW089RJ5AGIO0itDMlr2qIby+gmCTGPoGdArA7zUyT/ICpFWZ2E8TVN
MCi0csiItY2G/e1ebbQhmQaGK6BClOqcOGImbtfttQLZTrIm9dkwAkECVokidGeJ
7CPlce+yet6DdPTSDdm0TlOgjuZRUO4PXpqu8WQCOoI1rA2rwm1uAKsADydaU6jH
fRV6+1ts1MYsrOEyFKNBb3nKr/bbhs2UH3vRA1aAd9xe3DdrVFb8b+8utmz5QVTN
bb08Y9pu+jKzeDUgVkOd0wJUpzm8enPD0ve7ybiGxsMfd51EuYcBTrQeEzFbEYgm
rQpDVJ+5dBwPbKGby3LBOC4g+TQA/zvDe4EmWnjQbRy0gN98KwD0PPs6pW0TDEd3
nVvpWYNKa15EBtNUC+yHcJvxw/xiOJAqOcCxjBjrpITpKm1pk53f4QP9zT7xZ2rD
83BbwfcsHEw2rzwcy9nnQQqRTlCZShedbbxs7lINg7jhCVK9gLkRDIZ2QwF7T24N
lLO8Q2iaBUME/U+xnMVHFp0G9fxn86huyEJIf5H6/oA3fmQsfVboY4bC7tSNhouc
BMBy7UfLIuzrwrAZCxm42BtJVJZJcGIWjpWjdwoMoonEYdc5hnVE/iP4nkd7FLrp
MHDa5k/aktukgyExlwlqYy2ylNlQUXJtoB/RZ0FtNia4UJCdU8xag5biin7vjOMS
gLWHV9q7tA0F2WFP55tyWkJIBPqvb0q4RaBXixX1hjHVLRdL4jzOhz3KwTvzGsCY
G+QDCoQ4uaKUJuZZntp7zqTJ/JAeH794YifEDymp8qiubv1GJRycD2QNOTfM6Ssa
HcaxQXPfrnDJGO5P4LTss9xUwIHXjQmj1gVB5Lma171YAAdTbGZx4V6d/knKMXpn
zjSs3wusZmo8vfjfb4qgt1pwASyJPjtI2MhugEGLsmeHyuGbaiGA9MBH7AAtUzUf
Dwt5LC2WEnyN5UviUBb3Fy88gKe8+aE5OJPQs1oJy6M9/G8n4GAzQoW38H/3a9yV
MNyYtRPT6nRuwXdhieXUHEcCIvTQ8fSVbqY/bJTH3vHwEYF8Yz9FdfTBF+Q0qGIv
4K4xdxuvnhJiQ0WBxaxDfrJkT/xejSAxxn6ZCBPRdvw13Zn0LJdJR8AkIdBOLzm7
Pp+yO0pOU4t+/NzhmDBSUiWkk6l80SQ5g+asKWZ7n51s/3hGd1ce9AkxeStGRkF2
67b5Ncmn9sIsFsjxm963Z7rLtfhfL1TQiPEU75/f/p3vPVD7V+CJMUdActJqoT5d
26VJ5jlOv5cx8Qo4N3POvlJVV6jTfA/+kvxL1GpfACIHEQhq+7MGjpz5c0oGJAI4
xIMXE7CozEsBtotg9/KeYlD4d9Nwcf3sYuZ5pbjK4G3WurtVR/NkVHGIZfTF+6og
hcU2EXl6eJt8eenug7fwTmci3XkYBC03bpT+SkrhA84z/VGui57VF+dd91X3HwEQ
aAxlPp1uQ75EV2VgLHmeO1z1csAJET2l2X6J0fJtDKyhK5pvQAn301lUEpIGTn5e
myfb2k0YYGPIyqebxHog1gF8duvJv3UH2utI8F3k3nX6Sguq1s4MMwuxuzOWO6dW
JoF1vEzExPVkz/R+vbPbXGrsc5EiDxQrka8l43pAMc0cDSeTR+mGOTg6l8+seCQG
1nGITLX+Boq5cjqFIxt33lV3ViSuW6NVMCcNiA/GF7tAKG2d2vMKF24e1+ssKLN7
BumXZsvJxzqVKXrskpfNPXW2ZiEDAqdfKaWJV+vvS+soiVh1dVrc3OqaRQn629mn
YVkwCZvT+Cj0Joe9qypeTCpMcoJcjfe4v+PaC3AgQzQEF9CLtZWv93P3yC0WXgYv
ECFaMWfPJRebKehiOSbZjSey3ZDaH7TPHNR6KBBl5+rfcY/6Ugr+srk4bSK4K5Co
KfjOBnT6UAoLF6xLnEy4oBi1HwbCcGbjKkvd/NAsfMb6Iy+c8a2fAU03HzLTcspQ
ElTdheJVNlwK+2xo4C1P53ig8V4uK2z35q82rmTT3HeaWNBdHu3AtN/c6T7xBD0N
xL3zctTCEtfLIgGrGa+EFRCmwAuQC93/SgKQtpWbYsNFyBO3ecKdOsuG6JBmQ4i/
KeyCQu2C5mp3dnp+LoTGnCg6rE5AzGyjMAQ8SneWpCjecVpMFyFZqXbwURRe6YYX
HZrdK26qVbZrZMoLtKM86k5465KTPc3HGF9Cno2PFLXckEyydJP7lA6xhJIYKHQo
FKMP6TUMwW0y3Ve+lS3Op6DkVZYQrpLkUqjsi4X/oK+ntSZa+JsdU55tdkX3IAjS
7VCPAdn09oYbi0W6fWdn0k+F+xHvrarTT9fKiFtJFIXbZo9WIxonfiudNNJgegd0
HHioO7RhtVdI2KnNHky0Hq4rCwyL85vn7XCHoI0vilRbIMmuUkmYhUNGHq8yQqGr
FKHwjkibWPg9M18OP/x4jI7kKbSvNCeAssJ4q8N0qlJLRh0DFPtuIe6qG5xH987x
h/KD8lpJhbuq5ZcAxjr6SS0u7o6NltvkcJClv9YU/4y8U+d/6eJE0JEkVusA3yve
fZgtGhLlV8Z/c0eg0+Z8CNAFSdueng9QPTIjfUXujJI70T37ackpaEgyzAo06YCF
t5ialr6P75l7YO6auMm9IggfvaNR5PXSWZKglCf2FmweXyG//pZ49R9F+2i7xPSQ
TgXoGQddiLIOKcgP61/kpteqLemiBodXkvwEXjhu149Ceys0YWMR/CL7mHUwJbK3
IEdq6KGrHKxH7jYHdgC00Ekl0uLc8Tj5s0qFJMV9TmpcHuj/lHVmf6p1lpqFnxoW
BBQt84r1rM42GTl95A1dQs37GKKy5nSKu23AW/xEJR3nr4W/N4h1egY6VY94xvm6
VzInPFksI/0hudQV+ZPUpTV7Bjpd/U6uQqcB9H0mM1IyHmpNG08DRCkmF81UEXia
SogDac29dlJI7AKm9jtYegdzxOJmmb5Z+BBobo6D/ek80XR9ObqXWsBopaG16+Vw
iL8gXEWBMOI03Uqm6ObRlvF83UA34RVXSU3JusT8rCWEinYobUEN7zB7ChgVFww+
qXV7f1LU8zCl0hLj5fV4opdd1JVky1zO2ks4dFw/sMxWIH00MhzVbwP+7EaIEFLf
D19YSRn6Y+gRXnSBLsSZpC4MXYzXP0biFCjlf0bgqQzA/8sdEoiIE/LSCcz1mTya
t3qqREiOQMAtQ5A0w4uPmvZ6sXh1jhdnfONUFGrm1bpkmbqP9mA4scdB3+4XkJlT
alMbAdRv3kONG8ugWsCz6V88pQzeWfVqNo2aeKcyMO9r2X/j+1GIQUSK1p9oEM0t
O6Ebifk8738FabqsQEU9loMaSsH7yEh09DfI0zTBevkz9wYT9shgzj+y1y6nFR9F
n/sSUIMkJgsMU97+r8olgna+8/2V4JCIXv9Whl+YbPAdPbC3kEveIy1SHJtlfzm8
X3eujfANQ0C1lpk2ui/LCGAzspZ9YJImT3vX9KzL5ykmPNCnqynX19H7CIkgK9xp
wvvptE///IKxTQydTtMECJq+5/7H8pVHrslLWL5qko9AGflG2kCcMbzlBpE3h12D
zv3Z7OyBcZeahmwn5IoyM0nEQ9g84D8l2XffyDwCL6yMlUJNlFR7qUcPoXSpRoRl
RjxsDCcnfWTPFZW/G2FnkebplqKaDJo7zmjH6CZRq1wVsBOJGx4TAtbFUtNhR9d6
GB0dXoiB2DJ2oY0jmSwXGfPmyZvPXq7ZT7bMO2OCMWvCV2gjmyh8VAZfqtpRG2ND
gg1BZMU2ENf/8Mxdr1ABN7WlZer8IDIzVXfsaCKG5F4Nlmji0FsgGmpClmqkwoJX
TBUiqJbNjDMrCJEC1p8qixPk19LdpCPQmZ18gtrkWMAHiTG+R7V50aRwn+tdZEnO
QVRPw5zmtsJzIhHmFH/8jf2nZrynelQwVC+31uIwpwiU4GkJp5VwswSsqjIWhgTg
AehYcVo4PkIWLnYf3jmj35+jUEPm2rv3CQGRZYlZ1ca5DM/rNB6KyMDojL3YOkzf
0rx85eZ0Hlt4vsNxLKU3PmRgGzginRR3yhirvj7bSkG2NpuiC0Tjm0os79iOSOeC
UCKeqFpK/95K7qRqV17sC/RSBYO2crncAPo7z2+T/2j58Hm4WxOHP8AHS3i7pwtG
X7Oq2Q916lHadtCTY508AoKetgtctZRCHa3KiH/MWaezd5zJvHmFMVAlpllV2Yqm
j3hFu+4A7HO8U3ee2lU7dXv36nGixKcCyJgMTgx0vkSc8Dzkp7x9aztzZHjqRNqt
zQdKYyUQwxor/Q+uu+dS9waNAXx/rBegyeCXOZz6xYsTeM3NqbvQmaaBqwVIsFL5
jg5fh04aUcHF//gt5bmPtVKcaZRvcDwpj3y+ew8TOBs8eZIirKvuMFCRtB9+HgwI
3DA9XfYJUtpBt8mfcnMUA9MLz2AaJ2TtnWFjjKE0aiV1PSHsvmNarlVqaYTozea+
ZLDO+PnKl5SFrzJd7wlb683R7FwGMwgHhnw9Lo0syu0nfLyt9TMuqzEuZm6x8w/8
1JO+0Fd7dxmgZIfhxX+WdihGUTLKCdOT1ABRWWlWoiPr/jGhmAnkVymMLpWKxZcY
s5DqnAOnLD8MNVTZjPSFBiNmubPbqvmJkRYAB6n7k4yGUptRuc6xOnw4ExN62fPn
eAPLHJRpCnC3KuP0ZjLvLfIoaUJXy0Qwt5dIIyfIdTVswWlKeRtAZtDFwTtclYT1
qwHjMt/QjCV3ZS7Ng2hw6oY5ObW7PaxBxl3NkisJ9/1YMDM9FenGbyAsGBlyzeIk
UYdMLE6ijrXgCMn2p5LCUBJsmUYVQ3yETU4YfDflH8B6ATI/pJR4XFgqO0PARKD7
mHLSfRqORX5s+/1WE+p9SAA8gdl/mDWax0YHy3dHXW8F5aJse7TYITAPj9henkqF
/HCPvNZiquoFYBK3fxyBIOJDFjRQVmqbrP9vOZNB2Z5Za+nfleUELfPtcM9jaT8y
rdFVnw+HQ29nTmkTJUx268eDV9SbeRYcn4QDlsycq4LfEMdbIrPUa29OqYiu9oCk
kIVrv1sMEX7eutgZjFJYiUpVjgui6KkLRVUKgRIPNEsF3wD5J5LF0FCsiVEEyjgc
7t5MQzKnRGZ3/yOa949KQyRRkn7dqTogjfKmp3tI3YF6Re4Z1bLKt38xDnG8kgqo
39GIsprs+8kY/FkxnJoPMYuqG8HJVp3w1hQdDpTNFgjw361GDZy/gmBCu/a8svyX
skE6EFl4kpvAuIgKdSZq05oDd45QTys0XPpoNDPPD0JwJpOEBctUPmaMLgUuf+FL
2M8kW5ZmePk49FlvTLxRCHg9vqb1gwmJ+HBqa1PWLfQVj+JbSUXAnBck5Q/cXdMO
yUu3bQpszKAh8vygEbPolFUfgTHivf58YNuuG/3OlolZ6yhho5vMP9+nAHazJ33K
zkVZanIkAzsP9fS8Z2BUtyKlaCfhX5wEbhDSPZCtZrVOvigcwsK6iTKKHiLCNwtj
z+2sSmTdfdWaQpzUeawQfzloiYqoTW6/8VOK2vfX8Y5QwNez7sxgzMNMFlk7lB5s
xNTwO4ZePArXIacuKqmsGS9dkyl5Kt+v6rvLwlDIs3b2ByinIZ+pZPm+27tLXURY
tSte+v0vlEJlW6X1o5mPrYvP6AovdGs0RBrsCHj+adK1+Jd/2zCob+fMp9hmVeJ+
T7zYPVKiyalbqsQcNuHFUBsSUwtYWJRbiwsJc5kojbaDKw7FkDJMI3R5dhbMeC9P
Gc6+HX684ruzed+1De09nKXoR/6TOSPAEYmUrEdO8XfCvCnDcnyi6aDrGkgw6t7m
K7XOBnjOm6Ep/Ky7JLfEgDdpuoU1IuwCeXsT1OXx+0c/FN+790247LjIT6Itvyzo
kvzsi5qJCwMBF4Ohw3gHcvDfPg10DkE0yDzQxXq67qElh2CY0W7M6HXn0R0AczXT
KOpxl2NFul1ZVSQAJTwOInCIeGj8BPtS+IE025C95jW0hMceV3B7tqDibrg2EbGS
OkcU05LjkYBwZEsItVI8aucda1/Xu4NL/DbHYUrNFszVwvETs1rm0apBOvxovudh
91s+qURNnJLQANVwniBnt2UW1rHyS+uDoHhXNpDNahP53BjujRA+SqHAV+TBqUAd
RTaF3q5Bnb0PLgUe1APVJHmlWAgxmi3zgCtWAJgPFC0YaiRC43UvKnFF3IneLEkS
30UJ169Bs2YnsaPcK5qLirYtbdKDh2Ii/QHir3sY0QKYXbsrTOm1QZ/Hfgo1BRJo
R5ecPROlQmm+J9gFkBKcJLVMFQbPlW8XHaJZx9pRQwyI/fU03RrHqF7H5Ec/0ElQ
KleqvDNwMKUjMnD8FRXcJgWXiRC7+q2Tz5G+RM8IXlIp+M488lcWEdfFyhrwIgxX
B65Tb756+IA94I5xVqjSXz8+wyTXHHkE2Nkp/jkvZkSQwJOaGmXULzJwGfMgI3xw
V2uGQeXcblPGnuzgDSSZUunjusnOLc6PNgYaemy7R0uXbkrFrl+Z5ETz8swM4wSF
2vX7aDwgtbz6uH0vpB6My5rvOL+OD4+2JszB1S/buenpAT+jeMdNWsjr0Poh+Vku
wPBW2QQXciLAmnupBNjTJgVk2ZvWDQuUYcBczb1nSf0UVJJ2izzoSiQW9oooMLwk
Y/iWCt0Ed7Dmmh1fvKChN6nfEReK0CRSwM1gXuRuWMSBEUb20pot5/a/+IdLRAIc
TCfys+QUibjn4a8TYDU+HN/F7WMAn64RhnmbR3GPBYyofZH8SM0wzJ5YVZps5S4s
pQlWiKzBG8d/AjnFZtqtSPRK9V7KGS6tdRaxPm49UGK9HsrJNkoSJ1uvUb85Q+om
ds2YSUAKl14P8aeK5LaxbBq4nQXMsGx8dEWQGHkxO4giUC/j4y0HNuoAd4eBRWjp
cHcmp0ZGjcMkdDNKxWzsSCN0uaiLFWa/XMc+F/Uy3j4mFA8IWveD+0lf5cuM/AHQ
XpBDgA0Rx8NORUe2UZOchI/n/ZSbyxKFgxjMkSJn3uC9py5eb/an8eqOjwkjdXom
Ieh8a/h9+MEhEA5830I0IO56AdbCeS67xkouW67utXobomeWfPKBOJRwB6083yfC
sTDwBNHPD6hsTrXKTXvQWpvsJVfPnGAfxdM/kkpJNZ4WOXEcddrC6InBcigk0uko
oRcU/kB3ho7ml1a6yN5OHBnNS3CVdRuFFTVR4Kd1SBxR924Mde4XARB/nnQO4EOF
E8fpGh5vUY2UvJuVd95IfKw6t3QFm44HQJCOGqQWUuhiF1zNnyh33+QDkjIRF7wC
ftMxHDQ9MLuPKoJnUy2i5hIWa5LGe+7RrNVpn7pGTGQ+/u9lICAAtrD2G2lHjhJN
98YcMP9adMkr1iiFPieTYU+ty+LQqwwDoxVJfVJeg+tbWPuW3izu9QXkEPOw855M
De6w5QBXa9cxGD7EgoxEBGTpmqu8enNQ/cNfjfFCPvMi0fY/0WyQUtMKX2TsS6FR
r/zbSFFpsUoTwcqh1LFEISbpntukT3Dn6THhRZ2Ix0AChoNGvEYHCHznR8rKHiyo
CeR4rUkr1E03ZvflxqKGYRryEx0ZZCbwNWnHgWpkrBpYUgMQ+/swHZkehEm/XzbP
VmG7SzuJDys0CXuJZ+pLb9vvFwI67D93v1T5mBzLFevsKVshWZxIcXKVBk53WdNR
fjikcG9uVbYQxNBtjAM4NMNmhsyNtXqgTGsm0DrosCyPuLOKvM78oZB9xwXQ1DXt
ERj02M8BMTzxvMxQ9sJn8eNyV7wZ54VsRQwvabZ2vIzehg2DVt6vcKJCtwxsNe8y
xjFVG+emDr+SvXGTJj0Olsb1SQckVs4r+C17ObcX6v1xqOk6QUv/9lcTYmq+Pf3v
8yyFHoULdJuTb7CmfPu/iiWKnmqR49vfZpp2FGROggq2xNr88grZFQSE/sLsqbWn
u5p799RVRyVtgMIWYI5xFQHh1k5Gw5+zEyCpNBjwiCm58NMHjhBCyG39NLKEo4Ur
V4afS7c/EQbbRI+qrGf5QyXWck31wbLqYCZwAV3ytKiiVeb0ZEYLPLU4uRpLARbf
ZQ4o6HokSfm9Aw5qr1bUceM3Vxqwh+zSJfIVxoTQ4xarztIHhaZPu/6Kgpiqp+v/
m708Ci9j8JyepywnHVgm/KONTPNX1CgrPaIwd3Bk3h9vQX5MtBHl4Jbwc9Gukjjf
rHETEomrAhydp4wKPEwEDdB+gXGfPdKncfEupp72F/B/HKws1Z8AtqEhlRUNhNtt
whdH+hOvEKzUaAXjYXTyl6S2lGQzuityijm08eM0tJKca1cWKyu/9PiVEEGAPGOQ
xUWXGSHbbFidY9FTkTvH4k212bclpMS9xUGN4HIvC1HIBjtWV5y9Y1FEgW1zmN03
SWVdKNGhvT3CdH9npnsbkz/tvG2As4qzFOdXKsb4xq8AJa5gugMT1cuGiwEKmZx+
/IH9UqMRekN47jHnv2qBqjnY7zbsjBeZSKGhklWXvqgZ85SMNBRXfPEiK4UX3qGq
pbDQZVuN9NVRFdzT3letrYekHfsbwqPcKWkLRp33q0DpIc8qicn5SKqMB8O0lEUl
dtRapwHmLRekLleisHNh+vqZbQA6kOy3NEPEslQGuIfr/Qkd8/sjk82S3g1r7Eoc
2jV6N3gDuE+opNtKMSKY5F9IZO5CMHJTZl1dafe4kWH4hqusBW4pvhR6qvBwSYUu
jruv9o+3IU6Jb1/Pbfjc1XBvBzQ10PXVklOPA2PkdNCeiq6Dc8J9Jok/KwuPPRme
0N/B0it828wAQ1w5LhJelyTvylJLPcpBXaFEi3zhbhXT0xZ2J3rEoVBHPKjf3rU6
HyZq8UUhGfvsAGQZv1bAwLfgg+NMpzN46GpWZgkpIw/4TgbApgzVGhIqA+VzhOSP
qVscEE6i1CZ+OLrLrf31qmWtQ8CvL1dzyDzTucXmVuKoIZHrWF2lzXosZR0QlOgB
OsD9rNM3v4Qt6YCuJz8yEvffMdrsztsrN9OD8cwfazJOb1kxpLjKZgQyti4a7f6z
EK0TF0ZdJGq3Ew0ZSOooUMTdfoFEoeASOKE8WhKzi1otr8zxzc1TVffIGVHRGWWr
4PyQvMjzbzS6uLQwq9LsiWpW9shrUELWa7M/FrXmjvoZS8J+ITzr3fnXcLCA0/KU
WSkIXrzNS/Rf3V+9dsyzK9tBnYx/6AcQfX/MS4C97fjVBoMt31jAslWRPwzlnlZr
ZSUAnPZ04sDFloAZBQcPZ4QLHP51UfatHLoQMZtHQnvn/QLzCZRxsigkO4RpyiJV
2BH9wrV7c32RlZb9OjlAjNNNOHM8PHiASr8pct/LDymLTS1jWN5zqhKyJcjSMhJb
dtFpSUTTE8wndmD6KFs8lCcZ+tMp3/QeZYQPZmDmzIxtBMwOFXyKDJwdMyw4seRQ
FWX5cxeV+slmPAPbV1MxxQhEEr3A7pHsAMV7IMmGOXckuaJvXQVqYbKN9tclQaCA
eKa3pAlOfIS7o56xVoAA7fXVni3vd6sdBA9Z2M70vmoXkGNlKHYvQVIiainL23RH
/a1I3qFSC3flZuYN3ylEzlLaWb/MznY+WxAlneSDSp/1pDVmhMbj/B/MT4hucId6
Z+JoyOHjrD9kcMRqW+yV9ydE5nlS5Ejf3HZH5/6bnFOmAnSgFUOuKj4Wn5gwf9Pd
2FYQhyJzbKp076P7dO6Qu/xoM3xoirq96UFjWAijQ53fCxCHup4ZkFMZhJ0BPsPz
DU/vuNXYwE3rF0bblhttksiL4NiDUQzE4qtFs1yj29YPkLaftgb1rcF38dGpH9yI
0vx+al0uijMrHl2RNhTPS6Hy9a1aRJUr609rxm2hMpgvAUT+6WxqifjyuZilluI2
4QT/v9sNS2pzRyfaWqkG5IluXqlkQugBUOpaTeXQA5ccHQAKpc8PJBcGeHOHaBq5
GEeIleMMYcDX3uLlT88OM2hPO16Fp+LeGGbpz87PE59yIm8g9FWwSkfMAHVuOOug
dVlQE2gqZ0JSd5s/iQeUI0c+CCHG3jRIfH3+ilrHbBe/LvO/4+felvLgouC/x63m
IlQgC/OyiK/TFhd7en0UEfkBUYA/mcVwAAcxCznAVxOyXwPHrN2Q9JRSH524c2KW
zHeeYy245nnx0+zQ+e2epSNmIv99SBbPxhbBVq3qUgjQ7Mx5pVS8/d3qMey2VHF/
KJ9T3lrumqPkc8HfAOOj7tM0fbMKPx9t8ldrFVm/Dt/i6QY1EcJ4GtMmpgxUOxav
LzfvWfaAHbBNQaZv8ef6vOuo3vbpFXATBYRhX3M1RRlu/lyLQcTdxcnDiwh65LJO
jYoe3sc7hrA6W7RJGFgcWnax/aS8YXe39z2DP3j+EFcQ9iVe0tVcvqPmwOGKVU8Q
ozIAL6sncVLd3RD16tPWGCt4PSEpWG8XxfW9JWpAKXUWY5kdATMbLY4W833BpvRY
AVp5Zd1c5tosp2s3RQPD4x/juP2CMG8UeAQLnG5JuoaPhVydHTh5oXx8HzmuBu+V
8QIUXrPkaIMEJ0tgG+G4W3hE7j4frjlAd3z87B0Vyegylu/w5vFLvA9839p0IEMG
WZ2Pa6VurHBde4t2aQmPVizgjihVvvcC43qdKib9PIE6o71D+Z8KynmEA60nC6nV
MzaCfUtr4YOi03dWrsVVfQtXNkh1x6h4IDLyUZaSVW2uGPrlTl5hhxnKtbfVdrwN
CvVxpdB6dp5OGcBf9LBqndH8c0caeX6um5Gk1XTz+Xjnsfb+vEAapCwRyEjkBGDM
IoQhkX5veOc9jxkgVEUbBETIjmBtnVFWL9Jrp/jOfqies2+KU8gXKUBYawpaseoZ
aYrIoQMJxOyjNRH+2g8EhtwU9VJ3V/5t1IV6lQPtw33nsewz5ocfr73aCtYp9reW
uv1hZnuGG7X9CqbimFrstmWTfv8uMxZGZbMAlyOyfdUuKpzOMaw4gRvCBPEiVUHx
9Dy3tQH2OUoij8po+MF+SqWD2W58qin0vONDpepwqdNUzP726X10SHdIzLOMvsUy
zG773o7EQxnBtlU/7xusmLD9NyHXcdY8bphWO8UT/lpsLHhWB4WRgSYQkK4nsXkk
xu0AUJr7yBjctGx1/6SA80fBHh2CrBRst/KvxfRzLiyWdzTdz+Uzsp67TqvlnuoR
c2hVkzmgmyR0o4jYWr6Du3r4fSwj/uL5b7El0HJ/WA5Fo5wPuAqA4ZW/UnsrDmBD
T8gqeL/cN3GFul0F228DZD+WO44JHbhrQNRrCF0fHvVg8Q5vJbwZTjYPJI6lV0ML
5hlJik55YwAJdX20z491P6PEkXfzcRwXaANd7zTpmUd0HudfPE6/pJV/4gaLnf4i
swRxqDaFQhWgBH6SlWCSCcvtqZpNFDSiuskfl841D3ty8v2hiu+0BnzqyYAV6lxE
IXLwKFIQlTSbRArEMvxqmQr0PtTa/ojsbL+xwfJ1IcJGCVwk8fK6NJjUy3Se5vRB
kniMZMN1A301O3a4/P0TsJu08Kmg9iKeb8CjiLG1N2UTbTRFEVFqhQH4E8DfOput
1Vd+arruZEPxgmxDPIAMJO1qvdxr3fOb3h2T2rUOFDq7HkIYYNYpIb0o/hdkhz76
FBXzclpgkRNyedjEBgPmoohcPIULj8VrdFtX3ArGLDYEQIriHa0qqCLCh4CxTVYX
nRkOhC1KJmK73oN+VbWdEdqRa7S9xuKki2/QySE4Z+VB82vg89kHHiYg4UCql/mR
QuZZd3Nf7hiyO3/fdKwHXU3G6uh+laNBzaAvijRTnYPIxyDQUCdrMSsq/WhxhVM2
0Q804RgWghXd+zzLUoCs6QXUXjsXcEtGFTdEv72qYKd0lerr1ULDQ1tkXoi/0Vh2
Oy+kF0CR+4csUun/JlZ2mRXNJMh0K/i0YHKtaRsC7TLy18M+T35UXWmx5ugy7dyw
BEFwAOaa7IiTwMiwSctgTVdTcnoPMyaDrF3u9XZbZ9q/Ttd3BOJEOOS57vmFs7pR
YtRTBCN+O07oxQBwkMr70X1MsfrrvVlmx7LsoFki7zhDPwPN/TzZ1uqrdOu6MpnJ
aIaO40eLNNvLbcejbb/zM4YYT8fMh3D08LgM1kgDszXd7S0MuGPnGkk67IdCFvHc
tRn8SMVRjYxUWdDTuCNxiK1GLH+GzSBL+Oiy1lRuHIZkpwb4k0G17lWv7yBUuLjo
Wd8XMEyDX35pso/at9lGn/5g0+5kiSpepTJc9zcUz0U1QjxEvODB9TpdVrj/WZWc
T0ZDpFh1La3iGEOAbC4kAMXI4Dh4Lc5kS3wquSxYckNM8wt7rk0UewS3CkvWAiEc
sXxLvu4fmYzf/IulFqpNvEBo52dDtSZYqZUEM/4S2FuBPryek4TfXSC2kJy2JxkJ
nHBSUH5E9UP+JrIGyOyw5J1DCATwB8XsKU9Yji5KQ6b09MgAaBOzfs8S7ye3PV1a
KeRJjdh7fywghhJPe1izvMs/sJpbyzfJQpSz25eQuQ/AzBg20BYmnOQ28zLv3z4z
eM9Uwwt9weEauvp67wDmk3c+LD5Wl0DuoiKe8ui7I9e9lwCayDdEuFNTp7vniy+y
59zE9vW3HUjua8JQjy5gG3PWYz5kGdRMUvtDeuiCzR6/uRzCDp15j/qmYWgeMgLW
y1si/tpzuHwGvdWDgOjHZp3TDhsJUBfL+iH754scQB4lULMvcHpGSiOrnWd5/4zF
mc65Xu1k/yFL7G1xl7q2gSc4Aw42YZsV4TbFtbK971Yj/A3yN71B2UQq0ANp7Lis
oad5f8CZuJ/YvRdV22DjnSfUaFGQIuahJdumom2Nz6Ps9fil8i1YNKRzS5LAK7lH
gaiiP51kIpJqP1nyKdn+WaiMewzeFUjhU54K6qAgkJGWNgSjp/SZiaWQYnEnUI7a
HVPb94KecsDsBSouyfYmwfGwtp2fdwKOSmrICIgkEClqTJ+3+PLNcX3n+x86/qVd
m5TaDTPx+CYK5ZThsrThaofilirXgeXehZMCuzKtZGWLU1EjcqAqKw0w8AurXHEw
jhHrZOShXsMToS9+VZc6ouHAlnRxc0rgNn3s9v4v4J6oL3/aG15AuoGl5JYq7z3u
BmcOkBZVyL3m8bvpI3rj06i6iOmvsd8v85+B49HNC7zUTJbmuVqPA1NlmMmv0q6B
kAnPIFL/QZ7LoRoDzkad6r0f2a159C+IBLCpxwsuBFQHigfVctLqZlhMEs4mzFLP
b7riJGYyPC4xN25ZZt+o7Ru3+xNfY3uSsD71OtGxctUPj5ZK/8uCBdt7L6VfWNKu
52GZmQEOnUXh7kRubrmZZ19dWHBUATSIoH3foCjF2iwq28+mB73QFoDO38F1yro+
AetN9DwczsGKYWAa1ud7uQ4By5j/L29U5XHmfnFWNPd2yy9h6iRUa9nhv1mXseJ3
VdVfzZnWr7zNF4e/DslLpB8v6cZjttsIXs9RyX7RcHjg6/bS+cIhq7LvHbIZacQP
hZ1Eiw5e2ENByMevVYtH+k4NivH256K7j1vtxln3c7QAcL6oxPJ1WyCmM632YUaA
Juqn/ap9VL10DVAdcV1F5gn57GcgicFMUa0MNvecrQOR7ANG4hFd8uPTmOJZeKkA
idUxT5+CkvW49AV7xeFx88TOFR5e2u8xUalszMZN8NSzxjH+HoonW9+QldvJBkJW
dw0TYHggwkcTxYoy5eKdLQ0j4EQpLS4oO+G1THfo1kEJqvCCj5N2cZQbcqRnJppj
WwVcen1Y7c2cv/YgnqfOsbTv8mSix9frdiZWEJ9F9TZcIkwdkyhyMcQHXHUq/Pqj
RP+u8mskK7mu+Iwz1IW0vXwncz/j6rZmuq3GcfOlTmOGG4CMkfypjfxn10Ky4QRs
UGYz06qPf/cxxrA/mJRo+Rn0kY+52U7GX5+3QuivQoN/W8BYrOOGfQuW8gAcITE+
L1z6gBge5l3EAuvtWbZMDxI+SBmxwYhgAAME3cccEssy6u+NAm4KrhXQ00n7/UCY
rAQkzoYlqwRX7hM1ZwPyGQ1hU14jLiwUwGaZ+FzGWBvK6iWHT0BXgFoqLaf2lObB
iUbMq+AJ7m9IUVhi++G3SzcedLXLaPQMx4yFGPLuTRCwIn2hEdKCKeHiXGfFKssp
wVt4egk3yc1bPXIiT5S7Bf8HFfYOkjZOG+NnGUCak9ZBTIT62H4ObQ2bllBQZLC9
ZraX5qf61fTbMW1c6yJqP/FDDmzR/PpMHpAshP23SOlwUCxnkz5FgOioo1Bmifp1
QaXYZ4jeqB1inHIP0uX/vyPo7fO0gS5/Kfstyb88wahE61NNzlQ+JsAAMxCeUAG3
tJaS3QUnPQDJEUbhI+RsvvWNW1VsZOj3F5YtAg0n2/+W2KiE1see+sPncE8RIJY/
c7u4KzAmXagf00x6wGWz4zzs+VPRWiMmEKWUxi8DOACNFzIYspfZDo8PptNgKshY
U2P/ftdpNckHkoKe8cBB30SGfd3mmlaww66Hcvy9meEwHMTFQIoaGmTOe4/fe7fM
rGsBYlCFNEERWUKVMqvpUxOSH2dFeIxpm3+3rFD6yaphcH2epau8hR+NNELts+BG
NQ9f5gF1jCNb6PCjS+yW6GY98liNv0TI85hYd6Y4rkrLpZ0dxZpI8Fo40bEAzNkh
0niSQUT1QGb/Cnn7Y3mw+7s3GLpruIS2xb2vsiJwsIKBTHLaCXdHh4X05G6OGkih
mkqJS7XnrvuaNAwZJZDtDN+iCb84PFMVUIohH3HLAp8iAxQU0SJng9p0Yf1eu+nd
6ZDI89uLrDl7yaNaZa7C9sIkODY81Tdp5M5P6nknib1gisjjdYz+HCL96o1ZMHtS
rztJz5Q3ZFyt98fKI7CeNq2CJu/aHb8n57OrrGG4pmR005bx7nAtySiMoOoryi8/
Qjor101n+JEUG1pNO1VYTqnbPhMWjtHmpuLzaacBGE759ah2oe3nbEnC/E6rfpKu
RHo+Gl7746b7aA4Qv/iJXKPObiFk32RFyVX55APeNWAIRpULCqcXKE9EFg7xsAxv
wx9vi6z3LDUtsuaADUwVxNQqi++5BlrrOVd17BBJkzilyYwdPD7oore7dDVY1dA0
rERbcRzZPEZBdJ7ZjbJ+wST23AtB1Vju3SvVivla7yoN9+DjG9R6NZ66QLZ+Juc9
+iWB4c5e4R21UJKaaebi4Zpe92ep4JDI0nm7RozoRqMz4UI2LENJhhTuBDUbrv0z
KM8qERhLKIjigBFS5ph94phZeTTGE7mC62az+XuOI79uqhgcuX24cLMfNrSrjeTu
VQWvrWZskCrVPS9zxvNaDtnbLLbTCICHKumPR3UkGSzmZUv1EK57E9jGtuT9sk1g
6sPone5T70Vpjb+xw0+2KtoBcQYnCS9aqkkT61Ag6i/p6FZtwTX9Kn2qTvrkyfKT
eWz6QP6Av5meW/5fU8Xj8U/Q2a+jCuJ8j18p5tujVvYiP/NUxYrbm9ZVfZTBeHBq
F/FpiuZV9iocm6B2NcIA6B8SpwSWfnPc+tLJVBtRvzNT+Pg3k5Dhrxqr9akmAYye
Ad/ezzn2QRgquSeQiDXQVl6ztnrl5RQkHsS/+Ybhoel+QE9S8ELrDu1DRZSpz929
ZZPnAvrb5iQk6XQArsugD9RGknzkPwc3S5Yr+HtK8fBInJAqe9yuuxBG+apXZ/x4
DK/HQadgbvuoIauygoizwuV2dNulG/lSI6W2jpB+oa7K68dHtFGc/TjtvOkIcstt
ceCrofAkKYNMqy55C0awiO+5gJIdf7eviOwdxy8tW2i3tMacUa4r74l35K1GlFh+
OONtR+fc+N74H/agvnENlFjeHiJn/KPqlw2Rxox/PHQIGbLfbqUJwT/Yf+ltfGVL
8eJbRwsmS4Y35px5JrTO5jEXzGFrwG9bZZ1+CLD/giuydPP+DrWgNAmPOgNymrVK
JlAOOwhE093zO447Ow4tj5EOFQrXrTwEiyyk+k7obuSXOjrDNz26UFRYwsn+oaf7
Ic8AOjtMXJW+nTthm5w+blyHNKZ2PzM9sj0dDxF8u51hEp57fcdEYgCOkBrNSG/l
BedvGk2tz/yzUpKwwJ+rVM7NGrM2hJ5kCsQxNkRChfL9eR3NnnRYYIcS9najXae3
8pnEiisporPP56KlD7r79bgfvKnrIl4b+KPYgmBrw2FHecP57bH4v5I2pu/8gUg1
mi915ZroHMTgK28MbpSijXbMz4ov23IrGEMYCshXSp+BXfo3wxS1mF9TJFuDHJMd
Jh8d23dib/U+wmgQjWDYsLebfnDoW/0CxyE8zhQM9wVgyJvdAMgXRn1OC02teiCP
QlvrH34d0KynFEOcXPvFrMIlRmLZicMc73PA2voLkjJSErWqebuwt6l5zkxdKzY1
PW++hR5ydlSaCNK4P1RDU10ptUhNcb051n83dkvV6vpjxP2ckaWUO+IcZZEIoE4l
rp4nMuRgzZkT/3JUwrTNfYDZtIbuFSV/cgtLTtDQJ91FZTD+8rpOG9Q3+g4WWC+x
BWTvgjtGBeLjxO3aHAbkQ30XZR+CMnrLVek9SCSi0iXETky5ZUZhrQLfy+cSIY/K
yC4YdZBqLhHnD1btPgdtijRFASdg1y7uH3z7lziFWqvYgaT2G0lmLpqUpZROzBmj
I2W3SUhz02ZSeMdVj45XJMz0WDRpICNwDri3MD6xAvdidOtjnCdR3c/UivTj94RL
VRDKRW0aJo39wbiQWuCkY+C0xbXWeLBm4YDKBsAXnfFnGwqghe/ScuF89sb0GK07
XEeI3NWGDWWDMe2tujdUsi5QVoxrsKPZR3jzrXJP/sLOvjP972UOJ+27g2g5PgHS
fc9BECE+5Fp8cA+yeIe43M3RyN0ZP7Y6GNJKYln4PshQGBe/sCZrKedyQuIRMqAa
rSfZM+3ECyOJY4O5qI2k6fE6NFGthrJSEje05g+6IpPa4knyPfIzDmP9swUn+A0H
oF+6aGWwFwtfOkULHKxDLKj4YT6HhOz2ezFRGlcGk1TUJ59SDlYUhENHiAImGG4N
Dt9c9QHpnefhbpzuGmV9jvR4i3lNINK4tTP0B8AiG8IQV/FrwhbHskgsgTNMhK/0
9hOOcjhZ5Q2oWvUnx/t59fFoupJ7ALAPda/s6f5iBSawCEwvqfdm1qFdXVXiTASp
yeJQYlDoad269QK5MeLwgxOzx4qSoFQOal+agH/Mbr0WtVHPdm+j434K2w9pBCLk
BnSR8ydCT7hYjZWc1nhLucL0NDEo2U3rlLViaEThFgd2zD1eUQdS8VDOehJEoO9P
zZrXaKD/91QoYwa3dWjcN+20a2qrh/MCoceg7aspjwqINq222iggaXyoyaXs/0no
Vb+9+zZiYdEBMrZJM2tLhsaxo/0UDNb4dY7vVweQTpbRoZO1kEZd35P+Vn1R2CZ4
Ugm3600nrxKUZEv3tQ458D6ANwySwnIJB69oRB3vmX7AFyiiW9gwdX2pT/wUMWC8
eReF87x6jcA00S817xhpz57oZgjLAMfKpLkib6nHFhXe9fLz3vBazFKkEuA0s12U
Z16EF874exhmTEDHSpD3JUtDH8EVvwPAbe0X7b97bsaedTyugpBsF+0ptyJ2yx0w
m1B+jEKbJfvTf5GjP4sHNDnxOdYpMteXa6aHCRhpad7tCMJ9XYH6cPsd7fNhPzvx
nHZxcTvZ/jdIgH6F9jmT7SqaNdipjrq+f2mDgPDrzT1SDpThhf+pj+YK7LJR8F6y
o/nFWtmkX9G21vcMAmBSwrcLW+CleMt2sdePhhkjQnbYK6P5xgxDmzU7/JIYxfRX
GI7B66bLWHjBR3uuR4lvm2OlaNS9J2iPtcs9ruOnyfhiECOEG7hXwkmieUrUNI3w
aLfkkosdvpfbKT9l4dOPUNIg5admhuKHbKpQIjF3Tivm1GrtloG1akQyyvZrwdg0
NIlCQ/3xiR1lhNFavxBdY8FpqsDAoiMQfCoX3XiOdX8F5HstUGQlXqj26E0Is5xg
Z3jsGQAHCnXZy0SdKvhZCFm7xv1v7DwKoLHMy6iJpOAslUiEu7mDXlX8mBRVp2bc
hS7gQ4nCXXOaMf1epv5uC1p/BUEuhh9/3upLv/FyJnlSwVaqARsmmLeKBSfEJQwP
vDyEdiFg9lGZ+ulgqJpKn7dv2MjqtBTXIFbKb3QDhlPSvwRqIiOLQadBQicCRCz3
SMwyC1rfIhOAC8kqeZh0bi9WJBXZcZLWnlpDDJry/uGHfZ5+ImzasigGQh8EzxGA
cBOCO7uAlGA9t2uIAzixhJtJo+cWqvuM6Xo41vjHOsYyDJccj5wjN1dHWreV82+I
q1GRwBrtWvTrXPDcu21zJzuaF3PM/bzWvKolQ0RTrZO3N96XUrFcq6kkjb+QHI1S
PeLGD90BVr4+6CYqA8R0hyh5eTHK+BXyK2/hN4Rls3Q62SFRxSE0pb4aKg8c45B9
pwwLtEwVWb87X9T5JMK3qatm5wfvv1uoRfGo7xP1m/M/fYmYbioAg8xUticSn5J8
N1C3DHW779lplDoKNzvCcNfulESEmsESicyNAFBIKP0MpXqx0wUQQy9lpDlesS1M
AduNmsooh6oqJ+88sKH18IfoZCAImOdbd66GWPdnOh6FN1T/6bk5AmK1SAbhAT1j
LVD95dPOY76faSp8V0VzxDK8YwTDFG3cl8GSIworVCCnEjD47ZrJ22IJRdDDO0AN
mRoytTNOngWMEZvW+8ziZtY2MoMt4g2KEKv6fFk5edcifTB6O9C7Qc+vHLu97iRu
ei/AuEwiT21XsD+ilRNrs7XSf91hy8ow+LCTuozDyq0ampkOglCe3mH8/OH/ez20
AU1DJUc6/pBA+koZzOlQD+Z5DcDBEmCY6WSk9sLAhJGirKKkq1kaj/0e/5X+6XJa
4WiEZCbygg97JRNWttvN9LI5XV0GwmomosxXMGxYBwtBhTnsa/v7OHhc3PEZ3B4t
r1E0xXB7fsEcggErc+LVIMi1XsfWsP8z4iXlFEvszrbEROcWBKfJgDlYZRaJ0L42
6XZs3MOtbSkFXmLznwkWwfo0KNCwWvC7iSaq5YTAUkKmDiNQrAIdQowf1niviEvx
ITDfm3q1VufKx6Px2szCjuJq4F0nFpXhvzqGZ+K9rIP32b9vh3KQg4EQNrHGXZqk
Qu6Zcq5MgmUEOptHAPjj4AzUMjn1BvW5pg9wYWHxCACt7A5yfRuz1ECG/MPKUJm/
O9co9LX3h/kkDBlu4fADUrkj0e//6JRld9ORWATAYRlkZd4EEFOOBGfQQBqpgc9H
57mX3f/YXokntxnVTqIHfG6raddZ3JpfHND21of8Hjr/b85i6vbgtQD8kyg3x9Vs
ImCyLSV0qwy1CdtIFOkoZiGY4ZK+6vMIbahXzUqu/86XiILqjlELm/E5E2W1F+D1
LNGWWEL242L9FnsJ33/1okrC+dhm+ABR/kkNGXUQjzyu65qwFDnWUkjQr96tUaZn
DIFWrteLQU+j0B4qtbJs6OJ492HrjR5dtEvI85jSDH05QL3FMDVZgwlDGeX5/ArN
M7XVIXvoyLmTfgmZAeKSc9+MQBBDGqcdL25640rXvZe98x1Szs4Kgzh7nhyffNPV
urmOyQkLOOpz17tJyIrmgebPUpZ/V0t3d1JF9gNFlJ8mJqkPEf3MIW664jSVEF2U
Fv43m5rFvUt6ZEhbP5GmMJ5F45yGuLuVq0yo2wS7s8bJKeD4F8ngn6Fr9Ey56A5J
GP4YgzkqsCvkDRWtbHMo7hDFjlTSqzimcnyc2rz8j0o7SdEpfUyb+6giTwrjg71m
p6OwS0TFIqFwZlZ0a9mtcLuYgoM0+yH8uAITHXnzXAQDvrSm9U9VZrDEjvZ2VrvZ
Z62m8Im3NfX6iFOR54Fwtp+IVMPpSYeUZgE8+gzCo/BqEyOdUIcU1Pgp4IKFtFrX
AXDNkTHQYPtcwaS45LTtC+rpvDyyZ+sALgErIfSL1rZytRqV1Nxqlc1PQaPK8ftr
ty9c4wHbFBZDUFrOweTi0ie2qlG+lQFq3kKgqa58nSJi2RAtw25bZDbTr95qS0ML
3wxPIdOZVkQZqYbZUDm2HyrYxP9F1C+NwG0HEceLyOfcuZjGcvgNyfLnZYpBayXo
e8Odeq/WMYVPadw1v0Cw98yEdrdeylqHPnUJWFYdrO7EGLoea9J8rlrg+ru+9pXu
5CRIwZHSc5/P0unBunesgCgWVzVObfifeDokO2neyLPBYzicISEBJ88auYKFMZS/
BDZO+oRYZnokAqhEQwBxwBADcO6S5Xi40jfdgVu6RdXlqskTzkS43ulXj+VyblI/
f3YFLrs2gIcfOtDih2EfYqCX0BL3/HlaH80uH8JmOjFjGgft3t6Din/H4I24uABx
m7jsxHwR4h/mJh8IW58aV/xKrH0UCa/NE0tyt76XH25yj8BvPXaYquEJM5BpzRb1
BKBAGQgN0pN2vZn3GRixME2GLmmVurdTOTiUN9BU/UtavGBacZFRVJflydA8ZNig
b4yJxsJJCtktTgTUXrQc4K8ECQiq7YAsfc7PiEVLLQ6xY4jLW+Nbuvez93xjP/Oh
d7TzYOCQdT4AKbwxMwVqFe5nvFLoGIFbnG72O63QwT4QzK8HYIZRd4NX/PuOB61f
h+K5ko4bB7Jhw/Sc0IPhZutmnX/RacYd3sE2YUhH0KNcBhkK8iLQM48o7F91uO0+
dAB4BC0oOZz0LHoySB/csPi6hfy+gYN/e5sVx1v/YBQ9wz0Zhjj1t9v4xGlY5Mpc
dmntIsQdpvUObqd18IEGXxOxDek0w72ebfEWUnQUxZqAbpbg320W3MB+OFJNOemX
0403EF9YjIrmy/47oVbXgfiANyAa9ndXp38poA6OyepG88SLbV3oj2MmBjLq8jBJ
IR6ZHIYk6g+l4espGTXMz9y/re2TDRUsZ+/nCsWLi7DHvY5LL97EOvOdQP23yGPY
uMQ7a3+QScz7RHMCEhHgis0UkMLB9XpJxsAeheZYFjojsaps8NPTw+feOALmBwKZ
ggBkz6gUucJljpCRRcjj01NCIyXX12lsuTQG4YQS+r5jAYt2+kE9J+lOmsUEkRrq
Q3u926gDO5UIx3qTs8F9vRdi9DmBcc6TVhD0GzDX4yYVA0bcIFa8nx1lMs9zn/R2
n3IT7iFtNf5FYr1oP07dOOwCkxTyTivNWqw5sa9G33A2MAYXadPGTHuLhThemYbE
58m1qY51CqIjhL7LNr5aewnIrAOnrZH+RWosepgSDA1h710ViNlC1h2GIPYR1UVd
nffvuZkZdPLA9cROSNoWfm7BIzN2rZkDzT70IqfCP+1hWybCjAdZkSiTa2KgcJhD
fJ6UyF5WgSuneCA1vTCykp6FVYo1hEU2dOmmnDUxplbp8KD4P3wLlKsHOWr/Jd6O
aua6+cRDC2OR5fgtM0kl4faSFJ+ruD8VQsPAaroWdpvj/LsPtGh/8DUY+SlCVUp+
ZiSxuyQeolLkT9JeI1Ofz3jGb/CdCVzEMnW05Fi74BVtx1eKRRb6Wi7TbxEQn+Vt
xHqQ0tLvCHfFpXu4ROuV7CMyyRUHeWT6zgZTcJI4QH2ykYdw2lcTETMgmRM3xq7j
5FHJ522lD1asgEjoN/drbz4CJQDqGf4Dg2nnZqHQY3LWXWcaWcgpI7UjdHh5jMIX
ZBLMJHPaGoMcbB8uRBB/HJ7SA06oMf02jFwqgPmeKBKvx+Cy5Fak+SkhBz2b9yC7
i7xVN4KSfh+y57NyMw/93Rvm5a7TuYP7U2C1x0uQ/+3LChGhEsDoRdBtf2FmoQ5w
3cEw0ah1mMupwxArvYzx1fx+Om+PYEib9mEv37935PlYtl6EWrfz3a02PYbEB7l8
K2ibBCIdLc6iwoddEdfePUGHvRTfjVm5CLtY1KPBU02zdEOSQUIx4U3Ox2hSn7el
5sed+qXDAxg9RFSQG+kOow7leEMulve/t57iVnBDjtvDQLzCPkh7MfctwqVWL68k
C3LF2vIooBwJAeLBsEZSNXoP1viUMcV+krhiD+7OXIwF5dZbZMWffe1V71JwsAqD
vK0f9XwTkFFd9JD1GlY+aIVje54nhwvBga0XDhe5Vu6ssUTKnWlQFDAqdGxhEV67
h4EpI8ZsLzgOh1oHnDsIFO/sD2M4ItUqjplS+NLM1Qyh6IElGoXVdJ1rYyO76igq
AazBHpQQuTY/8X39DRw5P2ccqrmCR2Dfj1swWPJ3ql6Mv3YDQ1Qk8ansIH11ft2X
0qcHYsjiiNyK4p4hl9CT1yYkc2np8rsCk51KmgOHKJtMnCQP3mz86Fa44/drVkwo
ug9fmqkf2NrFR75By9N1kXjHLO50qbcsagTc5lfYGuO2WSdMIER/ddXV9fJGZ8C4
Miuo7H/gHq3POuY3UocOc4fOUMIIB4hR0mcfBGTt54Xdan8OT4au7SRgWX+GQdeg
Uptdo+6gRXhl2UbfaPCWIAXDaSBsw7sj73nsHkT/cTwV61D3kUo7JlMhZ1q51tZh
zK9ztlSCNnMD+Fk2DBJ+5McId88zJEPSd9jrRG0DqN+SlQbO64enYUWSjugNkXnt
D6BD4wq07ugFpfzj3s/KeiJFRthwFXHCOf9awflu+FjwxtZ6h6inaRkZehBO4ixj
wdxV1eqWy3dSnVrTvJ2JvGB0H25wHIB0eG9Z0T1B3oEdVqsg/I5jGL4RXulitTI6
MB1m6SGgg9Z8e/NyvL6GUhckt3P3jV98+HkWLATCoITXdnZKk5/cOugVf0E2lQOG
zAXBOj4f+Q+SyPl5Bd4Bh9ipGP9nYC02Zen+z3Z7jF0nP6M6Pbydk/fWf2Yen8Mb
rq4qBThPV41i8Hwd4JmLR70daJn/JBn/OFnn/i7Uprr8nvMp+rb8lsK9eXCfzCTs
IzdDwgIlFCqRYf6rO7SU2c0d4BbelAtw3mVZw4vV5gOra4MRPvTFsvyiwi9kNAK+
KUyqbrpFNN59/8M/iecbMK2byD1nGgillxl2olFdwXGVgXiuKz4IHibtkD9HlxEI
GWG70NlmAezHHZL2FNCgQdNrlRVVnPZcsK+q4yeNJzvea4MR5M7Q9sf/fTt91iP7
kgKGGsjMLpE7wcRmjLNqeuFGN+NJ8dyvekD5jMZ334FU/C+J6R51i5EB7shhDbVm
AmcXrOxD1BKekuyuPbTzRoARQ+8hHeqR8wj+LIpm4uq1IBPkiGcJ09wZGmjqibLw
m/HoiA5JXIJ4d3ysldOVm3tqm8dxrMBKwhz+McGnwQdmhRqp1VuaUkizuLihtwhn
t61XSbGlzVuoXqzz1kYpAL6IPIizGXlVwVsyNyEWfW6Pl0rqfuarDB51dC1a3Rov
NLRFv1Uai5wdvPLfVJuP+B14UzAbRC9ZjMSUdRdT0z2bCtCcmEQhIQt/5nUvRP2c
WXobkL6dQYhuA7DFKLBadV0MY/57q2oYC6wAVSK4CPUDXQUg+GRB54Ks2fFG6UCw
v8YINzXIKJkkjCgIuwvz3BExhRpCSuiDGlas7Z7IZ9ihWggkkssW7DweUqpP/K8J
wotbYw5fU529UCH9+6/09I1HfnM6d6bmIrHnjTNhbPyIc0Oc/Ka6dLQiTBJMEKPI
YmPKEB/GHTapnHd1Tw/6rjPn2xdMPtMnDHx72KLOwnAjPjWH/N7eFqOAEQSVG+nL
4CqF4nWByVZkgzlURB5TSyL5oYimn677wROX8N4D2RJXcvX8nUGaAohn6pBPhGrS
+mgvTTzjMDnjaxJHGlFEGC0NPOT1D9YTsCZzJAqf7AU2FXerp/dp8mT6ClNXWvus
9+MtpdFjDu9KvyQwWAbTWYYEfcsXBF0+twvjkDXoqJpbTKtWX1pkxdzxGkgB1wa5
CpDcvO/GnEFQLwUh8RHotSfZ9K+iYtWacZ3EqiGgcmJNISVOU9JRZl4gUTgTwpQY
KrjPwmGU7JAtm3T1/QLVxKPfp+vqOudM1P8nz8wHJHpRJ2LEE0MQMkWiClBe5+vV
trvdhmPgItyrRhuAZpZfefvltgFQX55YdT3QV3LwCDYfjMj/F1/MX2uC6pqMOsXZ
sbE1zuc+ajDQLmg9MAT9LUIQj8Um/eTBidimzzBUtLdVB97V6AEGYeKhYg7clhSk
PZ29Rgluw0qd1xDomx8RDj6vqxwInt4ywOwdGRLPKO5dn27MM3xNQbB68cC63Qxd
el9IE/vps6bITdhoH5NyOlG4QHbLf5+Mi9PAglfyEuNp3dznh5bw+3R3czh58rRI
VS29sVu/Iu6sl/WnNWnng3OAbsH+LAcBqL0zCD0aqR17x0pRI66SRb6V4f6vdU4W
DPG1EBKtFUiOWfYrxaekhgkDTNMxgcN5R6xEZ8bnKPLBLGaNZ0aEqwLCR0bx7AI0
GxJt+8kRMhC94rgUtIexKbUi9A+mR8rrOM7xHxLTsCsr9iI1fN7LLJfPSGb478Ah
Q7xV1Nq7dHEx+Y9AhauCjzT71nJ/3Duxz/2K7bxdY9nwpn0wn0xlYekBURsGHh75
08xvqvkvQ+69Z2EzOBgnN6jJrhSG35SSN695roAyNDFAspS+PsUX3uPBOTKS9/bo
bZ3lEG+dAWJTEb+rdNzsgp8og6rNDvfrtZDEu0Hngu95hDYQJxyFb9gscqJTeij7
GGzQFIKjyDiT/PgHZfrNxsiV8mQcI4soMPjiETch4heXzcZj204W5KfETaWsc0iu
1WzYeQ7ehViXswwrbUHcqBN5x5pBvpfkOTHL0jy/bDehxatC03SgQQs6R3Rf0Mbg
mJDZlG3/u8FC/8sOOL6RIMvLIbjnQsQbQAaPzoVIK+88qQgJl/NEVfOJCSy2Fy37
4RvNRrjfpsBaDsJmCnG/mhi8PTHkEbqPSILlpKkJhQaEC0WJPrA8sG8ELt71a3l+
ppa6iEhZDeyYFQPGVx8vwQRl2h4NDB+/1XTN/WWz8sb/PIRqOnKyAQ3JqDmcbo9R
/BhPybauxObl1zlXsbnBj1WUyFepPHlnpBFP84+na8hwY/HqbC8cSJGpQ4QGmQfg
xh4xEzsdQr+hs70hIDcHJhBm0bD1GNs2dXcXQcF8/Oz2zsvCAoTv7V//coCoMqjD
YNBeYt49kKyYduDnZl8lXEMqm7qFDBj5cNV9lXWpx6hm1V0TtPHxteWxodMcL5fm
bigOmtxvjcHXZt20fvZV17MqQvH4pSRPSXFXeO+QxXz3n1BHmiEd3Aw7DUIRM3vl
Mq2vds+gTmNEVu9GIRxPlJ1T+MMxUXUvDuBgFPeaWxd/l3lCPQCWppUAOQSsARCk
3g5uMx04i3K6n5e2pWhCP7957QF5i/QMrjcYVbgmgjoMKSoBCdKrjj9l55D1vnLV
jBTSkquDUZkaSlDMLoqI+1DneYZRd9p0ekGEE318Slcc1jWiPCqS4oY1hWf5mKLn
1WsKr1t11SUeOAAaZq1Ju4IUCkfgcLTvrFL1XWxvVlMDIgUWrN4TGaMO+thDZlwn
+ijEBXvmBqqJmcYQ7vM5+hcHxMic9u1lrzdVkhVixxM0RXFJ/DgEFpSvdXLzKJWN
7NQdcYgueEXOf3tnfA6/xbqvSeDPFnb363BJTcGc079RMrCW1wH46jzgUFME6T/v
9UOeXZIzFhotuuD/tIP+IQRISacOkdJ4CERQ6ojTH07hjqZBdUNhpfyrLWXOl7Dg
X8u8rZQLDUp7+WH+tAfT3ah5Ah0UqitT3jDuE8EUW59nZ7mqUqlqvnJZmwLKDVWA
fnR7l/0QHpKq8RkvzFOpKSqVbewE3btybbMnz0PuhjK7iuDs611OYT5aD/2qfb/w
kujDDne8fhjvnFZpu2VzWTkKVYhyB2UlBK0K2wAG0uXmm1DI6QJeNBFd0SJm/7MQ
zLb1q9M3O/quQdOgAThxtandlBbF0y8ZbRsrh+7n5RzHaNOtLXxdCHoI5oFTm0PU
3kkTdv+9l9o3LndVbO3iBO0ENv4HnlQ+jRhg17i/GashBIUN6LJzuO/Fjqbl3n+K
yPiCpGQX+TdXbwicdIZxcMiq7HXAvCDvYt/yK3zGctHaMt51H1exz6SnrJnB8nbT
Cp8M+OyiEMhe037SHZnxPjzOF2OaseVy8nzHh02acorXDikI3AZTzn+rF+Gx/yi/
A5dUnOoMWvW1AuIPVWs3cs5QfgdwJT+IcTBnDhssHDkqfOAhOxNqq0+74nIWeJlL
1fnnJZp+3R0lMkU529NzDU4t8pTvsXnZfdM4lwAjJ6+WyXad33Fn83065R8ivGIF
KlieWY1CoJqzobp6iLEPxSMqNKX/vmEDCfcELt1epiZOx5Rl4HYg+WEfLcS9nOrG
qDej701MLiyAe5E76RuT731hViM5DEkSOvJifald80UXyWxc8YFS0Zrqy835cS3P
MEbjh8B8gD60V18n0X0WkjlWBSJGV7KmxOm1vf36PZThNHG7wnYHwWxcoEXRHV4J
3QR8F4ysbJFjl5XT8E2g8Tl9iIS5/L349B7iHDjzi2hv7CFzNokotPrWzyESAF+o
gToiCINLb5PXR+PVhPmq/i4hZcCWA2kSKKQwBLKN4EpuS0yfYiu5tebCRV0eEBCd
OI3ZA6elLVI6jPFoMoCqxVS8v40sXbxz1QP7ll7D+rPP/x8Av0MJQXJroTYYo+9U
Yn02Igh1RwpKetKffbNhc0PJHIOHbNp57Z6ncBmnCNyaWJM0jYrDOwrKZCfrHaGj
177usuM0HKLc4CLFc1hbASberb6ffBRJt1vMzfplwFQyMPb2xJ1tkr43w2333RtH
Pwywj5Ah9e3cLRs5zySlfEF8jbjDN9yrzcXJc5mCVnjRT1t7NR3inHjudc22lAAv
/GvSkk7Vsq9LNMhIqemxfHhfjnIAEFwu5MAfS9lS+bggvtGnKgqryfHrLAlCGt7E
16TYTPkeVN/56nBYL1waT8uJXgzUgSp2xC2mIK5aDk5oZO/GNSx2xEKTamMYDpJU
edcG935v8G5hLia/9Jjc7SN989pLiruqnceffVO/JlTOzpG37TjV0PD3AmilUAlE
tlyQZB1yK57H5bYQSgop/qXspzXoD+KQ8f85r2jQeHHzo/lK7qYYy7DWnu7PcTzd
HTRvNCOk1c9M1hA7kY7tvUsp7gkzRmTGV+a71fE1kfXpvYdjSuZcw8dSW6jpAZ/P
Jin0HeU1R9o5Zg7BJXlguhtkfmZGH5jwEuX3AeNJD57gr9sdgEz1YGoydZw3SAqP
cgKNtIzvuFlWikdblYqpPc+sCzHAaNAKSG8UNux0a1AJQwv28xsg/aPPAu2uVCZT
L5c/pZmye6RuMbqcDN9D1ooe8HqulawJ+wS+BH9TJefHhwQlaF0FY12JwLD3GWS2
0buVnG3MU9EDF5sUbFVXjMhztZSqT9Ehql/sA/gwcmM7nD2vAoEdLxSmtLFHvCu9
nJo5hdsntFxE0DcgpVqREJQPpouHzK6V5O3r8zwCKeKZsecEpQ/CFZ+fxLutcCPH
GBcbQHseoWol/8s5oaaV7MtcEFecR/t+BGkEjjaofcWZEUylU2LEyj0AsDpljGz2
9lV/Vy8DKm33g4nc6Q2v/ykBHUpL1YSiXrDFIPjFBhV/w6G+blthPeG+CHPfQfb2
injushgQ0i0Pb6cV2ZlZCOOCO8IFAk06nmkvjbJUHrMTP4Ea7+RDBd5Cj1YiZi4c
EspTmS93293ON/RORMgns21lO5hGGkWt62QvoJ6x+oQn6r0XSRXuezamvA9wBCn0
5gTdKT0VsVcl7bgTZYvwAWmATSqCYrH9ordtAsSbuxmFH3JseUpt40GQgEGdIpUx
IbTzkfwKt+m5Juaw8nLF4JAUvJvpODAeWhWzDgqJmLr+8ppnPe4CCSxBcdCkqKAP
z+KRnCOOQtgJmN6LyRqFdUAjfEDQqDh8nNzbXUZxgkAWOu8yAlr5eC4nE/v1O7ro
6w6OhpDYFBOgDOjTBSP2OpE4zk6hywGB516MeBwFc0z7lOk6Mallxkf48a0WKTw+
okFU9+YUSuo/HHtaKm3J4rBDRzNj+fS37GGQpeHjmpuUyLltx9JIhUXg+QICmzfK
86Gfyn1DhNeMcpDzaKalPurNwAleLx33xH7nBN65YMX/YHYwX0Q/fkJ5LSUzj/hZ
pjkKNkYHN8aZsCuCS6AvLsH30Gzjf3SUrUt/Ri4yBWmm7gRKJ24SEUwMbKLwkcpu
RUxfju+nVZP4tZQ/VBXfWwne66GXkcpl2bGIoTw4bzFClFmmsgf73yg892kPzEMJ
pVvg8wjzQotI6y6AweObleMDC53ImJ5xQPAxWZbm9KDqf/8SdE2EZ0ep11l/vC00
56hdjyVPvOqMd/2OLJVCKlTdS5BATc9PUK3cvAN0HCHihd/f7poiLpOSrle0dG6n
z6DgsLFiOHnjMPpubWPxg03o8gBwEdj5XyjySfMP4xP8vvA6yPUvYLDeKqR8oC9w
0Vy3uLBu0CFgLq8WUg1UPh2tchg63XAq3JNfsbspcXO/APcSs1hXI/HqWgrgjpUT
Gb9Aw8fcJa1l1yc9jTSHvQIjdhmwJHu/a0gn3g3DYOADNwiQ30U8VH91gIF1vEBK
E5LEcea8yPczkKmXoYHuN0qqqJe0sGgqRjP+qO2QrqXKmXCOz98H4weGjEp8RXGE
Vd9aFvzxNcP58VxEI0yIxjGah03MlCUH3xE/uoJ6Ql8AycXme3JPGj3FMbN589rU
BrVWXwYoXdly0MVrwfM7FNmxsuZibPEBB6Vi5WWXPJqa66Z6kFnTRRRd84nxpGAC
8671G9erCAXcWIOLQOblMesxE0ozrKejpHhKXG8lF/HNA8Mbv/D8UQfmCYAzztf2
n1JWvdsqIUREZ0JHEqVNQULJWfGx76JlFXrZpX/NFn7h1+Y9twH4mpcqWLtieEzT
p5qWWWvblCR23x3L90o50G9ALYwlDnn2l3qRk6rrJK7UdlAB4Mfn58yjnecjS9BZ
TlQteWmGE5zvL35FzEM8eDi4o4MjpzaQbsvkY0zFAAVyRJciwxCFBfTXES6TZ53I
DC9jchaHsmv/kfRAUJXa65+lHPms4FeC7I6JquPvjUDgL8YMd0QaGGZoW8HD1/Dg
8DTSh4mVI9N7eC0xnq923UGhOYRSDvSqxBGFm+235qBaEuMMHjyb8tOs88VwFyyM
3BCQtlSnK5KKmqbbIaOP6RB8EzcBbVwmoma3Kh61h1P/Jzaww2xo4ABIrZqeTwAn
o/xpW0iuWaQzub7HQoNYwHdz2xooe6xCzeJZrPcWkLCMEkxpoH7HXLMPZ34r1NtI
FvYTWi1d2Ah38E8pdMdwXs4y5xGAg6XqUEacr3+sdJlxU+udxFXl2TjWOAEDo1xf
/jx/gd9sozXdsAmaXfo4+V8gU6UIAPvtpmp3DVMlsghz5DlP2hU1t6zfG1ySHG6p
8bW4ss+9jw4ZEqcLW61jOGXiNw0QHxUGUt8ZeRrEhlQ1mUWHI+i1HZ9TsZPAhp/i
NgcCHEDPv1TdMDSf5YvgfXPmK653gtN1PodTmYahQUUVDu9VposkX6dAK+J7Q8De
PrxFy6ud1DG9xGTczguGrIq/SEy03Sbb6VeoGWteKVuyA4TZ5j8Hd7PrTz6p8SX9
jT1O2RwdNnTEgSO767zXLQ37BhfB1zevMXVuDy9H4hrTXZnHvg0yVuYqyqnqribw
gkAf2dEsGK14jrpTJT770ZLAwt6XLzB7f7jsp95f6w8gt8xAkRP7AYGnu10oul1l
YnmF+Ojufl/RgIZu8MpQXagInQxk/6LIYPe7YywJWiEncVUyLrpmXGUODENRdAmv
ZVukpe+9IraFUEa/hzV9WZenYTLQD7ELRfA9xvgfgHFa6PXtE0RIF/fTKUf4FhI9
SZll9iE/fh7OPOxt13olNerIbHHhOIIAtUSeru2V3Z00Onvx54wjLplYWZ3OWUQw
Eq4kp2EQ3XjZgSf6qZpWOWr8ZTsXOzrLrJWksFV0AnxfubsXvI3Q1pgVEKnRJuQr
+WA6ihx7tELdIiJzDA2KfWcqFxeWCeIxqVgihlWvc1MSbsmyuCQUPoZBXdZr5mCv
Rq4kFrzqs0NUbYyDDr3A/DvwgRIE5MgjgEs6tjUpWrAB/1KE3q0czL7UOAd9q8dz
y5EulIQEHXn+f0G+QC60rqvH2TRRfYZsWEE9XNK6EzADGXn5272dId2ukC0z2nPf
1QUWkMFqQjwPGEI9ItwDXLvXG4rZGRQLyXVTaTVRC7xfFRAaUC93po3+0sPbRL3T
/DKtM+zrwEOKYRenBTx6aWoO3CKsVJgRnn4CpnbnEFdDJf0rCgLEv75cXo9PBvbV
s3jrzQNvKzwKgDdsXhHL1Q7OyhFFbjaeyi4zs+ss+mvq0rlsWzzoMcrbKSFbvH+g
2V+vFf5PNmpueYpe7OepGJS+IrT5DERXPDNh8zi7XIxurOwhI3YvxU1TkriMhNse
RHam3aNNFrPwTq8YQA2qlGfnGfqLpCDn75EpYSRPPiBU0It5tJlLsyp5ay99cNoN
Eq3f8OEO/qupczS55ruk1FiphoeCJCC9c4AUc3NoPt/hfs8YOCVXs8WCNNS9RYJX
DsguanZAemPMPkf1nrOmwIs7UptU2zkNkasVt8EEz2umXWALGwmYkbj/mVo/DQFq
y+/hZMaHgH9l3ECR7JKazJOt4UkdXeeGNjv09YAuNqTR4KUyQE2Lm4J4/LR5WqN0
vonLCl3l5a8AjlMQ1S03tbpdz1CilsjSVV/LddVKoRExxL25wWmkzvQ2neTa0602
lFbTvfP1Ql/nYxB53GNUyJ7Xxu+yx2UCqa9SStWw8blLmCpilgzGuZe4Bx6IyI2W
MOJ7Hv4fM5ZomFjjSn0s7wKFXpFEzOVI6RQvufDZ2fz4WiRmHkVdD9Umb4+jBxip
kZh1dF9K2NgrTHVH75JwqxEte79XzKG0iatrMBNnSpuoEogN0KjRaoHopkm0As2y
oAQwAd67ekvz5Mn1+a1vizJ4zzoX6/BAtNFcInGYTpxeJ9Yixi1qwtAa6t2+eO9x
EjenZ4u0IIiPnaooANMmcb37AnU7P6wD9zXBFqnq9nKHTmuSJeIfc8Plak8xipJd
wSApIoOkS6FG3cBKZubnVZW8a2DCL48MCt0nezutzHu1M3w5nA8Mfd8Oin6eE/ot
hcoFJ4Fz5E5vVEOyTK2kI63TvFGyt9k8UmeVoxGnl62zegWt/yqRN6FeYDFo84Kr
sKNnuobUYUc+ngjmxRPK+UK/PehwTRUy/HLrERTe07TXh1cHGWVewPc8Q0omS/1P
dIOQPD68hpQlBYsk1Yte4ljeRumVtc23an9QPahQFUxYkoqELMXooJ0FD5vfHBmp
K0FMzk8ohcGw3yj43+r+gWTMkVBAw3KPnz+7BelVcXFZuG0Fnh4BRFBu7rTnxVVV
X7lkWlUfxV+WbnMg0N0qRQUXH07glGsPinUXZzPgzBlEAyRBaUFY9sug7mt7glm7
RlX40tTrXjwcoprecDk0eexyExeZ+nhWabSQHACLpuEK+GrFBD7TbCC8cEeSKMHe
HDXktyZsOvKQYzv264flbaFWxf6QVTOR4OCpGypJFmv6n+CVHBHkDCuc5KqU3p6p
AqlwsiAb/FARdnVy52XBpbSJsKWAMMM4ftXdsZGldWcaewGBVkce1XaGaWeC4AIy
vj3EAptaGYlRlUGIbtx3BDo/2DMLSgpM9Q8GSEgPotJDhX3WYZ3Eqa8AvPXO23Xe
Nug2qSq8xlDxahhX2kuFnoBMaoZmm4praxNod+JHMlCtitAtaPnNl9AHvbFPW//7
HO+hHNQFqPhp6BLwppgcJLWAWLVtD38PyXHoNaOW6CJD58zW9r5XTcRKBsQVt1kw
v5gtNnhtGiFEzNZTQg/btA7K7iZ2hc7GpW8o1GcsKgKgV8K6nTjMtHCzI/WreJFF
bNhkNckDXJeXSwX2wbatZok9jdyRRBUkeIYKxD9jhzoQMdKpyot5KkJWfGBxXvkx
1T9BwXJjIspIZOyHKEbbjnYZRZGUpB8fGRzwYiprDacnh9pj4JhB9DtRkm8OZbEj
+QO1pX/wOCjpP3BzSRi5yYD6ml6gcuixCYFU+VuahFuU40+4y3KxAPUz3U7v4nw2
vaIiAA+A+COeTy0VY4b7Y9iuryWMWaSj1ACrdKMruN6xJ+QvfAPZm7aRbvk28HPp
1dsdb/D6ho3R5bJLqGnrAkO2ToypdFgJMyDeNuLdsVdx7pYzleR6grPcEndKQfn3
48z1hCR0fuWxJHR58HaDSm36HyuOKeoPyP1j/GxFk8h5+iMJ5DtYoEGBNki+alg8
KBko5PDIBTCdHWsScN+MJ9Ul9n+GMbzuGp+i+iFp/fFOJXzD7D4vZnsIXZnyNVbL
OFe9h1E73fW7WBU7ZEjZRKuvbxiKzGpQHLMR/rQs+bmmls6EEZIi/9bhn3PMc3rL
21H2daPmu3P1NA/AbfkdkTbK7wFKkCgbRZ1TcGUn44D8GR93yhLU1p4buXiUDItf
x5lt3I9eGhyq3fMF4sDeO0WVhXTVKA35zko6eIpBFVfp+ia2qmpFNnPR9SAgvetZ
0Ow8nm0diJ+TM2fOirgpCudePSuS41h+1G++oGBTpHsOcCDbJLl9X8qetNBgttGg
VP0WfLU0NzJCGtpfDaVNZOdetavuEZn4gNKnW8GzLZQKUuYx3jGbpZp5v2g+xmkF
Egva8hEURso6HP3HSQOuB+DEMRz6Wu3UCDhwXVI/qxQ5q4C3rwtjJR/EuEgyxJqG
JoXwOs3mmYXsa+oSVfv35iR12r6I6Eht56VzQiq8I0VABZfBBmXAMDruTNbn8i/P
nQT8ZKdUuS0hL8pPTyQSd/c97+kPaqfd3a9/Pas2E1N2oQH0Tvd3v+N/MGDYh1jf
BdMeEQFrn+EXVZVNsAvJNpeAbmpVVVTyowt6la5Y9XgLX49vqVRRK6ijwJC/U/Gs
K2RA5aPoCvDVQ1VGuv/jI2Tzvhlbji35F6x5Qw2j/Hwi/44yXoUcD/0qinX7N6aC
Uv4nBVym+SeRCFxSfuCSCCmiJfS7P5XklUZDy9XnQc7heqUNRUTv8fvGB0b36UG3
q4W56LFmcv3LPZQmMz81A4z8g74KDBjItAzhmRp4pFm60ybzsyKDGjzdt+pAepRk
oXQLzHUy+2yCozf9NnJtTNwlQZOFuDbcaxbyzhMm73LyB2TO05jWzdC6fOSAbk//
ciKvbI98anRrbkfGT5rmZ80m4/ES2DDMn9t/LrO0KwQs0I0jay9HstvrBzWCT44F
M5aADDwaoNaigB0vlEJ/qWR8mTAQWOKmJX/X/kHLS9zCEI8ngZX1pi+axZ9xodyo
1mb9e3u7uMdY2bcYl280UILGyxhxYm80hBX/oXTnzk6xE7tvRi1bduROB8TQnfDy
X6QywIIl4jvPzkWf7ngAVzufBBuGLZ3zz/9cwF1UcBOeHlOWivxPSTWn+5lsCXLU
1CEy+vufnTsV9JzPEfOd1ML7IB0ZmxBNEUSD/MsQjampCxBzCOehEqhmQ2kpZF8S
Qc5ZnoMS3BCmFKaufLX7SX6O6YLOXEscN41xywDfI116GaDln1013ai/tUr95iRF
bGTB6L4oAwCrEcLasrPsPrmjIXdcYb7iyXNupj98sUaUiqSMGYoGIzbNStkrmxNK
n21qCOixB/OkB+cPpoEpoTuniUzjmUBviXVw4amOgqsA9ycouO/y7yf0/pGUVKNZ
xTbPcCH+/sRwVjR3BJ6SKPVzYuarpBTj/cDG/njtN3dR0SVXIi9+5NiOAnosCT3/
yGeMbrLtD4e/eUButDaCkvZ2F5ftIGzZD6PkrY/8tzy+9Sr/+Kp4b5Rs/2UxVkEB
u5TsiRuctFIcqRQP1Bld+d2/WA9OP07zZMlu7BeaDfsiRr8qJeZ77rqcptEGGPsb
SrQaDDmcJAFE/icj6n9UDcU6vCoyp1A9kVKQDR4TWtJ9LhZH3P0G8q7q09SxsI2e
Vt94tEJs1OlkuE5XnTdicnRLx85WcpZdPSjVNIpPKOTqAkxp7gBknuwjnzxeYxIL
TmK0Zibx1eCykwuvceeuPgKu5uipiROGrdE6EKxWxswt6UcX/M431QNMOdtNnd5E
zw/yuDEkJK4raCehpLhwyB9jeYWZJ8WL44EYUIwcGmrinnclALHfQk0K5hhhgddb
tMO6ZeRbpl6KJzuIqTKnV1Dnwf5KAXZ0NLf1x6HCmpijRPWKAIKdz1GifUyyVAWU
7f1Yb7ZQFjRirfK6liMglXCKxYXfpxAMujoQ0GUviNDYki7HqgtGTQQVh8sBxDe6
2Lq5HBqQeSidjfXOEr8BBDiH7fdoIbKd+Mh0tnNb//VyVV4W/l4Q2X9znu5J/XmZ
ZDqxiSQPjPmeI5joLtEAdi04EPo+axi6jH0ySMVm+XX5lRspO/xU9CNFcKOddBCZ
FneLD+fegfv4I4xDK6o2pcpBUucluUGCX8MXXFvac0oA2Nb9qyH8cdvCa4fMLbtq
mT0fJPQ5kUu3ujtlv9Uhy0A1zzN+xjyrDJVTaoZizBWW52inrysE4Vg4IhDuVsv2
1J2WKx8MCifjw790HX/9Lwopcw5Bz/FsvD5c25bgx78hbAdDNiXM2tOm6jpwdupr
Ei5JO/NCmoe7Af/Qg/8jm1wyVMMd8XyLPHAX7VqmIxmmYfNv9J4vkKRCar89sLq5
5IVvGWkR5UPl97T1B6ZidaEONH0g0BcW1rpD/OSYQUBJjlU2xmoeoJNxHgZOE0se
qbPyjvXkq9yLZ29ZKjZ6Dqr4iXT8MWpcQvpbwqKUOV1t73QZQFMoL+1Nsp2JE4iS
nbZRi0KMXoMO4Uwcp/WAwbBtNvqXHQ5lcpssyO3dJQsqX0SRs5ZtisM6MXZ7GWnQ
0GMwS5pdK8WJb6na6jjVEabQA4d7kZwwNNvCCELoYxiqRan/pugqeIberycYbRzf
iukRbf02IuXiqS+WPMw5qeRhQWIgwifd0ff+1hvU+9849ojp/IJlYOk6Rdq00UV4
PgJvaCuVYQ85fxlDviV4SlyVVRxxQcMy/gJR3rROOHRs5+emY2ImjDi9hu2Fv5Hl
JV/vxMXOnNx1yahqptWY5NbbJDgN42AqO0HvHp3exHF7gv9lHHrzdU3Iq9ZLyXzj
Yb/7cw2oZYGzBSxdYiTAXMeiaovn5x70DY3LFA2zm0nfTeNzh4/wmlQev1mkq/RX
ZY+/LUhxEGqf+cKxLbDP0h64CAtbYEXRGeoQYMXYjVTjTB74djbjoWRL91SYUKIw
cG8DkQnR7SrsV0frQhsJ2vHfQ0exnvm6BJxlFEari9TOYPZ+yZfUhR2qW5bpOTNd
S6+XZURFTT2ZMMjV6LMW3gGbCbM1PsdqmeLsVqf667V5tJTVKxxmI+WtxKpjlues
KayaUK1Bca6ToV2WZmVxVRNyiMc2etHkl+9m+8gENprghjvk23VjgdUbTxkUoaxG
Tpa7XSU5z3Glog+TMTfqQfOfNKGdg70jhoFzfeEaVxEqwXEwtNp9P9RAoypOiqF2
RRSo4Z3A3R0igZ2zFuMBJupivFgmDlcx31FRCBW5Skc8sg+t4f17SYVhq4VX2uoa
Fps7dIyNZBDBL3W6aEr8Zr1J/A2oRpeMmYx1sLRjTJZ6ZDNTcoUAGJAuRK63Iptl
JdVxsn/dfRff9yC7rcm4z1hhU/scH5V5l2xNgbjLU10XAcWC4zP8k8QiKiGCZboD
pnJ8grDULtsCBBRqMJ7nLauoF+RsFzB08q6MGOgqB4uSqxOLx7D2625PhaQnHJ4t
jrgoErfe6Nh0uQave+XhlZ82K/J4Mi7AxT9BULEeWLpetOrYSuIkebbEFCTKGhaT
uiK0nDygncAzzvbfh5kQF5pB5T4Tfme1upPGujUtplBkLOnbvUACaeYCnIsMK15j
BeBHdb9MHtVZcZpdo5alcAB0DKx61OPCENdEuYNrmcUZ37WiOl+zOatjVEA9MXSF
xccuVg4CEqaq8QFOixIfqDlOqLo9Y033JIxb1ehGatNU/XZB/YNb6xMfj0d11wGJ
3wsUAby/rPZ4tPUpfG6rWWlaz+yg2aZpJtpygtJ5RmE1rnILmy3YbPSIPdj+4EMx
TPsm17/4IzIpk6KMjwREgBoTdfYmr4V9zD7Hsq4Qz4CXQFHPLR1lnF14sTr5RIlF
vIEI2fIaTQEgQa0kRdNa+Zcy9JFkUq5ltpLEZNFTfPm6wGrvUufmS6SpMBf6nu5v
NM47Ot3w3ZweIlkxKXUMv4qbb3zl9qDhFe7lZ7oTlTjU1cJtZSRHlqrWja0iv0tl
W53w88/Pd8g+jQZh1qPl8XrMyRtYxp2Yj5QtMCCKrmCLBbTQr2hpCUBBPHwC4NAd
TOoetJymDWgqFFuRAaY97//t7j3zv35ghzatXCMe8FQHqS40L7u9VfNwR2bxLri/
xCVGAq0NLqHoZQl4Mkk4EYWJgSkQJbefK+ZEk93Zww3umRuKxODPDl74Ytu0W/Hd
dNQ5oq8xUE/KarxVkXwv4zoYgJ74SgEsxI/0Z4VEKv2IycHUEWLYENMK1MHcEIKA
OUtxhHapbsa3Y49AUYFWbkhPrvbR5Lvj7Prw+AWpsRl4rulr+1xkTLwCNfHfRmr3
e9972BRLvspuBDZcQRhPZjMpSs1ejWoeKTY67ZhbLzpUHLypWt5gCVXqnA46Yt8Z
W3lRApr81JqmAE1yh01OpYjgqqyedD4W7ihvBeRvuC+MJ6sd6WxAH4TZmnWlwo4E
j1CHUG/Sg3twNqufZgT5UxTvK22tipwt1gkJCm4xtU4EYLDh05LB4A5px2O9+M9f
455dz+5y6Tb/iphYXp9z64YorMh5h/OnxikYC+XbcqJ4+eEiry46RdD4U7FQfot3
FzQP9pS+7Z+LyLI6hihIiHqZoBDP2Xhrp45ut+uKvc4rRUyA/E05P8QLT1Kp4Gif
ctZslS+jriTMqrw1R86+PJbwVSwJVxx9f35seNAA5XGXj3H/zNg/r4O8VNgxbxer
SXrpyqRTfkuzxoROZZTPaQgBfBhUOgZ0vMIYzvnW2ZGrTL7RWspxrqbmgI5xFJ8b
ca1UKZJ+kK62jF8aDlsISVymMZ2Z+wJkeplmIcLTIKo3UAT/1sim1+NdP8FLHfSH
5xy26Bw76DClflRY4gyY/J29vrfNv3DdV6HrS8I6F7ettH8trPe8Soii9p/XWrjF
Olf1Jxz0rL2jyX3+5m8MKswKquvZR4U/sFvpmprkjgC7GFXtXqn3iylzfq1E/cc7
KSrssLakOGM6EqHYTPlq/jADtMh4N7beH7myE20/X9DhO3oR9aA2H71eKA6gUeZY
uBGS1KZOd9fyIi31fHoURYiVRWBaIQFEEqPKu/KRP+wzGinOjUIYM1qFsrafH0I3
UmvrAY8S44bJRU8QQZ29JBX47EKK22Q5lx/64Ai6OhrYq++kJN/qGcEwbCEtDGXC
N5E8oLSCPQWT64kjsd8q4OfcsRreTWGNt66SFkGTRNHgCBODdrohihJTFolJ2qj5
9LKMAvRaZ+VLpvNfn2GLmLjOVyZRdSyM7LYYZtqScI1PAQ6KvIHahZCFm2Az4N9P
NliLZWlDiftgtWqbvfJUX5iJjvG9HS6X0W/4uR7nsbzzOtGiQzKb3iHxRgZraKhN
GkR/OxaeHLUd8Y0LXitT4PFj37KPElBoUSa7ueqkNuFjubwqG2C2wnVlHLMQPhBY
YVMzsjdr0k/XTYiMgtniiV5pPtvM4y0nKb0Hp2Fu3nxCVoX3SgbrfvDDPjT3qDA+
AYoApfcP0wDrvBLvQmzOozwMsVVFRXqQ96qhiyvpT7eu4UWOUjnchfP0LtYRqcMo
5dwTFpfh+3wlkVIzX9jMJpmdIVYITAde7dshplQM4lCE9PirDM2W5UmyM0VYZs9d
7afuNpWUIdOxKj7OjmCpt8wzrymK+IVr6UE0ldCOcdtyQVDpiqkmQC4vZOCjTAN8
jGFcKGqQE09XbvIsu0TlljdevrbUt/S6t9LDpVexpyDMM1CzSqSmCqxQF+l/djcb
7Fn0yrNhn9j89qvzj0AhKfnntFM5XSXyKzvSuwVdTPEAZbwi9E1c2MWg6eGa14tp
dlcnKJvdplSJkoQrWP8tjzCxX6ruzJIolnUGBHXp0jA9u0pyl56lhcpfUXgpiuyh
aVCD2oNVBPN7PSz2mZjujaIBD+37RHSpMclrjJjHS054ilMip9hcIv6iFbLmvgty
iDm/SKx4i7UMKx+/R1D3RaCnfHghyKUMr6aXXOxm0UeykQ9aiQVW4J0IohTl2NSK
/IjTrAiaE42HE4CvzKy5pq1DP3Q8qpkHCh1Py+mfsanNQh0XyA3CeUnQlT8/2BcG
UPySnh4cp8wn0bz1/Va8VqTchG5NjCH84tFsrmjZ6gazwYc7VFBxu4KadSakqzXS
LgTg5UwFinfuaHz/bDXAxmgz29KOqBi5gB4n2ccrtRZiNRzZ0/CbG0kOrHDcnCg0
7HLEGN1+g0GyqnACwX6g9M08Tu4a0aPUw5lpmb8Odvzj8RV6X0vIGerEs9qeyb/V
fHxB08ZOOA9aNym5eypIHJxB4Tnv8klWo3ONaK4uknsYoaIfqpwDHwNyF4WxeenI
DJI6eXpPy28yZ5yofCIw01rhuBoNTiNRDZX2wM42D76GXJ1dOqlMd/ahUo1ORkLa
ElEzYd0zZ9ew3DF61/L68rgctW3ShvOK3DmNGY32xar97wgUZ2ES/namuL6iz19O
OgDRoiaBLEg7S1cbKOf4NH9fX2WXO4/Rz3+/oOrfN231uFRxpSHKEMNluPMSeQbz
0JueV8uKF8vt99kj+Lq780WHDxb5r9Y8y24bggwtjFq/eWMR1IDiLcy4jU2BF1RL
hkphLDIuB1EmEBs8b7ZA2f77Txain4gSb0dEILcJdWvM60nqdzFXvMS5ae1iy8JF
ah8TKjVNzx3LlpU1IAAqgZynWydQRtp5TTMgl9YUiPEz87XpEf2WI9JHyGDgQEds
JvvDb0Bff2UPNCUHKV/Wzbxr9rm+HsOVTvPnYOGql8TYinDRtiDu6LdAfLKK7nXu
qoZh9k1CvB5XomsnOkC5X5iuY1s7t0igU8fQp9gYBtAM0CTg+TuHx0ZUKbznZGAW
lSCzUbjLXQvozNpqGd+g6vAoobHGxsDXrWVmeMzd5fQ0CKX8CrR9K/YXRi3rBboA
fQnlFFQzugBqWscJYDsyCxiRhm5KeY9Lv03zCDSP92Nih7yDZzgHZ92VCXTqS4pW
Nh4Fzo5D4Seh9hMaC78gQfbpy4T60FSs8NRq/cEfJyFluIRm/ceQtMX2FQQCl+12
swxB35OdYBtS0Z5tPiqNBRLSjZPtDhASIxPj1t9bX3Z4YqeSwdklHrLsydo0mSG4
oq/bcKu1ErpxKjBNaPF9Uddxna4wVYN6byAsQ3mkIjLpbOq/F4ya0pdu+5h7XSmU
XL4rEsSAY4Ne5cMU423FecI1+f3wBZGkFJyE44/pW7Iu9MxG21kH0zOm38sJ7dOg
8Qu20MexbH6ZHf9sNcRatBxFaGzQPv8xNIBkDg6eg1nZCOskq60TM+X+m/JAZmef
KGLMCY4EiM5McrlZLHMdN7Yo4siDs64pRxEuY6bV7yBDG4OD/S8kiUsWxX0Ti3/7
PBOU+pA4DavnD0KeecejS0JGxaEb1yBvBuE9ux3W+ZCeeGawdeVRxSbhwHWxg0KP
W8bOJ4vnBrb8lTDW8SYBdlAtlMPhDZrz+ezfXS2Au56/EkD6XjmxfBmu+9YSF2r9
HpdhN/0MWmFSTXqtdkx45AWLT4VR8gleowSZ/ffF6A+7YWnlALqDRIeMMWhieAij
WzxYR0geQkaP2atwBikhUaRN8bljwErKKOgDD0LnlSpGJruzCAdNcwihtR5PpOBH
q/3iKEzHhUozoHTK/lDMlcqwNgHyJx1rvOpaa8noXBWU+u7AVBFrCFawpOzRk735
C6uap1zj0Ic5nls502IApGNv9Lzl0v+oXMXFSHbHIS4j3KAAs1JEGSkvZCiKap7H
YkHZ8FHFVEaw5EWskpf/6aXp2elpBdfmE9q6QU9a0AhS53qpkmOJcHHJweL83vJk
2laNCjnnvqaeyBX+KuYTfC+MSsNNxnW8oDzIxSsoffljYbEjKVmeUsqA+b8TZFHh
ExcZdMP3MbQacL28yoamnFaWxgSRN3N0a8wY2KVm1Sa6axknVYfEsjc2IXEHMfnE
IvPI9Zj5dd1uqCTijJatMQW07i3YVi4FwjqqdFCVfyRu47lBo/lD3uD2oDcNIJE4
8fgOAtVY7Him06A8WGYtGFQFEoUCloWvI4lA4qvWrQnvG5LERNxLuHk5h8Qu7djA
3KODucW1KBhKEM7a7gZEobrFtOPUZ/CNOARs3bQgg7xPjO8M9IR9GhFvE3V8ZT45
uHhDGxojEBeev283ajlfLd+jB8R/jmsN1LiF1O5PZX311mBWudFhTWOd24XWUjO3
pTgvRtzmBtYlc3lhA3q68y4ui41xJNX3KB6xfE+ASFjpBs7BXYFAJNHR9FIl66NM
qTfzQSJAI41/v1UFD+4BrXvAtH3rC1QffXJ9fYFMJZB/+szLmg+jA2YEFbEo2Qxy
NvyoPxerBEppSqk+lqzxY4wfl0X7YvDRUFAy2lMdn5jnQORViHzTD9neBGBxNOMG
mTgKkTsfx64LlvMpSsEWcqU6IKBMaXSUXKiU6byTs8EKpmaVnueQHdLlvyef3SOW
pbW4ZHMPzzAgsQsN2+LNLOshp4HGF+wU6kTh0+8UtfCY41b7Vrx1zbfRmRN14KDh
cVZK8GH3MX4IIu0H1OvvgX3O0V9U43kGbIxG503rWzuzKYv6UGdqVdqkUqCYN8WG
AXkhIeTUZ9Xa3AO4DAIqo5fthEDZtLIp1NldFZfaE6sENJgqatmuIA6Ntj+HAIyN
pMS6cuY1RESibpOFBiGOW0dN9NIJPDiTSxAJVJqI0VVEJ92bEx8V6Es3fmwXleeh
EYxLaIPiLx00g6VMok5AGPBM6UfZ9f6rQqCfaJ9Tm2SdcPuk9vZX8zzeGZ9r4KXe
TTN8uaosL4JKHpwjXqdlg7PQoIiSDTtxDGoveE+PtaEWchdFMTZ1L5Grr5d6pAKX
rVTjoqjpP3Y6FFfk8FtjUzOzrdTdLoxi6nKhp0zWlkJ0dJljY6cHekckzXSwDioo
0TWqWWZp7qH6N8wcOGLdAqapfX7yv0XFJQJ2XxNgviJTqyD/RjhmbiHpOL961GBB
EAnAITFOH3slnjxeudZ5/1mqdlFLfIZv+ISluWdDzmmrB+mPrXq8k37ZjtfYF1yQ
HdoS1SF4MgnBU+smB31oKgusqU9bX/Hpn4tfmab5N5u83Q2v0TYE3WrLjib0zCHw
FU1dQ+2gwAACtlZjz7S2g0pBjPnQ9Uyxw/W0rtPqP85aZef6X8VdsU7nJGTEuQjE
GT/guLvCjx1OneAe+Pu6o46xj4rRRu43LjlAqSFqtXWt8LqFxwrIFWNxMr6uJf1a
Q9Jh+emiNzQXoLFbT5nAzyS3xFJYDhYVSpYZ4E1j1XHlqwrPtGMgGdikU+fAP8E1
4T8Bo2T2iInvLK/v/GPDz68fehdEE91Qg/yUvmV4oPMnIpucK+CkEw2Azdox2bE+
c7Rc+IYiEczgr0rH5kJRUQkv2jLi4uKxB75mqUr/Ir5mSdh1xk8a6kmOLUX1umZj
+r3QzChKPz9yUj5b0/QAzhaAYQ3yDdzIKTNbz7/Le50IF81noOmaOsJFtMGuHBQg
AyaBrf0iAISLeNxvZNwa9Is+24G6UaA+72izzeO5vsX6rCUZu4I1rUAIaPl92g7u
+oCRshz4OYiJuY8Cg2jUQ6PgKbMW4XBPB+k0zRXu0NP/4qPcY+XaPs/9djVuQAZ6
s+hPBiB5jCtBagN+D6ICpjbqu82orUH0sczyxcMFyTng4SpgBLJE+Zhk+QDOkG0i
gXskJ0CBJWTtmNJ3F61JCOmaVb9g1ZaybhBOmezG9Ir5a4y1GO1U+n19LuOl5wFB
XR0cVDu8Ln0BjTB9xjle1bkDJi3TEnSffuG2P1iKiG62mEMct7lWQce9bYQjRTDC
Xu2JoiSPpSgf2QF8puyVSYIRXRZ86MN89/F9T6vbVCJEPz5fuwl8M5mNPxBbBqIw
HoBUhvDW4XuW3417+3riR7xAe5H+kKmdvs/ZajEg6s/ajXXnvLfQwRHs/SnHeIG2
QlxhUPJCRCmLBg6URKk3lRPgArAMj+reart91yVxsLJaLs53+621B+eJhi3+pi8i
8zC2GySfJh9p5l2bmn9457dAIf16WvjhdFH7/ywxG/seFgzW+sKmmXbWjItzgUqR
jqcwjcv7YECTg6Na21t5RKVtTrmHcbOazm1B+B3WejwMvmb8UxhnGwX0ybET6E5d
d+YAwWiM4KLG8oPwET1Ll6qpNvsaApP83gyCDD33MCV0He4imFWoMrnKQAD4EYxS
oBxpFZ8tyFffu4TeGSCot8mg6jTVUAGW3Ud4ARj4r8s34yPY0pWE/RC3lhlhbbph
2vnMSQSLZ/ebv+2xl8B9SXuvosfPIZG7ncYr14bqckyNtp7MY1gfL1RneRImPOaK
AEPFsNXNqzaTX0mHnOQPR4yokR2VupuydysZato0N5PDOs+qSlA9NyUzWyu2cJlz
N3CVpKLOUulHLOdKcXs+KHmzxj+ar27Is+KRlgAt67NgdFjeHsYGOkN0qM3BbHIp
S21DgGjeTbiUWbniFrTxVdNJNeKD0RLCrJKr07W+5gYMUzwhSF7atgp0W7bNqrI4
DaMAKXh+h4IYgwHfZLl2CVsWn6XhXbSFps0RnXW8Q16Xwe/oXwbH+Rr1RV8BVhfX
6lK0WVnh8fv4Uw7ZJrx/2YSvnATiEdDOsXmslL4S2XxENdI5tdVGapCUDtuXmJvB
LXgdnZaYjb/mIgHyOZYG9Ql4R8aONRlPjiEDv6EOxUmIqOQ5s+hpTow5/0b74cpa
3K8E4okNZAVScylPyN7DR0Km0oFEWbo5fgn0Pw0pKMv2cU5Sa/vyBnntO7FFbO2d
YL0Lcp72MceXDUsXV56hobYdaXM9ZgCtJnapcBubgJeoAZKTOSsxU2gpEstybmQ+
DePeH4Q+MdN1nqfPa/dMC3iMfFTThnCV/vckT+l2aT/n8Tv0gJZ6s6ry7WgIJDyg
WuFdj/Vgk+wCWhA0B/3enZDoycvI9rYuTvP5uwIqyiIFpUE38SFYQHpzZGA+6AUl
6mOa/MEygX7c+2n/mxGZaEywn+hYG+YdpyJ+aU9SVcTRxDkAQ2wpgzhdXvq6cX+C
Uve79143+hAy2cKVomvHeytHab1EB06ssFgEzBir572lE6/EdbsDebcgE5aZwUqW
i3f4SkObXiWnyfB+OWRE66spJLesXBpmpZLi/x5/uIOUAdd1cBN8F+GVF62VCC8o
DI6Vb1hK89ZA+W2b+w5srzyn75inOaQYX8WXXQjjT1309FyiufGnIaduPlCv5dRS
fcFswIwc5iX4FhPpQuuFIH02m7MgPLv9kb5aoJpTx5hnCBUdME2DskeQy6I2rRZl
fTos9067tuy/FhRgv2Igp0HjvPizwjAeK4qlI3OvorxcppL5eoIxJTiYEXp6rtNh
VV6y+/pCJAc+Bb6MrYWEVRL6q4P3JnKbzLdyfyK9Z1XnA+MnaDDErCpg0Olrz0Wu
bYeNzcNKFnNUTO8oAHpXQStflO/N78iXxrk3RWo6ZVCbSOtJmPU6ZobK4lpSdEFN
BrW1zPZSwCeWJ8isKW4DIln17FSQM24C+JVcro+g/EJtYwzzgosjLORZLCFI+DYc
/Iq0aBTfT2nz8p6uDVx+0MilJ0gSLAXFxjl0KfoHj2xiZUG0AzyPI6KMV5jGy+l7
p5Kdd+JhzTOPQ3BIN+7J6Me17xoEPLMTbZ/PjX6CLMf4/R+o/wrQZQgGG659VVod
8tJVeOsOKeuoXa6FDvfRaaFEVhJLw550Sn2uSzXhaN53izoQAJuGMhc4xP0a2s7Z
VsrkBB1L39JMlwuDKdymvGAWToqG/E/wbvUQgXdJTJX/93cL42LFHVMRmVLt8uaG
TUnizLIaTpofvsWWzRhqWnpahboCFlfSTKq9XO7nbc58v56tM0qbj0EsY9rAUe3O
kqwlWfZbiw04PFAQhdt8fkSqT7wo2BPz8ipzYRr+fH0WQJJWIN+Z3xjyUb0RJRqH
Yq7+JXQJwP2WyeGa/VcYMVT49Ycq1gqOMEfVlcjoqhjNOrirSy/X1DY0Z8Ngxr+n
/sFUiYSXAgADaR/eQrmVMFu2oTZWwnKmbpi6LMzoWnlcqFVJw/WXNkCt4EGomnaE
wKxl5YLg6BeeD8Cde0VA4h41VbPgbSjIR0UGgIhjnEdDxW+wvKqinT6YNo6/CXud
n9oS/Hfvv9QDGUcEqi8HPBK5sdvX/SNoL/xsOviSMU0SCUwRtiQ0MvUXAtXJUT7+
sleddm74bvkZkmC6ivDBThoIn5gp3P9T7SoX5ZwgW3vCv8LdA/d9yPBs3zFA67Hy
0VHE27Hp9M3EOA0u3fHoG+L+V38Q9bIoduJoHN8D8iEWKgb6/8Y9gaChCP2yq2Y7
bCVCaZxr0+GUVHCutB/tf3iNhzNv3FfBCT06bOaXKmS7ALj6lqEs3RGVPrSophPt
gIEX0AV2e9n7BvbW4qzEJAfH66yB3RY4is4EjZF9WCqBkstvKR4Elq0LAVe+Sp4X
vI+etfoVsrJ8A3t/WfnUOUjG1dnzemls0gXqxu4I4ZrVXICswdD6k3iya1DdyETq
5pMZVdblTzeqDY4fP0P1ByCOrrt1j1vhdKRRDqnibPRkUIWpxIfXQ8u5eXVVYqWA
e2W4lL1o6Wou9LUnpa+fvoKxlqt82J4XmCm90b2KXUIb2Sh6IElXWFfLuYNQdLvX
KiK20HXe4Mv+/tnpTcJgs23ABVT5pVJJhdb6WARZ/Ey7bUvYZZ8BglywiLaQR3x6
Ty4GxmrLTdHP3bS56vIIfYc5aO/98i/OIVJ3/XGGvl9fH+l1JHl8UaM3rTF9GZB1
OyA4+zwdIzTdiggJ3ZNVXtXNLuCuIDO9+7bEeRFOxSrkp8/Xnu2Uk1q3BoG7D6W7
Ntil1RQ4Or6xU79TNpsU7wUS4GpyzfUznDEzxETDkzxXzUJBo2PdeYlS9/E9Z5Sq
/uajrsEZTmKfO2hCUjhJ1pCGeio2nPjM7OocZm6+Wag3k7V9JUP7872sWeVGe3AN
jv5gzPT5vqN8fBARMx8hMAFaFBfz7O7Xo61mUNQqfflZoTM0MaKTIJCCaGirc42I
VJAOeUyVeZagh8RSsi5mB5iEzirGa75bAywsJU352A7clrO4suHQ2nsKRqZZCqrp
gtb8oWUdNssMYKyxwMSdlcnqC3LZPuMxFoC0c2DDcTJtdXZFF+26G5WaAOQ2Bdc2
GALoZ14zoNMmJiHS5rVSxPsOq9cdZ5eYrHYMX4HaqUsfiw6k4smDTCnScLXr9PeV
W9wbdEfxHrQiiEK6m527ochqG0qgBKjfPaCscWrbHvcH/MSsT20WWOPaBrYlp0sN
m9gOfKg6SjbhJeeJ73A/a+6IbwsCbQEw28w4Ye5BBeVyCdtmnTmelT/3p5o6sqsN
yB2t6V+DC4cKdmxac4RabXXccpFup0SXQDLxjSqs7JcL6K3CsZIzfQqcwF94oTdu
1dRUeGBXpuvv2QAr4ndjEU+bXMy+RNVMT5DSYbPc1KWaD78mZAKScn7lZiiWwaxy
2IZMei7rIGQZ3FTPdUMpkvR7YnWM2PvgBXcDT7NzcUBmMhe6E72uRGdaQLuwTBsg
WTvF5h+OMl/+6f2b+uL2YPWBlgWRzBZFMftXCniTmNiggFd8hOTFgwRALR1rQ9Ds
R83CxFkIigVGx+bvtZFzWM7zaCkw+lnH+1y5X+NXNehjmLsvHJeqg02xJnBJzfZs
BnkEJvxOaXyXuXUssH3P3M7CUnYYsTGAXjOo9jl8XLqEIdrx6YUbvNwP781SG1Lv
aBJWbjSr27s7WTcAXFuJ9E4cRDzX0TysyohsGFSGIaCrOYralfOE1dn7DiQyruSe
iH/aHOgZNCOQOZkKn+3vwRM1cEhCkVTBO6KxdrDj9F4ObP6zGLLHTEtP7sgr9Db3
0BXxXuzpfEvIW5A90hJSu2zNa4iOwML5iRIySw5K1L6LyR9TME+DZLLSdKDPeGdh
cmthaO1jrSHokgyDBy9mfCpAIBSTTBQANaPSbovQGLdJ5V6yZ4bCiJIt/evEmlPK
2bZcjTOsHIdfsTOj6TcvrUhsk5GPIef7y1G4p+kFfGzVU/k1BwexahB+uOlE4G/q
iWwAKttrSVoehaVyyBoyZQp/D7AYGa0jwYYsKZVxv2Pacc/Zlf/yHDc8Ge3BRMxv
joZjJkD/Fcj18kdjMMcvDTmw4Is+T5iVfGg1xZgG9FFTRTma568+h2JLosf8h620
KzutHnb3UKgm0nvnpm9rhZB6ksylskSrroWaQ4QFRAV5tVlM/OLjWJ4y7gjnaJXs
UTYss2PgEpjn9588Sduw6ZKcmTD3IlqP4NVigC55vcCy1XIQIdRDC9SSbknb01ec
ZypU6USmtJKhnU5nDl3rhUCImExAX21ZPKRkoqEefmhOyr23ZD1WrztYE/zbAO9l
MdtU8wdXuAV9ENvHQ7RoalNYNQ8gT/XQwmJwGi/VJpSFbtsb8+DGCcAx+h/OBspK
iIGnFj4afVaJP3rxNtWh0ljLWvCYRHx3BJGZcgxyXxGeU9t5a5A+pZwXex01ktjQ
Lp7zURlTald9oOWZeWkVevoHwLiptZscjcoZ7KFtLwH1Zi4PmZ+QjEaaSfBM1wjL
u9PrIBL/yyBRrXdzqakFuKAbg52ZG/tdI0b1EhySfGSMQm9RbWv6M0uhwRhQGK4D
DmqmS68wStdh8fU1BnlFSs3GPAEYMOHhNE6fZRB+UnO0dpEtEY764O0lRo90Gpli
79h7lwJ2jLSD/Ujq9/ULpC/1QycAUj2T05ITFXtFDFHbSEyWDtuzZEQAz+aeMlAJ
htIlCM5hDwUWRvN/NiZXZETHhztGINEwfli/AMLdmqLfsB1A+xo09a3F7vB7wG7/
dgaQ9z3DmAOeYIBzwW8WqjoNY2t6Df5agfJOghqFs42YhVlXNGAWbF0RhTH7ee30
8r1DAyIOhNZeooPYiZWV4calJcsl8anR5uR2oH5YKcdrMN2js5HLNIsecDndMLzi
hZySLHN+fW6SNmsewoV1YzvPE5TWRpvfJ6Rgw0BmCnXOVSrS4Oyap8ULfkoFZr5k
IvbnRpcsGA+WYzwE7fiOWNHGzx1iYqe28DUHT/CmVb1I2yoqSv6sSxk0A1jBdE/y
1h1regbYfSmwzapdsEsSNc9Kr8b4bjbGaKS27NUbVnF8/d7QwvaauJwl4PK36g5v
KmCdPe4e2FW2uNh/gMBRE4IKimiL8fMT30JwNswy0HqtgL9ccmmM0QiuDY+nKLn5
+ytdqoOfpApAVyKEaCWEyGptTe5OqzoJk2dfbqGn5FSFJmD5FdyfHtTkTjhsUZ4P
Z9cURW2hu7Kl02R9twaEQjxlX4bY36bf52DPn6pEXZ7FzcYFxmCK7shIMcFnL4mh
EXW1Thbeh/LbaNiahBDDmkwyoS2yUvWwJYZ0lblOXnn7YXsyTjr7XcVJU3X4IVEj
W4HCIPBObvmxWrgbkGdbb77h3RljpDbLUBLqafP9TwTtw3V/CKkjHjCBVZAd0CIO
s3LQrU8al5/2bm0K6BwTihQ7RFOULvkagwDtHfRArbEQQcgrgnYkH8M9P+54IzMQ
NzDCRsjoxFk+VfB/UIZPRKuaXL7Lr3MQbihrC1QbQEBLVNl8UrpGez50nF2ufD0T
Q9QOGBHuHqRtqd4TmuUJcIkOBBOHQwW4Dobi6LOweLgORJkGQ/WDhZDJ90KxKptI
7+suHjYhVPDqmbUXwOP5O94LvTUPOt9vjixsd0J21NhocncXNfPta7DCyyxsNLZr
LW0/oH5SU7OLsp9sGZJ2UrNIE1wgCufqq3RqvH5jF2KaZQ4kgxNVXjfsZbO0uRfw
1iNsxFpQFOriXC5rEKl6a85v8oKiN3pT2HZzD3HIZrSbUDwIWTzPvzzDqGfcd0mz
rwm9qr6pyBvni55Mj2cbHwgfWw8yXaNnFBVIMBY7wz+e17wGrZDRVSmUz+5wPcRo
YwgelofGcqO9tgT8yIsYDIRRJMU2u60HrURYlLRkCZuVqoakqG16/DVRcMY+9k40
hXf2msEilmnkkXECETBx5FrdoMndepEl01S6iNtTvUXfwdn5lCcHhKVSN+hpgjDK
YsWNb+zUqwQSe+bHp7/oTQrgHzms/Lcp3AJ9DZqcTtlsz2LxkQXZruNfFsUFCoN3
XZA13IGRuHweYjRhc3Pzo0HBP9a0ejdhxO516LwwwqG40OCcq9nbxRQ9dE6vN7Y1
6gS1n73/++QN/clxdmMxrh9a3zFB3OqvUlbbvQrVMmrjDYklLQ1Y2TENC35HU1nE
KXeKZTTSly6gexXqMf7aY36BRMqZcB/JqZz0zH4WGtQ7OmaYsd5NN5tJFV1yvATy
d9VzlQFy52ve4JgpHKbgSCo5qR6eJRKdbN1SrhI34v5enFucD3Tz8ja9/i/Slydj
HqLL2XvhIddKq4wkbSN3CDQUZF/ePM9ZhCFoZyjU0vKR1OOLLHswtCzUZvFeI3Xx
13V9MKN5FIMoacvjAHOebQkOrMJHV+Hhqiza/Nnmjf3tucf5ISvgQwPO1369R1/g
u/l92pOPsojvlq5VEsqmZSVgBuo8y2Xzawt1Qw3ETiQXro/zA2jsko+d0ZTziOlZ
wTV7VpBEyXZNtcZHUjYliuVlDvcPWFXyYyfyZ1Lk5b0vlK2TyenATQ6jX0Ibngls
A0+NXtnI4IIeSQH1JqUIS/kYXcCF7hwYEGmpHg5NN7njlMB5S/8rqR7qn0lD8nq+
CnSdbwaVdOIYqrupaMXaFi1xM2Akx1Pt5F0DdUm8rcFrPnY6TGbfa7DSOOdBPBQB
XoVSQWrfJsEtbbmnRuQkrKF0eEi9tGf9em07Ij88RFpkv1VDajD/jOVWLA3VBP70
PjoHNZPUj0RSR9zekpzK3R7FDzzHzmYsP544+tF2D98c16C0aTSesPD2bXntYVaG
SsIlR8ACxCvzDh9yxHlE/CdFwK3OYULE3Pj9QoDVJ8mpU7OIBRJ9G/KzRvtaLUzi
ebOIwtvhaFSyhqqBJNAqMIfTYG99RzAB8U143eFRCwnytfaqN+iUvSnF4tRR8fAL
LDXlyeMb7WGTXAWq5U1uH8btLrCK0MvwPWiT4wRnY6eT8lI9gGGmCqHQyDbDfXF3
QpI5oLazdFPre2Xt3Pr+iyNBNFVPcK0MNzRmxQNN8c42TRO4x6QHvprRPvgnpKwg
WO0iQdYbdOmJbzCK0yqVsPV9y3CL0zHqRHAn84o+KapMqqNCCIEqm4HAa0zfuWvW
dLjkhXQPU98CUVPgJDT+8h0kovbi+bWu2XZZPklURKm5BkPrTa3ut9f+EYHcCY+i
lH9LMW7WKsWEnygJszHVUzKNYLekbbMjTnjdFPqSlXvR23W/eI4gn/98TpH2V0eg
BzMRaBFEvxaPq3ZxjQHnR++i7N3Kk22wX1rATdKxYlzGM8rpP4QO0x2YvISNtoGk
YYhPPinqhWAR4mHGoI5VgDUcUBheNQLlABOrqvX1WbptB2nYzZi/gUpmrQJXNWu2
XG755jPZhQCJrjf6mgWz2qYyfycKWmtIIaGL3qiWuj/Cm9rUF3IkctOJxAqQQ8Fy
IJddHcypSmbTAwAVFfLudYESgTeoFyemEsVrh990SsZ3E3mWvoC4C9iQZaNIy4JR
X7nuhaTbv29tIDKQVxffxcBDuemVu9JlmLKuktU93tlxDwxqWt2NygTMtdX6uE5/
17l/a1pK+8KRlCfVaH1lDPsOnxL63O57/dir/Ula22ajt8f27bbahV1Yo95oVYkm
nQF/TbNNrStc4waALfJHBYA6StEVMrZJDyJIifGakN2Hh+s+yRm+yst0Dh7kcYlD
dM3kE13sdYqmwnGEEKA8TfO7PlnYi0s4A2m7fx8AxUnsIj9vhkQBOTO3AzAD7qI1
MzdkpcTyan3XAvyUGHq1cJyXr0kNOJYu8gtjhDwx6xhT6wZQqQxnA4lY2XCLoJPx
IOk+RM6z7Zh1ZGMQl1Bn20z/+Bo2DgXBYbCdgHOFj84jZi8dytzWX6qpml88xjru
nGtSpR6XOdlk76BJAl7bALprjOpMwodFRz1+0bRZ6KbbJC/NWJmNUkWxelaaFIaz
DsIxOoY3d2Z2Mb/YabjncfG8fbsM1cvomy95BN36SfxEto0xv20AMRKiXG9cg0EC
UXSKkiPrsriopqGQ/h1J4+YAn+MorLKwpLSo7vp6nEJOiW/535Tt2Em+ItyFKN0G
Ty8YOyXULlyCzevAjLIxo8HEY/XbvTBRWG8WYCGBsmEOL9h7TrwwL55An9ynAlA/
5/1QzW44lPquN1yVSwPmPxFWuY+O8NCEZozjfuHisB/SVgFnr3m8a7klvegPUx1/
iEimgczvjoLiKKjed0xWTMvVB+javZG15+s2br3sIycxj8WBmC7q4KNetJYBVFiO
FlG8SP+jsCG9lCXlit2FGk0FaTq7WLmP8HY3xP5XxwFwPrX2WvCgKLRVY/xQxhS+
LMh6qvaSJRvmp68GohfNxzltMHvSKPqdRMuDfVZfNC0chNNyLVE+BoqgQIuGz24v
VZLBRZeVhtdk9DzDfCpjdzTE9eiFz6oMceog51+J9YFpWwasTaGQztY8Zxh9bxvq
HWG+TH9+foFXPYmOvVRsThJr1pfVtRRxnamSyzUdyWPzFykqVLw1+k7Pd6eksDaw
hz+y1H4qgvg3YLuRkHAa0izhYoiXXAY393ow+Us3DcRvyyMBDTwxMb47Uyxv6n/k
3iLD2O55OB8HQBqz3UWkE5qpr8zSmFirtBg2Z7it9nAokljc19okQyHTbhbDP0D5
AcKXB3duWnklpoPzucnEAkh6tuKDvPCQSVGZTM65k2XmsmCUkJzvj+Fy+U1lmD97
wkaM/eqZPbmhCO22fJOSwBHXlKFQP9jfif+9/kvTgtjBkWye5HVZPW1gzcFD7nUO
zFIAAVziFgBmA/2V00KMyB2TDYhrer7EL1pTFECoPefnCLdHyc65vQPlZsKfMwDn
G0uFekhHI0KYDcM6tbUDnOncI0U/GdsoyIPYFpf75tdt1V0UwH+/F9uWobw7DDES
eAZFRgn7fygHXKNrviwSSK+l26NcUut6/5BX6cC1N72cOe6hXKrXgS5yS4eqikEX
`pragma protect end_protected
