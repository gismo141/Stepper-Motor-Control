// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
NXgZUUPHRJi+7NphD7kn/TsADXNpXzGtRJj8ARvzKTfATzv22Yfs54vgBIVOzMiuSVz4BA7v3r5z
zTA1Rw9e+JeUVUHdcCydxZ+j+xsxaYOzhfr/VntQ1Wer7NmVLE3oCr4VjzX61sWRkCwWST6HvTi1
lmChAwT2q/n4/DxTXsV+MFZ8ozrVFM8jQfBuBIqdmpRfHqy37MK/xkUf05hOtrcD9htKBLMZgzq4
Y2TMyJ61g0bEuswAxzA2yNR1RSIgrCGvzYhNXGYOTccAe8l+mg/K7yqo3aiTtkH0GarzT02Scm/a
FVYMkrMnbXZvt/Jf9GpUBgyAyKxOp9mf8f9jXw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
UMYuOnszWAH15RCNiIkPtjWqQ/MtYToJ6sWbHYIapHFGzvJVkjesYPVT6FXdNVV9VQKJ+sNWKH6/
H+WxDGI3BU/vt5hFo1zqPqNsLgy3VX/eG0GUZj0CRop/olqiy/mcBWOy0XruwVnXp94noNljUGJj
7Ku+M+yv6QQhv3vZz5XsDKyN3JUadzRv3EwCwRAiy4cFhz8bbYIXqiKILA3hq4L0u6Vi00dwQxo4
5Wh8YSVJIjFFoeIL0yidZLBsePlBhUsDrXJ4IogaWP6uQHRvkd0RfMv43BsQlVinsseU9b6PagMr
UnOw2HQyMbHKnpjzIxWSovGje8WFCTWJYfqUUOtQaNf9j7uPTvLhLhanSBe2A2zk5W2G334de5fc
NZ0lOK1RMXm6QXSQleywy6E//TO0NdTJTI2hxVoNo6+6bqBL/guIbWp3ntAO4vtHZibVPjHuyQd/
9l7DV1pidI0yNjVEjMKzDyT5UTHjzYbL9Yp5QGbDEEIhgImyEHRXo7Vge5oBiI9BTLocMrjLBcgp
NDhD3ruoE/TyHdc8kl5ceHK6SUfR3briUNOR2m5MmCQQ+/sszldu0fnuWXXntSKBjwRDC5jRYx0P
YI/gcgdUklgpH3xyy4znIDqJvx/zxFhLok88lBiAmZzFw20XCBMMNSAIcjaVeQywYtK5vPO0BRNI
Vnzi1+hww5IyqrvM1ZJ25U3+cv5JHbV+yatcLjNjzf3JMcwtEcodCMCHjwlQAgw4G2T4t1S55+cA
0nnC9GSUwJfo2DdXU1CqyVQQid8FcreSoJmTiXk3gnVJEwVt2ai6kCj06o3M6WucBHDRzPZ/c8Q3
qXF43ceZVC+FeIBaH9gXhMAXtoHyiZJ/iJ1RtLNY8Ksv0u9R220oMNdfDgZErdQ4lpdMht/pS/9x
fH+twsmQSjD0G8tvjdlNGdssMsZYSNdZNW48nC48mq2L+LkmjymGeHEkY6F3IQUyFFzFhxkUJaJe
sIn22pplhjYW1yOIdHnVKApXOx0FD9Os3b3HavA0SvTk1JA4gHRG/5atcchkymDt+pqxEY9UhP9s
SGFjQfCiUEsHO37u82WmRnBAR/92v9t3O8rN5yV/oO1Fxpy76VvFj8bHJFadeYSa62j9YjMKHI4w
WmcUqMMUiXIY86OlgtlAQbaB+h1ikSKTDVIQx8WHsJOpT4klLBuI/bJ6AbJvcxhug6kEsxfXIQW1
l3PGdXbSuEkcP/TxdPD1foOWuDR5ovs0iEufh2KkTHBJhCEYwKmVyeJXSfNZ6lBckNZQbEosvn6Z
vXI41JnJz8K4Fta6KLrXJszSjkvK4DNGfijPGBiJhFOX2Ik8kgK46/gM/KElG9Fc6V9kXaD3I/TU
3x5xjFUQEBxczAcqjzO5naE5F7uBHJDJEnhQiX7SuoA7qwvy7taaVOJNzOfHskW+UaqEFvsGiiWK
XIRFE7iJpDw4RuIsY4DJzR3lyjCnYiY4ylsVJiotvnvr6bBC+k3qu+IQt+M5OlFj2mRPtjXYqFtA
TDmb0fTRDOi2NMzzNEfEbQN7RxtnLbZ10zJrdV2zCDKeuuht6DIcB8y7ZWmURRFL5T0CbA0MysQi
SgskhIoDSGhvKFawjfLkriSKdP5sDhwMVy0cLtcMZOFegnKNrxhhZZUuEdwK3KKeQR9GQSzyXSlJ
AljSYBgLdUp7OxXVheOORPH85XYaYbmiDV+NbgWYIVViBhVLIjVcvzZau+CfhLDKjhA9wRDxAhCF
pLcOTudzhTTcFQCxUfmaCUuEbi6D/UrSmwv9DJVpSaa08ZGlcgKQJE1z87FGSKMltPbvRzNpgJ8q
TiZmoalz4XeuwZbvgAozjf3m/00QAKXTy6DJ4NVd5MqkFFv3n+Eys/FKx0NKa3t1tc9nb8GRNwB7
yDD/r+wL7WNh5TkkJR4lLiF+yNS4JyK/bWkPPuNKuiUNKsNidhloaSrogMV/MTqX8OPO2LTSnAyk
C3mWSa5NeCklYDQMk5o9v2VLlI9xYoAomNG+8x3bgMg8dv+SzLc9ar+KX1A4f174YkI2JUM0XIre
zSM4PtPnMzXxjCTle+qQIEhQfupEM4aJYswqFJzNdosM5Q3gA9COnnTuP4QoSv6kdcfmkKQZwSKD
MANSViaz0QikuqCgLeOvh+GpJ05CDJXdFfJv8Z/+VaUytsiz0m9aMI+hFPs+WjnNCn4HbcqRwCrS
+t3prBx+0fiwUjH+36bllmONV84cFTt3gOaOTuCyIuzsVya/7GftBrKahh0/VMJEIhzifhuqMgtp
Ihq3hWGMEXh7CagKHiXsPC5fT4B6J85J3/v06XqzbyGaOuJkm482JbJDkKroEQ6SRdZoYY116ibK
PK0zoTRkJeKHLYzjjcKc1yVL/ydcHqF70taigAxt0fUro3j+KkZJITu3iMbgOB7rzRpbtjEC2LGd
AtZrzwLNn9wRxRxJEPb36CQoDPaDwRHBYJXiiKCgr7OcAnMAnC2G72u2gaIWzPPkLoPpnuMnJfSS
sOq7TGfXek6uTHtd5/WT5lrCvhjiqjYLZnBYigOFUTBJvor1kNQZyvwL97cfTGg2EG1SBhnicwBH
WFfF1mQtNvXaG5zkjG8g3Jw/Svv7hIjh0p0/wdEwXtBQ7sbczUiWccmoAu9gCBpuukWChL2DerQ9
tQhr5IGJ68upj9k40YAyhCnF0IJR9jWPhjtiHREAYPV3Dklo+XJG2XfSwyQP0puSFaaa6/YbnOYl
tcVEsBj2VjeZoJdzLYOHXy6D/CpRumJB1K7MBfpPYNWHjdQZ78T7s6TTqPZWKbrQJ9JzhrXHU4Zk
CRiRjjfPjSkGBOCBbNsYTcu2DRHQIjUibJaN3/rE5GplhvigDXwDOKpopI9/hqu93eEgj3HxMibb
ZbtbnFWfmwQkkBn5eB1IEXt5v+3GM5+eH3/PNiubL6JZdKnHMBqPWVrmcuE8dYOoFst3eOgWh82T
PxyXyP8+9ZNoeWLcaeAyAMpST1XS966naSa+1AP4dKCOC4c5rffwQgTPM0RXXW+Ad2rD+ksgVbVv
6BVnAFJlsYHa2k5JtlUI6ZmLYnauWFosG5ZWdFlVaU83GswGVkeOUaA5mqkqX8FpjdkwtxY2RhZ5
CpmxB3AzHwu16BnqkIwWV8s3ytTzUvWLsL28jhBsNxwkhY3O0SKgZ4auiE83kaLa+u/QxUKlRVaQ
M5CX9asaJye5ACsltIn1ycfGMGy9EpB883/KTM9542H2xZDTO8q1JP7Vg/tn/osYbyJ1BA/09aew
KNRqLpvFuvoO2GaMv/JLv6w9DW8GNko/dHUZtBDU+VUizj3ObyrB/XPR/ioaKvq9pudYSL+VE6Sf
aMeJtqfZ5tUaSekZbLcRIhS7woK+E2hwxfYDOUE2o979qn0/LqzP/Meiog7UxkwaG/FO9IpIb1TI
khSDDQWP3XNIfwgV6cbqJjhftMwTX6SnRRAB/wg8v0gML4f18xiDuus4LfymFKUTc7bO7UGcS791
gyhEnyBoEOAjCXNVdnlg+R1wG8Lki1s6t43bAOe2+BmDpjwZs26Da/NQ6Qro4z3nDJaNCAiQPysq
TgJwbVBjCvRpEoMXR0+R4b7x292Klnoe9xWO+XVSJ+zNLOWRMFOTF54ty+bjistzZl+rQ92sr/Xd
k2hEgGM2dXLMUVIFiyrOgIhMgC4Ttlfu/20Wxhj3yc7zRA8V1OCpjyzZ53pWMwCPetXsnQFtLv3m
hutvxs1Z+gFyiL4Xi0Z/8uPZr/dLar5fRVWJ40O+1w7YEB6XFKBZ+ppQy/47NTfoFdIsxoKNhcSH
n4RgAsJPaAoAlzmRxC/fQ2RTC9kc2AlMD2UasvkdXi50X2Xaygxm26h1BuccS/wQ2HQhUQJOnfRI
PHv9PaXvzgtOhhYUECRL52eKTK09/TvHsKEXmElm2nNaFpV19NGPi3LuECSUY66+vMPJiYyTVG4v
XT7eLyirl/wDmvGXzklNt3DdFtK0NJOzENcgrYxccaTIDvC2BE4GJR+96ytBmJ+vOgve5H/miRcJ
jGgXVijB9C6pRw30hDSfmIdXNmn4TWCy5Fdb/IDgHl4DrLigjrz3WUxeQhNZk6bxQlHyKXNb8wOG
SMwRc2bX3z6GyNKwMPeMzwkjB2H0Hpf+7Rwrsqv5iXrjnxKTkHnPKqOej2mbUdxwnd+NDmdHhRRn
KiKrkrtOOO08EFFKykiKvob4CeqA0Gf0IcI6o9MxbxhX4i0Kx11ipB/miE5cgaWq3OkBfH180FvJ
r+9mtPbBRLfUP0E7Kih2rgoif5vF7iqHtwZe7O1gGqQSOMTBb4usDOVYKBcsJ2jZkUGkTW0kbt3E
oTzzMMSFbgKLVmURDM1R/AiEeOVF+yk0k3RVbbbSmVz+sm4zOhbKyG4C5/piJx2/mgtWKGc+o2Da
gysbAt04J2L53fMau7DlTFi4mCXT/pdc4foGG/kayuLteiyuEFlxY2OatN5/6bWZAatJx65gcN9O
cVjSEP7ABbEFfryKNzj3JUHOA7ROkC/aWlxq4AUgobAc4vAxsTVHq9mALnvIicVTBFY8IGwdpwzE
EOPO4reFS4c5Oubg2KVmt4+dAFuYIjUbZZ0DrUu7EefU2i0Pts/8YR0uS8cwbXM8d/DtxEBWVorr
silbh6nKb/lVLu67etqDUfB4ByCK6IvobZkej7t+KnkHjpSlNlCTozY1NqFesCPhb5/dL0NE+XgE
C2nwvpEg5MSnIOxv5DKUPezqbs43Wwdil45f/l4PFOnCq+GlcohPRqz8DEHDBJWFn4B0w9M/kwdm
zWQ+0WLkvVTxdMLkBCbgz6msb3JSDxQpErDd833ULX7MP6bwmt8MIutZhuVCaZT9QU3AeXUBuVqy
HAZ3v3ntdDVL7/TMXmOF0lE9oinjZtwaOPSQ4Z0XARbg6FLdsf9LqT3g6lTsv99A+V2HIw3i0Ohn
5G09mCGQ4+MqQsr8IXwVZY7b/naUGXib4qQBRGqXO/ZZg0O3z1vOokeBwWCklwGvPotf1rYObRJ6
Ac4oHqik8me86qbqa5FqWgKaLpPf8fCZlskMuwfS1o316TPOUiLp2aCqGIPWuLWpwLNuzctl1bv4
RQuTTJ43G2yY85WYE2IOh/vmFJl3ZvDPKf6BvHf1fC/BtDAH5QNDF/+DzxB1cwK5JCP/WnTIEh0k
D3aoG7fEzHtB5sdw8q0FjT9qdbmat0WC8gqOUvJFqdg3JuM+eajx5dcQsh//j0NBG+rYq1Swaoj+
3AaGdPLUutcU0woHZzqaQjfHqhIxIJHo8qLazrqwZZaQVqotMzaL7MH1ekuQsGWHbZj+vzvsMJ+H
9U1+ZGhx4vlTX1BS4PO5BpKdtbG60Dx8QVU7C6tdpLx/A2B0CvYpeFr9pAD4/VZ3gXcE/YyU4/IG
NDwJaYgay8FdgcB4mdJ+9csUx+ShqwKZIPGDuCLkCi2V5rTkfDPwJFJRH2wpmjGF+BcsesGvjwI4
cC4xPzHCJmYX80O1Bo4BfrY41+ierPWqy7CDwM64ribTMhWn+87KlSwQMkFMZiO9ZDgM7x56sp+7
fSfM1Nspu2GYZvXRKt2INWYGd1kbqbhiNBCnD1YcULKLPa0IY+ssV3J0x5JK/JD145onFNMQ5K3D
4l9q080thgyVYBild4pLoiWLaGjSgaRoRmdrnHUEh4Vm5bgcJD/kldpnsQHB6l6zlTjFDBdOHHtK
5M/H/+nIp2aEYpNQGmpJ7h33AkgtjA8zUQtGRao84H/dk6lPpWqvE7riUgP6DZjOHEpW6IjAnjgy
7RjJ+LyIBiav5V2er/yxyFKHRFoVBg6irmZ8LQrAZRxsLnYAdSgy1tbILrvw+yIn9Booyw8OOdP5
dve8Iups7wSOftdCDKeeIohbTfEGKdW2EVEXLpCP7DDGKaWzjjCEKNsqPneL2spP3XCzDh8MhadF
uBPAw7Iucn1OZWklrnK1hIZ/9U21E5EZnGhFiTZDKDVLvtLhtT+ecKXCJvVdiFBsmGB06fXy1E6K
2maPZGsfBGaAJlmomTuuNT6ZrfEBfHi+zSohVVtbuQNEQ6SGhmrQkSlh1omh+DU/v5fj8frhpGsB
mY0o3KY/T87ucmQ7Sf+5ScdiAOhgDs7hViBwEyq84o/hbXAexWqJ8ClHrwN5RFHb4DQznUZBwBCV
0VSr1nQFluyGJmqWIeeJ2pDrueABoNMCKd198F7g50fr8+4PZhV02NLaevzzQwsVTxQFJeFt9ax8
wDDLJac6PkvKVb0Sac4QCQWfYtbMvwQB3/WuarFYJEjSpJG81B8vgjFMA8XfVXFryVxWyICC4xRL
5SGjM5ny9v4BkDeZBDitSDvEujvL6YORS6M6c1Di34z5SKZA3H/9GeD6bGZhig8VlIo5wY1c+h7/
26NT5ZfrPvfQ+2c03TZ9nMJPl16kX42xVhfD+cB0GEkVDp7sNLAc+0xqyWEZ0BmddR/r8LupOELS
MFQSfWDVxLlu0RSp2ZjFaI1wh2vxSvReJv6oj6HISenDLRo/E0uWlpShs2zskmFd9yrquuIkbLHj
DQXBXAUaV0hpwKOXMHEIIfmY9/kbQjYlh7LAsbX6vhKgfCWE8rI0Or8BWkY6xb6S0mBeFVeOCLES
vUaxZjVU17v/V8l5JrKH0Jbp+w8fe/x60JXZN0X5W++Otumfegg9PDQINyYyZLjt7gx4Xp5R+y/q
qwjosj7wTO1nvz0bYoPYpqtlJRP8xyS1dbpgaIQuLSzvhurc6W8oFiF+r+aVfd1svKVSQHNfFthR
x6kGzdXKtCqBrw5fDA3U0/U975oJK7q+GZ/dSaS6iqwRuFA5vthcGXTtGd+InAlbxbxNXxTRDlja
B2r0VzAJcpUUZL+u7so0QphIv30EXLKy1rHgiy6KcR82IxLvUajE7hIeQUmO7cXfNMw0sq7IwVNA
bLOJkF8uZ9mvmcEXgb/buiqX3QURmv2gPj9ITCJUouvL2PtKMFy1m4nN8UDG5VwjyMzqA0aQF/XJ
B3jYWz19QBNj73Y9UU5d6fw2ysuB+8/2fQ85d9EKIcrpi+eeOQMSVXESiY2HZ5UsGW6b1s/O8n42
AXHaQTOt2VFr+N9Fl4o13GzUjt8ua+CrTJu/gxoP2x333q4ovaK4YMmFt/Ky/zN0UcQPKsddbeJv
rw0gCdYduW9w2wPlOPNhTNCPvFG8IZLKaUS+7pnwsWQrBk5TofnDuvODNcocRt+a5795DqylkCrW
UgVVIFH+R2sZLNZiPe2oe1A0//3nS9pvBVLB60n05FE4qYGZ7Js5n7Wrm7Vd3Wks3Jhz3SNUt/RA
RAzQ/O0JLcVJQfA2Jnzyudh4TgvfO34p7gsEcU+yFterDGuUZ2R4n+HIHlb2afiwHp3YHY1u+DMR
TcW7Pv1X2y5hsf3Jr221xehY+YXbT1bY0rLuMVou/ejNRGSU09cSb9yMNSdLjF2bQ43pqNzYkMsg
bGcx0pon34ivd1ZRcRc29H0CR8INwGx+cJ7GYlEs4bXVdfmtV1WGjxff+rvVxoTT/PfErmn9ylFh
vQGcNnenBCQF7JUOrkfeKqlCY2ykzveTiNBqEcK2IK24SL09Zwdt+qbpSrXYk3MY2lpEZALmWXpM
jcZtSbV05YobsbAE1tAOZUjts3e9+Owy7S1mTlpwwwaGLRgCagE0qvE83a7diNvkxKzipNVvfltO
y15PN/LZ83OnnSODACvI5JiU+OZB77xPNKj813QoNCZHCiMaSbN9AUjxOMElZSFq/BXb1Dt8M6eD
rRalAWe+GlRgYzP4qYHUBIxvVIbluSDbK9XEYhMyEZdxgIBxO027ZDn/DNN4SxUE0t8LgGH5rj+O
nNqCJFgc/kW6LHWLue7PF9RoY7FTCB3MUUxi13yVqzoi/jtRJO3izihArTWjY9FD6hgU0j6VXJuU
WCy70Mlra3lDtpwGJD4BfthhQCjwPxMw9x7LZ3dobGIMZHar4qsJM/CzqLjkixXxXXO2XOyuEfNr
plw49gHFANagITWVSu4COW9oIfNUROxsiaefXxN9JOsWfThWSUHoqvqsQYV3Dh45GkswAVBuBNas
hZYzdL8wGQjKOWdM4GQNqBBMQU8pWjraNg0NTqED1pfsM90p9uEmnSal9bpwTTl3437OOyW6g7UC
jGutlvaxGxTwn0zoQk3FJZ+X3pbLrTohAfKpm3Q8PivlTdDAeELo6F9bb4PiMK+G3OPBaPtFPYOo
1+qfzqIheE3wXRYo4CGlkKS84QfUKAmMp7QJoXnb2XdfCtirl5L0F7JZ9xLKFXiZqtfL+n22HOPR
RbPBQQNtx0jTAugFp1DL+GdBYupqZSvXGnz8KP/HWoG6pjh3iY0RoPfsvbffyVMXbznh1thi+oj1
4t7/Oy3qrcuzFSnP/bquotFCodkesbse9oupLaAzAbDnpT7H2wqb4fyGf3J+8hP3OIcWqyOCV9mP
KPyDu2PtqlmdyXL3YwBTarhUlHx/LoAG+pLVNO34gXUSJ8LNMXfKI1B+yT1/l291s9I+02LDS/j9
0JvonPJiupM6wf6F6SmEe9b9J2CyIDcE1l3vgHOSFk5eL22NmX0ldVW492Wu8CFt9JKA2pfmLDBp
h9kJM6IDWDhRn6vV1/eAUZsORPTnEWTnFvtYYaAdWzTInHAqi5AVpwgSsKBg/tE8+JPlbddjDj5f
cAppJWqZEPSA3A6NjrGwizfPytJiqe8gZT5zTM7xM+rqZjFJiyJipw2e67SQ0gdF2pPesxq7Kaqf
wANjCIDcg0iEpgb3DxQbqlKG0HYc50HGq0myuoihsXVM8Eyt/8zeCtiXURyJKM0pcngd0I7twgX1
kP9QQrsqIw8XOeVI4rWvegTvgCZTCtS4QHlhCM+BrZ4SWNuKsEXWGksZUcXh431sUt4qk5Otl3FF
Rm8S1uLLvvKyS7ZBd9H8e0AJ7fsSzFn5TBycJ9tNnqSaoVdWmiimsdNzNvTBLh0VijLIydt8tNYx
oR5iufkxl+BGpk6zwAU8M121f7qh/4/vrc2lhEfyL5rO04dI/ibDBZG90bkUgzKgQ7eUTzhoOXO9
2YNY5ckzwaRiMQ5SnarqddLvaAYE9c6x65P2KkcXEONsrjYlxoM7N3cTAQzQpivzZPRI0gloAEgO
5Umn3FiOLvO7m5+rOzp/rAPw8E89C4Wtm4+LCCRS4oRwj83JqVfoKtOwUCEv58K7ExATaNrImkjL
JmtdzdqZSalAPlg1XZKvx78kSvkEaPqbTCAaU0k1l79Sh57CcpkjgKMxGxP2om2FEF0N5cph7pjM
3P4wZ9lCpT6p9SENzIE1tyFoSJK39dqJp97qM9kRmyBCmozyPFVhXMghkOzSLxn+bApZXsSLJjYl
ikp7ALZEzXQhfrycRoYR3L7eds94GN3mCl2UO1ZPqf4xiB6S64idLpcUoB/T37vmNiZGpbZr975A
bZU3cs2U0IpISwzv7jklat9ppYv7aEme0xpLv22j7FARh2nNdDk5GX+v30ZMKz+1FOdhCCWwjq2s
9pB2hP1R/lPbEwry/G6YOs/Ds62UGee0jElR/jwPQQ8cJHG6o+T93Lmt+bLsUby6qmx6/+4/NvYP
gLc6B0vJzVKp2I4ueEXS9qNgOEnJ60jKJe7TihpWG+WYPQc7Lh04DGBjusfGP6IC5SwrOulyLOJA
feW0XupxVAwL/S7mdd4BQ3x0wFtrb95UTzV7ud1XJa7kzhkJOBNXKj4lw3hD4u2tI98OnIciQNp9
ufahIx+RIt8Idaxd4vFcxU+FZ7BoilMbJ8BNZ0P3/1iyts7B6Hzxlwo70mC0M7Ai0O2QyV9SsDeM
9uGKD0XzIEcq/i0vafmcHcDHvCyTMm0H9b/x0NIs18Bo94CdePrgZ9gnIOP5t8wz0YToY8huyOc9
S1ToPTi9jjmlX7Ju/BMt6s1SPpHT6+ML3TnqPURplW9/rO5trZ0Tw8+SLkPMIvKhFWsnXbC1KyEH
X0goZ9FQLdcDPTvzp46hFJt9u5zqLy5KZbBMUr5Qo508u++sdmt5Fi4u/PAicKzGfKAqyWz9eCzn
QbsqOoJbptfieAONqA6a4x3hnCmHouxlpTrPRs3Sm4Vmyp63+fLgrViO5DC8afWDbo8MDLNx2wXX
HsIqtJHVbB3Hml84C0wUk4zQb/yjjj/a9+QH5n4LIzS2Bgo3BlT5M49viqNOXPAKmWbR2f1bzHon
CXbDI6eKFRWAZeBzunByw2L2T7mbuaI1c94KaRrQCpT0idjlRE+FbRz06e5eJefou1Dg88sZ0/Ce
8DzCzOxE7FX4amBwQbOl1QcZNVVcLvuo2Q3JYmkfXS4sBZH4kEkYMxZsynHiDtwwWI0m4DyFnyOk
rp0kXUCYJvPvRTPF56jVrRR1chbwPOxvxnZD5aOBO06oj9BrLZu6W/GyievC+QAYTZ7Tf+grnQwJ
Yug8bpL5k1EpNEUXUBWxr7prUjAgXOQ5WAJiKkWrDHIoRq+KPPr0XXCE3MwxKb/bPkxB/1M/lfkT
C6PDZSLgCt7LUUbNCnhGNOlTaSdQPoRuVMYOJopKh+aRyw5lZxwuocMY33BGF9OYjPczu/peRh9T
7SA7FKcY189J0iAJ47inOtSP5cAZ2mx3Ed+xegS67BLLk6sCaR1Sho7pk1UebWaHdlSU0bfcF2PU
kF6zos30hey+jHCJU7U8wRDXqzgfFSZyAoL0mq1oEOiEwvwalquzsD/x5HRtoBdsuPfCdX/NiNfW
cFgv4TJaQ+V3UTKbAbt5HGFeCCpQyrz3Vzp6RNg0f3cb7zgel5ZOSzgq2S1GViCu89JnKaRue3TO
WzVd4ovFRmSUp/XqnvChrIANDgtXz0wRTbbj2ApS+g3PZVFqJez28vkZXRAiEp9UySyaHbPFYd1R
1NqhXYLRo8M/IHUjsSBPTsB5c/fW5tz3olEef2TFKbU1CmAQEEPOIdVcGLNLEmYIvr1d9EO2fqhK
d3R4yMbuosFgA+Mh0OUv87fPB7KLft9nXIcSLuChZXjtpTyQ/I9uUsW5dRjNGN8/nocpPxsNyaax
T2tFfrfAeUqINfPvk0yNAchWfK1HMPxuQUqHkPcV8LBiSB1O4PG7p/HmV8VcYdY+piDFlVfjAwpG
nw6WUC1P2je3jjf0gzzj92uZlN5KXS7kCurtOZEEG8hkhQxcO2Tj1DhMuDE4vSuJUIhyBCc6eTvt
YMmY1MTfC8lyh0JDL8j4bSRWtSPMkIjkGFPx/WvUPW+GVC5Gb8ps8lZR1KWnoIOACxs+gqoiJsGa
llLvWG+gZ3lt0t6xSgaNWnTLUaFO/RPmuQu/bbCNVohE1qGPQVw7/fbgP0jkvNRC/d1yQEVmI1Ne
xVq6a9CHzWuGLe5jdGt3Jh490+VGcdP7jmpRxzlaLIa+pNbiF+4nY6mWe02BBXGD9En0jTPbLeKe
ZSgi9VkIiRBgNYPP0umDw5y2q7LT9FHICu2hNvJYT2egm/S42rjPEmJoSDIHXsdcg44IEzPj+Zjx
YM+ACQVN7lOUnX+13vsSVcBNJNpmg9qHpPk1MLiIkx2BZMzDkIhEJBcbvbKOR3/NWAbeMcNyUHWL
/jbKoMjKFOzyq1BPVBuiuNRpxEMkBRmgbrU1kqm2fxKspZK2En+WLGXzrJB7cOEbqJlju7lEztcW
Joa9Y5iV29W0J4QgWUYTzemge9C5FtgNsVRXP+uztBefZmUwVGYrqRo8drB0RIm1+c2uANW29O9/
g7ggxyvy63ufLVw0EqbOtURODdwyKpPeBdSyLk92O5Sn2Jduziw3L/aoEXc7PKL4FVE+hMLJact5
A0iVhushcAZppcRVBi78Trs4z/h4sFPSKLqcMwV8EO2dVSsGn1J+CjzL/UEsMH/KS+gwuN+KddBi
zul8QGspdmZrzZrguAtx9O4ij/ztDxe6qILNr0kLCxxinTIph3eNKeuXS6bSuZlx0AK7bNFDuReD
35LBcKMpaks2IAY8tSU/cWyf4R0hEAJEQOeYtbn+/nZIAxIGhHZ8bN4Ejdl3MumWlM+y2K39J3Ta
x9bKKtj3elDKeWJROso/PiRHKs4IGFOaOY4qBcPlFv43tnFU+UvOFPRhb0CCMNwy4uMAwlDNw7OU
bju98ZIIk7mAjPop3CK9P9Q+/HiItifFvz5HaM4U2kDxfSrCfrw+ySYhPlZo0miFlxJ+tVUb1CpF
YOeyh0qVtkp6DMYjF1fuq7PFTLhivpKljZenuzr3U1jHHcbWO1E81ZJowc3XQ826xgTrd0HeVy4R
v8CEOTOW0e0wvJqGhQFmQkCFWT4zMQlwAWIAN7aG5qVYlrrzoUgZ6+bXEg0SFByHrWNVYihBxpVe
Z3xWCOmUAFRKZMG5BQ4f1UZNvziaBmvslhp6OzpKi3Jxak9glppKdfSvy0Xe6F6qfYOqF2HPJrKv
YqAN8PHN35CvSn32eOjJ6hWD/4U2Arvs0n9gOZPFVCl6qAz7ZTJ7lVdEvkXldC42mC+IPpd7wvMK
t/nkESHmtch2utx/Is7wslftksCL1xGDJG5vSvC+lNOg7zT/WzU0wOBSyne5KxTtdBfw511Z2W4F
ZY/AnXDKv4sIFVVWKuFHOjA5/nDB9xS3WvrMZmnleKVLO/wjOsfAqXGS6gNnFNYufcdO5H3n33X0
rAsC19vym98CZLhq+q49OvSTj5B2H7WBLtd05+giotP9XvRYDdZnonB4lCq7hQk7e6QhivWE8fL5
xYghlWpiOEaLPplKO2Vf1tDkGaDmKVPHLdoj9scMP8OB8uBuDYs+VKUddJi75NpgVcPLMn+XbUJR
ZD5fX8CqOhDkumAJjvQKw0xt0idSWtIVIkojeqKC3zHntWjO+a2QoKGwtWMj4t9fm6eCvfhAbgD2
++g3nonpHm9ptjeMcu2ihdFZ5ednOkJ7PbLpj6p6wnHyGbNDXHz0a1ZX6yXM1phb0OYkCdDJSFxa
+xQ8UGQ7NXGFY+YEzXZNote3w+WP9+svfqPNCAZcbKQp5khxmbhRViwDoix7M9F37iHxJvdppFrv
FI3Am/v5YW9AD0JCZ7kwRex96NRJAXZHl71KGUk84j3M0FUMDggwU2MP5XMkeVqCOcHW8XdNO20+
+3OSJNYOQc3hj1viNBye/AH9Cfpsvi0hb0TkWxb+xTnJHaosH7AtC4/lLGwjizkwLeKB4FTp7oMh
Scws7IvKW2HEU4Se1llGJgKo7EJwVQ5h0+IYUI28mZe5UcJd85AGYd+6RIJ4cFXVrrIr3AH2/+5n
h+V+YmvjjZ/sT2EK4F8mh2FeJSQyxVQZTN9H5AQJy8csky7kz5DnmrAN+385t55zdHJo8eXP3N+s
gVD8O0LbEhdS6IplgBThbs9VdQJhgJBGXqqzYX/HX1Q3ZSiioW56tSn/gj9twaRyUlkY3t3tYmMn
EgO809UZnByL3uUsZftFj/N9WKw6AEKDr/Xy/bchGJq0MvNaDfT8yaLRO0PEI/kPPqa/+r5LSL9k
SOuR0nFbGcZXhfmJQV8QpEvhoVJcLrMpv1QMzFwfnLTVaLeHWysnHdo8Os0iRruKowzxpT6bigBL
FllrclnjgT5Cszr1yqBePduAabC3FGHI192DR8k3yLJXgGxHLEKyf5G/GZ+7n97nPXE3HHQLl8wr
LEpSlhOLUOKJ+tSmkvrR1KGcziy3YPPpNDQJNAXmwmIvrXfG5yWYQZSrPifvEliEZVckrjuyrkdN
CqQjLY5QF+1GI2hxMhDdCva1Iftumt/figzjp2jpC/mmfmPJgs3KvlXja0TWq37nxF6hwUQYjQCK
r4IY2eCmE/oP+poZ4wG2naqot81ZsjtSdZX92K3RY+ASmcFRtu5gJ8UpDJaHjJV2q//Kp8rEMfhs
dLGk98FTlFW9Nct/vy4A8y/k9mKMLBqBTJqiFfJEEyoMLd13Rg5qp2FbHCi7h/x+oSI+ViWHYA+Y
HG2Vta0NCPWHHprPo6KsNgXd8fgcY4g7TIcDTUk0SwvmfMIK4b/V6cbluQMwGDKF/56bmRCPwmRg
X5pDPJyCgPa1VZ9Nz5KyKDZMXQyL+2yfq9wkkRe0U775tokoaJnHGGaeILFz6hzC/j1xHgtV3v+o
eg2si8HBA9OfiaGvnruMChalIF0F9cKDEgIZ0PMr+IaRPXnwETgSVtdGpj+nC2ZXUUDQnrepAdTX
AYnyoRMzlttSvh87W+b6c5Ju/kq6yZScdLf0d2HIBxSmO+Hww/hL3XnAhTYu88dNOz3U6x5avTDy
qSynvsvX94Ee4LwaykRezFRWTFe/9eVL6A5Fy4JAiT2h+MaGCEtsybameRAoMEsJXW3IyDOruXbG
3OWro+eN+xOdOPtJhrUgnf3O8GCoHaBHw+2h39nVtRcRJkPoahcZrhSYo6TIvJTvoQPXbQrg4D3S
RtjNCCY51qSb+elQ/iCaEj6MAUp8i51U29t36yx5C5QFD9XjBtYX7hpxoTvNDwtiYXg04RCr86xy
H6NFF4xYD+hmxPsDoQFjc3JHX/sOYlvfaMrELfPYtpTQIg1JTc4Ar9LfSHPHbyyjUI8bzc1goHPk
9xpzyO2vpzuXSPYmb1rVo8q8F5OIzBSyl0I/WkRH3uSH3jaa3FrGNHjFyOqTAeVRSA+w0zkFFEN9
CB8u8wOh4DNo8HikH4VqMOvfIkpA29VTUtfuhHNqG8irbUdByqxCO3l+kbR1z+36K0/lWaLWQDqW
qUzgAXhEmJcMmLz/ade8DlcHlDiE3iJ3Go7SWIbpu9+70Wv0idFytArf0Ar6cmSe0HJLZn3bUceH
8C/SKh4pyoCAmsvb0O9WP8zMvrgRBg3xAWCb43Buy6xF25jNNiV5z+iHnzugm2pu4Pl2qcgQnD7G
wZk8GyofJqDUlGhTsAtG4+onJDQUkpEqV4TV1byO5cvN8FvHSAwLk3RWz56Mz0rsE5aG+8vV6D29
/YrqHd3vHFEYeHgcjiEVYrhbAsujvrZnlxP/iL9uByznzbdAm5OD8ZK81UEupH1fQYsec56ZDpNb
bXHO9Adyg9blEwvSJbFuFPeQwEPyiicM4Jv0OoDVbjPc7abhiKlx5KJjCzD/e4O4f1yeYXtReTzp
svAv8sI4FbedDfAVTX96+cSW6mxy/N8TkZ3WlsvluTqdQV6rniIrIo6A8YdKWOFMOMmBVaLf9eMV
K+F6Hkjvl46zN/zUAUfOoB/0T8/0cdoD3L1o4YO+szGWnh4B7flVWyFPOI8q9tGHQUnXfAXipz2N
ffbL6UoL3DvjETkTTWbVgARGm/u0Vm7jGITR05whtYiYevxmb4XpCNx9VkL5WkkfcnxiU8nrfVOO
nB/fiiWunKOtHsDAYDCCr5bzjq7hhLCwkaJUcjh88N0E1x8i0mnvTTceqM0XLNKdMvDWgv9jm22c
TNdnReWX0xX+F+9O+xJ9zEQnSjP4y/mj3Ywt72Kgxe1ic8FoWn83ZPjapIO5dcj9YpzkdN0731tn
l8VZL++0oLlrpTXk3IxKg0I6pCMQtLbrDAMoiMgZLN5maQqephU6uRbS7hqcOyLl8YHjII1ijQNz
7ZN8cFUyObS6Pes3aFCFaYMIh7ZtuN+wmn0xXIGa8aAUcLmLDi0vg8dQG2EWM4soHUQyYumyGAY4
K+4bgqLUJ8drMBl9AlJ+4UDdZSmyZiUyMtQt2ZpIQXPXtngbBKXkh6L1nItM1EffkSeLHQAKHJCw
RxSRgwOrXvnpoNVPMl3WRt9db6czXH8KsoyzY+ifekarqP44lukpTFP3+JEHZIJSjaugUS/VetMb
rpQxx/A1d8edcsxsyQISkQwFyX2z5S7cFxigWG6c5J0y4iVUfJe+A2NuObHe5rAHw+92ubQH75Bn
ylicDcuoJMjNlrpGbftE+VRJVFhDQ32hvSS8P612pKoxFzZ8FlNSLDa9m9IN7c5o175cwQE+KKpI
TNkB3rRSUhBADDOCKaXDBedQzRhK+926/wlV3NHhq+v7jmRn4N+1icxeTURpQpL6nMQ39ynSDAC9
UH6VcsktbMm0HpWY/NQy/DSdZ1R34XlQJZgN9u2SCZMWVmkBBIhGO2oRM9n7M5D9MgQ8DLxQh10r
dZN7JLkqjJN43OM/qwkKR1EWRzZGSQS58Kv6TANy7OZ+trOAkdhZT+zCkwYbUOwYnq43N5KI6brg
8R5Tr7+rVFZ7KBiWHX0LGn6atWTGMWfG0TdQAu5IWyTPLM4YxuD+XIkZh2FSZRT0dobCGCewqptr
7TLKACCInJqoL6mqlhhVz/S51PmEStVbU/5Qu9w+TEUenLzYoAcq8R3zMsMLqrBAg9Kaf5efgqr+
Vz4uqiyq8p20rcNfyp0pFZNnJ8l9i960LZiHFjNIx6qQor/CId1hBs9jwEvqugA9krsJ5bF/CKr+
eJZ5UkX/j9l9gqmQa6NULlcjPjttEDGncHjEWqwuKlmuDaY5DP2YWgRusugPLGHLWtB31Y4fX7nv
jgpggGlMudLgQV2g8CKGBnA56yuB7ZqaVgEcxb4OCz18uQOnD+ZclTiVQ9GG9rc50sjl7lFUtIHS
scybaUFvrj05i26oG4QoYdqw3BQlNGKpXrPAYKXAixmTJy9W2w4cTe4MOh3LqRf1D7W622bv1DrZ
6oKjdRMOoybUH3PP3Z7m5I9+u/yXsl6TbnmQr7GEYU3Z8H/NoJ06GXSBBXu4rElQnWNAZRhwv0eN
V7LqwNGMLqXHGmpHg68OPagoIXGn5zGM0TaLHIdL1btkSPEJATErr40kuwo9o8jbCDBWNvQDUY6p
Wu9ymfuruZfZDbGIgIvRm9sREwC/qucMsuzknW6hJ2fAUFF6hYLc/Sf/0E2i9TtzIJPYR1d3MfaN
BXKPBjQ3dA/Jhc2AzL9eNCfJR4kPtpKUp4hniCudttHlc1UkeFClSXpurdvsRmjR+x+AJchXWhSH
rlY6ZKso/6XkYm5dA1GVeSykXJOsE4Has4J+gSMhpsjMRRmDj29q2MXI6tmV7AKmrcmSRHu56cxg
OtzSCq5aMLtruDZf+GxAwXj8My3fEA3kBdl5vX3RMsBfKWDIwWmHhe/b2BKsfTjxcphA2vGGOVXe
ap/wW5aoto8OZYBTBKoSCmB4vklh6aJKgIWgQzTYR/XxnBSzq2IELF3opNTy91Pe4jP/csMeC/df
cyKb8I5vN9IR6PKuYTYkGG8+tNQKjgJlef8tMvpgZUMWmtNHuLKW0RKOafkpz01Uy0CJrsYOrhNa
wv4l/J9ksZQC5UfNyRgau+YG0QLD0HWQ1rfiCHWxzIG5qfFeKkzqZ6dxtKxYLMixuGYl4pFDVZ85
3lXqG9TWWQDdMs8GagvbRJ+QN0rgtsAtis76JKCAWzOK2fTSofuqdOI/KoI2p+A9m+8zu/z7A+KX
CWrw+WNurf8EFDqi58r1QW/InTYIx4qeCp/tGMUNrPa8T2MyPCn3reTfB0pPBwpFdivwQ93BVLTu
LBCbfT4vD9hqqc1EsSbs7ZJeBTRtjXK3cvu6ih5UFK+7gDFjn3awNXp8wfX7uLMKkhX/R2+N99r1
elHXWvxSCfT3NnhSyGodM8NhPbjDw1ZjrIuszElUAX+brQe21MHzAArE2s+XOeXG0MUeeoU0w5Ci
auEeffNmXMwjuzWeMKiEEPKRWDbkiXiPOTI2wfDBu4+cN/cBUxtIJnBn61Ug4GemwlfeIifSGt4V
jRugdZ7aoBIRYQKbtIJp+v9kVcMzyLMHonhyYdJVcnjuY0y2J06ZHwCKK38M4XuK0DQJfQo4kvQJ
9Z76fYcDhxhT1W6PUealr+AFiuKvL96YCMqpRrPgGtGqiRtotTrTQk15HgfN4XggwtGaeXQWoo8L
UopqEx2CUyIeUdzk6LVSyzR8hSXMLCe8QMiZUKXQ0ZJDcKZQ7QoOogoZkPhlsfYiqnPCYl+WUCFm
x7CEXYt1UjK2/LvqycV+YIQGY5Qm3Za6Xgjk9aVDwJOe0LgllnuJ3KdFv+IkT7LQAbiK8kdSs3v3
XTkHGxThpd7C7HqnIE0sNm4sG/bSjzqgoFBoc5XbTtOn04yUm2PM0OHP37TxWPRKuRGgjZ0qib7H
0UdDWjI6sIZWvutx8FaUIzg0tIaVCaBl2G6wSeXmWgweI57mnbSYg5gIY9+F9XQlc8jU95APzp31
LRB3ZZazop3ao0XiSWiUJawrFnnasRdn34sxTVypBWXNYIUPJ+d3vOuqB8aLabrs6MLR9VLTBgAu
kJkvf+spo3Vlz4NUxSmQU1tkuHvYubj6WdzzrKy3NzwSa8y/eqWfeWLVYQ842Rh/e2dCRN7l6WrQ
8SAPkWR7zeMczJSoDCH4C/ANJ/1uZPUU7B9LN7Lkf0yVmhbb0S4PS4wfNAYt5lloAJ2Oz7DLS5vV
qHWamSdBxp3b76Dket6a3nPmNGVPHE8lKMdgPv5WLWLNSxNRiBCkjl1FRGOeXyNMKdRusOWnlkRA
VouUXI4GLoppmEeJwvz/XxIw95qsqKAY+W673KPuz/dOEY3GlWs1jpOwB7PLbXkk4xoSWXs6yMHP
42hkoKAyE9jRNvNv4ah1BdQcCpk3w7/3K8LbOdhEs/olJok/jQqBZR1v4tzVFDtZyehE7JhuRk19
Vre3B9dRpzW2AZ0bopjS1Vc/xE8Utqvr75k4+Yh6fe009208IYtaKiZuPb5m2Lqt/eOuBFsm87pw
A6xThvYJhwE+xM67uRpnm8zKTgNNC2y3PV02u3bY+q6zoRJvtvItFzd3T0EjykQcGkF/4wtyA36T
BPRZGcGJrUeHvKiasK4XhLE9Tkx7x7UuxGqwywsQ5eQm4xVgsuuef4YrGvCnZOg44GRWxyt7g5ns
1a4zrcYu1dESX8cOuVtC+Jn+fSM2onm+jWa+dbIskT7vYCA/NUNyE3HlcwyMuWm+UPwXVlNNiP+3
7G+iGXi/DpjW9RHm0HmJpCxjGFoSZHXxDLRv17t8sFZa/bjsEeZZb3JM5fDO3eQ6/fQA+XuV9Alf
EUsKVekCEpLb8Hzxn8qsDMiAzzu8wUYbCiI8Ry9m4ZkE7kuvRLUBtCwKIQylAzdjamR75GD4N5+M
EvmdNMryaCDW8fURRYqKTrbARJAnt7uZ2QVnUG6g+yjHBuPx6+OxpCXz9rdx6Ft76IiuX9hesEOH
5QbWThmFkodj2UUQHPA+8AqlSB/NK2N3XEOxIFs/gZN09BcaR8zPvC/kts79JZgOCz0Oz8b1N7bk
HqI/skCOyhq2YirUVqhp0w7rkrnYEgAOnygSiNpOzNX529lvOVy/8lNSX1kW+DrMmj0Nr5ho/3sj
3Pua0t8Ct8qNITGB1Vc2UdaFrqFMrJEQh0jgVZ3LB5+o9MDsl/Iam4Lwoqje7zg2JvVi8C8gUTFB
bqH42vQXwjViww4w1q4UYNMOMQG+TRGMGi8CCQj+aOuQ798i3Ve0R+32azlw01PzN/C+cfEP/kTS
j9/Xw6ypig0sN1cvAq4OFE8LZVOXWCA3a4lFspmHdEuJl/V0B125RTKdvm1DZcACRBvrRGD0j2qB
bBpXvncWG9Ilr98vBGFSJ9/5985uT0wzifzHL7/0KaZT7o3O0g0+cgzFfa5io0WhnhCyMLq195DA
MkxSx8ecy5+PfT4Qswbz8nL9uKRY6ke1GsayS34vWVUy6uJb/tIALtmmOj9HrP1kil7VNWS+Zc6I
Z7uN3Q26xIVyyhQJWT433kdTWPuCgWNC/+tD/8q6jN7YdYbACa3TdU7EGqUxuxpZw4DUsG5lSzzi
QtHbjXW+GXq50UXqYHnUSUbGjYFO/AWXB8IYfzF2DL8bVAlppC8wa9D7BNka2jDgPcAOVGU1QCVE
4xtIvO4dzxWTqcintp0VYWTvo20Y49sAgjqYwIWST1mxIM78g0V+J5iujLaQJhukw2XiUeAAEiG3
iOBtXU5gF6zObB0ZBVUCdNv5xzhsS1HPnO8iRmnwksydTPCVh72g71hjzHdedxY55YqmMr5snljw
bHnMx8x5fmsilFvA7vk6Q/2nXQdr2J3VNDrnqpbX0Z3qlvlC/M137xOjcPr7IaVUUulDoTZjV8pl
M6cHwU8rKIV3fbBUONpX3RIXmMUx7SiBeMsxuISkFW9urfagxcUhWYBhWKyLWnQxb9TWqnlYgepz
iDgM6bXkK6vsPLIU1y2nfQxaxgtYQ1iIDrDBTp20MASZs0f3Fl+rHYBVgtZ+dfkp1blh43ZGYkbn
HJV7CdwAF8BUqca68EPO64GsvdkTelI2YjMJi6IlvnSppBd5JAYtBME8/WSALakovxcaGAE1Umr4
wEDEUfnTGzSBIgbdETgiMRNYYqaq85KhBnuhXXdFdm74FNPljUTCJw8WvdzikHBugzEwGLuzqFe6
TNWKcAs+RNbq/e8dM57oJYRNTe7zgIMax/lXaf9jvRTwYoOGKVd9VF9bmxsw2xkp2CY8n9fpNm90
i5zLd/cLBpVk5iRHLB9wUrnczL6SUNHa86r/cLIW5y0wxUzmOA6HZXF5LTxQgmIkFoRKgzjmz6U9
NZ/V0Z+AEQNjbnl6AaO9EB1hfjIlxkOMvYmGdOH+9Mm8RdQdmcjxpOrActX4EgtymzAIdLT1Iuqb
m1DSC90ijdyweaHM51viTC1/fL5Sodxk55kBzy2WZ9OGEG6M+Fo0pXc+sIHSGYrASBhUcYbB/WG2
+KQcFWocfN7Z8roZMJkMh1aFwkKzQEwJulkUzaj3aq6Wqpkh7V8YufafkVvtjhNRzdoKnfIN4Wc3
DZPvFp5sO7U/zwX6XlUNoZFTutXlzXDAaSZEcc/JCP+swykNDX5ZPs4nTVnkAd9dLFXmxqwdDmYq
96BKMbzBybMP+1+pc5mePdbqJgwvDMaLuzBOBgswDmSngvUrd7TMeTKEqHzSSjb0sEWl+Tp2A1MR
ZGVDSakJxfPGw2TzmIvcsc5ltN+TdlIWt9QuFxGX99b3Q4OdbNxLXGhf5C2ZPsjqVsXL+2Fl9W//
jnOdHbVbnClVkZ6XTU3QaPbGLJR3T73MTCJSQGQzuQm/3K6jgxVJ4BXmFxXEFBB8LGZ8RZnTTjWF
wIpMA27avYn+9Js8Q+15TeDBWfwsOqOLDOrmAOxmfVI1N8GdUIkqkFsPXv/yxjHeai3LaAML3u/c
K8qlQpiywChDbrAQlMekK23v24IDtkgifChJcrWdrOgme7+973xYeZqxXyamCsT73BReROc/FW2/
q4/WFYY1F2cfUa4f3PXTUBuC7x57TK0TgEGYv7LKdatnSvpWJ8i6ezqoWH0JB7TSHkYFm8kIL0OT
ATBwWmJgy5oqlGJAz13GVgr6BbFyqHJnW6AGmnlPgswMT+1jHlQZolBSU8gf6CwIgkE3VNN/SMPB
2TlOmTXDHEbVXK5X699A6zER6I9ZpYJWgdF5oCJgTc7SPtT+98mkM4E5fchh2eDtk+FsFxR2mPNM
+CibkcUFqGuKHfkylrBXuKf93Ehe0m29W8MqVIOzyA0OQTOvoPmWmAJawUG9Ixz6Hlqc2n9rbJjd
N33QLpG8z7cB8ya7j2Lr+T3+o3tfdEBsSvfM8huSRML6zG7dQpCwRBuBdgCHxd6m8FycShxcVUEX
iVNLUjbT/59g3/aUiWisoNl9ADjVsTN3/P2iwaXFDXSlLXHnCe8pBZLRgu42j7N8UDthIWtaZ3FS
iGkEVK0C5lyQDO8O+tbVAyVZDpH84tgLihEVM12fEKgUWvOk+NsyLEIWT+tP5rfDsy+9PicsAW5i
KxSpPzJgbzuFG66CJpkaZuxke479VtHZTjPfEkScSQG91wa0ItK0VzJsf1+gvmYV3jtE6/rWBg/n
rS65tI8mI6eQdDVI/hutSqYmH1jGHdCSfgSiWJUIfCr2F2LTegPgzk5ye34l/RLg1XUsnrEB8zqX
nHj8WQBsKKuXbL/7ebKhDB7P7kGvK1GZhSswbamPJISkhL9IvmF6nOrjLQdp64rs3fn4Nq3g3WoP
pToCs0N5d6bwUYx8njVFd8S2BHlLIKwsqh+fMdYoJZqude7SWu8QHeLq1lj0I5pRkIFGfYNdEAvU
tRcUs3WXgDZdUO31iehH9mIim1jW5Q23fg56kpS7v7qoyUTZpHgp+AuaH/vte2xi9e0MNmjR19kb
/sRXb5EEZx7MQL4VOd53+hAHs55b+n9MmgwTDTs+WM8sUXdvMJ5FzyBW9fQ3Hmhx5TYPUmy4sGOa
Z04XK9QZXwsI6PHSr2meVAQgqA3V9iGHsOhsdoOGZ+dpq5KRN4Pq7JztnEG/scGHJnllNkLhDODE
0iFWxiQ3NQ/1wqwwpW689/AR4YAEUWWj1i+W47rJqsczixuAGXUtAi6EVpFh+fMRyiwHU3VkXgJP
sJy90tSaiab7qJ+Nr+RdUGQ5MgdeLgC7GqqLC3BtfvrU3PFsDJDw4Ifdml2ux/45C2058gdGRxxr
xyV6KB4NSK6u772cylpYOZ/7TwlZnL35tRs4s2YtrhLQYOEOjfDELMCvGzEx84NdE2Tpk6meBTT4
4LoWk3kSX7ZNBRzukVwtYWN4qXPAtVD084oh4l1fb1gNpdtYhjLA5hEC/Db9NguIl8Lh9tcKAhJf
F59JLUhson960+XydCLyj0pQY+F/Q0+wAWDSj6yM7l1PxelbWwkcrrIDAKWXvn1zc5TwJEBAuUm/
DcMzRK3WI6UzNg/A8leNxI46OFk/6BE1AcpLS43efU2QtSNRW5qTWtZbyYPK6z1er55G8TeLZhO9
HpX8QuUfkrKTQmuzaXRFL84CICCnvOyz0Zfd1Fn+IT5Xd7PFuTesHathqN7ZQxt64isT0dtOJ/Ee
sbYkxhU1RzlHh0LnX5WWLHThLIVn6LsSd/0EdQOian8wnzR3x7snWO/0vLxOPeExj46vM/ntsaYF
ASVsKbzyAboLBg29xC8bJuXZlLZr34AeiE4lk8b0vSAPWqi4mwbvidCXn2OShJOL2o1cApVizaDX
plW8+sdN6r5h4NvBP275kb7EqPDPx4qErv/4GM0zYW1WYLnnZPQ381X/DtrCKy6mfK3KMl1eMmYe
634=
`pragma protect end_protected
