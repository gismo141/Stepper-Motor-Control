// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:51 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l4yXLr60Qt3LX2punhUzD0yf3N5M7SId9GNc2e3b5PTvSRbI0mO/HFBpmmJzuglH
XxUHlVBX7wHR/x/YYpl/36artZEAM5C3Fb/TVnmdlozcfucpoTduBUg2axdYE+j6
U19lOUSHC3oy2oB6As2G/Wb4rKeY+2c/8ARadxGjdlA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11840)
tHIEYwreSJAlBzTX1oZGxCG9M7glqRv1er8N1ohCz6c+77Nw+GxNmuEtEWADilRm
gN1wTMxZeBkm9NkOfSlIIVsd5kkoNkxcSZE6ymixdUIgw2sK5ROzWQEhUsmgVgmo
3lJYBSdX9ULS4mt/Gq/bp8PsS0fiuu3i4FKecj9FQdnjeCGsukvzBjYvxbJjPqcx
Z4MownkiWj0UaItLskTFiXx1/AeMrixf1IClIoo14shhD4Uxz9n+JXfjuPgGv82S
kPYgtCar/ask9eA9WrzUTqeBXTqJXeSQWYAyPVLKi73DzchhVPTmLO8MC4dssGMs
y+GF5XV0U9CppQq3xcylZODvBWfuRBYhbK5Gu+VFRTjFDfwieqIpCBVE8dqB5hnG
MzFMdWlaTPpKQsgXKyUHQ4IY49TBPXoF5A7khlE3nMgxigRucVrLlFxo8hBclq1h
hy4uEFRueVRMc8hWR+80Z8zM56MXCbLfLPciLzg7IJDCcTMJoAcvp0b+EqJbfVp8
Pvw9JNAe2TRtKkvoK8U/MaNitrFdGuIYcHpzEDQ6/6YrkeFBoYautttnPbgSUWdo
XHESpqqKpKaw17CYenVLkGdBfnhOiSkTwzWtQY+ODBZ9WvvcpoOHTsm/mcVoI4vO
oPYvB/lWKVLwJj8x5w6H1l+/EOb9kbcCdgKJ9mvQ1XRDRHieTyAG59UA4VVc0/s5
oMswgn+YDWEtQUIWvC422aLUlBiV/B9XYtLJ/PUek+fFpcjK7fW1CZruW1AAsDCw
ptBItCBlKjfbw7tsCvcsLbUg/ynb34Ln4bw+D2sKFJhHfinLuaJ+QeA6naiFKF0y
O82/q7nvmsfiR0fsaFscEi/GbGiDp91N30e1eQ46d1f1ZVw5CnCqDCqp0oCDfqS/
Iuq06CdmMhM/Hx5gAJogrkrNUX2P5gQeYrLBlGXsogIgCdK9DbLJUHqLWMMGYKGW
pZ/JQECNAMLz2QoHdoAPPxMMiwzxQh8i2QZB/C5/o006fDG8YAW7svixMVZ8or/J
NZ1CfqYk92qoswQz40soIaLi0GwFXs5YJPK9on/nB4jsjuNk6F84WLvGuSz4r+dD
wNea+4DW7Vqm22zaxrD6+zt0HL5DI18nc9DH/gjDx95X4SPAvNLpjiuVqYJ2l7Jh
b8nHvst9bQqBP4sQCPFEa/9PB9wf3epg1yxGHn5I46JALBKKq0amKYAUwv7oTglW
Uj6XI4pc2b+PvU6k5Q6q9IUg9L5u14E+eVSgKwtz6Hwwqz8dGJs3e26xuYImbEdn
RKpWvx96kPzjeqhLifx0Ea0UMhDcvqOwevoEOkR9pv0pP4n+K69G5upIuv4RQHaH
64nXWLBN74ArvmY8Mdlmh4Jvn3dCHAoT2iZw+YwSfn3ZzN0TLe77NP+ICaLEgG73
dTst8mQX7QxAGVkw7UxsVWH2yyn6yKRgfHa/DitMk7Dk1DudP9qJgTrKznX9MJuB
KLpGt6C2bjqzEykbCxgMJIQ49X9r/wxeB+wONkw7C71+vZmjVyKm/OhMfGo5ZU2d
SQSyBWgi+q7/F9rPC0buTg/NSgUNJaeSg8bd1W7J1lk8y1dznukJcZkWR81CIP5b
MNf7Fvzadt4siagmjiQ2EfUAqJFsRsOrnFwwZOD5NNCR82vJSXODiMWSaZyIeqs8
yZ6eAu6RGydh/QFGLkXmkh1W6lYmFkx+K4ogIglMRm8isqZhg4/6P483cjWNByo7
r5w3OdmMpNTwO3Cpfpy+cGwGeHjsck5wZ6NdQijZxAP4js65epsHw8zub2NT4rzb
WySNTZYSkgx8xBrt99iHLhV/AFjikA9akpjJuS7LFns8iXrhpQYyDBer9iuwgaT2
3unbmg5RNPNO60OI96B0GuGBJlF+XmF5upuhGL9Ta0JClG459VEA6G+szfAaSzpQ
DJpJJuIsREhYgOep6f4LwqYnjdh1Fqathy0YZ5mreHtJQcJhhW8QREnVkuVXhoEO
tcQLOQwbiDO1Cf3fLFAvsPx8emHIrIUZuMXfpmA44bt8uyYza9Y+KD9Sb6bujQlD
QDX/yseJO/+wZzoYzrHvzybZLeENflhEbVUnmcRsQeMBbXWbMIG50Kb6I4dfcE7v
ltO0ammHdV8B5gTvbe13+hmvytQOKBlT8tLN9lGmtvIFXnPPHxhidnH98C+e6j9q
UjPjKK0Y5ShNUbTPo04ONG640uc4COGQmeUKdX6nlqinK3t8a+62jQPo4u9uM6DI
BNmXxOrcBp66wZ6ROhqLf+gD/xKaLmnicmwBsJ0x0Udi7LZoFVkHcaijHgRFEhOp
7Ac9fNMEr3HXuGLmO/e+/qHoON5nbFnFP1zjZjG4pZXxzN4FQPJ5Y6Icz18OBJZW
CWSDG+LEkWdQoBlgl2ddotAHsuNz2q+zmLIEStJsQlBpKWn45TgxoBFRiTCNI1q6
q/NfRqoO71K3NW9NWZ+Lxx8x97ILkUEbtGmt9lgd8tybiah3VeqXZKFBdf6Qawny
uhkU08L8LZry0fAwZTf9MtVgs4YyNV4nQdZO2vDvKGtNz+/sFT9x7Y8nl02RPDwg
GvGmbQabx/Xs5X3esHiDnucDjdcpdMromsc4TkGce9RVXkQZg9sYSE5MhY68B1m+
jeK8F4XNWK3nsCE9GqkDRZuvYXZ1PHqowhCwErJl5WRgi5f9/513KwyhQmI8thOv
+E1wtPN1p1sz40qlFRQL1d738HSg94Py+YvThXbx9HkDtYY7RlscUEBzj73T9O+4
CLaXvfm4YvbJbJEfyQBYtbJHlQIRRU9OHhVr4Ao+xZ3cqmEASEHQrI6Dh58CuOuL
EGmPexRkY2Pe782fK5+aCE810oP94O0sh847BZsRbwby4+CqcMK3B0Dwu0LKqsSk
UbJEPRtPapj2YBW6vTIoMWr+UKe3vysr3Kano1PqK6l/pt6CIk2MJpx8pYd/pIcL
OQY1DF82NlMDRcCtR9Hd4F3UwwQGjCfwbonBUXeL8uy8toVR60bH7hbCkTMGdKEz
+YwtYMMhzA2WAbGs5neP88QEUwkvzCxUU4KzYH3+KbThSSyce25zgAIMszl6jAsD
efakVItbu/p/b5SVu9sGQtp8DTJrTbcHu8+/Nptkoh7QECf0p8qyee7kLWP+R/5d
ijFmV5ZUjUQBj6pa8XcJ1oGpHVb99+JIMdYH9G/ysD/UoWzEshgajsHXnAS9SddL
njW1v6XrNB+P9aTC/YJbTgGDwUSVIt0CWCDKE6Wp6iYdORdY1DHszIF1ar1WFCaD
s623JeedHO9qJkHoFB43QYb7AdZylCAF4XRevPbLjQFQAejq5mqzvBNnk1iHySIy
9lfyy0iH4jvWovGSFn9JkjcI2+Fh0uO22CcvcqRAUxqMkM2tDhR829ftxwyBiZdq
Bx+VwRJSQM0K4CZEzdlzzowg/mDuAt5O3zeFDwqQqwrdpBZRzc7QFr8SoC5G5AFe
rUwzZ6W3cQ2vwz9ptAmVEO2Bu0P4TwF64OJKnPJnDRZxNBamUA1fcATRyaLqPwj8
7bcZsxWWdfT+O/t4Hq7NOiqdRuWPdXm+/Sj54Zvg3L90LZKG80XRv8VJ4c6WGmal
zCgyn7VpXVWxtEXOG7Ea/j1/GtGRpYxUB2bjGULPz5DLMbHRJ0zG/+rzn9u+vPEX
LwDMY4wcP5hul3U2XAtQvYt/ZKTuNl+k73F3UNpi+5tu8665V/lQP65NKwlAe7kE
9JY3l32/IjSBr2n+hg/CnxhvzvBt6aXPGUalQjbQwMqlsSeFE+aQviU1ha35m3YQ
2C2ly3+QV5xyiN4HIoDVZjklXRp3C4FwFHR84wY9m2cQE61iO/3Hj216VKjJNUQR
9+Urj/PbDy2Q/dPvnkSEM3Uz75BjrowZSHNjyCULfUkSudDSi7sGs4HcOl3o5GFU
jUli5Kn1odSPmsyFAc+5mHruxkF+ImH6SMe7eEswxEOGXYWqdOPZaXdHA6AHIFkO
98GzJMcufLRCqC5U1WQ3hoc0R/23lSgheO9zYFwSvPdODdGEeFflEIarxUmAVjCx
QN2qmlNZg6azXHml/+u2s0UpizkAG0Io/MFEHB5EcKEuOeC/gFVTfdScpR6ylwHk
ViwXCFIMG1Ee7ObRIIjC8twqAiVe/int5LxzDcFiMd9JCKlnRbqZBqCi9XsqPBey
/f0ftfhaIXgoXWUrA5fAU2hPtHEXxaF8j95EdDZa+dUHl6feM5P3OUfTxFZ5bfN1
n/55Fbqsh6+y2rCmyeVs5VzE5XRTwJPYjP2GJBO+6ZlOj+qwdNeSu0u5ILN9O5bf
gLr7plmfqHmWJsefMQtoPz0D1m1p3SNqmnDaxkNCSu0G5PHNUg5Xw8zjVaaK1MIU
r4HAWDlcPO/FYCQc2NWYihycSasiG9tvjNX6nnYHMVM46PEoH4sJ2X22UvbUSmKE
c4ePZCh+VuWHXjQXqwk2cJvuloEXBN1SqcJTIZIWPdMoIE+LyK/e4FZMtqBpPH9E
ogYcXkyXdcH2SvQ01tZg3zInxj5gNJZraYdZHSsuPszVElWagMsz9yD+vP0g0DL3
riiHacKPnKsQBIp1NxfkdyGxzyzk71qZ+ECG/CJNz1jKUxWChBFYH5TAms8ffQQU
KtZwmwd+ETj9CLYit8d+JIHDjOpJdhTBiRJ6MrIIeXfRlbxjouR7CpmX1ccAFntA
0EeXuzXVs9SALmRttOMTcu2JdaQOMbVKaYEk4vI6Tyc/RLRRXqbhKhYZ/SUHS/rz
QP0hkqjxggQa7CigNxwbwVIY+U7Mb68mEAUtxdyCFGkN8JCKNpRsas5Rgt8YYFtA
ZOe9web/kbOR6oRUdLJrCBJ1/X9wQ23hTt18WTjM1VtZDuYC/2NsR/Q7FXdDoRwU
KgKk+ADdGI5Lz8/Hu/wqWu8+Vqpt4TmXBCBawaomKEsD1sN5qGzWg2xf/Q6cVcbR
eK6CAphjR4TEf8kvan/ypmBMSF3F9uQe9EmmNocrk+QvEkkRQib63gt9LD9Ev2Ea
ixpa/V++My5Y3oDGJRRDvgKZe9KDUVeJXWTJuMhRUbFREp2ZKXfUxBkn+kqOQo81
k6wk2g2+7akVAd1gTy6SL4MzGSDW75V7byeTsBT8baUN4NlYU0zbzZoTS2xIM5me
gTt3FiU9qyuE02y236kJXyzMH68si0hFOIFyyOx54bXfEh8Fz87wGlCPZQzqYbzd
54I2SmXqDqRxgoMlXwemGK5cduaFEp3uiZxWo2/TITXaPEYDh+CcDorUg+oN+Oyl
+lkN5a3t11LJG35nZSNHjd6BPjJaWusMmPi+jVkidBI/VEkmOJfBMLXXTi6NWnrz
6/7uNmz17r6y4GBouS4S/5O5NAlF6gPqSPeeoh6ka5iW1TLndcYJQlrC/XauKgJV
JL62N9Kq2lUZPqDouoKHkWavV4scqwehrNCgP9peAspv5tpGngIg5k+aqpGH7esj
XOwC/NySLmod00+I25ZHc6Vd5vgjY5BO9q/cnP3/pqquFQ6gSocmGQ61CHX0GARY
5N12SDxIwCU0L+UvSUqUG5ieLsqaBhULjRiDIf5AbOUl7QjuSV6AYEFc9KqeIywl
z3kI5rDXlMJt7OaaQclcOhrZXjrrevSKxu3reyB30iqGqyg7LQ/f5kiuag9fKdkk
KAY1dICbChf2rOgFsvIdiS+buxsstWl5vBwuZy3mHyk+bTD6h0/XatA2TuDb1JDo
FCZug+uOdaaNUbBp5ezxdCDaFZD0gvvM99E8UJye3H5UF2PbYEQpIk8g4/lfDLyQ
SjEclifCOX263mwy/++LZcI9YGWzyItNkX1AVVOalMO+X/3ety0YtB9JsLtFbf2L
wOO+ilCLXEKT8mm0ox5OS6dAd0LAwYX1HDNavTWBBkVsbBRBSScGWUOP/o6OFfsM
JcYLN2VQVDQzXUDSpQWhCEj2KJf9aii6Z8WcuQTLTn+rZTfQgJZ1T4GHmdeuqEiu
7+U5d5kLt2ARieZZYuTU5wgowCq7fta9cuebMpGAiSNqWKK0dr3au6Wlr6Vnpmd6
1KgNMcitUE5DxK1TX7akXaMXjV0CUA59QeiNDvp4Fu9hfHoG+dSXfORL6LWQ3TSC
qyohPpiiusUnwSldmZUITutO3bAxubvPzxj0PfcZ5jYK2PLrAteKtgZ0Kl9YKGD6
8TLR6mhpm8ZovSeUrA7IU1W+lVXFWGunXpxzNhEWsKy/iSLIYKS29MN9ichD/A+S
Q7osL9u9X3s9ILxAghf+WnRLZlI+SXsnerv+vO3cbF1A4/8xIivpF7k9bu4MCica
7NX/5bR7TcXUptrz67ImeF/oV6NrCFNjyvRAhUaJCO6XWEHlFdD91gcG6pOBp8+j
DNhPlhjYUehe5Skm+D/TXvr7GkWzAMihQUwT3JwJbbJ3JZKrhWAoMg87I1ZVFlUh
IlrUpLwv0HUXiQchnDxiGAPZHVD2MU8IHG5Lmcq2rn4Rn3IIvvlLndBEn/zkd2Dm
4eCeQMk4DrocHcGBKKRiE23ZNSovEuurTTOmPUDfzr+/hsoQTQgz0A85ciScmAaL
R8fWdQlEDz+fqFTUDCuygmbDUb60xTCn00Lh1VcUV0UQ3J4CfgVd2YOcT02OZLbE
UpcyvN0EW+jC60zLFQyJqiJw4a+x4Rqg1mXjVZjCr3iIykzlG9SUxBivTApOd6tZ
XWJ1QxLsG0KIStz0GCe2r579Af3Dvr4h/0f64IdgsQDDBVg6eAK4zg/UVWO78HJJ
crSpShvupzs9M1ygD1cpAYIyq8Pk3PWH7bkM4ttVThmHbFQ3UGO6svZqgMMyO8aD
X/xtt+sW4wDNaKYxsfyIevQpoOS/G3KASAldZa1z8FEoN6N44TjVX+gL9AynAOS4
h36w/ccw8cWkEiZSH6JfCiKAsfy3Zwl0qV+xFR+g7orrYL6eM9ZGCE7HT8pXhYdu
hKcjFyYtuXgysiXcN/MUZ0VzdmkE82wzR5Yb0rFHJCs40v30cNkUCQmocDfthu/o
Id14lEnfSsfUYFrOShE8sSGDt22+XdLMK+cEDsj9eFQPOzQGYJbygw9QBOVDSR1g
BRqN/pt7p92NjWcaTjm3inXeHnazJcnYyXWCyIQonVC9/Yp1M4Y9lm5vH+TNWn2e
SrW5ubMLE95gug5/7T4IT1L/cHrLMQYo71Ta6oTrOpBFQSCVqpQdmELbL/23JhYc
NL6xBlkmsnSjZuKJVatoUyGxGjDyZ/cyNwE+B0ckENjOkg1xVtgAA9L/Cuv16SUi
ILXoSlX1Ro4Vhy6QyK6FBqJWQlqFxIrBY20lW02loO+Ko9At32Npgq5cs/WHR3lY
TmfQcVQ/SSFskMdvi8xDmKwPwEFDP9xgS1bDJkPnQU4Ytv5DNpMIJo7ek5yW6/rV
IOZahPxV75Yq6lxMyEBTs0yyQCdQlDVlddRB4MWtTK1l79dV975SXG1QEorJz8p1
7m5nSLYDdO0tyZ0oO66bQCHcgHBVIDWio2jmIggQPmG46KCWEyOiMiwjJwOAaHTP
LSGvagNjYrqV2Vcv4/RJrOKaX9E/2EUIxmMIbSnzDbS8WDO3J486SX6ZrDe7LIaK
o9bz/I7qkfinQu4jl2rwYRoi9A91Lx69N6TYEV6KKPt6feypEaQu8Qwur/aXFG5a
d+KUVUqfq2ynxWD8/yA5lm1eyt6VQaVT5bBDkC1C1Mltz/Puln5oi6tt9ThRyDMI
tglFFX+zE6p55+Lszv4/dJSdmDmmTA5N2krFeuu0GghZYoP4IMaTchpPZyiLJgll
Wlwip5nKuV2j8axs5qOMzcXptQLmaDaqRUN6G9XbA7/wOz59D0W7qSoaHTtDHCb2
QOG5sLGOexr8OPFkVzMMRpL8X3gUFvbAsYc7zwLpbKWK6/hYkzOzJDnQkSBMNO1C
6ljhu2vg8ifD26bzRviMSr7EESoByBAzOFFkWDqsMvivSswOVIM/57IjJb3DfgWg
LqtrVaXbxxQKdjzkJEcjjpo0EGnzD19gfaNNFAqLjODpQWh+XIj1RfdwNep+hZ8Y
kcu/NYqsPiOhYOLn61mIE/SAyxQ8BXBhYpcHABaUlTtCs1RoCWatrAkV/YhlxS1m
GbWnUj4dViRKorh6u4Kr/MKS0ksV8pLRbC5vhVZWBWgriQmOXFABwawSqd2cUBtD
0zPL9jM4YasxSxE8Cz/yvTHWmKSIliv2RlUsWP+jTMyAsUpiSubdxuI/cJUfzh95
5rq7tGbJLQv7sxMH7VWBjVZFKm2K2Yh5IjDPDYAqxxh8/xg3TH6fOfqqJ1x826vh
eSj3zXn8FkT4v095Okj8Pn1OTnDWdDMiaqS0n3CrHjLaSiOkvVUdZf3WzWpww/My
BSpWORNuRtrYeZvVhN/gl8mJ7nV8s79wZBUPKhlqQj5W8tquxFvGUZ0xHyQA2/Mt
xQJGLgqnImTtKvQN/7jr82feC3aTcPL1f6AabOhmnv+vIyX/5qivNcPrJ110nLNo
tBd13KHvjkZBktQykt1cZLypSghlDVXFsQfTwqyVuSgvdlSRUi50lSIrCflxYVax
VxikRA8jxnr6oMfLo7Mk32mI0GRXK86XcHxhYwXevx9QaXKjcnfvOa0JlxhhUT79
yIoMIozZNsQsmKa7dqDA8bVoCXWnuVXFBLlFwMtHFEVy+tmKrqaMKdAnWqR0FyVm
tiLMsz86YCs5AZSenotkgedfbOf9lpegOgl3yzai/i3SfxNjG1UezXkPzjJTRcim
iub7J7+K50z2SCtzZGqoNOwJfVlg8l9y/UbfpbGOZxzeJDaZ64OJ6QFPr6e2MFb1
YS+JqZ5AHPFP4u/zHukXA+6p2tgz7oOCltq3vr4ERWHDhTNbc/GwHBf73a8v7Omh
Fq1evWxcY1dmRz4R1bkU2Hh3gb4FikQP3l8Dmbm3SH2ImkbyaSPUNNFAQCt+VMlj
MtmEOQVA4uHfa0cmGs3shQtcElkoDJGpGa7oYWecqzyrLKG96Ksf9lmyukrYOUhI
BDM7PfhV5m5fJ9bctqwMn3k72xR5PMPiL1IZbi+ILN1EZHLC7mmNzYSANoBXEywO
0j3zjAVe6rlxZWAE0/fVYOtVZ34SOVyBVk2L9XUKx6QQ4zHo0AaseMVXrGlqwAFq
6dvq3sRy0fytJHQcHOS5lFRmbMdOcIKz1gZN2cbIzhSOmc+XoLJPldmEtoOtmKYG
+bq9nawTHwS1ns5vBq3vSHjtlazA110g8YRZVK41JZr4sUr0IXnwsvphle50WIAQ
eWhA4S2MOLJvUPgsfhySI2RtBh6msatTJSoWtLBArh9RCmyujg2nnKSHZRINxqW4
XrH4Vmwp0i6hIQF+HSESC5YWzowyJvqIYaHC3BSa8anpkTd2Rd/wS/EI7ZsFxKwN
GIrV0JH0ITZwpqofNyamtj2f/2Zxxq6OIDlIPyveybvF16iLz4VXxpTr8zsx+JvQ
VuDffcUOASpLAVm2T7aYZ1xudcdhYF/HFGBmPDVj/GfpV+xHGiVpgquZ5MsNZhzX
3E72jQa/pTAjS2L0HMWLqFraIFXkU6L6BVBQN3UD7tR8V4WsScIPbdDbGK2bVK5r
YMjgYSk2j6tzoSw0Q8nKHGoC8+KZqqwp4xe/0i+2cxVpCpeQ0CcpqzsUnTFW0sL7
z6Cr7gtGi5ShW6ODqCoMXayCkCJB0zui8z+0lQ/5oYww0cW/rGNYIboVgchwapNZ
2ksRAdVCRUsdTQv9vydQtm/x99JsTSFzuAgPQOa26AMldp6s/PQxES6m2ku1Q26B
JLiPi30Udjy/D3Jjhyk4LvpH1Ws6pALmeqHzLyu/ndJu5rGcavkHDD7n8n52Lz6S
UL411ZMW2acGxBXydL/d0s506MyTsvtjhZpG7fcog9E5/NQ1DEcW1KjD0XIDdWyA
ONvBubq88tdey69kmdTURTGeVOOPnjtvaqj+DzH/icEqP49zuWFFhJJQZy5rfo0C
qmhd9CUcdFP/sCVZE8EhWHCdxcmKxb8oN8HO8EatG32aFor1xkIUmPlfvRGIqaFy
eotcxe0ZDoizektEMfXATho1d6TjUQFzeXOVooaJy3gd/CN5MuK43rETrIkux1rI
8pFv0S662BeQxORxW1YIcuWlVl8zEHZm8KwgMF/jgp3sCmOt2cxs7RJwYtrpus8l
vKbd5ON7Ot3z6CivpPCMH9a5DPJc2qqLtGDiOzdtaeaZx4TSWKHWqdsF9fha4Jvz
38MzKrkUpJgUZ1U4kQ7E2CkkXqr7bspvtGsk37pshGtfOcpCMzraf4Pld6hKj4iY
u0GBSgrRIwKMhb9fSWXiIgrVZjohXR2sBHH3XH2FhdckKBDfhIbLgFsWkkmCFT+z
HL3Rd5T/gvPW5ihwGYqqy5MtNiHQ/lC5EsRAYF+uvxXu0u/0ESY+i3PBJcVaYNEG
gcYRpIl55ZZOKtxhbjCgkBuQe45kT7qGP/BPP98CzQP6gATa+jmCnkoXVWz4bRZ6
y78OeUCstoyAHfVc6JwMPx7FwNsY8xteCSL13O4gHDoagjIUaGFysSUF2xQly9EF
aftETCzlIp7oJoNc3Ya1/FgLdVlIZIUz5oLmwDa8eZwvTd3yaV9KmMvfevL0+g8g
vpR3vP5ibzhLfio5O55YOcZdUz3ysAEwEz5wmCge6UU727V9ft08NvZnbujrWfFL
iB1DP8lAEveKFBwTapiOhduS2HsQPV/bXu9qCnG4oH8EMAaQo+enDTCuzqB8bbG0
N7dJkWJ575iUl4qneDvx45wqC5pztGI/VX93YjXJJJlHPSmMOyj42NVe4MWamb0M
jsq6fqbKHggljXj6pcx1EJEnc39JSLcZCB0cLckMzJkaJ9WK1yPLXYvwEyrDINzc
ZLahNdkeJVtkfnjWlyziU+p1rzLBrhoDiGbFzd9tExcIbyBPyal+8xh9SNx8JAgn
3m6Rue1Md4SdEPCBGsESfSJLBc4kd+iU2F64inp8UX6+CFQuTBN40zmRdPIkY1pZ
qbZtzfHeG1ZsSCT74Fa68KdYdwdvfR8GycM/EhWhOqEgrB0vMhX451gsB7tU1xkl
whLBvzjxF2sPvz6Z05I5CeCFZr6G5zQnD7jW95faLg/L+URf9osWbOMmTsex/YuE
N+nQ/qTDjq/qGQ+Yyz1czn+CYFsGN02yGFkWBIi6lyRpa8cBTZa6m0Ced3iu3t6k
LBCIfHKb02Jp8SWyQkleyBDDKaF9xR1ryhPKITcQPVWBhKXH+Y3LtqKzLWqdh6W3
ERQOfO9Fv3CD7KYceVdoXJXOs3bmJTHvSiIQf41zM7uKTZk1EzfEdl9VMArDsIQd
KxyHMh8iVTfD9MMQ2nXcircFWUsbRnR48/vn/afyL3h2fMYkcLWaMxfFf7gGu0m8
jL7pHTJv6ZI/bJ/3XCsvDf+F9BjGvKxgfAl/otg3qB54MwX8V65kDUhSxk7nJMpP
N6GdSHADAijJnM2tGBrOOOZOOs8nDVh+OTqnbxTvzv2jCK5f5VUFNtdvZDSDJTYH
7MlB5Pv1EUe0ODKgOqzN1MzuMuE6RNcuaT4F4y2Bi8+muUOgvfJPnUKqsICIVvNc
Yo+VdAyExF83xwniHDFM25ZrHB+J3vXtIHJjagImzgwusUSVcC1cSHZAFlJx68HH
//Lfd6+MFIlz+Y/TuKUPP7PcaZmVnR6Ww7QrZkCDOCcL4rWrnQRFMc5T4UcPRaOy
2BdQkFIKs0qL8stVYw90hr/UdWsTa5ehSMcwD6XZ+XRf8tpCWFQW9Qe1km7JcPGS
lq7AuaZHjAnuNW+zLeFCjrNeLMmGfAYjT7qXZebCX4SqVqqVQ91YGkJ1UMJyUe53
S1ZAXrqqM2+FUhk221VxKIqeCeavIvrJ8VSfPhZZIqM2HdlxJ1+eTDS03ORXZ5Cz
UywCa/DRIgto3Rryv7zpx4kpF0ONWiHMVCBjaHA8ann86zWOyvofwvXTJtVkiXgY
uMinejYB7AF3s0ARyAGpITvqEi+lEn7asjWd02rLNhzFj9a8nwDa95ae0bLSm8N7
JyJJQCbLGwINSpAwyGGOqXiJr0kL02pesVVI7cSzbYAs7S010Ihx2pKYHg8zh2Rt
uy57Q+qJMYZZS7c2pm8okUqupP0p+4uiwyVxO4Q/xAESr83nY9DA5LWV1dP20mA/
QDFrSIbrJRD5v7TZ/KOZ7FtSmeL83nIgg+RVU551J+glYP05pz9VuK7A4Tj4jWut
Wm6i1J3JWMAOcFX+EwNMzBoMBBeN9s7EdXZpPN9riTCdju5g8QHxNWyPill60scm
wPkOq/5NLdCdKeSLIcisgBXrhKBxSapPNjbHjzn4WWhYFiSvHmRKinEyWFGZh0Ld
MAklcU9xapyqo29g+MNvID2R42JXkb5tZv06WRWkpZ3biYRj8RMJ5SL1+Y6ldrs8
Yii9Ret9xNPvvtzDWLzpQ1EezpXeJ6aAneWZUYW5H91E/+o8Ka/aw5TMXsZ9WAHD
XmfJTSF4Duple68C1Xbg17fNj4G+PkJ8Hd/4Q5VbVM9DwnIhDkytVVzC6DSfIT7n
LOBXv43rnEeDhvRvSeiAFpOS4cq6e54uKi3NnNR6UfdnDletexdxWGOybnbaosPF
pPFDWeNpr0pIRUVwNDS0cSC4ZVb+5tHxcs3MNnAKpBq9Tki6uuehiAJzzBhqNxOl
FwrCLMItaCyuFo9fJFCG//JCc0nEndSDq5NyE/RBufzGcQa9ZQHu1lCfqWK8hLts
PpyQp2ryA115CfIHfz8T0B10O2DtDGAGIRnWg1zM+K255vQ0txc03eE2iwsZTf+O
vYngD2dR29LmnKBSccYm8bEWBkzbjYpBKeA5UNSfg+ocseW8SFDNu8WwL2cApiYr
aa8x3nwZNPSxqKnl1zmkwiKFQSqJ58BR4zeLcV74H+4P7SF/+U2TOroK9jXPPjta
m1qP7nurMz7u4Cn1S7miaUacsN8xzq+VJ95XlpZYuC39u781IobltNU92xkGzMom
zUw/tJfcbPJQqpri+QiC/riB6hMxn0BGtz+rugQYouZokoZePQkpFfa5jGQKv8Yg
EzNSbhPAej1odF/h//6HBylEQUQT+GGEVVYBnlAYKYp93ICoia9zhuR8A0wn9f+l
HiXKlPSFAHQcqtMqwL2nAmmCWOi2ZbDldEzchEFGiNK83ib0Wqd38ee65dWxfDgy
zkxh+UXjGG5D9jlR3MgotNLTOu/GL38z7nRXHBwGSjbfbStbhqLBkFzcsjCAmzOM
ovVh0XQmT65nxHmMUfTCE41Oy+B8s5fzfIkq28ITA5zanQWP13jYc+yVmN3DIeiT
qrAlXyDvHsleCLNFPDo0CWCUK4XRuJPNQKfPn06x5HOr+XFTXF2N+pOcaRVRh7bP
AdbPiHvTJlSkDF8doiXQeqr7ZLKSDdiV3s68j2aXa1S3aJ6P1PDXcDAWQ88owUn3
d3MZwfjL9UFOn8nOd+/hFfQJEgRnzxgtD7Tl4z0YbRMBFhw7A4YjV1Hg3ydW4lkm
mlkhTVPCaDAsK6PZdkZW1i+Y/IwNvxRPyHioMLi6X5PAbAuJ9iBwyjVMJr2YfT14
I6cxirRpch9N40GFQ/5vWr4PytejijejLcfISVNzYnTNJoI4MkVOJbHkz8iC58Lx
SSq/dXvATf4qsAm9/k1MnhZoQr1Yh/Oxuhm3uP6XJR0rnSXc5LfWaPazd8hmX8bc
Q8WDdmmasP4ouSOBQyt34e7uu8Wnp1P46mJ4rsK7ZgX00nZEgtBNVq/CFn2LSgpg
e5zMauOM32FrHVNeHMjDFpN0ME0/Dgo8v/fals6EWDQvSx8IoC/b6be5t2fK1UOo
cQgs77Z85P92/MXNx1JCdjI4JmLoyeb2fTPwlwt0LsgI3EgpAC12gTZHmWNAR3Rx
YdeIxlDsYOSmWXKjRADnq+OSGXSJWINqDBK8oXieBFqla5gXB9HIddicaDgt9qnx
0LQtvSOG8QtEWJS5jq4bm1mJQeL7RCh1JDxQbm5M4BGPczA0V8lPc6zdcMQbMpD7
M4MJ/L0f6aO27ydX5bbzgrQqk9Vo3Opow4SHh1xprBNjTafysNFdOlNY8X0sAED8
OuK+mdlqeKLIkFkkIv0JNXxxVF4oLPSPhDCIYi6YKFQvRwOY6p3QHpoDyDHsnea+
q65J6aqkh2DaHcPy7HWjDcwCNjA34Ym1sV1z05GiBHH6gsR34zUtoHISBQQLdS3A
9op8vM0o6pddNFHfkVeFXMbGwW3gT6dicdNo1UhD9HyRuWjcwnWVZJhdxyhGxmR2
3Ye/EUuetH6OzsPXka5tcsBN785M9aHVSzfV5lVM0ygyjaSZau5D71kO6Yfn1lN1
mh7Hut8v9q5x0rMhrBdKEkOjM9msXCi7v8Z0bJ1/YK3Nogl2fuLvhFafwBPs7eIc
SXI44NNX16QxGkBO3NlenxPDqDFvvZeprf91n8C4RKwxu717Av6+MnoZAR+gVl+a
RbeRjboHmNJJXr1Fyd9J9oHwWQr9P1CA4eS1yZmYTRx0vdHZ8phOru7hpJF/7X9O
eLNsd8jbGZP8WkrPq8tpXXZXVfGALSlwqcdL2xRYCulUhElZmNAtd56QqOxZceqe
uOFXlq8OhyvgP+yVKi1BlHy1+sAhTu7Lg78bmnv3v2Yz0U7Ao3vqiYLVu5WnSwaD
5N3VnAs9YPqC2qRqi44BjUQ7lyk0DZyp+UMx9MDs56JEfHAZo8+BdQzgKflgJqHn
G71d/51Eoxs2jKuG3eqRID6wMBrn0KyzsfDLKAJuqC+/CcTVJH903GM/R3BAE8g4
oMukUR6P8NQ/VQjLD68Zb9pR+Q0KjnX3OItkIUDg3TNud6S0i+jvzWYXw5188rBe
1i0rqccY4kKcZSdVSAmD751dg1lRr6BNtbt3znYzpwOOouz1UTxq8tqJb8Z/FXpY
cd8sL2Z+dOjHFkYmAPrf79t4jqeJTF8xYtJQjJRPCAqcoEiKM4nGd80Hkw1/eqk8
2wqmDn2TOopul183eMAVvKKVj7bnAb2IiTFanWHRhe5QRLy1CKLdZvxIArCq4Xax
WCrZrV6Z8o4H+klqPCBhTPRp3Y5hgniFQD95XcgOr5j2z8dtDmSCSBGuwy9I7gCC
+n2ULmb3ZgUe6Cm1bFFBX1Km5M91lTyeu3Jxmel4g5m9WYJT9tjdf+3Mk9A2OFZg
kCVJONgMu6be2Bf/PG4dB6RLTD7iIpDDRVFMr2KZJQLlyjx+0DkY4ZVBWFHc227N
9KjvsnStcbcLVGKoKgJuYoibEd7muo5CWEudQx37dCMT7of68VbcV1X7tEUQc4HT
zcHaQc+/xTo6b2KMA0XJke7Yh87RHLLqV2EsZXIwGPNCG1AJwe0uAdUJNBkthdrF
at6iMHYPne1O+NexxSYpUi2bwuexTtroa+d0m8z1xeKISTN9uyZo0JOGyZx254iO
K6y64GwGKcz4AOjmvo9O4kPppoOlsP0wIP2q4qY9soOJTp3eECTyRZrxCfsgKkNB
5x7Z/Ptcru7VyDEws/Z3DMlSnk8Bcu2HBDs5qOjMHV/HNMBQWVx8d0V38jYzxuKt
KaIkm9yxxj/t2RZc6f5mIYgnhPtVZrz8mSLCZ/u6w8KhrDRRRgrmNQh3BOPycezn
BloEZD+W8tSbJZL+0UoiWbUls936VMQwCYl2mUXbmARSmUZXea0w5oZ4+RMpxNvO
h2eWkqXlTb5zN4SVhE1PR9vsaSElcMxXL8ACjYLdDloXOsAALlrfRp8BXyrGxYQ6
0BCGU2aqMcJt+AocZE/n/44aMnWPlYmWrhwoVbkE46o4g1Xci1qdk3/2ejm9Ufbn
bhyWzH00OCAnLp9WYNeMtRapstXgGagKplRbP3T3xGI=
`pragma protect end_protected
