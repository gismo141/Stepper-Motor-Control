// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OS+kzy9mAwAOlYzkftHJFcHcYSzpNDWoq6mnoNIV53HsX/l7PfO9dNEQhv34dNn9
yOUimcfuV01GMZrIG6Zs+v68xWPKXa97qIGw5A83vtlXttEnl1kykeJ9I60rtmaF
3FiWik5j/TVlGwo1B2vzX9T3SCw+gLZD/oP2wKCniDc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11168)
q0/EVxn+LuxY5QndIBXZrMmIHKogcPlMe/xszL0QJ9+Me7tKOB7NhpOhfwZhB8XQ
GBqMQ25VGT4QdLCBKwgy7R8knSqHyxBDq3Y07p8GZMq6GDupSfKay6Vc/9pxv5sr
SzTCs8S6yUG4nTQC7E62DdEeTJXoaHc3EBMD0kAOSRim+kRXuB7NE+PgKZsx3E+C
Jv1+BMuEeEG3sc40e0PnXRptk3kiWZP3nji2bp5b7zDvR/2csxEkAYguB5YBls8e
Mn1VV2Mi+9/VrIKbJHVyPWD2WrNp5UnFuKN+pbLhRvjYg+joWQ64p5scqheIau6S
f4Zo4SHX5Q2Mttz8CdAHQ2vDehKwn0ZgchYuGAemAPn8TsQEGAE6CuqwShV8DaZs
vNBXiA18iQ3iEUEOQIuVf1d8DtDhgdLs54+GDAH9yJswDgeXonPx8KcKR4Ce/Wfy
rF9qwQvwcS1wPYW9tRA/li+O+uRCRioNgm32Tbr2c9bIZsngP2P57LdujhZFf1iu
b5jxF1bROWmKYQXM5mYq/RTdVBQnfXvmRzCiCtWckH2YzPNPhVnPHSGkrZr4ml31
K0x3zbIq+bQBadqgNvyzO94HfxU7qLv7fZ1I0pSa20c1QCjdK0FcMLMENwXDG+Kk
7I2TUe33jdtvuHSb6fivkKW/jec3IuqijpZZAB6L8JGfScav4zFfzFvgPBFyT5QS
pzoh3Z2ytTyk/wV7H2LPyredPQlvGqyH+fWa8Jk2ctBWACR4F91IiT5sotU+Hwzl
wnuokUqCNWHW4NUAApU9sxJ2pMwR/O3/2BfzQ+JxN3TNVf/w3XaLXwjtvQncJQdA
3nUd1D/KI5APJdDtWnQT0X2xaQ4QEDenrGD6cn4dlv0RxNkmd9kBb5eZ2O6m1ChF
D0rtB7LZWE3g/zsEDXF2lntuwTpR0J7Y5QQcbiLi32/TwMRXR0hF6SwmMqWHiMd2
STWa4mh8P0mLRpCVhjyu7or0v7Qyw4a2ILdAgxhyrfRDNwpeIXrvfAS38q/Q1tWB
wm+hdZCQrKG77tP4yhQDD23Drk+dQGFmtwaK/tnmfmmBwkGFfoT05IzN/hYQ7A2Z
xy3nHzkMLMfnTz4hDZd0N01xhpx/3C83hb3EX9GASVvcTfdHbIme0axCbPibaWQT
pQQzgbzuDWYv2GGTacnoppmwrdpS5b3BR6AlvIx3kyms52s1KJ4xauiA9FY6o7R7
2EqbEoSRr8xlwR7kqoEsOOjtl6F2JA1TVnzfiNtKG9jBhAE3TBD9IEWkSGlXw1ua
rRnQsMfYbauz4IT4y5E+buSpghY0xHhJeIedeVwcGP6Xq9h28GMHcn3/I5Qsvs/K
7yXclfXcFWLHHwGV3oTQNjmKR+yk0PL2mFbCgrH4QVNGIi6+xdtD350DY2tqUal3
wOfJuvW2vYW3UYFt7BAzMyLLAerb81xMYdfOziUJkFlmTlg7eR98uPz9yIr8jc2J
qJZ5gb2lS7GxsMbL9taoTUhcgSA9Ob1fsZPh8qQDZFH/Jp/klNpNCwcw0ag13/17
0Rtny3HU9HrH8AdsurxdhX3bj1ziSHFpfoQdUcFO5HI5iBiLGFHmr5E7Lmio7yi+
f3lNi/4dgW0UrspPsI89joDLlAfhSF9KDNiIbI3prabvCdMTTiRLqRDCwpnVUt9z
NEB7HJ2gRYZcI6iEiysJjdLAN5fAh9NbKSUkxRBhRgHJRfcacvrFOp0jCl5PRW43
cEJB70g2tsPx2V89Y/tN3ll9+tSVU6pbTdcSX8mvMuFiSkbQ85fOoLgSK8bOBY67
jNvbu1C5bMWUDuSI+TP67lkzmXkQHRGxYHV4LufR5XCNy2a90wAxlwKyQH2ycyOm
+DDT4IRpobN2RmYMlWwmRuvAlzVMlyg46/b3oT/d3F9ROcJ4ScVWAFTj5Pw7oM3s
hqTSUoq/9blK2z2uT8LFTvdNnic9l6S/DoOalD0oOzbaDQQ2AD/eEwTtht7LuggW
SYeM3SZYNoYXcjQYz8LTFlGXcNOCZ2OoZt62y6HuGAFD/6JcN3XA51gCURbLKYJP
wBFYNaC3W1Bypsym9nJMTyE/VQYsvb4qic8BATlnFBXXpMJuv1kszBBLHVYDuKgC
AjpK+pMVHFfWZbhCKH1sISDoX/dKCh9rU7Oe7ROKqxQfRu/zByOXCMlrEDzcpjKa
tY29pp9R3qMd0sWrj/0WFlmDZGlhahrkumqPqF7nYvETHJFzvAOmxopaHhRIcoVI
WEQnjv1EUIBpYbH1pmS6BLyexpyhnRLMKYybU0kIXmvJXLd16Zf0BZPEngdQFXQz
K858n9BRev1JfSp0LQRU4l84j89ssof8ZkS7cKtK8RE4vGbvrWl9LlXsoz0FJXvm
Q2aaAnZMAlWIJ2r/y3t47w6IDN7GXN8tiersw74qvtzByVIOtGXtZlR96egrOhgG
LY+JO8+NB2OwshBgxX0a+RDLhhElKt64B1BXlBvpTgcQA/4rDdvfVB4HgUwR3RSH
uIGhmnc7jhGMRmjh4jxuxSOu16ekGMnC9V5dftyIIOyqZQHn8HufduMuwqLZT0SB
a4BxFhQraSTS7e5nvJxbrCDpSsZKR9uXnjAzY/mHp5DYyEbLqKtLXUCJssmR3UUu
4cLoDTcff9WQFC+WuLDe8ufiRnvljVXmQaHfkaU9RMluVreQJhePr7btL1QXmNAq
AAJ3ZehzZGX5oidFm1OVDy0dcLCNVu5cHzUIuwqpFQxYFGCzVgVGLBgmDPbSVmNW
054EedKDkVPZTWqO5GN0jRSrPEsVdmeJZ1KpGfYCFZlnwfDNQ1LF8dhdhjF17/pK
DrXXoJ8Udev/I7vejg9WjgbzdJq4+eepJNIQs7taWuwm1IqsZPzw+Mt2Xdi1irAQ
jreorA52eCla4Cr7dCvkcy7UxAeCSvEakKpVccoA2+6nNs5PUt68mY9WIo7pqEkX
DMNxc7KYZaQOpcZ9IDZnpuNhm+8Sn3M4/4aVBjG/4F1rw98flb3FZQ1tA0cWKDVE
l+4NfrIIeSrGMeAreHi1VZuE8Q7kcowd2EAL8TN/Xf/GsKeC1uV2uGTNzB6H6XRz
sOT+PbtrH0yf7MMnZiSz41j1Q+r2hoZaH0wDQiQ2CF6/opVksZ9I8BiMppC2DXgg
7xyVe3OKRcRMaQDTSGlf1s4+J1fiGAtI5n4OqNPzCo76hHJO/ME7U/N77iv1DTir
XYpgvo2hip5T+FuL3r0NvQ59weyOsJayp0l+d2KDy3TYznIC+iIHCU691pbWeQGD
2nhj9AbSh5BINjGrpoY+uOsx9mzL1LPgYcz345lj3S7uCxURyUfTM7EQ8UHcvsqZ
8LxkYzytxSFNSsscTvZwrwHZO3J3w2bRE8N856lFf5Py4X9Hzok6+coFN5Ql/Xri
B05Iht+tgqmWI94AwmM6UcaM6gIxvw9yYOSlVru9Y3IMc2Ym4QupHNty4FSyI9Nu
dWXrboNYEpsQ2GR18/mOQWVLd2masf+1+ACB6oipT5YmdfY/OpkHk6eCWocl2fkh
8zWmf/s/6vqHuTlh0PaTWdBAe2Z2kxFoIIIsJTIXbEq+5NXhzZLcJKyA3ry/ck/k
Mvzay2ljntXyaMZUkdl46pch1OHlQdRxhlG/qZtHC/S4C3KX1jSr3OEt6QHUieDi
bAbf0BVQUtNb9Axi37P1N1aKIQo3D4JdSsgBBfubfzFFF7hgxegmvxqW3KtCh4Y4
xI7nfwUjTIYdsqId4l5hJpetTx7wpc3gWmQSxUTjG5tBF4jf4IHzRc5pk0qn7sn7
ibM3zd+UPOMvPvJK1sSv4b3Na+ZNsry9ncI63Jnb3oUAFmmo91i5pD3MfTmzEpwP
M8kSTBCwBxh7PkJzqpY5bNF6N1h5R76kQopHFJyvdk+0OH8Pja26gi17LVPcE9xS
NToCEYBSx7w4oj+bhKif2L8uGx/+ZmkzHCkn9PFn4vNfYWPlrKdMgCgFK3lo+EQf
x3H0lvPflYhNnquYVqltvdRPV2BlUDhImSy2NnFKzODu6ouX+GqkaKbp0+Rv9oIK
s48ZICz2aGbtWTe4ppB6pJO9zJBi5aUt0Davly91GVhdN5Gzx4bSJ8QDTGArcaj9
GJw7TiLSx5odacHIjEuYGqGnh5thODVXKmN9wGlKkK5KjH6ogpX0/leGPdr6Mcmq
BnHs05rifsdHB6x+UKUrAqQlAlf9iWEqVRCvUp60EEsO2xsV0xXjO7Vsg6ft6dCw
HJKlCh/HVcD+Rqps6kjyqQQJ0wJFwJLRE76mAdeNOKYhgd3OBBOQUeY1oR7cqh++
4bv+wT+7d73A0zTYEv/tHgCuW/pWiSbTMP6sTWR/o89kF9E8og7NfRAaOzimE6BM
UUJz6oLAFOGNfpy2oP0ZMeH7e7ragElnXYHjUDgDUnlX48ROoSW0AnoafLQx42Vl
c8Pd152ELES+afHZhe+ZrNKMmfYFB91empwHvwymmUN/FA6nWElpp+vJc7LS57BI
q97fvEh/BeaYx3u0wHCKlPUfB1xJM+nvadnSRKEg2rkC60ldxFaOZ90GJyFINTuT
cgDqTsppXuilN66j2ywiLtvT84jT+rtzU33ZWMQIPeGtIXSaTClo02/xfhzohKXa
QwIM6fHg/183Zjc/kfpt+iYIGBQIq4G85iathmsQsri8yioeo80c77jHiVB0jtrN
swj/WMaOGGXzQsocnYFK9AuO9g0nGU73TqJQB6qdDwTU3fOb0cECgTlVxuGJ5a2w
Usjz6bvhe989l2OsF/CH2k4OZO/hQpPGLKNXayxaKmQuGOz8LwnIEIXU9R0OCAhU
QOda62j+RaZfUbxYBzLZBaAf9LNUQ1gmGJQozm3B9g62tyqQ1CS/pNek7yOXrZxx
i1pygXKLz+zIIah6NY91CaYSd12MozZy981QQluKkkByiNI6OZB7bJFtRWxZeOot
FF0H+yGantuy0nmM2w2fGQNrFc53P2zrktxKA8ydUAdR+yJirBprZQ9AmPx2TuUx
dSCyJXiwmPuWGSg82abee7FKSF8cq7+mBQBPml1c8lBlnOQQse4PriAqsFgemPGy
6RxnRcO8BpZZAnhhzjdVmkjIbJiE65Q6PJSPMdek103BSYm13Em/4/0VnDYfRmmI
9CvcQXnAHkZqqXecoiU9FtaPxS5gqUuwEHpszVEzx7ETvCohGWC1NywwMcE1LA5s
ouuPwyTm5PWm8Nx7WPVAbpOl14V8hvvyQ7W5bUYQwVx44d+bC2ULM7PLH61H3jW/
QunW6e3yy3ICn4M8nKl7E9+rl7xf/PY7gfprU0VJNDrUtvgZjzQxwbUBo4nJM+hv
nlx/Na5hScqFmZaCgFMJiqDlEeA88ZYIMV8eyaXvSJ50kJjW6xly1FaRMMctncTR
vhthoE+MmMYr+MXHGzVN2LxDPVkpyv3rpOGE6ZRLLQN6/3Y10OvnQqKahjotmV3M
LyOZgrgHBARF/SAsRKw1WabnyuUHcEGdkDYcZNUR3ry6+y732gc4tk50TojnjgAw
8jYDfB4Cr9/ftnV/xKIlVW2VSijMf2MhbfRk8nvZGqHIMl1I/3ZWYTWzTCGGj3tn
EOq/UyDUFp97udF+igaHB5TZuHxUrChxpuzch1nSMjNn2Z6Fu5G2Om6xg9ruUtM4
RiOE0iWKUZEBC7CImFEyebjpgh62U5g7V3xSNtUEL0L0snLmltgcEf13B+3DNuil
1lfCj2yoy72SEsffc6xvPnzStBSQqhXiPXqzRKwu7ogey8rkE+uIKRD5nHSiuuTu
myX/q0ED68v5sggYPx4n4EdkFS3y04c/iXOPD92Yub5+YLTRDDMOddbTDxaQ+W62
OfFRtYqA6T3JuRaoo5X4VR+HetQ2myW1TV9w9xcwB1YgLqgs1PBS2niq3L1d+BGV
R0e7eIqNaDTbtFqEbX+uqKOF0QLwfxLYFw/VGmzJ1oGkU4kh+gqzcXMZBtDbxrVw
9brEm+lcVvEzBUaYV1Kh7b52i/DXnBB48jXhfDWPhls0gfdql5VhQ6FhEGDMS91T
Y94QaubIEKO8JkfFktHqY8ZfIjTJB24N6EXii5mKjGJWDjwDHTLLQeO1t7fjIECO
ar9lkx3okjZfEw113SW4TSptDatJzndjk1OmLFo4itrUCZdPQpD3fW39vK0Zs0f4
xNVNP5e3YdqNbW8RZUIgt0BTFKVP7mu9RTZaa+frwJ1Bbcj5XwY5TBJeO/Uqc9Do
mkDhnnzE4hhOdupXPVzn4Ho4OXR3p9XPiV1/qDhQkaKpCG9ctYffBwx7/2xMzUqW
6L+vEFE3TZ4vvbz8DIZ4PTScG4fkdxuGXpwEByVXTiVpW9RhDPFLlxUQwOOkX0xK
9RwwU5pAMznxLo7uZF+d+V5b3/P4c+s16QVklwy+KJHime7tDWo5NkBv84jHpXUN
CV8P/d94QtnSE7SuFAvN626M23vi5wH/3uwIuRpvoBPPpXzrGpvLSwYeNupXF/1b
wKBtExhFtApLOJVyAZrWtYWeTpSI6MdPZM5i8l7sG2mV1MWb4dzsWrF1RbXbMiMw
wO1LMl6Mw4sKtK/2Bx8qBC2Lnieron0kdqO8vlPMT0txkVEj9BBcdfxVuWkOMvQt
yu2NZnNAoXSa65mYClhMOZP0jArG4w+US6Xkxqo8HY970xlBh93k7Bb3iwHhdyE4
dWKlvJbFTUG+mHm3CIYsSiQS4whSZ8J/MkS1ay/W87LDDIKKH0NRS3wqFiedWBoe
jMAzA16bFzD31pAGNXqyrPEdAYRpBfBNtms5DI3gBeNrORy9sQ2A3mj8msxJMrBZ
svUT1fUn+5iLeF8um3+/pN+18cVBLRzEYwilemfABYXzmFBnZj6oBQF9EairaYOB
HNHSpwl+hRCy9+kkYSBeu4qI34a/G1/h7ByrKLox9KQH44vJ8ypcmPiXT3zC9l59
myOV0hXyL72EHcKdShZBDkQ1ACGw81y1+XmKJgGQnpSwI5cnvYSyefmnClWffNze
18v4nU3lGW3VzaWJa8HqZVhhh1iSpzI2WWCjGO46jCkM7HY6w6F5Lv3CP1Kwdgyy
8DCiNwVYtyQfMy9UT/AckXIgU5MMRP1n/kL4QKe8KWnNnQ0HxYHeqKEwT9iSahxw
q1zEpM9FDv4ZKL4ZqkK5qYu9OSqSwPQvdhzqYxMCgVk8Zzbck8AmHUw+vI8X+Pfi
krZ7n+nG9zeDIeRlxuHQe0WE8jpV0lVNFTDgyzqKTmVST2v5YYacdVKZFswouCkT
em+M7s98dCglIoqtPEr5J/cy83/QrOfpa1DJN/JuxQkBu29jsg6+9MAV4pMX0t+8
Tf7q7pq64quplYlFad5DTsr70xIOVcMBj3D5LwjOEWFpiYmESQVHTJlSjMdO3+uG
9gkbMXf3fx2I10aLgC4SjxW8e4DG81a/jvcddcB1VvpdWUx9qQ6vf2y99RXGft/A
00kRLGgPuwqucxNlOIxrkHe2lxaXcB1T+41JdtHAGB61ZRBJT70GmD3IMvIMtS3t
F+OHoiaKwS/aVnOmQF5syxfyTQyUcKu3dplqpJBZtxHXihRJ7qaoP+qWrZ7c399Z
gTLSrqVtdZBmy2yA0IZGzqR0GwUKed9wqFgNlSpU9V7w8vfluEPhMmhUusPzfep7
a8m5iqQV+siMMllfVF9zY/WcWsw7Qr6WyP6tFT3tqc1DLbWk42c3Ob29NLZgqcDj
rGOibeQJFLfmBykbBgoO7gjk+olt5JMdFFTesKeigk6smJSNZGjqvqHSbNN+Xp7r
PjvhZ9F1A+xYDtQLBCNlgc1ds/aYYxRJRZy/pP//zjDyiYBi/kzJYLLPa3N993Wl
JG+TVPfN+4kG8QqDa4yUTG2H5XFXEUqhitjhxi2SsB4cY0BDEgS8Xc+VI4/Z7xwi
gEM0rcm1zo6TLY646nXH3g0S5AGjqWwyM4Z7aGaj1TiiPi1va0IGbRICqck5gfRn
21APrp+SEFDdjnwbRpfIBec/iKVyShey2gAFhCv/IYnvMR5Xf5RKFdBJaKcV9/qR
2nP7Tl6BgTulG0T2RBSpJ6rQOZ/QYreGOQNEMCx2XoApybk+8d2IN2zLNsVRTNVM
sHE/vSxSedgadw66oLbvxarOYdyHrArcWBUEU1R41HNHmCfXulZKGNYrIjgv7Icb
tgrmfcKU9GVDGluITCMmuVPBRZFn+ljZXVa88FbdicQfpK7300HZ15P26e5l1Jh1
ppV4pt307Yf5C5Ke53R1fuCFEjni51UBW+3NtFFDHN/tqJmbrCpbalz2BMu+xt3o
aRqulyoUWpxftFaRJo7VS3EPvK5XNvsidyzqkUG55sAlTYtD4VluX8qP4B7DA2QK
O3aLqk0MMotev5iBa3lDvreQXa4uyaUn7Et6CEuFT8S/n9PNkxP/FavEpswXXMaA
3+jqz5SEwtjxaJ5bb8ZJS/pXlTGBA7nXyFylYh4uQ7M9kmm3kLbzEaFV58+qoZYh
5+dv8AqukWrnYTFc/0hvSBzLVb3EnxD71oDEysZsdTflDQx0MwF5WskjCnMHTycX
wBALkp1iB9fCR0tpOBsg6k/strVzdUgsZDlf92cSdnEg+/ZmkIPnhOXzthL+nKZG
aVvKbBIhFfJjN23Y3AxeFlOJTAMkvzcMXkp2ELJQri+yTrr2Y8H+kFMqXvVrdrJy
5PWcTM+WImR6uXpKXOjeSqMT24K5wgyU6E1ygSjWTLWxqBGOMf+CBu13qPYe9RJn
k88x9bOesTtFsPgSpsSG/cY5WqYtKm3VDBJCrLNWicU8qftAHfJCVys+5rV0y0rF
buL8FEfPIA8w2kxtutn2xkvgvxYMUZ5tNQ8z0Poy2IXGu3xwQbtxATTIVCh7OCai
PrLZ3j7HkK0Hc7P5h2CRpozbDEZEkAdQEJNHMMw/bmx+6ahDk2BIET62o6K1hxk/
Abs1iq8AmGJCtsxivrPG6TdQB4bszU+eyATZ0jHegFgH4vQqNrWBAcIO3xJmuJf9
cooDM1+H02gHw1/plVRXKSIMS+reY40mttUtuU4555bgBlfWX81LKP+BcsimGmLH
XGzLLymQ7Jvsn6wx/0ivSUSakXyRUQ2J48p49HjKdk92j9jxwVsLOD4uhRTkFSTT
JkH6hDOhHSdXuQLjRn+T/jdt3cbbxWl7JBahjf/dB1p2wNe1KLUmvoNotLP8b0nO
UqSdXbA7qfgt5QXg1z7ZJEBfnOmCxmQey82szPFUUEyaFiKhQpxV4Q4EutJ19vMl
nZvkWSTnitwQwkrZmYB3SlfTTlhf2uF2k4QktZgoP/Zw7fnsliLSf21HTeTuNsXE
/66fdfFzQw4R9KCicAs0XZE6fV+tMEpu6hyLkg2x++oXySkzqb8QYn2S1k6rVnoT
Mm9qXIlMn1NcbghMINJxR9y0e3AF/bQwH5/S1R1+ZD9E8tipA4gSpNuucmwla+Ln
rIraWSmoXT0U/Kc4pfkbepGZ9D8g2SMQxLjB7OxVvFCiLZBdVQxDZdNwtpABW40I
3yNo3LeEMwcwmHVRkgJDg+Wghk+a+xnRJX5H68NPAOeFt5X6rFv84/kA4dq3IbN7
0OLDF8TNSqiQSH7zMhqKdEaok37+VPJ2zO60YZcWYz+vJCnrUbSaFoD6RDP4EbrO
eqdIGMM6aTCR+89RjlQaW8QSAv/fF0dgFl1VnNPpMCxKWtV2LI74XBsDHW8AHivi
fDOhE7TVlEeSkU+w7xzHoWmIJ98x8BNq36tT8iI1uqgxvm526m1nnj51OhlZuRl6
RJP+vUXcWkzqfMmonINWhhAwd+8OULeQjk+4PzK1xOBS5U8Mcn29b0a7KQEIkG+p
pZNvx4/sDOj3foF+AmeE8qiLZfHOLsv2a2xQxubIlUgRloM3Du0zLBORWPP6Ek3A
ZdgaVJkVMyGuVeEdi3/IHXnLGguo3244MnY+3WaEpt3rt9DJbJPw7RV12VkdJOgu
qlnjZVcehxTC2ImKV83VJA3RUvnffZ+x1WQqjbuFlhT+Hu/UvHDPppUPA+jT05oV
84pLPN/vLawyXozRKCeik163N07p0CuhgljOHY4BdwVNuSYi/5XCiqXH4yzTvZXl
LabGsm8Tn+llkwXWAD9NvkhoStuuz+sSWFRNPlj+Ta6xzIr0yjIbvUp+NC+MESRK
Cy7kg+/10NOMkeCiT6YnQTuDMdf6e4ivRcx0DWTFnNchv0Gqme9wjdoUATj+YrN0
efMbhU9V6iTEYqugt9+Q1nJnyuzY3opKy+yx5n6hm53TiyWnccKpOcUrZ/vXOEG9
/f+vpEg8K2OdIb/trCjglbZd16qkPmUU8PsGEArrBlNXm7/eMPu+xbqt3+Y1Zhqa
tkQu96uycUP9tXioaIp8v7WQsKIk9BY1xxQ/ys+Pe/3aUNTSGnOFZGFzl9vQtEGk
UCi6oQPLBkWrdKxDEO+MXtJsceQ3DwPe7WBEtZEWKWf/qNNB2ehXKMlLcQIH9kxB
QtHZ5bUAJa6XB+TJTm1I+ZrztL1ri4qkIfqKywgS9VEKt5A0Q9X8QxO0U94XXLTM
z9mGD2ycfrQScy8h3WDFVhkbxvqc0aDbcWYC4zsAr7VNNTnjBxmxfGFMpe7lcROx
t817vzlfzUbKAWTyHBIg/wJ0FtoW5/X2kN/BUvhuUrTqJgyE0aDBV5Wvq+6FZG8P
eNkTgANN9SHNI5j28yd8JnoO/GqzOdb1AuAusm/wNdlMwT5WiWt4ZPCZM/Nis9vi
+HguOechyOXyfCBbzopkQraf1gcE7sut0D0rgeAlVROACXzwWGVc60ToAc/UkI85
AyQWfaTxmJG3doprokTUiE8ROhwybxMzxWWnkXtVOAT89cS39zsG2GhwaGzqkPTa
pX2xdRPKRWKpiwxuKfn31f9FqazeDW2lcmOgEaPX4ZfA1wK0oT4KDrU15yFSIchH
0ZqpcIbK/gBXn10bB6viyeK2cbe0/lzHQOW5wq1VQf/pJuWAkrfVVRydnBs8SohF
/aa+0qRSVyr43gTkVXctjnTVzALIIGwKirZvwBI+Oye+sXSlfTSUaPtLobVl4tlM
XfG5Nh3+92+O60u1raf0SseebH519nYedoAe7LPsFK2x9JQWXTjjcDR8z7oM/Qae
BofDdzOQeNCQnww4pQ6HSAPhLkaOsuqFYqPcFyiEbgTTMuxH6GLPczlsax0M/dYa
tLpxAlgxAyVecSmsCjDpYcTH8iKELLKItBpQ1m88fRWReAWs2jNisxjByOOYlfj5
iICI+b6hJ/EEQhBTO/0H6HVadxfJaDorrhhtvFTy2OAgqjn80iCic6H/gcaCyY/v
gWQvp15xSwcZX/QkVnpUTHtoZDmPSskL67qzT95yBHps72i6FPoxEDqk8t26RZ1I
hvk/03fTtpbW019G0NxAFEznTYd8N7Oebofk9dTUWrteSIZ0zQCKGii4FpY/rpgw
dwFaGx5Pwwb4pJhH9lhYHK1x5yNz09OBfeBC95McwlWimooml2INeANZl9qkZSFX
lup1OzjLrkIarGiZcbQ/hjaK7MXGtUXDQ6uXo95l9A057R56FuzkuZXlFqZmFXEe
O1ojT1TQWQaEUjZBr+2os6OTop2zX8nVg4K02IVd79x9eiGPYMjhNYijTs5oWReM
7bT96GsqQJ+ydVKm7ugsGRpT8aiFu2nkpgfyGKRhCNpQY/G3FmzWC3ZEVADK2ZHF
YVQwco0GkTV/sRB8OSgV6KjlZ4Da3mwhUrwSyUmK1FnsLCnsPfLs/hHi/TIflIkB
isemN8bcfQZgC+w9+Txe0/B9MlRv2QuZwG3IpOYa457FV7pRi2gF78mKGAwwCA32
OOIUrf6vBkncp9JCorUEb22ndHE+8lMDvpSRrofL1R9Rf/7yXP/KZ1XHCQmt4Md3
VFieixgueUT04ClcQ1PHpVnFXnNBU7y+bzdTZEUrHbNy31uypNSFzHZlYsmO4w9l
+EIvJlke94OY3rP4iEpDgltwxHMuOpOmi/CUCBVFgsoQzFYT26YHo5V8KnIjWBRx
ytV5lFKDQhWJfnkMD98o0qdoia877QRYgOXOMWwyg3fyEeMiDn7JeBZM0Y+52zie
7xO9Sgk0ReLcitiQUqMn4trHK8odEGky4o/OLd2td5OWEdbvGhI4+S6DOBDik9dM
sfGECFkXaBES32kMcWF72QdgSS1gVdYqIY8Y4lN33+TQcxKcJuKyOvfu5AOVqQi7
b4ZsiikdZXOR1/WNc1Rpl3F6UTh5JKcIoJO4ALFL4fCKR3GRpGZ9KtejiNujh/KK
qz3G3+elBdNZBw3Mf+2rVEC+QcLDjNXL9loNsuObFraUB/RNwmHFXrTjZg7F75+O
Apn7wLGqiiGOUuvhLp/J+r07xJpifu04SKthLCtu4TbHS2l8mAkdlGY7xUXA4anZ
synAdFvH/TwHoY0yCimXkcQVSF2r2AOrU5K3u5v4zvi+qNzSgWpooOVnCc8jVQFu
7mgW3v4MqGj17Mh4AdyYKpmkUB6e2fBDT584iP367Wsfcx7cDvihp7LGERDhBOBk
5X20oZ9WoWXUbHadxOLpxeYB7as0sAn5tfr0/mVBXBvxGqLQd3ZUPg/2iI5GGseK
0RM6JOgQbYNiZHkGN/P/Vo3Fqz9mqN1UmX0r9HHafdb9jYez7AB+X+CzYQM4tJPs
tjX06ghcYVS4y9NLsg+7oP7Lj+goHTwZZ8fc47fRq0pcS9EdtZPNGJWuvxFnAdO+
nZ/zhTeDAAgGl4nQZqELvSKLWUWisYGzJMZQwC3uDUSRdH5AjlW9xnyXTSJ0bE4P
utQTtiE/ItIUTnhaxuAjNmMXS30TN/wKo/Z4z4aQMZ2EhaDR0S9QtwsETANz/tWV
RF5eDRnkYZsu7nOIKC/Zf+tIFCPLdANaBPsiJGpokHAOjWD9omoZ96XaW4e6uiHG
enr1ktrNS/1HVQMkpEG+pGAPJFgoysniVNHGJmu5iLC0dAVjnwiL9jfriQ0/LKui
YUgx/FsDCDuZaezTQxqNdq3T2GW+KLSLVZBA8ToUHlylp1zICuh9ZXX9CLsqu8/V
ZF/1yAqaC9UklAGUbEvFDy+cpNOlrqJqShsYujLTZIXG1WEd6UukHU5+4vmuPlXJ
gKFJetVUpNL72rc5u8UxEtRo7uUVHJ8qQ66AjZHU+PC5T4DmoWapDkMVMEv1zFc5
LIaW5eZiXEGT4093Y2S9Zp2A3/tHAcWm2VLwGeXUgL0aKr9vAXG+tFctK2oM1zVy
RiVh7phA1VuDyc0WoywWeAhrcbZMyzHkpb2Z0GUKHulzRD1WjLOReakz67pZvu6h
YQSrowBU2fnPzFao5L4dblVDpkqcwFbB0dmwVtWJrrNZj6aj0HyoL3ae6F+Y+sAi
4poJNwZFbfBS7kb1IyoP//Vjim1T585nnxLLTxF9wHJzoRoy0GDQEvAt+JKovC1u
Dl+Q3WY5Ym6Nb+YaCuIIw2Ksnv+p6Gps/522cssh7m1LcD+BPGKrvP7RAQ3tmr8X
q2CuKF3hMn15dKiade813YlaqUGhQ63pPnKNOtLgqi9gu/B/p99NvrGEkZYVn7+J
ERWCAukyZzU8OBKXDqxx9yA3Os8gSEy19ETm4lLJYpvAR0mdrsVJaoKIfr+4D1Qc
wntoEhUpHYY9lcvO0SOU5007ZD7NDp/uU152E18eplwQJ4XnkFt3e7r7P6hKHotp
xrIszqlhjhLTzy92PXG2L8AdMu8IA0Z5DMBQnqbBWcFXJunXWzQehMWyzFy09st0
IibWZ1Q656mDlgcHLBcX7zr7PAImARGT0Z35xzg+0co+IKTLRs8Xwzld40TxAkt0
osBwZtYRnlenJiZKUh4zE2f7aEKlBHcAUsgBWYzJm7LdTbZWdEDr8+7r4kyeIad0
mU64+2lgCm7Esk90R7FvW4wvGnAF1AakRcq/G3GR5f3JxfaMJUs2CVvG7mmBsrCu
A12xCI4D04spbTfzvRLL6vIL1Z+VMfOCuR8fswd82bFHbeafnMGzuumQGEolBgNI
qkwKtpG2CL1aW0XKjs3caPGkm9a6ohyFTlye7iTQvPW0zmmpEB8/kMZnRRb1uvp0
yFMUBA2+h8TTjnmdbWqY+PIxrB9s/RDhnFBlOHYPgw1qJFHR0RIih9N3HxgucZlA
WvrFo8wF4e3vVdyzI3D8D3AOj1is90FQFHQogRK2Lbafd5KXWkApoPTWLxMPIxJs
HQOrESjpFXEIWZDSsp6GU5pwMwKIrkM4FIgIQ5dhvfWTqSx5Cu7VFvyo3XXtCT3/
vDFlka+sSa0mOhKRuMlxYVcYpVd59cmrAK6d1BGZhxd7SXl1cDtLLaMGz9qNOiJ6
sBj8gtv6lD51usG1cqUj2KD4CEu2pJ57s6ZAo/m0KZc1hclmkZ5QgrZWOFw7L883
IRkghzsFUWOwIrXScoDlfSwqO1cK2ID/IgHRJpu3fsSZ0rlIqcoK3RdA0WGFx4Hi
qH9DHCJJOtlFwYJ+YqmUW+5mpSpunAN0GgkWA6f674bd28NFoBLZlInfc7FQsEIh
AYFRjLrbMBH0wpQLS1UIXpZHBXSgL5pvxZOJN1kw9UNK16lC+aFqkGHUdRe5j/8b
xyeKK7DJmWw0MuT3gTsIz+P56iNNPQxJI06PjzG+yTwjVv75SYIRWauGG/F6ub0J
vGOdEmmUKNT0JY8XBZ3ugUsMADY0YEise9BtW6dgJFh/fUKAd79ZW0z6QfmbY69N
hUkbHt0WslPKOY3MZJmju9oweqPZSh/gAryyQMa7mOkob4uYtGkGSohyGm8X47k9
xR92e7R2jXE0aC47++Drei0GIsvwuVZ0ajquMknLGwsOJN1kr+8DV24+G+mNliMW
GDtr516GLT6XdvliOtpCF+B73DA1yhR3txHodxpu6HUSkvVHVpxKaLRcjPvApxh4
nScpNwzJOlBMiYiBfP0IBuT4RZbo8HvqWk/sK6zSrUg=
`pragma protect end_protected
