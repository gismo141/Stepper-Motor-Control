// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
M+cjxkCSVoEl2a6fr9EWFPsiX76QS7yzFeqzTCezQKDVSz5SLvdeBjkwv0cvvUV0
ZL5LZ2/T0zulhdp6ro4FrAfLl9fmcQfxjHbQlPi2HbwRuMfi57Nhq8UuxvV9cMEo
xUjnT7eA2LFVdr+q9MGUH+ypG8tSQU7i3zgge5StnqE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12064)
MEKO/jxsHG6NITyApWzVIqJYvE9Eo6UfGwKz5cATx/uTIbRAEPYlUAukkPGDq3+6
XQ4h76+dS2VB11lrfXAKodsM0BqebwbrAC/H0ffIXGWM+GMePxUmpJdf6hpZBqkm
t47ga8WBHS56FyH9Nq29ZcVcgvXkRi6Cx/g6tA1juEaKNx0FxqaEMV6O2D9S0w7D
TILPxVL89aCemA4pGKmNdwEk1eZsiXQhv9h5JSFx4WxA0PqJHm8gBQ0pfwkInzXH
S4aLlBXbKaV1a2gYG1wILvPabucTXLef+vwNEnfPQUKXhJzfVAs9TOxu0GDP4Ns/
BxS6jTtmLhV1N1eekMZsQYCioBO36I7RyoYRkM3QdnDQ8w38dAaPCe5Xwu2NAiQY
ROvmrXiPseBJc7MNmdLjidDDlkYEUfenAaeNhglPUQgQ28ODD0tyc34E7jG+mhKS
6D7QPGcj0cDfAPz3lGEDbcg/OXYfBI2ukevZ/FSKCI5mJeow8U5rmv4yFblngoQU
q0GwVb0YjFap+vNLTlCvqkWIp4u+kA4+UOQRrBVpKnQXOAkCfjWej8K1D5/MYVEV
q7u2lyGzRDbamWXQO/86eAsQwQkYYTsRxGKeB7KQeo1+YFX+pI+THGw3uCpUDiYi
Q8umk4Dvx+ROlbMKWUKf2WUL45SSfU2+zJ02GX9bnmglsKVrmOL3/Kzs13QOoSd5
w6P6283I5j8pRTwIH0nKSzYOv/j332wCT98AHEYJg+KuOwcvgszH2LYqA8SyTgWl
2fdujY+BwNXr0Ab19NWOutl42DR0s4+UZ5O3OZjDqbAaEOxB0u20DObxCfujPS4f
4B8zou1Xj49Z+quMuLT27FktdMTKBUqnaeKdykOWJjI6KtWvla34jZls9dE4VFq2
Hg8vwJyFS8LDQAzKv4MFAIrx4Wd67zymw3Ksjrv/p2Is4n8qh8yTDpOciBowCJ2D
funjLbPxGOYm64dwbp/xykIGlvTBJb9WIEk5kkMnHuEUvJ0TeZxAUro9YySnJ/Xl
1dsDW/9+PzTDyqL/NCSsFSBhWcNZv5hALAf/CvVM16wd5wkYo3BMSSoFz8V1EbHA
zG/f4OVsS2UhDpt27Y/p1OmO9rEFXZ6OTnXgUsYxCMBuU7LZ77NnmElQ9J6mi+GD
hsP2JuOZoUQ8k5V1TIteOWcjae38Fqv2fbdMS6M26FppDBUp+La9lcE8qYZ3Cfaj
Ypi5/Otg3gPU9ARTA1SrxVrLLjvJXy77duU4pTqR9DYUFWvs7LHDc41ZpzKVVVRV
5ndQtAeZNWK0+0/BysMX2FQfZI/djd6FRMmZj8U62N0Pb9eOxmKrWD/W0Znt4UTW
kkO4U15ddaNpPfSAls19XAsTkU/Uk/O7vOywqMehb03IhSxhx60N6pBw+c4CN3sa
//VnwJc1QubmvEXYIsch5hx+vkL0AVNQAKEDuHe1qhT2xDYHcXOhBPbMycW/imNx
mkFeF/Wg2sLc3mtjq8s2imdLb8J2twcw8VlzO9wZmtGsQOPJ3Is7iyJ0E3N3SICx
zfovyA64Mq3hiabEihfUrIF8kCA5e+JKhjjvQRGajGTiNAdFjIKYj08aksxN9OD/
dfDrIifxhZxyeYuQO6T7Hpf6Z2F32GFn3hXA0efh+N9wyNp+eZhWGarcR4M58jI/
K3snCW1qtJvxURG26aoKIECZ8RjCh4n1CVi/d3QhJlfQWGkCOpeCmCPWGTzPBIxU
Dd9NxHQWJjuZU9+tPRQ4k/GGQ3sqVhydx5gD9qEbQssdanvwIQGHpYEqflCAu10v
+xUwTnpHnEHiDJ09Fat7O97RSwt6T/vY0GhUlxOVXHT/XhX19s5FRiX/K3Adc4U/
G1logmJch6EQ/ZH78oftM6ycp+3hVx8uVzQb8phoB3gNr8mj1ibQYs4R5sYTSKY3
zPqlb9E11Pfs/RfuS/qFuGUjfj9D6KK1+74JAfFvPig6LnvnZtNuPdlEsaOSxiew
VKoqyg8Re2rcVWMDc3ZsalKNwnPyttBdqMqAPeDWVGnJ3R2/JyGNiEfcviMJDD0s
Yo0PZXgpK+wmSHun/Rr5crFcV7Qnm/wgt385gz9pX/eZKRq3nRIAxqaPwDjcIBXQ
JAQ/05W1YAKKg4TcrmmHUIaGokzPlTC9e2YK1Db+r/wXKPB65PcCzoeysN4CMnOF
oIxRwcmUJEnwe0PW9eYhsiXbhixWIhE6iIskilhw+Us+P9JPDCMWnKULfR/3IAQW
OmwApSzrY+ZfdcDHFQubuRvOf6ZnNqUVEFDQ/DyzVY5NrlJWuW78kIRN1niiz4mr
VsAh5dmiDOOIND5D9azIl0dZqqnx8/SBK63P4WXUwXfVG6YYYqlShFNE4BG0Kok5
2FhJ8d0O2MawYlUxKQ2YxpaDiZQyojDmxPiP551halHEJPGGTgUMPSmq1G3S4gaj
DaXUdU9/VePYvtQ6kl5rChcNQHI4dEmnvm9PHbXE+/sskxgfIrNWg6s/4BHR2Wxp
JQ8ZO1a0cdrdoTr7QZZinzb0wrh4rNyepxISK1mg05C1qSeNLVBHJH/k2YC99sby
Dykq92Udrtyj00Z1bIZgST3NYqteBMFnOvbdj532JHSWQJUCXSbRaKMoJjmb1+kR
DcBY3uotyK469X5zJ0naW+TG0PPijZS2EDvbR/1SSYbXmerlnQ+hnEoFYxfvkBZ4
IBKwU3RICP3TxWWIPlWPFNwx4eUjchzk0Aa/Ie6lINmmnewqLvVr2rg/4KHxOFqz
afL3exHVpO9Lrohgmc+tjQ2vQalIXlpzWQZVBImxex7P58J3ikvcJO6j83t9N0Ol
uFFRqB6jRq+UIMC2JWKgZkEr5IrhPMiBzRPBnPN5p1Y7DyR3hwES5c7U+M6ZrG4X
JA5bmja8RJS2spjFWtGJ4bQhy1setJGtX6zUIIbXw3ZzFFa+1A+w40S6nD8cr4ZE
Z5ubDxVd0DLtUYO6VriMpVPvP5KvBDU64mDrm+f5FoUn63gK4GFA8nx3cyuzPp/U
b9sRaZp/Hy0Ae8cf64u4OiJdMV93BrJfc3f6N7/93i6CRdnjJN3jGEjWDICLAEGG
+vu3EpoOk7wCO5MHeIh7Bafi3YBdUvcJC5Br5p6cxvLWG/DFPcvlxKf0NDtO0ML0
X66y9J1mbJhIOVJU2j0XxuZQF6t8ljwC6wfckFcG1+MF21fPatRHK2aON/PyPt/h
x2OTNrHQUUCnKvC9k8u8fdisLQ5l9HeMAnqIEQJqt1N6s5WTy+n4Rf2XruBare6l
RVbpicqvSLRKmQrEs8udD6cFBhS9iDOqLEzE9nVwBagVn4aMcwDdDp6Z9BENy2xR
ubOXjtH2Uti7Ta7Naoo3LCsIvUNp2SEfNLbzPx5rlA82C7J5W8zLpyb50wiVMzQp
dxk9nC4pYO/ATXybkLBL28DASUmK1UvWgzKv0lGBzPlBromlZBUjUSFYKOBvx5/V
u3by5RXFMAPxmJMj51IlCsijc9lJvrvdrdg9RS7hUVWdWRAAYWoF0ENkKg5A1X8z
zIAfl7TQgvTYNxbikLKLEmzhsEZnavKySasfMIHclCtJ385jE4VnK3wz6eyvl8L9
Vy+Jf7hS3dIBTa7OxArUmAS+qkXTkyr2g4c1dXzr+7tzG71clUwlH2PB28ZtcKXo
el75X2D2rLUUPypOoIAjxYBCUz5ogxML+C6n6jSlPZQ+irAoVa3CKdqVGA3Aa4bR
Sm+Nohkqv2/bDy2anY5RUeJmhfNOFCOiWyMPPIzYzxOtkLVxffBKgGMA7iIfkksO
nIGTDjI45GqMhTrWtp3jShDPo+8K5UHZG/HGlobP8DfYFZfVKwyxYWIh7+vY3f39
usOufIOMS4a6EdOzGFSPqDfOFf7mPh63aju1abr5Cbnj+OjEzPB4YTgf/B0N2DY6
Ay8mvo+qA730KqD2hsbc+ED8dFLB+U62pDw/npZp0cPY80d45VGQy+0MgHG5En0g
4FPKYGgmOsYAQx45n2r1fEhc8lAW2sbld9fuxNwNXN3Vuy0NR5WcWT4PEFIw6PzH
eH66zKK+dVKwM0C7sC7UR8QCTPfSPFKG0wNmyOcUbAabRacVgfJNTH5uPD4pfAVK
aURJY2S2GxkQybM6N8urOP2Sgp+lcxEsDr2yZnbMlBxUzEq8ieklrcQ/meOg3Jua
kK0bxct0cVfslB++vdPCIDR2YW/jAjv6lj82OciETM2DZ95WaPQ4IQRZQdGBAeBp
9RXKCqYlb/GmeNhgcMGY8k/hbfkHxYZNYBugUnUmv1gHtNbZOlpbTybJXg/1+5YN
VVzaa+9LiAxoWR+EykIwN0Z7Bv+wL+6MoIuKgvwiUMGpfo4zeaMnK855J6BsGReS
W/P06FZwezgAfHtUVf2oaK2DD9PAD0BOMLmnfdpwWR+PZdiGOXe+JYVP7W2naZX6
84uj/QrzxBztgMSDf/OSuW2kQhUHyuTwbfocbfQYPrdCwcS7XBJBmB8tQmiGCMXD
gSObgKD8hF+mVY2JSrehQqztH1gmM61mTXHvoqcp6qUbJpuonf+wTJ264tD1WKLb
2dnVd0vDeyc3H+8mDNZY7wmgsVgse8SBJriemutLT9s5NcOaI15ClCJe+TkgzEvJ
TlzPec+kFbMNYbSSZx3Wzb3Wkz5dqPky+v3v+QFVkp1ARafEhT1xpYvh5YxoAxSw
v5sMbih1qZCn8nQzmwJonMaGOXIQmxEx/0p8U0LmDnmGc8PapJdYi1y1yhM94jfv
9KklLjQsMxO+o+M7WZoTyKAfMrUdfNK5wdryzXfqECsQY+46B7NBNRtFDds1oEqF
/tQPSu4HZi7OamY9SBbAMFl2UqZXAQkdnANtCxp/M63QZM+1D5VXQE+DSZ7Cm5wg
OOxJkR1jLurxH+1T2kXTnszrSqTrr09x5pOlbQj04X04Sg8qCKYXnqBXAYf1VWbG
xKCqe7/2VN83cs4MnAIQ5lnOAbXfTszDqanm16JLj+mGCYn5JVOrSyLuHYUGrvIa
tafibkWVn4xlowgXgoHwp9NU27ide7CT62R9dQFt9wu5aBuQY5gK49uiUUmjQHc2
DSP2X/9KTKfW07nhcoF72HWxmg8V+ij8DVqAQV4k1MQbMEPLxc4Q1et0BmcMfF05
P3I9U1enyiaJUT99Qu15GkG2FsOvgtnyCbVEFG/Juh1TdVpF08fWOIZXz++lPtYT
QfAq2EEbikUuzsMC3zcrV/03YuNveaMlGxX3OUSXNuoP1TgX/6vP+fuzXwMeG9I6
4MTAOLm9AgRiPGrXBycQ5b4jMPpajsowm8nJcaVoqnhuhQi8E/yihwSmQVanmUEs
oOZV/2bcXDn6NRHa8jvR2k8nKt/O6PD/NFP2M4oF/TzYUrwQx4tbHhl4rHpdxaJu
vLkck04dB+7Su2GjLT00aPIVQsL4W9sZR0v4oMz9WLRoFXvvD/Fvn+ZCe7YR1Mcz
L5vpXVY+evovuEgULxD3oM357MDKdy+mZg2tAaLE7vs9DhfucbetD0OgUENbhHXr
0uNHcwt1uqi3XeLu4qPSvnA1jIQmZeJyVjbZOMnryOjXcQhO3/AIP4HT6MPEa7+p
kGXQWKa31SDzeJiwtEgtrSa4DTbeXgClkk+BmGs5Nw9XP5K3LKnw8XbuYU8vc+7Y
0NyIpSAintUPFbwUM7+xs5e0S1idnsCrLCoYPFiVWl80nTRA6NHvbCUfOL4lTdul
tmAIuJIMV+KhnsKn39M/XXMFMAVFb/QoeLNsvmn2f+yvFzxmANWsI6tNfZDN6M7x
stWFlVzqFaEr7xGnN5pxRz2XHU2PIRZfxreioNBmrR+oonT9YmH+UMCU1tskCe7L
YF6cJjaErJjvOyME358oz/6uxv1UTked/KNXyF9vy9f/L2EtFQiG+TyBbjop8Sib
h7Dq+D6OCQEJVeqq/v1bX2YTqR/Ek/smEL2S/0q2HEIxOd6Ar+k6p+d8np7cZue3
T6F5n7bMrrmk3mDaYtriIWe33pATGVtvLsCP16/eOV6GVnciiRtV167eqOoe4REm
H0nZEKsBb7n47cz9YMlGdKXdOqTzt9/wpDzX2BWvFXhocgvs1CGk53Y9MQYER6Py
eVQ7OZGltsvBsBIXiq8Ci0rB4Ika8qhiU1cCqjJNCPadJHASdpCz2lmVAZX6wdYj
dZROvZmuNfp9YDHCVoRJxIoK/nq6Bf7CKvIhm6Lt0EqE/FVkuNHM0w80yNTkqe7c
sPvbBkLi90P02DOS2uJwwMDQUsNHxZqRRMUue9ZrWhBxSvl/oaIffMLnIIvDDt9o
p5l55WOke0S7j9Q2AtZgF8YzeD24L0NEfqlX5EzvovP5fQ+0FmBjfM2ZNqDuGyu3
eVx9wpflW19QYnWWIy9gNjfGBMFEY8QBDIL7KMCMZVPfUVpYR71W++QkXbSNGUbk
VxBA3TGwpsnY4CCdHxKL/q7dbn+mcxpU0WdL2Rn8WTl9mbx91gxP48mRRlWDIakq
5hQj92t1g4wwjCbCGi/FGZlsvXZm8OZ3Eg6ySACNUTb+17lpwoECqY8Z5hF7lbHc
TqP4VooXurQU4PzsfeDNmpqIR3Tf0XukL/jvuWjEZDjdHCZnA8VUfYfOblJc123k
0mgh7ZcYm0qOEpPbAaqj0sj5jaUt4vnA7qWGq8sVEYAv67IMGjWJH5MQMNlakI+a
pWOFTYSntg+S3G0I/pmQvEJJQqGJr5Kzx4rFXEDt9bnQSEmmexmYRDTKvpfbF7fE
OjA0PY5obCV/sEu0blbcFrXuYDu6IlcsRm+pOraWIwuc1L91IRDXhDeok6AR+j3k
A+kRqYkyyJIaV567pvgNE/xpFij+be5xHfUfFcr5zNUcwYlwjqtmF2j6jcduTC1T
uU/zoWGDbmtHTaDtD1EKhmFBOP9xf9aj6vMDQMT9UQRxAVbAh10I9p/WnO1MASlk
Sfgd7wNND62UK6Koc7Z7pdUh9G52bOl8RraFu0l5UFMKUxm3lwMp0TW4V5i1P99k
q28J5PFn7xXeOrwyMPHatlfiM+ugsuXsAuJf+UPfIb75KjHWTOpB1KBfI4MAmaXD
fBMNzpDdZ4R5bu8PKYVMtFM67bKr4EhH703IvR4LvIlO9w3dIbAGxqbP5CfD+Ydw
BT3cwQ3VhEk4nRY0uNg+H7xh9AxywszfoBEosjo2SFA2Mz6v1fHuqPYWIZhbxDxZ
3JdMW5R5ZuO+cetiPIPOzsDJyYO2JGcrG5vkODlQmlG/uERZa8lx+/iP9e7Hr28k
cHWhnONrUbYuPojVE83+t7giOTWKdDSYUvyACgSpi7JJMJITFt4QWK/ba2sr74n/
p/3LcFDGWmnSHR/WZkt25nQhWx36kt/0n6emL84ugBbRQAntpQ2DhmTnM6h31GAE
+dzRmG/0pmqcmp5H+iI30+m+HPuU/7Gg81RrTT6P46qttMP3+8gkTFNwf4fxrPTA
UHq+tV9y7bue0/JnF5l9Lzt6KRkTv6Ia84Dtp+eVdE7Jykeh5IWeBoqybs1mKulj
IRC4jaEWgYJxEsxJTwi5AXrokBAxo2qfjV9riW55F5ZxcsFi0FPwq4t2D+GifoA0
5POUChwhGDSP/vCWCMIua05EbkS7wIetKcAcIyUFE9LcJzztBRyV0hU67pQN6bfR
qk6nGjhPquC+J7WfkHfcHWiw5vbmIrwp20EmbDr8H7SNSX26MBZPGwDxGygc+u+i
IchWYL9nzu2N3xTFD0vQN8yN4C5fKhtR7U6Cw0aSvFXEZQypr+jqJX9DyqwvSlDH
BPW1Qq7Snqk/6rG5LmIuc7NbSMLxaghkRBdVNTyK0rkUa6BMluySkBzR00mbjgLF
h2MBHUispvx3f/OpT6srNhB85TbKD2HSU4j8VoLKQYfQiePMgh6zH1bdB9blTi7e
C82cvB6FSUzatdMcBLvWNRxtgII372MBD43lMvNMqaQ2D+soDkYG6xQwsY0qTKij
KBbNkEPGFx9ryHJlber36y7utG++G/svm7CL+kLBoHTGAd6P1R/Nkheungg4RaD3
dxD50rT3jpwPTRXhoaMfzFGpkcNX9NtmMH9gc5lwqCkHqVRyIEU4l4ba31f577zP
GZaq+WQoWpNGc/WKxQ3i4B7XuL8/ApYCsJobfw6Z5D4uG8IhtjhB0c8xyBrCps1Q
4v0ALChHlyRaZeax23hxFcTT9fwi+wufna02a4gET6vcKhpDBXkzCINUGnxngXMx
ajdJuDPM0HwQyendX8dvMMoOUOscwAnZgbbYG1/eUZV1/t/+YQU9qDHoUTWgxyO9
7hpYYW/lLzZ5y8XUkb2DwvuUDw4WRIUk4KSiUNetAaM+jXgNOxQUfqHXMconhV8C
J+bPlAKObQOj/pUeA3aNmk1ydiKNRMDnY/stBwmMmtcq5Nabo9WtcpSsT6j8q5je
RkGks+Ye/NrkluiB/gmYJgGOIep1/BAWR/wT2OOmChVR4EmDGltTaRc9e/TZ42KV
WwKTAlcn1zX7w6/5b8dqjZxTHfxOfBTJ30mOM3crNcysScfjbIPcrOOJuC734RGn
NsAZEx3SPSllq03E3+HPvqu94eHnfZow4SW2SsEy/XkTQCocPvmMSmQSyVJW5Dfu
YsroMRdtB91dnxG14vCWzLG8vuyArmZYydNmjv96HTee5i8EbWpMHRYYSOP04jXu
6RKc8pM0D5q5VeW6A5gg5OwnHtO/8ancr90GUuAWWTjBC/PgdAEpq/AL3y2MJcvj
l6ZppIUiTJzEjwAKenExIFzo5Ty0cGkrKGeB1srmZBVoefXtkTmIcSDNAMzWW1H7
w+s8GpsVuui4ohum1GAkeVtLHDWZwao5zIfL5UQyXj3itMUsin3awr4uH+abhEh7
he7VY5cMsg9WhCfISHlkfoooHlEjxHKJiTSnezaieEbii+E4wKsyWC1qXn7wOa/D
dN/JZcMQMWl4OWTnmMj68xUK84plvyoKGqTgJ+THFtTyOjY2iUI+WYuFj5+Ux87a
B+y0fdw9cMpsjoMUlcUk2JkZkQ0Np7wVvtqsWFAOYediqpi4Tn5XjMxeUlUuXZiz
6QU6iNhzzaRWc+cQP3kChn2tRBFNn65P+sRr2SFzUOiopW2GizxWJVhwUfXeuaEt
h0F9Zb0lbM7pbZkFqu5XUW8pGWTZ/ALclIN6VpJDsLd8tvx2goOf0zT30doQ7PwZ
7TdWn3g9EjCY+Rm8sJTYq+EmWNv0NnLLvjnLjHRE2b4RPiZPT4CYEYkU5gX0W7sJ
C/DkWeQ6MpWYNMHiO71VZn8qXr35UJsckvVAHLGjgv3DSdjVDma3hgfkel+l4oJR
rYO8uHaIAK4zZB97WgaZ33K/Fw+ROKcwTuSlymcBllAN4tN9XxT20z77nxJAw2ES
w8DU+L+tSkrEI3mqFJA4Z0nq0WpqWRZgQgMuu11bqUo5cdr213ckd5mvUU9IV0/V
+Tya4ElkpWJThDvhLPt5QQo9sGcOeV7j4DaiU4csfTwxaKOk4GHdH0ZoDwYn1zIA
tqIxXH2u8P0VcaDt+XJ/U+JEF4+3CymFjEC2b9ZwlFMwrRZYO7g+R+XePyzX/XlW
jKe+a/zCGBwZXCR3G3LVII3R3V44dNMUXFT9pcar/BRd8y95lYwR2MTbro4MVIRn
RXXo0XeSl+hV8AjxXMt4ksDTehzAdEGd128yYZJja+8CMD+H5kG0Gid7GLSc4O7F
XZa7TpyjbMfQzTRzGKvAXOTw3qwDKW9h8R46YQ0XddGfutMUOP24dZrhqgBf3+at
NkKdwKnmzRpsSl2t36+Gp4Rftbsrif7vNBsrWjvWgZYXbWPppBnEi6DTTO5Hd8hO
KQohI+srNhAi1OXS2OiXDKQoxDeAVPJfKTsTozWpFFr6WdTAIoATjNlsFGPDBGah
Zez7F3N5J1FtFtcfdCzJfEfGBNEbaIRtn/JeMoN4VS/Ssyf58fepbp7VypzGvjEe
KgZFysWMzygCr9o2zXhACW6/BFUgE/a3u9VxiWTNwsruTGoXahknrEBj2pO5dL+j
HX3r31ZwRsRCnx05yRlK1br17oHWs7jF6L1rFiHIGqvvW0Y5D7uVfAzQBNozFZrq
yctCn257L2qm1XFUC5MuD+Hk/pypr2dc/WQoTZFS/OaojKEqybIh3oJF01Cbidzm
NKF86zNcZs8pc8W9ZyEGUEJolMAXEagBaXWwseIf4mw1jMzjUtI8ME69TeB6ToO3
TLVhPT+N9RrquNEFW/csHP+nWA4CvDHzywy25AEBcVwnKSG1rfZ6AjvOp2nZBb4V
PRGIFZxfw4dpbW0a6AW3Y+C2lEMLkOJy7A/cTe+Hy9SOYTRFcah2Ev9ZthNb8xpA
ejAacBLDxc/R8T3VWKZGfJgFgxPMm54tYhyFQ096oH297fe9mmftBJZKEFVx6+Uz
k8M5oHyzb67c1iTQNQKZrHw7SYkOO4+KnXjVY47sHkpFY7jplDkluiWrncTbhA3C
SR6T9Nf4TLFSt+YOwRUYyl0aV3Q9Lns/vqA3BldaZdSvR4ZN2HBSkVui01cjG3Bw
SbZ0fe+gRkbyI39ZCuprVAII9vtzur344tYNVL87aan6tR4L/jnEMWt2Dbyf/KmN
VB9Z9PtweRBLhJ+nh2KVeBXiGN9FOhoSMLiKLEO22iLGUlzg6s49qSWekAu90Tji
pPBDk8y6gJbPl1P/gof2aO+uy77CbeOuk6dZdh9g/yq7Zv2onVrJlKj1RVJQhWoj
KOGD4CjReRtVnZEA2J/f4ip0qfA1XRjwSlUho491jYgNfN2GzFiM1daavR+l+qg5
6SLnwpSWlkju0JiA0ByL9UnsqkbptzutEGAA3b1Q8xnSv/x8mvoHA0sSSi9r3IWW
6WWUmcy3W1pnx6vxbIVbA1Dev4oA3t645wOKueOjdnZ0nDLfuiblIxu6rzVgawx6
tnc4qHCIDVfkfYI8sS9vnvKziGOU/AYccZDujMII8rMnLNieGW7JHAis4u/SKfBH
HiAxldUix6U69AmwzrH+r55idZdisYPqXzSsAIOEVwwwQF2TbDKluhfXnTiFADsQ
flLmGyx6CinrBO7fMAQPfcQh5v0GHAiIewxYhX0pwf7EN1bNEy7qgqSzR8LGLgbo
CuSLpbDxFX/8kbJdK5eN+HCGzyBv4EzVtp1kN4CCAX0/aTHF5U91ROGONfo6u5N8
jcMzkcSKd2NgvPHPuAjJmWAthkNa8IcPXDfPRGzSAux+Xr2pCLTe86GJma9JTCaP
0O08XB15fPigXLkEE7z/u0RFNYhGSHd4XcNp5ZgoRDbZMtMMefRi0U4xf1xTavep
dDMmytLIkZ72dCELmL5QcK2sZ2fEp01YpNkJrMh0lEqLr/SK6M+0rGa8rjfSDlSu
WAbjyBak8LpMw1gQhvchppxypJrkoGoJ90PK0tteAD5umSv9vvXbbBYztxuOKW10
djJ5WWCJz5Rbj3rVyWXCQKpWHYZfby31Z+8QIC8KiVdBT5OnqxlOG9QUjdVuIvCu
wiGkEXjrrvyBGhqVQhqA1rWyD5fraIFrPGdFi0fDIXhWzUzrDHUqXw2JjERV6MIO
JYhLkayKbc983DJzq78v59gJFeruMNFK/k9PwTxGTSBuu64gXhX0VQokxcuqzhqC
0C1EStvn0KGaDEU3xf4Ke502rRxLQvsYjr8EFHqPxvM/cyVnD9T/iqehFfK+0QAx
Kt11BJi301XJmALcaf+zO1m6nmb9ZcdMnMLHL+no9XeeVdMx3603XPbpQYzfXTER
bPrgR1vDyh2HFftOh4/Q+xE9diYHQsoVBCpEzXJadtUpUxYidwmFkfsagBZaQxx7
hyD8i+IcoZ5uFHOCvIctS4X/ESDe7J9JpGNKEo3e/qC7oj+9oB1mrFAFCsaOGf18
NCH5tn2ByC4iOvR1iq9MzsULA0Ec14MXlWb7YeWBoKBbqHin+5M8ZegD7lDBWvJO
Ue51ceaGobDksMGqoatquBuGPV6/ovxoHEv44s+OEO+Xw1fLmQIXX9z/JWk1q+Df
qv2sdcdSktjcQYvXKjBWAWJwVmDOTCGTxgbZsx1E2acQ2tB8jUOMs4eKROqqC30j
TFwbl3Be6vzt88NBeTGAoKFsEt5aN7fdAetZ/PHkoGPGoTRg7va0PdKOZAEJla+k
RSqZIhr3ETtS7I5t411lcPxGiJlLrWAzx2KiLx9OOlGiP5733YRe4HG5dCEUWkTx
PKnp0oMLrVEqTh55NktTjwVBFFhizT76q9RYypXrz7IvDFEyc/uyeAhcr1h6pgcF
8+DgJ58QA0pn9wmdDAMAij1U51fTcsYF6wPMmVuy0weFm2XnAO32cJGMPbgKvQBg
7QtxDhD/owL1JzljbbJWlG+iOPa5B1B6S88LqHmVhFu8nfrYXaWOedBZtwSPzqRz
EFxCU8DgtdvUib/6peB7+ygAuDHAE9m7iwQuudnxMOdbydcOj7pYfCUJGuDRKCqZ
e1Tko4pGMX4vIjgYJ/2UI8sQ8j3pASJ1Q3KYVT8Jhg+M0g85czEvqh2Tot3cHAlk
1Bdbk4YjC4Ak+giuAFbB2ONP4SkQZAUqkK8J04+PAk8DvyXq9B7vEs99s/efK11b
LYmfRo2tKrMBOYEXKGBz+dIqjSactaohFr1XMEPvK3banOdfiVY+kFtU1W6cDqGe
OxVGybanRJj6ndFiEqovvfC1lvJmcgdvyBbGiZKapjen1gUAyV2OjDEzRtrpaIlN
limBRLkQSOmJeIuQG8oV9Flxm7mk0x9vx652zGWnLQWOlremzppuyxjeOJ9CABca
6km2rvmIvpogmqm6Nt+kBQs/Pm8GPaCW7U+3/04gfJRhX6yykNpSFI/oRF2gNo4N
D239M1r6rPc+FyYBwS8+szM8uwsZyNzb4I7j73TBlnqWLjHk26sjrwZ74qgpOiro
KgHk4++XNwkBm+wNmgq6YcRxpoXtyN2DvaIyLN5bydKgs+1694oBJ1vlCq12Tkh7
Yk8bADQIzouLmrgA6482TVBxuxs5k1d7WE2p5RkrWQYiYj/0Od20kQtBH+0KB7A9
vCapH7uXtkW3JECnTfDIJgb/hz/16F67GRSridFbnhqfHHINS5Fdpg/dmvo+85xE
YUafsGXRe6367a2foEQ7K4WuXM3CzvxhzYYm5F8ZA/bsFKzcJycTMYPA31Gy1f6x
pvzIt42TE9U52GvX+e4boh21825U2LBVf94+2h+xdZyFYrW31LYTB29WivcS4RRH
IQpWMutooXnoXDcnUvLF7RT3BlxwzBtpGPGZylhNvne/s+5QcXMyUhfxMa7eMR/s
I8Rg7+IkDg5P4kuF0KirYvbe/vzACsPw/8pEABgT2c2nNaljlAQANwvt2/0EAHuT
u6fN7R+4AUZnt8XXpqiTVAmVkVmVooOYWtoUsaDbd0Wye6cjm9zXHsKg7NOrbZHr
ZKWcnigqlkQ27IQ6ToxoihkKHeQgGhZkiHVHCcp/XXwZB5cpbpFf57hT16yn83K/
+Xr+ytAJpiL2/yAkYm5zNvM22E2lf2PdlQ4h3kxQuFQiJOl0r52r5bTIvna0J7Us
ui+DCKzTBPe70aLSPqfRI2NoiT7ILsUTgWQGamu5j5v4pkH4PE0/EHZ0Kw1oQGCG
3pR+V1Ud7G+u0UHQWsNKq9mHoXEWYy1U7QVLb/7b4Y6rzSzJtmnGp5/HBy0Yg/CQ
qYKKDH7JPnSWIVA93a2UFSzkZU5Bto4UN3CfohvgsUULUeWpr3XUk0Z6CMi35iYf
VegsvwvviYMO44Xa1hHyPL3Y1EQg1UUXvTfKe0HyB0rgvmqb2UtIjDuB1oXF3yma
0jmmqc393b/Zxfxjb5OnbE1u0sbfEzbibxiLPcs4YQDsVex7jk4ObcZK3oEDCMhB
0cLJiZrR7JQTOBCz3ew3gbM9HT3wIOPs1Q2p70mV73X8Xe3prfx9V1sAsvT7c4ER
iaQyM1SWZWiHcRN3XQFTk9jHqEXNFFjGOwHzBLzSJgryY0Gik3PlURET5c8BBUDS
DyutxeVOMIgzB/JzN4nwJSauZNvkTshP4URhP56IZ3EOIAJ9F1V4D/Rg1Q5UorG4
hJOiZi30L3fezSWvSNSR76NB6LEWCOQiEH13BA7DXrKzYTjrtzMV56w0uNkNdRc6
phc45JofYBgVtfj6BcYnNzqshb8qP8+RFbFCSG+EOQIC++Uh73C9zuw263Xp3GxR
rfpTwmpCGc59Fm8AkdiTW30KidcuIqyTaqMUflsgEsy9cTtk7fNEjtH1tkybWqIO
HF/i0smKbhu6eCUEeMgivkIqOT/xHMznlfhF04SeOfq89lu2zvhHeTk9NncQPXNE
1JJMH43Q8Vk645BRtg9E8YVPvxYIxFRdWxVbwAniY/hZ9R8s5MarrC/4czES62vA
aIAPlW3zY99fAgxrTLK0LlLGzBjwVxF5F+jV6V9UV+O1eb/rR+qQV+/TDcuSOWqs
y4t61uh9Rs4TtnOc1IkqEUOCvfRk09kly25OlrjecUtCpvvK8UYYhRlrl/OXbluM
xqs1sIX43kRCTFYMX9or4SrIHmmP/XzHPtDs/9SCGzjoyddwATVSMeP9yHzxP/6v
vHY3uxojfECqCZLWhFMPsTRXYOF9Mqt19rwe1sxKyS8fIDpdqkKYGzmnyq+UyuL9
YXNXytmKPiRO0zZsYSYEtt8DdpOFLgT7vXwFzrIL/bY+SbOGsy2u6/hV3O4UkJz8
fv2SdHhgsW+siJ+JHgVNAe+p1GE1TjIQYob1qlvO7tWWxlfHjyIWPiyLt5vL/0zt
jzTHArLIW+maum13sFa07hJP57TDM8X2qWSjgTDSbOS1FXjZA1S5ZX5IKHezIA6r
PaBg/wZiQJtzTjjouVcr8XfmXq8ZITbuBy894yDwXdDmA3grU9lcwi6UZkn/gvou
DVIgS2StnR1PnoMkPNG8ZqIBjkdGU6ITSbDIGhRzr7G2eozQYlPf8Y6P17NKCy4v
AL7TiC8KHfZjvZokcIf7etXNM0kpn9D8bz+SpeCBmMdLdhPBX5ZQShbDfPBSFfnf
JLKItGS8W9RsXoK59pg4BYBFd0+X/MDORZb+ZLsI1052A1lrTWVHUZ7O6u0rl8kh
t1nx1nUV8cc5kWiV61Mn3+Y2eVss3hnFMXMoOTBqHXrVirG68sNXo0ufwNK1GrQV
OrKuwKBbVUlGgiUqAsImSDym8PoEpnXIkUg8KnjPyRz50g6x+uRDnCZJpr+riagx
9vRYxcK8zkC86MiPsRVa6oXifI5rL4d5NbHgfL5Eum3F4qgSnQThh8nGoDMt2KoV
bd1JX5De+BQRsgHPsx9vw6qZylNMuHuBBuNBEbkSklMW+XN3Hq93sX3eNQmqsCCl
4UuvhNnKcWATXE/O17tKoWoSqX5+P4dfiBuFCLE8fPNQq8vuIUdTWkgd1Uy1qemG
aOlNNi8dV0ZNsgTycs9lXA2dXKBIKyy1X15euK5dF73v+SUDEED9feEG6LUEhfL6
mbCXv/0kd9b0BYPzsGxmcSlrxjG+VB9MzC54XrWIYZo4PGt8gM9Z8kypI2hQC9mC
GMpYd8bzWsMjfBfZ1HGFl6q5LQL8Q1Qy3MarkE7evCZxY2ZvxobpCu/dwAGNw7o0
HBTUAeq21ugo+/it2YaajetwJoFYN9MClkTPhBdXaCUo7MNQt4wlteWjZNOs+Zas
saor9pM+KdlaN80LIsImozI29B5yMsgi90n163UO+GXVVrTApjbgCLADVewQwPcE
dXK8908CTcTWA5B76iats2GxXla1z17cIxQKhYivBUybeO2e947FtHNYC1g1LmHv
BgMEAqUczR2vzN6/QkOBR7Y+aVvSeLVota4mqtXYbeB0Z9VTGUZg4tBFhWhuRNX/
rc3up+3qPJafjFFCU3F5RbIyLMuJk/js2bt6r+vKoEYce8+RdDenVC6oQxTyK1pE
B0LWm7kHcDsKHABAfLCD2EUnZWoE7SDBpkth8SDheNR7sPwEWiXioEmTZs1JSOKi
tH5qPrdJ7Sa5zHITLi7nd1AUUREelMB4fAub4zYqEwGFw9QrAGrA9GoNzGn8GNDm
t37IfI2dcVUySC0ajJyPBXOpOpS/knaAKMz3k1x6LftLaX/uSA7RdezL33PK72nu
/bIJSXyZ/bXgho6Kdc0coQ==
`pragma protect end_protected
