// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
VZTZupf/dembtiP0Ol7aK5owI+GZDXBfrr48051HRRMgUSyq3h2FXppP4TIEtx21ek+GgkNpy41Z
GR+7vvwxSMiky/EE2i8VfZxDo7RYclh4gOFBPon8w9ypfkK07HQn2+BcFbbiqeE3mXsaI/8hpaxB
9QDeq73b7Ikv1Bhufz5DYGDgixpGZKTmxEZ8gnw9qO+J2QtGl+MIMOr9Bau1hsVNSg7oSmfJE5aC
gU+RwZyR52QbH19gKkNnLBwP/nGM/NsBY5zrYgUTpilb23y7vDqQ4bl0SUlk2sDdvXAyL0d2+n8g
DG9kitmSkSQAZ1QM8kWUjYffLV3rRBs/OGrn1w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
qrK+rq2HjFTbXP04q81U/MGNSOTjWHOkpShnxdz4ZjrVytGk/jzzGo7L1hgtgIUOUa+XiRZYcV6f
OZ2PcchzOidq5svg6MwbU4JKw7VUFyS2BaPvm0IXg8XXfdCNDordnw65tGoaUZv4PySbptptq4G4
e27Aeh/61JapTY40CHbDtONBUA2jyckxTJuwwB9lCClAzyfQQa/kXSMfLT9Vl3AveEiwFmPtJKaF
6ELpvf7AvTrolu7U/8n1+spMZcFOhrdAT6R+dO+dYdqy4EhoDgGTMs6INaUsZ06WyhNRV4inWgJo
xhKaDZNCAwzasRepE0ylSkGbHvv1uKisJY2xLPprdqf3n+9oz21oDB0rR3aP2+Y2yl9rATOWaF0E
5KsSIbZslBcGBVCYsKeQVaERuS5wfT0OgTkaWVnFnlcIQCVEnvIJl70aIBJ6XOq6v3MuGJ18aBbn
wjL/DZEPVytWyKL1hWxdLu8APV2cOxZ9gf3uFwkjKSsiR9sXpS1H/CqSTcq/Uoj6/msRXu+X1zQ7
3p8beQPSwHvLYwmT1Aw9hG0ysGiAuimU41Xvn91mQr4NEbn9cnWRJdPZ5M1/Fa7P3rR0dIbp0/ML
JBtaZf6gwTADOmh1Xb+cc7EpG1SEzrC1gSLzrhJZwpoY845vmausq9yvmiqruFA8pUYUwnaY07ar
c7Wyw+l/Xa8JodAZBhv1isFkBB+mPRb+I4KU5d+fkTZLKJk8/iffbjAH2ddGdLL6TRqkhaTWpOHJ
uDiXcnRAtwfxO6MjqoypsSOyWeBMLUGNsI+LFmzy0CxybTOk15pkaedj6J3/exluJllYB7D578cD
Y+YJNns2iyL2duvS9j2V1HY4MTZOcTFxQ4KTfj+3d1tTB02iqmdN3nQAbiBhy3tthuBXlrtOa2bS
93ytermQTUlVve68Eflo9lYN/xSzGEqBn6JQNrvqrpOhijJ8bXm7DcHftFHMMSXZs8uljhBmdxUt
29g2hqyrE9WCF3k26ZtKbJUug2/7q0EaHR46yc2607/6fGEf9Ew95jZksnk6QQFvyfsz4HNw0Uzm
a0QdUBKQVjb3NQMFKhQ/MCDgvMRPjNXxIiNPCiUIR4RxNBUI2dVmpRjEjnCNusg8TDIA4AJ1xTej
VkpbQB9m7XOXosG5aJRoemaSsjjjqm0safvwF3/fkDrmy32edCeD1IPvdhPVGW907UL9KIr5nRs/
vIRP70UgfSwICwjJeanAxollSw9Z+K3GcNvuyKnnJr1VjfEzTQ3gsLOboCQCmJFy/trFRRduM7s4
fkcSmP53DjYEfaRysO6pJz1+AvZRHk1hvgJSUYmOwRBgEtJDO3xhDhMdNqR3jNIOr6Hrwb8ilLpt
6soQ55GlSpo1jGI0y1uXuAwiIyA8506lLzuxNw6tWWKIFH2kDtQETFhD+F4ENSqP1DMd+OxRf3CY
IBiPOWxhdlvjhVL8r8GjpIF52ALv1jlYlLIG0HYQtql/tceROnRcCjScRM5pv/wc0B8GNSKUDzxI
acMdZVmZZRVSnwp9YGJ91r1UJiMZbg9KWKjSQcqQ4GKXU11qGN54HCXm0lwraI/aicKD5rceMJGK
kfoTIuND1aHE00tBL+Ob6ah8SnSTBxKL2DUnlSKIUzhTNkqjbUmO4B8OHG2VXgpBpec73jv1Odgh
YqYljqf22WvYra5n/ZTKUDQRsW56EIURBNToo/JbB4pZdB8HIHu1jpz3h9YUSmy4aczcVyjl0EN+
jgRb9BuJ8RRY+IxCiVG19YPnpBaoqO4x97uTpyBoPNqBaU/yfzEAiiRgdiJs/a5omlg6E25wvWDV
Y6XP0afjJR/nBMA3KotuatIjglUMVcZoYA04titDDFwmbjmu5J9w4dGtO/gd6lU++2Wzb4sxpKSP
M8v19gcs/lqnNI7os4yBlh6gxpxZ/0BbrBZS/hjMj7/+dQ6kSP2dERhkOa4xD5K4r6Kr5asb+iyt
RsHZueHCOfH2Evov4Aq3c0PBKax6cWCCL1f8UporP9r56J8NT23mGj47AwCSQ09cQcz8EOx1d95M
ZSKk7DTQ7AKkdub0QFaMVqLpWT6nORozZd2cvnD0p3jqVIwFZ886E9Oe8kmQqzNubemeDC1Gk2gT
CF1V1mY8E9iXHDFGRs/0ZScQvdqofeKKa17w5Bij6APULEY4VSuplHMYV33QLRgpYVjcGTHvWK09
7+gyp8ui6nqR5ivS83lPE0LtU4w4jYn0fnr9OjO0DbvFmU0o7bqsysyC8fuXbP1xPe6nJzvbxaEz
HtvXOxGXElH/1yVszzTZZ9L8XS7UQu2a5FTR3d7ytQXR7B/xQjnDIPZ4DN52ehEsz4mo3r+hMIFT
6z904VWpgC/OPvKxbSykog+GX+AVKYD5x6zxAnyqy6NkuW2M7TeA8pz1Rpt9tIoa41Lj3t/Pb6Rd
f/vwahfpB9pS5CZ7/3VbZw7zFswRfwrboFaRWc0u2omvy+aV8vTlaxuHxpKrUig6kk1Ipu66pkRU
qKehT4utHMQ33Y/hH1XoKdv+TyiptuhZTxxSeQJjovUJ8bWZ3xYc5eDbjTCV203hB2+QbJB/fULk
GtDMpHiCGFUAZOrgJam1xAtZlbELo1bgxgpFrdjh9KtHR+lDOKHVmcRXBmWkr1+faCfBZsHDFz0+
eOfIHejCrkGculbhDoLeg+v9v4pxGkSQuwWCyguzXIg9Zhkns8BTiC1Jqr0AfStlpIX2o/BKfRnH
DOi70CBEcFmH3W7ST1sV1ZGRN53ZYWth+v/z57dAVDA53IEbnmp18wD8are6BibfeRaZFsteZSDl
/85MfuoHIaboAlhbEMRkBo6/8spUR9JiWUMUV34yHxRNNXFBFsRQEdScJnPyAIkwcsaCBlTkPzWm
e1+uBToGJR47eNOwfHwGD+56VoCqHkYawMlGY8BQooNgH7yAVCYVizlP/sHRst1cbxpq98drCeFy
k8age2ws+qEDEGdTGqzwDiSAAHZT2zraDVNL969VoV5pZyjR7GaQPGRH57YwQKBIrqODePw09lPP
1o+WFE/h+nNNz9OmGpbSkQ65j9UGLOA+u6JImcU5oibkNKmkuaknp5W5s27ebP4UDjPD1+bV54B8
7l4GHDSHpLWB9e2aMAaGmt+P66F5HPDoYqwdzaxbO751jbCgt8EJ+PpfLLj7ho6s4PdNSSqTVnuw
cmCBIvevYXSS4B+Z5jil0v0qYhR59WAxDQUJJzX86Y16bL6q7OtvGJRkAsvBAr6q6yKRIeoDp7gA
x87yBXWs/XrOcyoAWH7j8f6OeZpM3JzHZogR6FOwcwA2cmUQ+J5lCZ5CUysnAyNqVoRl3Rbcf83U
ANYhd9Ujr0v2LEDkr1sOafa8lYZO0JrUsnULluRoiYEMUy+Kookg3kYycuSdh2d82izrIliqDkUq
bZ50QK15SNMbbmh/wRlpVucVIy7FPUg1JhEfqETaFpt41Bmuw0M33s9K+l3P4bswsUJULl4ZTFHX
xn0829p7xMuoi2F8EN3ol3lO4h+GpbhgPCFIlYfapb+pRl25evhT4q2wYRrUb0fi9tkbke0TZX8c
pnAFrHK2GsWQDFr+L1hC56wJnwW1pkqMTlUpRHzuNt9OGM5/y2el30sofrDruDG/4ryy16/RTiQ7
bT/YLOHiyEEfqnKaisvoVEb44Lk2VW763/0N9dyR+/W1eQWB7dD2FLuU8iridChqOgu3CI7JdyP7
lwRzI73WACO8eNrVClFLaSydnLraCsIVvm2334wGMxoizWLL3eRsAUXmsRt+ZK/Hv1gcMPvEN4aZ
juJXD/ZhnRYkki0/NpbdLHB0tkpZIXopkor3PI9e9SzXU6rDFb4x1Dave6iGpwl275J9D4mp24Bo
c8LS+B3+Y3VUryytUePV0IR+RKvkhIx9N1STvEmJLMM44hUvKjBywG0qUDEOGZeRh2OldHraPFSf
9bv4ivUBEZEn+tsBqC+9hWrkMbWTsztkbmSEOzSz+5u3X1KSL5TgRRRh+fzZDrQY3UBFIt1MUsM8
D/KQE4ywMQnxyTjDEirvT16OyK2wlbOzqZo+4EkOqWbyOKtxVcrn50AYuLFWwiigM16q+LYKDZNO
oK8AIxvw+ZtkoWAI0cdfxl5EVD0mdAXoT3cENU7zT5BPtufv6y1vW/s20fmXJAszp9qgsApnrEzS
UcCBLSYotnWXatJk8owb/p+CiT8P2MUCCTJfTvf7ywXlCRqLp2wdgntFndW/zFHPvcB+3iCTLdjK
zxM5jj1L2bGvZ18n0L5DjuoAeBQ0hkRXAxzunL4MMEKKKxAIAU84XeDx2CEIm0HEelUa7YxXFSI/
aQZvqSKOg0c7Wm3kp9nI9dR1ouM+8rGnjm5+faaqWDG8zL60vLwpN14ILGyGNCv5UlmGxxkxZlfd
Es98S/D9JImFiksHO9OYnFNkPS+eexn+7aDNuNLTVvL9IXlnIc9ubvuqJrEr2ItFz/Q5ENghRwQm
gZzwSx7ryOko0M3BlbqFkLWO1rotlGpQ01Nc177nOXoP/r0FzF7KIVfqyCMhylXSbVxPWaeV0LXd
I180R40+tUkUTc1qJg2V+6OJvqUwWy1aEmaoAlpADT4ULR/Au8Y9XivgEON+R+0FrTo1gOmULf8d
mrYkBv5Q+aLj3AgLEB4yNkgcJxwbzUN990Zz22kCc69s7utP2btybI2m+gL3ztXiO0aIxOXOG2Nj
NEzUx/E21wBiarNqU6iselFJ9goumwNx+7RhVALw7NAOr86fEhiE66CZGRWBFcKaLlQkGo1/Hdku
bsD07NmrXWjuspko6xcFY7SBl0Xb8as9kO0SU2ssi2UPDDXVY1ksBUrY4zE+qSgXrTDU7Umcq2SJ
/6ygDndn+UPaOS1dkwQrb7Jwxr3BW0nj8bxo7Lbc60bI2BQ7c7sVyIeTNZekFCpap29vWYQQvxFH
GB2uiwjr2E9VSLOyVt8AtZcqSqOSdJKmAU6axcwsqVnv8MdEKDL81ls0SzXT22mfaOV7mp0fKz8H
hXoDBAHi6dxg2/ESUpVYy9qdGJ+vsGsvg13u6W6nDsgHWb8/oIWDvUkJA9ZqUs9HcdVV5SVv17YZ
67jBtni+NqeLBa6Mu0Zhq1sIek5BRA9M4oRVvac6gpnlA+NIgamUUUA5Osgc47+BvfH3hMGtZZd6
J6iHqxg3eBBXOy1Tfmk7g/DjZKmE51A0jRGcPPhiLT7EuVZdCWNBEKxzBux7TJa22B6hAYs5xZCc
Ma6PX6T2b+RhQdJgsl9phA9E4rpQRg1H+hqDtfMA7Vy+IhZNZ0/Y7ot15u9vFc/U2RYZR78PpPbd
5jwlXg3gDf7Eg35xbbF/ilZbz42Zkgb17vwhWslyAJGV5AZyMFKY/22IIbVE0/hv1vJCB+TQIzY5
L+SfKgf9nGESMw9/ploXyx0CD3D58dKQiVSN39GZNEhBksGsp5qRcpD/RcXZTgeK+iZV2iJGYraH
HsXRfLjPuW1E+3JI/aybq2TBMj/3xkKzHtyMr9zMEYhUZaQki7Pq3XA71RVSNZXpB+InsA5gIDkV
uLjKwUJLNM1QxIZsHdMH3ZeqtZgIXASS/mRitJUodmHy9Lx23TGWF9OnGfAFmjzHvVpdIUXtTbiR
QFsoeEoZB1q2YWdbTh/SH4przqjfgaxnaS1O4c55oxedlvq5XC53+JQdGy134YhpDKzIKodJkO3g
GrrXVh+k0H1PXqK1fuIC+AJKy9P/GdfDNXGiuZp7peb+DEHyg6GtGUloUyo6gwZmQZhvnRiuXoaH
8GwUlwZuaShErXmpaWPuDrUU0ALIeBf5ntRnCBemQPtgkQGpe3qmom+rpAZMnjk3ili880B5vBH6
j+BtZxQIf/9XKB5Noweopt4m9m7gpCLvCVepSdhRvfw9JzJD+Djh28cZ6OGcS4+BrHe2w3PcM6Nj
51ixcdDgk/KxAG1zvVY2ezh1ZrL+OLZQJTXdOI8wfxdEMw/ltQawfdXQ1r93Tmnqs8mqnZFPD08L
TmMRii8eTxh4k7Tiyuiz/j6lmjbDAgCspjeLwN1qUNJ4Ese74lSk/kRAuBM/GUnlw51folRf2oJG
vRqj9QEgs1/x0mAOOD8JLMIzVmyJ3cuMHylVlKyIvrsbrSv2E+/PujyQ0/QEaKBzOVghCB8dqvbL
aefY3QEqR0iUZzba+FLzyjplOH3ZI3kG9ThBFZI9ntZ0wm+FVElqbv+YuL7piAKyxPdpnN+gFcrt
2mE6lgT6rIo7wyKPSz3h3F4kmBJxBYFxeEzBDIIAp68DqVVx4p+A2gYlQsb42JG5qzz+X3ESFeO2
wp0yhfzQqZljBhukhJV3aGaKJuegEGb/qroFswf5CGm1Kk6Fwp+3FRQ2TAcG8GWBfqnJ+KukGZA0
P2mSthRtBd5lWhN0ZPoHimuxZNxrdnmEyeW8Laq5wmztqsAvVHWVYnrhEiqF/CkNrt3VDb4y8cSN
ScRA1+hkDFxYdUI4Q1bcNdEtmoykSAC66rFC/Sl2gZ5JB6CRCyG3pVlbck1N5Q6VWHUgu34u8w14
/dfC9cAUVyaf7lv4Zuh6MCZXJEULidClt5HnIfScNvXCaZQ6GENdGtzmMeAvIf11o842ZYgcfHEx
gPascGhrMKSLPlR0Ovj1uVkOz1jg0YzBNK9VpJ+pf5Jy7Im6sPT71He5tK2Cd60DPh8I2kdkt9/u
MIQENUUmWSr/LsOKXeIJbl1i/EgOGCo0KGS+mTRHHrwavAoYMFxoM8D4ITSIThFWKj0SIonJKBg4
mh0qoxmOyssZP0p9r0+sWppSU7/3DxsAz6J7hipf2aoGc0AEBCd71lWWWHDPyx6m59qsZdUq84u2
3wNY4QzfkNs9DUQ59Lf4JZQyBDfe7hQhhaVkpQqb8CCvjMRi5uXWTm37qlHWwGb+HM2Lur1IFXUN
lhC/d1TWxSOTfUEnKrWVFhQohe1Ih4pNJ9BlOQhASdpK4KPbOle3CAffYCzOVsj5Ei0iQ3U+xDxG
DSVeAlbCwTwezR+iPcAxP0HriN2jCF5P1DuCcik1Sk5/h7AKKCTkc12Xw7qrXGtHkBRusMZatUBy
J6STkCKHFd7n2CtHtlNFpN3fZEpXSDE5BR3HhhjmnQ97yvmKOzD6yJRmjRzyyjahmJAGjwkZyBzX
zooOpojw0SRN0UCZDNGr8Qu7RPwrzintU74/fTGrKphZb60tAgc8gnMfxSfIg7ER9ZjTERcxljhr
ojarBw5trcgmUlJa090msCtmDzHCS9BSTrxmbesOlDpp2JzN/82/j7NHgDT6bt05dLad3bDPZt0H
zy3dYqFmcwEfJUTwmmHsaC0XBP4rFnnu1F75ErRzEJpQzUWk0yOO+WQR/hvyiBdlkVeYFlrNBxxh
6JyFXPfPy/FLu9IbWaz8HL5h/Lh4AlHKFD7tDcJgFYDHHBpv3ON3JP+Gd6QUFdxsj4v7k01TIh+m
a6VLR9Xw+sKXWTLVjqwwjkW6UieZQlOMCoNeNGV3x4F465omf/xNI074yMfYMEvJeFcNIc7Q+512
Xwf/p1qD4+ZPfPopj8I0zsLm/h9rknkFjeZpizu9tK/GKoJSB82WuMbZ8kf/714rB8Py09ioa0gR
2pB0LUn7HIFpIRigyaCqVI8SxOEpH1+N/K3gsj7rRv+o174JZUqz9vdsQ8IhsPrPj/VbcgFuvfMY
xkYrGRDoziG9VnkQIFpNLLKRv2miIh1+HwmwoY+ZpTEQ8nhvfyLVIQLEKBEzx0vvU8zvjQxr5CUu
XiaqXwqwHZdfY7vF8GBq9N3QHpLTnhZ/vSlZTm9KhQHvHuYBiG1W2gSDdGqxuGikxPyM0RB6wMuB
7jpf56JfYeoeITTzNdC9MDeVPSOlqx0B9TD1tvfPAL2iGo1HKNEvPWdKMlNvHQvZWPTAolW0pf7u
DCtb8R/WxRON8TXp+Mb+jztC/aao2QsvdjQXlqZqvNtDCt/LoED6q48d+vVHSLb3vN30AIAXh4mS
udJ4G7XG10fGSGCcsbmlN+hSPmWjDG5NGVdmcppf1Tvt4TpMmcv878TBpYVVj0c5ucHPR/FicPwW
RolLe2i2rab93vbWQsGwoLuv39iymNnmqz+QqETms7kmcAdBSFMNFwA2VJ350T3lV5rulxwbs3WD
7LWY1n+xrXGFpyF8bhMkDf1E7/ROM0yzycUcIdQkUbApDuBnqYdI8xir6uv/AqqhTfEqnG2DCb61
8oRZIgFmjtfd8MROIR5tH3mIbCdflBMdwF6adC+tRKoLorQ98XRzqjmg3BHVBFqNkVNA2/ILehDq
txoK4KS3R2EVMw0DcbwhkEa8GwjGVXTVdC/trV1T4NWd0Jro55W+jLfqZ3UMKZCRcGms0lnPoaMD
m/uT7OZY9f3G6jHe4y6C7HzQyjtJFUX0RH+frmEdps8+ACPz4n8f17zm6USZSFfsEt8c4qzXtT/J
+mF2Ua3UFXH4+lGKcI6/x2VhvqjpwDfqQbsrpR5FaSpp0BISSE9B1inVwPKcv1EcnnhXocf/IsLS
FLT/T88wwVoxncFgKD6OMy/rMA22vlJdAqWP1cvdXxk3eB5I6P+XR+7K3VUoVY/Fp7dvC8RP30hm
osLdTQFG3A/Cgn237CVupP6R3xxrV2MqN5pNn3FkKJAEeNDxp6c/xIBBEnnu2MoLiaoIu7oEfk20
6yKma7ERgSyrblVO6M86T5phnM4+qBPn2tXOlj8TlH6WieT9drnLOGoAvivoRUh49NUAVMjy14Gr
o4pfl2LD5Svw4sA2/dtWhoEaJtj/82p3xLGOie7YXRtDgzayi+weepgHTlAy8DTeWkIcqKozHxKG
zz4ytQeHXkzrfik7ACCDIJ1vho/N+1sBW4R/K7x1Y9/1i8raCQKZRy6m94yAue2dgA7IRZBk6uXE
m4BzVIDzU0gsTFgWndiRdH3n8t6barowp/6qA+S96kNIjYecnaz7XX7WwEtLnCOPj16bERIUHeYk
vPogiN+UKYBWJu06PxGC5GHbqoL74IzyqsQfNMbJDv7B0rwCBEIMBef3sKJJnb4r5yJEyhFhNuiL
3e9uwLThsOQ1sYensYwsYvst00bR5SHwbHA17QmlLs9kWcj9VmyixEwAf7JACCk6O5vPdsGhJcgr
Iz5bfR343yOYAcBFByw40WMCNSPG65UBcOzo/X2ONp1nxL6w6hmW1MbudBu/e24Xv2//nabsYuy4
KipwixKKdvHddJC8V8o85u+YGTAqHjmdZcBxUEqLCIc7WHTd73rbSSYCSHwGKnTKlQ7gt0xwhxZd
DNhbSrHoew4DrWOlF85wNYLz/dgAhW7Iu6n+ZzRbaHSv3utohqzsewls8nQfckkDgWkwAZWwCfiV
XyWWbPzNNVwipLMZ8xeFbtlnNqgymsH2SBAz+d642Iptt3+KnDpfUdlN9jkndtlXEAOrbYl/x0Kw
F5hHf+0G+qNBzxfiXbjWuyezeNgYQXJap98li6qlaEzvaFLhMTCQliXzzY1YzZ8j/swSKEzZA1gf
SPfozkgC6Hq/YJJHpNQxsoxuvG6zgv7otfmZbQvLV4pb7gOS7kLTRSVNRhajdAqoLyULhObNz4eP
kfTJ+ncjxahvMM6YluZjDavs6Ygc0vBYKmeRWekMhOMtcX1N50/rUKOzpAu1ns4OyDlEwGqP3e0i
1ZH6RA146cl206n47yU+ZgzLU5OAtlF1Vio2PApcYYFiuBXi+fmOH7qeZzJNQ+D3RHH6jAEgcfwh
XCnw3EHXSe0xR/Cc3BXtd6poBkMAj7SrylGE79kswT1d+dn3e+oxHTRs2mfDugwgzjuVaJ4CeI4w
on0v7kGa547VSbByiNebZ7VcXp84t35aJrgiySUJFgIZnt4jt8VafaMETl9HM/OIyOBtPwm3UtAM
jTMvoF7Ay9Oxo8wimADvf6z3VXtQjulrTQTinMAPiF/tTD/Pz8nTlQnnXiBUIUM9DMAvwcJhv52s
T4Wpzb0uuLZOwHT5Pds+qjnB+oFCe8+O/73xzz8OPBh+GWD/3vOJFxSkEAkUXPPPsmbyqNVG7PP3
mLcXq/huhn+Qyqmo8fOWEjxufFQlm20/O9pEzOZAREGvEL2MQohgczOXd4XuEPg0vbpKPjzG8zTw
IeOKoLHZeJC5/TKhfUzrrTIPFw6ZJA12e34vk72v5To+3NSGXFKDtzKzwean2ln980i4VOoFYrHB
rDOIR/uibIxKioZHw9sfmZtZL0R2GQupCIHw+aF7ryUbexZMZbLzJJUAvSZXJZXPKxo9oV6TuFOs
jukFSmdOYMRia1gV3n0AC7Qvjp32b4k/AQMf2xYQDLdgBf+wei22NDVHbZ+SqATRdhjDmKm9u/3g
/T6sEFJxVl2YCdp2NW+79MACYtkI4pVVzgKhwhJKx6fE/SIDXLyoGQjLge1juV0cJsVdgS689M6y
TyztMF8cw9v54eRkZIFoDSIhwFbcDm3l12Na6NuMEzPBcwFZnZKq+Fud7zeQQfhThlNH4ylrOVWu
kau5peTXJGktJUAVqYssEHxnrk67BiAO+Uk+NX8SAV3hWh+FhPPn/cYKJY3M/j5DEwjcaOfHEwNH
LwEbkaFZ9hEyAgrbreI5g7oV+WlVthYHCY9fHj4uQLcp5i72Fo5Yg7UedcqwgR/NS1Cu8XwVU8/2
UhiGVnh/rQ2Ea5F76mma7nyOiu+4HNlEYbpZ1aX+6dredggAoFdmjUmjxUVwgltfn1+iUiSrxzPU
gDeYF6F+TCynQb5QJXa0Nu13i2QlpBZA4MDYOlG9ny0Jjof9JASB5DaTsNSMzekxXw9nk1oRc9sw
0+x4AchctNFUMaITceHm80eNzGoL0C9D7tPB8O0c3IuY8Yk6QEQVcppbVHjx/hDPgaxwn5jq6bAe
lDQayg99NnxEWctzDWHJ1U1OQqMRMUK8nxG3tBybnokjKOOPqwHpi1PVqnda6TWJ8ggeOAn7eJs1
2/OWjuohZWc4fTB3IXNaDRvBLiIWmwkKPSlLn1bMk/BsVR/hPfQDIZM3wbPyqV/d9XjHS6EXWXH8
6SHcIfLjrq8Tdyxpr9QIMICwO+Ay+zYhXh5JwyrZ4LCfFATgBZuXdOmGWPmamuAgx/bDvoqiNaqg
fV8YnCjrieHlHG4mk9nCeZ2B7+HWId5PIt0i87FUY7n9h5jd9q5P2RjnxZObbYRepUpYFXzvlZqc
WMys61xTeSoq2EEPwAHtoZd/fLPUcmObm0diHEIslDY32tzW2u2DVwjmIFoPJUs8td/cTPkNIRpF
ySwIO9MX4ROmtMFR8i0cDiHop8avpeLgJgrsAq9bhx5sva53tCMcf0EA6CJijeAN2NRHFsVWa3Y5
mk0u3CDDmKEUS0RdO0C2/FI0xfpVIGsBuJUHEKzP3F7By1SnaaEKNIM7E+EDXUduXXR5gZZsZyzp
MdhAakC/mvwjCl2DaPnAS0jbbvlFzhSeNXRm68BBZMfo5GdLRducFa+Vg8ldx2Q2z5bTujVOV51G
6NLNU7w+hpm/jul1dQSeRb+asTdfwIxoODhmsYbyEzA49FMajxjBRKjB/V31N63lRE6d0scGD0I+
+1B1ErX5GotcYmk/G5L1c10648U4AEnNQba6rZuiafCTdAJSOq9isY6xTs7NWmcUaKZ/5dcXFGkb
kNNT2eBqoxOgSMOOiitAPLSsFXu/LxpbZix2L4arKEI/Jo302+g9cVt4COaOl5tyESzFLzUuI6+Y
m+GOQwFtfi98y5uUL53+OXltwoHNw3SgHz4rF5rKtwj4LYyS2rs+ujBelBKiAtkY0HaxPaSB2mvU
/y1VowMoAIbaBrnuh9tQ+gEx990A9E6Q4r4kVbl4t0yCODDknovo1WY+LsddYP4F1Rl5GQdaIPp0
KXaxALz5bFiZX4X6ffzKctpYQPraKxAdBboQKio3Z0xffFWOFkXS0gDDtuyvrDEjU8Hzpq7Epy6p
9B/G3L6HW5krNuz63lwPLHj0r/VL23MQysvEHwsWbjk+st3GIKZD65G2sGnkwPIPIKeaUHvpHWm8
Dj/rlIF0RCrCoOO1conE3Og2e1d6p1LEP5TcKuK09x3FxQq4rCJGzqsxsLjGoc6Ne9VXVT2hk99F
N5RhP/7iCGhnx40u5FW2f6r47bRrYVMbE29YkrY2aq/TgFShppfyjBJOg+09pG7Mb3MCquyVr32g
/cBOrdGSDvdSrK+SqRXkDCaLfYaB8YM89IcQIMcmtZq/ZYvkn1cahjjukEbng8J+Ge1JGjnmbti5
U5rEzYIXA3s72Z72HDtORfQdehO/Yl7GasAdcisPF4qIoGwrnzuINJ5S90SkZFwrPyZUDibuqyG6
5IFzC0F0ZJjVXxBIub6oSSgMpLfwifzsj9FxtMvdxajHzV3FE4/0o4SQAQOTiGydULS833kVtxhK
Nb0egx+G/iYh8OyWjjRpWAKTK92jLUiuT+CV/S4OaauxM0YK1N031foJjg0f5e3cW4vAs0ougF/X
xDtSV+u8IJoX4NdYv1GmUVNyCzZzOePBLsY6oz9wx2KpyMbEQJbYSngUQzVeL8mpaQ7R4n40I+Ez
PUJRutGple+RlWr/Bc/MNS0dDwWhNFrHKj/AhCKh4+4X/AgsLH1PrxP4mYH9NRaqXaMsPFWbMoy/
po6z9UKi+wRS1WItI4b7HXi/PWWo9UYOB7GsHZnQFffExqoRgGzf4GLjUFgeKsqWTwv2ZF/BY555
BDDy7/Q11Chpm8tKVU/cz4CHkJY5pwLftG6O0X/7M1Gjp7ocrlEqNHRsc2igWiQm8Ztspa0ZZATo
KzOQFcyjTmYAQZHk9rx8EhaECoiIl/2yxqYGZAW+v+49UXOf5vQIhKkt0vjgkn9sSpJw4vyeZ+6L
zgk9DlyM9Z/LgW1+W83LYapz5vYBy5gmW5JZnBUTYcDWeeLb69sEXlp7FUlS9pgP4pqUI63+es0S
0EY45HiRFFRGf/A3x0ZSEV/XdeEml+xOwVWKY8nWcBsFo06zvKxFrySzvRPGirwzl4XoqpUkPwje
cxpk2p5/SwtW5jmH9LkAmneyugZ3/BIS140f30BZTRrH5MGn3XQZLqNs2/yWt1xnWWj+1qdiZPvD
Vh+ZWPlcRUCDQoEbVruzDH0DsmVEzeHgLOSKAM7IxqfNTSdMphLbZGcWXjzIgtenMHyXv50cjPQ3
RXFoCklfPsghp3QcTWH1khb9g1pkxVeTjr7o3hlqSe/hmaRMZnfpAbzLd02OLNr6YegnoyUFa6WF
HaCLWamQR9CfVUwfFeZwGluF8Bxb7JG2mBslF2sva/rP71IJtW5oOfAHo+AAGJ2pUX+ZTVrx08F7
CBzLHqj5vMWFg+hE77mXDbSid4YiXZx4SUU1T4VXxO3OVf29IrlAYJ0OkXcVmMNZ/4BWV27skmq1
U84A8V602QhFEQLPk7Hk5+G8lGmviUtb/5NUFYPZVXZ6O40hWJJw8w00qgQKCqpJWmqe/2lUdFmK
BnH9zhKxXhJfcEl+6I5+xEyoPTQKTWixriCsZEPCmy7KIiW2GXAcu4dCTH62mlJC6bgr++IxZLEA
f8BYKFL5cyFhYN2Btbaka7FyTPqsQXxxh/zircx2tCpP7mBksZiZicnpCHEc8a3SOnc//VL3Faus
65uq8fxF3dO+twIXhUT4zL035wLw8G0ndAaIAwIpy9utCglxLlg5agDbCV63dPcHc8qEC7ztbFn1
CgRGR9AgRP7gpxfU63omZcGzbYlx6bezHGxDGsmpkQwwOuX/XW/hk2gIh8FXIIIT+QZ0SK2457Ln
nS3ASxRl5wcKyeNOTGQJt0Qn2A55gpz7pdBQ0PZrV9NszkXIbrntp9jxSoacMT1dIEu4oTzI5d0U
LdOBacqyEmeuYElVMUmKGD9AwHCVOfxOYFSs9nhjs0TcJL95b1sF3GKhHJ12egfwmFrNlIqPC5zG
p4CALsmlbdImA18xTqnSRq8mF19bMo9ThzhupCm3KBS1WTErdVjSG5xK1tmlPUvpKjX+MS+JKIra
OUyS33XZRjoPlgeIJ6RfeUlxVeXHxjtQtKa70mzfcl2wveq2baFdF+jbJkz4MHThJA1N0r8aIsL9
rfy6LC0KmYj7vf3UOymV8pAiuTSwBndRhJSXadXqYUFgE1wEIP/jyl1uixEqG7UZasAHDWqi2H31
rhg6ZXiCzsP84xk0txgl6m2ewsv2cGiIWSfTLQNKQ9KqXsnLV5GqKqwgXduO+yRx5RITdDiHjXy/
QDdEsGEkBDVgJdK4NzEPOq++SSjB3c53116iHyiiTUzhgcEzrRLsHGC2xhQR7Fgkxoz6uTKGpwRs
wYYeRXsIgoOMx8xZRCxah33Cpmz172P6TZuXmu2uhNfuG1t+y0df2Jj0ShWRNMf2vR1hLbCUBvzJ
K7+0GC+mSpKsfELIZAE/xMSg2HFTy8GeOjwYNl9RcduWhk4jeQ9S8jazAA==
`pragma protect end_protected
