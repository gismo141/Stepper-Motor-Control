// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:51:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
l6uQBtX5a+Aeoyb8cGsqQkT5etE4V32XBAigy4rdSavKFSWsQYcsMEMDbwPfZwoL
5CTIzYMniI9TeiFKc94eAGugVf0RcObqtLUSS1iLma4Olv/nXUHLw69ucEXNXyQJ
07t934jullqLil0PFp0KBlY1FseAUgQYJaVtVlovfS4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5696)
tBv2gBlvRiIl8nhzfFJA4mL3MQLRZgzCTMU7UfawiZZnZsGnxbJwKab110QNtsZ/
BolZzKMCuDjBEXcBVZqTTytFEV2A17NbpyPqNHhjaaYe8Zc9Y7j624TdVndUSUuW
h6LnKZN07TgTSPb2pSOV4ENLbpFuwd4y632G/swgE9XOis7ZFsLEHLe9Lv5RIy1n
YhVPQr1bQWqwXY3HquG8m2PiixwE2c2yNGvLN5/UzjWpqcPUARReFOYBmDBBsP35
I2nF+yzukomzxzuHHpPK6lQKbSFUwlxeD6XiyhQrz/t2RhgonhA5YtygNh3BK2ht
TsLELGhqvScjsiOB/Y7a5WARxfaVTcRqO/Kfr1XA9tgWNkEENCkfwjsI4SuDi5uK
LNlRNH2Gh6RANDy9n147AAK0M1HVu604qF09FTq9grF4SjHK4eS7CttHpOWTq3mg
JL3kxrErlaYXG7lKhhFj1UnIW4z96m0QNagGswxBLgrwCMc/7dgJh2mPIBkiFGyb
EJa3happSLK1UAL0eSzBU3eGK/1x+hkl3uewv5eOq7Apg6euo1f8pmSM7MAId84E
+YkSKVW0dXaC6ezhgb0Dtm1c7y6DKLFPmWAP6a8Jz02rz/VQFVO9RRqWbiFtZEfd
iVMCO10IkeA9nqhFG6yq3YLYCW9hbNaksBaTIdLQ5DtufOgP/DS/XCqYVB6h3XDH
v49+ET0gOP85nJvYHdESyO29wnnDuVRvgyJjZPmVEj7vlbxWlP+M/c2FeOhX6t0U
G576X+20Vms3FdSVRv7eAMWNYToB0NoMN8cVO4LpcTBelpBsz6Hpsq1bL9zYDd0L
L4mJaNmK91UX4f4Jaa2kNUB0MT3CHd7ZVrnGEcV/CLbbM6WWrB1xFIHN8fcrWfxp
ak5FedRQ5P205Na0yT7nWypx2S5qaK9PYZn551xF6YpBRZqxGe4vsfoilSfkVV+w
eKIxuL1PhBacRVVkrgukk3l/LfJlkpYYKSvvdnGlF3a3ZKUzWjG3hDG9EarCsKED
7kJmrBDpQM/YcavkiHGOtUKqJez/2xZDgvW97/VP/UPw10VQ65c2zS3pHTGPvfqO
FoXNIuqpfV3hofd7AbsdE7JUYxpRHBwQyv1EJw9aAolQRnVHybI4bz2Qen5+yz80
PhDSpSZhNt2ShPyxADDgxon/N/MeGzVACT70znA3nV7dhDiRxAU4qXJhY1mHX+N6
bySJyOcvo1UQlDIESPSFkiWEdRip+ieJyU5W89FnfY99PUu1Rz/qZ2NI98pRbp6F
4l8HYUq3mpfO9gS+htKJkMD8J3rzm3CAQqdz0ZAv7S/qqFD5eOSEyEgJlxulEMp3
VWaUPXCSeQsSrc/J6h74PoKLaCozJAS61M4c4sHVRF7eq1H3N9pIKPQbncTz+Qzm
F+IhhHYmTehQflA/qluQr5bPMq+S4IiRQADO+p3YnHl6dbT2rX002Xtm8vB8DydO
78w6GC6bLneaeDPlfDrynTairHY83sqM0ZdiEV3bpfUmpegtecPJkaAD+MhGZLMq
LjS6/eIP9kMXQ+Yf8wCOm0k1wf3Yq1J1PlX3N1AbEbvrJAQaXaWPyI0LcoBcHSIb
6ghg6RGgMzwmUAWKxjGl1I87uMuaHJaIksCNvqWvp/bEUQrN36HBgY8xG6WGf8VB
OE3lk3t557aQUexgLncB6X07p8z4z3+ok8T+2RExVTU34N8Ober7lYrJ2d+UFjaE
TW5lkJfTlzFabvwSH+ycx/bIUxv25XQaugK9xLQgdqSVp6kQvcfY5+riwj+RMppT
neuH2WBNUEAUyCgcc/sufznwlQ87jOw6C5hnt0hhqxfv4yKv9ka8ptkFmh2e7FdX
GU+HI4U6uABp9+kdwp/+oq6Tkxq7kEpx25qSXlPTkaxQ9XlDmR0efYeBChXSz1bt
DFk2fd3K4GboDFFqFRG8MBUAr7ch3Tbnl/JQalPJRoCcAzGXinTznLz0kgDv/kfS
rpzHYv54RnD5aIajjDtunUKRxWNTMzU5uyg2IBiBtWM+1hz68Uhz0NTs6opewR9t
JHwoR49S2YnrBloq1Mekctn10uhSvIX1iJBCVOJyIt+jj0o0bwbpvV8g7ZvUiTNw
ROMebFJ+V39JpL/pjM+2VEvAP2CnwVj6yaymOHiKMhIn+LV35+CYXjtwU2slQBsw
I90kiq5fi0h+S/ayRqt5Nli4MLhfbAWYUCyc2xOsJ3jxHMMIIuZ31XVrjjzTzJ2p
w3xe94AGKMUKuvnJivnPJuQTWanK1OHKRZC18KM1vdc+iS64QUASCDBVZeVUjD5x
gDUSpu9xUQ9Lx7+K13/olmyiI202o8QddbDS38+l2QxwWddP56WM0NApxcgsiKW+
6ebFuudOMFIbp4MsAtYfd/7u/Hu0qEHAEdATvhVkeRtAuVXB6mONkNHW0lg1vurA
F+XdGs9YyqR4ZDte/1UWHjDI0BKn94dB1MZPeF8HytZ3qD75cs8p6Y+CYmEnTOLl
27GwgQGYEgx8bRGg8R93/0iLSXtLbmmUI0bkCgHiPhs3c+v4A4Fmd6pNe89K8Ni2
kB8PlwSTwz6z1vaPt2IuV8eD2V5saywl9+ZVXUNmZ3BkFS9vPxvysIvPdocwH8FW
LyTMQ9RQhPWIcMliAk8t0ocqrZ+Um8ujpQQx5eETZTTZvV4o1TARzOfZo8XR9OoT
+AyNxicFnSSkjBKM/tRu0ajkhqcFaYW+v7Y0xe+ezJFV11exDVeDz0pd+wlHbU6W
+oV2DBTOi9Y9vVTXY4WeaRbBJ2DQYE+I4gz9hcgX3bnDETELsu9xHnEI5cScrgBb
jBuyKgyymsEcuyiCHnL0Tn6XAPTEL4Qg0Oy6icfYZQ94b1OGoEqVZIsakny1XyRS
R7UE3ikHitxvsKn5x4LKQGqYSd1I9e8Mms+rMvXN4o4O1VjOPixrnvgE6Ouqnb+A
QMpjtfiOxIldnYkthnGp19gfR4uRyGvPqTkLz0PXSGF4GyN59qqJ0WmB6sP1E1cT
BBpnJWXgKxBD9XsHjdVxX3yxmCvTHGW4Sy382uaCNlrnp+ycnv4GBq6hEC6KAloe
0c23HfjCAee6Aqka5OsiTQ9BwixRXophFA+WLZqaMN5cUFl5uhT0KS3clhyqyBaj
VHFRoEULPrVGEjCyxPUaRvfFDgu/RipWOhEOUJJoCl4TaQezPS9myLT92oo7X/4i
q2efm7EqtqnRpA7NIa0qqin/ZFUHQP+8YwNgLLKlxR6Gxh+cLbSd7aaTm47LInfk
bYeMkDO8vuVKCeIduKRzPC2Ibi5qYgln4VWcoCMJdri7Avker8Uk9aH96e14CoLh
uZMq+fXAwY+Sib/a7PC34kfz6+02hiccIDJwz0IT+Q0UsCkaVrY2vZdUgN29RI7n
z6a3Cxoi2kubarhKY+o2pEub0i1udaik/d4lIAQET0ikrhG9crKIwKO4++UgEPZ6
1oblkH1eerBx4DRVleTZo6ZbivrWeMA5tfIZz+Ft005kPuwff1lRZu9pL+We5H6T
aKKD43tXrDLyiCdE6kYRLFJUxjIH0MAQD1m3py1rrITfVXwEH59/+aLJ9oCYeUYz
nXQc3Y2ZwOp+dcPrxE+lxgvQSHOhdQXZWVo0zWiplHEtIiUSSveBrZqHa+McgjIp
PFzyKY1SxsS3FWE4uUzQOCbJMqX1fzOR6XwyhCT40t8rtb0roVUST207rBn/v6MZ
SBAYjNQV2NxVogKOPlVlPKwaf4fvqqeo8YROIG2R6bhmEgrSVlahV14QOmpsSn1q
dYRw1+08bz189W+fWdBgTxddWsnJOqEljnJmceicbRARzXz3jg51je9qsakhkwSE
WzXLwJ25snSqkGwkkaJD8OdbVA50o/Z+GHK4y5UtysRRe7QkDXpHDxDAqI4whizn
9NfP2jqeowQI0lEtokjzs2TY4WO3s9RMXxzUPemAWaA9/gwhMN9hi5DSDJz2I7PX
7+SrdZElUQayccg6u1GwhabkjbD36PbaX84PU2Hhnkw1itEvHKlw+uSbvqZzNaVj
lsKIRzjwBVqvaOnUi8PScmQfVv0v95BCAA1oclQpMRds4GxzMv8iNDGiNWjF3CTp
fmgYkjZLX7IM1H95NrJEdZiwusdYj0ePXQzslOFFxA36JTb0Wx6QWf2NoACy1hWq
fXiEea+1lJHDp1bW0PQ9h15LqY/tH+KWkHiCu+gUNCzbThJynLyqCxenXveXHoce
0kAg8CqePPuulKQ+yr7yjiuPpt9VJAIs1+IrEKmWbO+KaHM3ASjU209l7VDISynk
UZspsBzHI6sIvSudAbVIbIUVRv8AXLlQzYZL1gxIvo966XFuq9w21scXIqfSKr4A
6Bw65wPTVoTjld35F4qYracr8XqeoR4O0JFoyD5isvQVSXDleUL81Xrul8htrxuE
nNMMELbcnaR282tWS7qgxERKL5e8E4krAEvSwRwuhVR/tmeiZPUnlkUUGC14iXME
rI2u2/Ys2lcoCTqR9KkgSz8fKvvzUyiR+LWxtcMwEo03P3e/REjZF1hA2Q3b5iQu
7YTz6lZkzXVD8WXzitphjHFRqlwfODe0+fauJCxH+kXIRz9rJtv5EWB1VixebRjH
OU3XgVtVDOIYL2x/dtpSQEYL0NX6yccq8vBO3HY0ssbVuVoPbjSEo3p3v0qP9+/B
ed4IuKU31hpMkl6Z2A19EVhsPTZWdKMEpNPDHb+GfbIiqWOMt338ihHADhCKGHWM
sorPSFHenvnNBVmJ579iXguwXLxAjvybSeEDrv8PZCXMNbe/UL5rLZJKq7SIoPZu
8ayDTFH5J9/QwGrArAWyeNtXiXR7nsfR8aLRhiDs93ND50fAuLoPi9Kxg3TvO7GZ
4eXyCegJTCLg+SbifITF8LAm16WGcprB9LBrlo6LYUKhcB7YZSg3cRAmIwKAOwO4
zDnOHCvZjalCvnSH4CIB32ppZBmq49MJKJRLRW9EdV5seDkZrVhy9srNUxANnw6C
PslrVSiaTZfIj1WQOjitn4CKsOYQsQbzgs9G58XHZOmkc92GbXfe8mC7Ah/buboA
egpf4nIur6AlvJxw4zFSs45L7PrIQKWZjupmkcSYoo0Y21z/PWa2Zl5tYo5qhhic
fFAw5vhvGyBELW27Sdy/wWcc9qlbDpDd0RKR/68mw6g7kMcxuc+Y6LWsoOI+/0Kv
M3h+cRIEEUN3pGWdYP3f+ofJmaoGgpjBP0tmFR0mBu8naL6iyXZ140CxUIOHeH3A
0kqLlozKR4iq5JJ/QICY2okwetd8y1BskdzQ+MITWU1sKCGHQuDEjNIRsghY9/ct
Xm7p6j8mTLKk5Ez/4UJU1OpznCb4WyuWSFmDzvZMIkQqbjMFMCowWVNHTnfxqwTJ
jzCjSOMPt8zisExcDyNi+MZH4UpWP1A02FIwqXQewBVBSlL4AMy0dMz6OM/J4XEv
I1vKDPbXorY+Yz66Yz79aUuZjMZAH5+kWy2ijjyrUdurkH1ebYBb9/vM++eEmkba
VFukoZisLoTJepBmsWk5/mPilQ0OisY7FqwkpNqP4UFap8IrxvOCWeaDN550nmmy
o5WPJyEK7lI5aUF5je4DlV40amWA9QVDkssTzNJ0gjrNZMKgYksi6ORG2iuUgk/n
T9Q7MHtd29U+1KpHYN5XZA1xDE/68KSjdMGOtyUTOD9zBrogXAP9a90XGwOeHGIf
p6Xp4SGfdda4kw8o1/lZlIlfd5puadmWWKDdCaNhK6Axi1/8+Z2kf5QdF86wX85L
cxxI2KxnrvtXLcFbn9TxFSko00SJkkXtwX8/TuzoqZIe+2dOW3ugluidir1Wfndf
Tqo0n4vlfJkA0ey/1ZJPCyCRXskSmYJxaSn49SiUce7Y9M+nhVLP/46FarHsKB/6
xzFujiMVuoJWXqHDxQQ6zq1/FerLfC+W8/vXCWzBFGGBbOnWWUMnP9OYPUhHjyXp
2JhxvY5NCtM7atN59zzlS1dFH5Bla9HIfhGV0DHKd0JoVH76QF8IjPxRT4UdBNtW
0C+fFaMN4VmO2XE6vzcbzdCS9+5cVT1/OlWoZlaR+UNTChtQ6Hha0CuPK3IWp3/3
1nQRwzcRFyLUE0wxx5ygJWbL5z4/+Dnkc98WrR9q6BR4Uht4m3t5BAkU7RPpHVKY
877OOz6siqCl+7dw/Q4rDmflrObh1THu9+j8IFoQ1WePDGJHWaqoagiVTwoTiQ/g
HpWipoepV1AEj6XPmd7+wUQU1WsIPKCMu6ZMmwyFhkC3KpWTcoZMbpI4bJzt8rVM
yoiW6KVFGtxsdYs+eCG3A5guH1uJh8CTr8KxdIU4zLhS8HCQdRE4xxtl2ukXHpWF
dTzs6O9K1VqqSzBPM0HNLWLiz11vs5HgTWEI5cAfGkzrUNdLPdPajPhiRjYDjO2u
Esk3GVXCE/QAjTiI1a93iwOMEAKDKD+GAtjRrOvD9XRQ2YxCNmd5jnsH+TnspE4+
2b5gY5Tl5e1rmAXJVOIH2yBAnIEyzVHreySIWZp2fw28h3HyLkS9zfOrdn0oDMWB
lrsHAeh+IGCxHK4nvByKymWNir3QGtLmg3vArFoHDkmuPsgU9gfF2mLICgy5UNKq
X0qJcxnv8RKJ2mSLpnEVYmKF2uRVe6l8d7MNY6HjGYd87f+we0hN8kw4c1SH56b3
tNkh9FMCz9dCp/e6ove3MgUSrdH0N329soMtQ0r8nW0v0JaWV5sOExDq4BYTa7cO
eNbLEV8j6rW324VERVhHsDWpgoA8/6FI2PV3XZRFVZFL7EHH7fjVjWMARO3KqOiT
aXZWHj4E743vVlZcrBg21/OhYp+CVdquY+GJqd4wYqIvUYy1POrZz9Hg6zsG8cor
Rxhi9S2MbQCSbCDGC6XW7Xv0BmO1Gpt/uh7mWeYtECllDECYtugWB/RDyjd0NI0E
UWluKiy6RbwiaUQ0PeXb5Cvy5qp8fexqb05ElyVZZsvl5uN8nYFZkSRZlI05/Q5Q
e0nEqyKmX2Y7ixV2YL1SIwqKgAAGoeN5X07TZHvp79rge+H424e86uG+G7EFnJ2J
0juIVL3UF0DGl6qxsN/Vpu9hj5eoJ9847IdpVScaBIeWmrurQIXfgtAnRkHKADve
rlLZ0hLiZ5h1VExZBo1DmN+qVozL0BETGZ4kvylKlC19tfXdADX30iMS61NjF2IT
X0PgeGNyxGYDc8fPVwnzo0B+moPJyG+WB7kvH8YoI+yDUKlONLQ7nBAiwaOpiqxj
tIqk2oPW/5raA5tK7Rb3Nq1jMihUklcsLM1XrpbU7Wk6HlL0IDZp4rUwvKtJmt5X
5veVfxhX7lXWB8znE4PLGmVFTpVJI6XNmfIYqLqF9u0erN/pHrr+vp1klaLA6eWv
N2ShIPR5jGRTG43L34mw/OmAYSfYEoaYzlMN8RknMAMnOm5b7EjuIQ8zYlG9tDwe
hIoBFTRYomRz96MVe4OBRPGkYWj0L8bt+wT2/uKw5YkQIwkrOoykvxeeblLP1TKw
oK8N7J3VbjQobc48nVCiw3e45dC+IaLygG3CODrxX/GKhcXUBlmHVhKE5s9dmCfJ
SUhbjac47mtHP+OT7k7DDNRAZDJ6kLVGs1pFPQ9LvHc=
`pragma protect end_protected
