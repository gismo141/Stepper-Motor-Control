��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n~����1cg�&Ft��ͽثc��N�i\r���y���AKK^�z��U��Z:�;��KP�B ��N��A�>	��h��H~,
�z�*�M(�b	������LV�laD=tp8F�6�!�~�\@NQzB5�1�kR8�W��7�����e6� �����ْ����5�}܇��M� f�/�_�p���Y۪�^�ow��PS�*'��,e�/�W^j��������ք��ݜQRiZ�-
�}u�d�|"4�����fTD~e{�I��ks�W�oKG��]��6Du������V���r@�Wcle5�t��"��a�ǎ����"b:ٯ��O�A���k���֩y
�^P��}cC5	,R�W)��ɑ"�C��Wh9U�sɕ�B{�T��'���Ч�k/Ƭ��7�kֳ�q��	�c8Y�&s�mCM���lZ�~>�f7@��(�a�JL/��������Ly���C�2g�& ;���ս�\w���Hu���4J4Y���!P*Z_|޼��1xA�/���m�������/&���Cʿ(
��,@�d܈�K����~?8�d���s�s��c�8܂��l���SX��G2�`�<Tt5iP&JP�2�8|�1*�)юa��А�t������p���������7?}�s�{��־���l����M}�)� _
�o��&pPW>���X+R�T��<�V������4�\-N�����U�g H3$#6
�q�֕�,Wz}��E��ۅ��Zdc��(���f�6 "4����a�O̀�R�mrM��?��Cgh��7L�����43K�ե��Ƈ���3ylc���}�Ū�`O��b��R�|t�����.���!�F#�0�}.*:"���|�����Z:E�\�d�I�\Q0����v�֯w�j����Ć,{�+b�Q~�X0�h�(D���p;蜁�!p+~MP�O��X#-t��f}Ɏo��`R>V>�����^��]W�X$�7ˀ����KҚڥ�}��7�����*�דyRQ��#[�H"Q+���A�ÿD{�@�
��LH=֜B_�,g�B@P�S*�[f�y�1�+b������N��l�e(<B��R����(�yu�)��?����O]��EW���(jʄ��t��G���K��EӮf��_�E��vQO�e�ƻ��mՀe��L$�$�=���dr�:�Ru��lJ�]��Ʃ+Q#F�o����X,�'do;���1�~����-|����Z/^�(�͒������B��[�d3�+��EO>�/�'����H�q[�lF*@jA�o�P��y%s������y1�x���֫T ��2B3����9�T ��'�9Y`�s�r�3V�l:|��,cX�(����t��2w�osG�q�U'� ���j�wM,6$K���.zsh�G�1Q��a����H���l����x;��\��b�\���7��[��=��g�茬@X����|��K�cg
�0~;J�쉫E��c�@��dK���NW9iZ&��������rdy�����8��6畄Y/8;L\0�iu�IE�K@:��MD�k��v��o:@�b.-�6�?�Q�`����Q �.��څ~�嵨�k^�@��e`Z7�Q'������Y��L���]���V>�x|�vR�	����N\�B��L�����_�g�:�[<N��v�%��{�s:_���K��v�G��z�c`�	ma���v�u�1�<64��:d���3[<6 ������߳�V�tX���4>lFx�i�d͏$>e�60f#��h�G�lR����s�����4���ZƤ Ќ*�b
�����,g�A*N7����f~ �-��+%*^*ʀ�d��z�#�Fͽ(��4���FYa���5oi�.<� 7}{�̼�P��/3s�4��64�(����!�)g%ф�bwG�/I��ծ�����]FbR$��O+� �T��c�Ég�S %K!t��n��
�zZ'V�!��kU��|��i�n3��;*C�:���ܵå pE�#�*7���CT��+��)G�$Dxĳ�M9xgx��
�B�+n瀧��N����*��HE4"x��/"Vu�������W{�z�S����}�#�A����4�tW��ވDy�"�T�&5�	�M�4��x�o4����(��#N����랉�JCdYB�) ���-"���L�.A��Se�2�UeP}��A�fM��U���̐;n*&�oR���{$Ϳ��,�4,[`��M9���dC�i�؆�$��:4f���D�D��9e��a(��da*<����P��͜Aa~5������r}5��Il�u�Ԙհ��h��o��lR��bs�#(��q��n�Q��[erU�Ob��ʓ�S�i^�%,�E?VWM[Pr�L����{ [�b�9Q�i'l1+�}�#)�푇�D�CK�_?���]P(r�7�UG~�����6�ڐ�d�j��wt!��~N�2�T�g|�OF4�ߪ�O@pz#�)�G�=&w��-�m*�o�n�2�3��?����-3/h8"�����<� �`߶0�pؓI��4Zwc0��'���hR����[����sɒ7�?<b��?HS�5M/'LM���1�,c�m �Oj¿Z(H+��&c��h��9��w�KՊ��R�V1���:�E,}�I���Ӥ���<-K�	ꖪ&x�)���5#�z�T/�{�Li9�T�� ���y���D�ӔQH�ܖg�=�j�&>5�H�wHjIh�\���S����=���0��������{9B�������u��+�J"��	\�%l_ZɎ�ѥn��R�bk���M񺡘N�X������xR�����R��|����,�,r]���0��`P�_]�@ߌH�H�[܅����34�ᕦH�f?�0EԻ��@��V2{���#��3@O��7 -<v$�����E�ˇ)l7�����st%�n�,lr�5�
[���HW��*�q}�r$�@4� ��NR������k���='�t��t� ��C����hI'�q@��r�q5�|�C×ڏk	���I��/׃v:B�N�O�|Dm��b��m?�A��$�A׉<��^`���6{�}d>+		��.�9��W�oq���DX���&�4_�.�;��@�-iwX5�'�<��p�S��Z��|��l6��C.�6��9Q.�b��j˙4b���'�ƚ���z�Q{_�#��hS��\��Ə�\X'��+��G���$�`CNFhC3�D$�ꠁ����.p�x.!�h俩�s�8$*������e̯[�V�s��':�OY�-���6a1�#�_���lhrw��5��+�ouj('�+�ί��+��²�dG��`�fS�{r��Θ����*]}�;��K�v=��;^�C���n1�������)��T������m�X�Y�<'Oe���
"�-bI����YB�haH�/L���:n�k�����7b@{�����+itk�Xʎ�l�@p��$Ԍ�3E����-����]|�=��4L�����xi�R����lqߡ��yƻ�@hw��A�J�TD�s����s����-�l�Fb�Σ-�H�F����
~��Ѐ��f<��x�m�Nr8K����҆2B[�B��9T�T�FP�QZ7�؅�䆻S�'EG-'T���wJ���uf�<��$�а#v/`)m�#����H������I8,�8���^(�u{�n�E�EF���U�B4��;]���~��r�:K��� ����Y��q�u�	X!��^�s�`�N�+2��*�ѱ(V�E_�lG�-4oF��������M\��/�H;z�L�!fGm$��<��Cp���qm�|�+ ��rw<����3��?D�7��..8�>l����k�ѩ�Zc�����(��q����9�0����B����$�`-~1M6���ƾE��EN�{�Ľup��c���4�
��-��S��<��YGa��z~Z��`��.�Q�PfX��҅R�w㧂At�vN��c�e�����ė�� �u���5Mn��Ӽl{���N����&ak�Kx"�xƻ��!Ж�q
ȱUޤL���j��0C,�R}+Kk�O?�(������%�=�v�pP�ښ���:�����F�S}K2�A���$�2os<�x�W\�<�y�&=�ߏ�k�	$�H�d�a��҈��Q>� T_xލ��r(o��H��^_$�w��@]��������ɘ츃�U�=mp�v��L�(�L} �A �)�+��&e�U5[�9�y+PQ��7ʙ�W��O��%�K���w��$��Gm	|�Je��6.��@=��T��X����]!���*f�}�:�{����8h?��BUE�	���'�k��@&��O�(k�iE����^�vW� /��id�ec�8,�2��#�?t.$�݂���J�[� ���%���I0g�QfR��L�ʠE%�'�����XBt"[#���U�2>2Jߡ��#�pE���~�+V@�8~SL�ɥ��/[20�I���l]U�c���ҭ)w��1�mY���;b���������H���T
`ћضp����"Ph�J܄T�Q��sk��7��jp���Z���/u��K����@����P�V�k�2��^֦|�Bq�����K�j����D͡���ݷ�W�yJ�z	����阐2�B>V�Z�d�ԳL�i��Q��z;Uo׬Zw�gŮ�"OiR9�j(���F�7_sh��}�l����	z\[�.]j�
����O�k���q쑶G\�Ϥ������9AH/F��v<�ֲ�����S���!1B��X|�(��~ˎ"��]me��U����Y�IՈ��Q��+$�]�3�Ոk�#_/L�uR���ߛ�ؠ�
������p;�¹4y^;ʊ��@tk�^���Z��6�gDp���ϟ0���S����e+�g����T6QƢ�4b,W��g[�u�W��J �B���]w�z���e�m�I]�8�f����fKԔY�^S`u&J��"�7��ɮ�]E~�����I��^�\�:�7"2���[���E��%�xܜM�ǔ�2�?I5'��Y�����4�@J�d���r0�D���ȔRZ����-E?���ss!5uw��Gm��d���ٌ��6Gx+��(��]��1��~��b1W��SSv��47��.h��� �Ns��/9���>�<8Lc*��.���ԊC��he��b��� �60O��:��>p���R�04��a�Y
t�^{A+�@~�9����x������ꆪ��P+M��%�bІ I��>�?Wb���`P���c]ծ8ڌl���p9 ��鸑���U5���N��=#�����;o�#g��^/�ʑnZ��ߠ�S�~֥�IY�j795�EE�:�vʍ�����J���(�h���`-Y��?Ё�v5O�@է�Tp��FGg4�Wf����qӢN7�=ɝ��y'	~��#8�M4���C�N?��{K�2�v�{�"����e�"���Е��H����#DH����)���G�A�ѳ�:��Kwl����3XiKu�F���0���5s��&i�c��jU��We����l�M��V|�G��r�o�/0�^끑���d&x�u�	�aG�.L��L�f�b�uM䈅[�Li�<��ymxzG�z"�k�~�t��8�\%� �9��\�e����4�bD�����)������1<�R�F�34)m��8ι-j� 0��@�R����7C�r�p
�q����	:�T����r�W}�
:i�f���kF|?;��]��-�;k�:����ͮ<�\���9;�ٮ�"�I�>�� ���-��]��Mv�./s������f���E?
�ʥӃ˥f�d�L�]���23L��pr��_iEj���/b��	,�0g�At5"d��ɗ �猾�~L�Y�ӄ�+�~r߳C�nHfĄ}�h�� �n5�z^�����2o_�WK�Aׂ�'	���qçoq����@�}���+^��e��,� ��Xd�Y(�9�.�Aٿ���v�ڌ��_����0�Nw����2os9K�����,|�e��b����]a kv�tUލ��!i�7&���I#c���%.��.i:�H�D����z�5�lHV����y}��`Y@�N���!�viP��Ǥ1�t��eє�q� �ቘH���e��2�I������w��W��,'3���Q����v��nf+���o2�BȂ��������D�������F�������x��� ��9���\�m�`�� �i��;�L���:��Z�r�mHK���)gj�Y�αp�Q�Tb]�k�>��<���p��uҼ���4��B7?����A��2��a+g�V���*k�s2�'c�:XdS����x�u덺�XOG����w7��������y�8��T�<%�~�
#ܾL�l�l6��Z�j��Ga�al�KWa�@ŢD���?S����X��,!|���B��UA�F�Y��S��M�H@�a�gE�H�3K�؏_���6�X+MY��X�����ģT��5`������i���K��ƞ'Q�N���!����ҳN�I��f��K�ńs_��<�[�B�:�g�̂�vh}�������=:��jj����0��=F.��[�O|�/3��s�o�|��'M�#Ӳ�Z[�cm�y�"Gi�t�^��^��14��Y�?�I+���<��=ϗ&�L�jJC�Yϭ��鍹x�W1}=���Ǹ��2p,C�n��fP�C���m��ky`}y�
sI��F#�g1�UO�X��'��F����cP���tƳ�C\�徥u46-�9&�|�R�T
�oT�������~�������p��
a�o��3ZoJ�����O7(��ə<?�0t5-cc� r'�+$�X.��4�FtęV<��Sf��kCMn���w�XF5�U���ڈ��i�կ����Qt5պ`��l�7��R�q���,�B�������W�Ǿ�%������:LU�X��J���Qz�@�2Z�3j�)r����;P�YeH���cN������Jr%��6���e_T9	O�8��LWA�zF��]��x8k�#�Q<������_�n�*��3q �@(��/:?��:�JM��8ק��y��q�U�:�M�WcY1��
�O�c����:u�\��� wKA
x��.���r�Q�	��5+\ēA��l����-xf� m*������o�WR��L[��;�4}?΃�U��[{�Pb��⩅�����}���G��1D9Z���C'��v*X���ԟ y��m�K,�x����Ѷ�9F=:�/��t/�u�Twɮ:�@������[p��|3Ԓ��� �2��`�;���Y*�E��p<k�VYdR��d���˕1��d�Ec�N�I����6����w�G��ٯ
h�S��,Wqt5Ǹ;qMP�|)�������9��n���]r�����=�v���G.$�g\��Lf#�')j�oH�� ��=U|8f�C��<�ڻ���؊=��!����)���P}���V��-*������٤_�<Jq�[�o�bB6*�Ac� �QD��/�_V
������bD����-X�A�0h8H�¦�鰈�r-���U,Oo����`�ۍH9H	[H��.y�_o�t�ݾX�U ��2�����>�!%�VT)�$@x�k��hَb��&R��>�z�P��z{񤐱!m��ң20m��P�Y!X5���4׉�fv����8_��
%u��f���A���?���<i��}���%��dh��o�/�y�D��v��(�NH��$����%	vۡnt��!���s
�y�f��6����*_�<w����x0J~>��fo�J�f�(�L�<�0�#��v.p ��0Ɔ�P3Tˡc$���|w��,	U��[��D�y�A�N��v=7b�ӶS7�	w�~\B�C=�+�s-��4�ܴ$�|���?D�L�8������SF�u۪A� ����z�>�b-��q��V ȷ�9��F�0|+6�u�M�h{�$pE/[��#���*�#ks�r�i�.����//9z�p�n���y�;���+�[���5�,���<��Tc��T� �?���;�:z��G�bs�<�.�S�jn�w�hD��1�|EGs���ElOu坓�G�2B��S}pw��!�PƱ.��Y:�Bh5%�Eߥ��=M�{$�D�[/�mê(�������Rl� B���2w`Y
����V�l�Ⱥ�MQ���kb��3�R��󗺈T|8�w�����ۈbT���t*�K����bO��<x+q�p�R�=reSϩ��n��?OǕl��9s�n�L�U�	TVP4�kڤ���!?5��]�`�%��+�#Ƒ���G�T�b��ot!�呐��db�欧��z�".+�1m�|.�'fD�n��96�W��N�,�٧�oƳS}�w[���t��_�6��S�2�M���W��7����U��kI��� k���(@�
�tT/��'5)����3l*
���Kf@�w��ܮ�5��zY��䌫�~�Wk�,�����8re�}^  ��I������L��.R�Q�Iǥ�Z}����dV��#��!C��h�3���	&��H>1Y��[:!,���Ȍ$m_n�"�+��'	AeBs�l)�E{��+'�Y^q9?�f1��@ZD���P>o�k����
���WJ�'�|�1�W��i�m<��C7���N��KCvs=	���\��56,��NW��K͆Џ��.�*�x����f~{��]%Í�k�I ^��O���A=+���h�i�vU�����������؆`�V��L1u�o��N��7�Փ�a[���`	��g�p��cM�v�	��p�(Q��q��1�J;씑ܪ�C��G!|a��Aht"�IN���w~Y����Ox��É���>���`�<�\Kgp8�n��ߊ34g���B"=VE���D/�}K[�4�~^>����c�):��^0֛�k�og��;�|8}�-&�D<%[��u3�<�v�L&�F�&�Q*Yj���0�� %3~��[�<�ר�e[%Z)�	�\�{�lUE?k��<ZEKbj�hіّU?�T�^��i�f�JbW���������i$�kE<�h�WB=�_(<��AM�M7u෠e�8�����y�R�W��ID~]v�Ջ��z6��<u�O�3�r�z}�
��5[��UI��Flp�ɅQ)D�ߋ~��S���F>b�l�8�R
��b�%u��`�ݟ��pߊ٧�hg2�W������f+RXQ�ɻ�+y�C�]�bН�O`��-�oͽZ
b��C����=�DB[���|�܆/�)�R��R#ᣃe�Lk�3����`�+:\�6x��P��s�Te?�4KO�Ϲu��!4y���JX��+ ̓��^��[ߵ�1�]��A�ͪ��+�B������Ca?P.�>���`~�_���D������?bk�Z5��py�N� Φ��`��C7<�X1'J7Y�ª���Ï�TB��4`������9��#� ���ER@�7������$
Ɉp�gy��G	���������V�I�=o��.�]-}@�0���Kۯ�â���{�R�LB�"KI"���J�����N����E�&ϋ�'����)�(0�2�w� wR�,��~7��*�S��8�2�lqE޴Qun�DiIx�D�^��N�5P������D#�l���������'(���F#]���QXv�Gr@d�Fg4�:���M��]��41'��QR���Nܪ@��z�*��lQX�^�S?��F�M�AӬ2(/��Y|�1Q����
#�z��d݂�7=n��$�;�|� �|$����ߥ_�ᐼ��!�񬦱H������;������$f�G�k`���G�#B�,48�J���ᨗe� F����(1F2/v�ږ�{Ռ=q0a"si�,�Z����.�sx~�ߡ�v��a��1Ŧ�bPd�2=a#Tg������'G:�D�8��À�?�I?(:��$#���u慾0NW,>h��+�ލn�a�j��a*��FLM�.�*���7�!ĠٺG���楅ԏ�SW��I�?@�z�[�TH9]
�a9��w�+p*�
:��ȕ���&Rjd�6�\o�����G�O��ѻ��W:��%�{��6b���j7����,��!�l[�g���H�ʮ�A7ëski��L�l���|=�#Hz�Y�����+To�AƁ=[����2�x���~�,��h����-���+�����s�V��H��W�Y�%�Y�SD�\s��%�M]��
�X�g����ev;3������JtKJv����J�G��X��Bi���Y���T8�DMp(K^G�6��A87���b��o� %���A����&r��]�_�u�S#YĢE�!�N%�ޮ��n@�h�OV�$fG)(�p��0NMk�k��I`{�C����:����S�w�O��4��%�����G�D-b����6�=	]GA$TC���9�^R2�r�����I�ԑϡ��glh����)!\�z�kjt$%�\*G���e���R9�k'ͷ�E_����0���1fyZ�f� ��X\�Ҏ�o�@_�#:���';K!�i�)m�=ې���H��K:���]�lM�
1-�� �����ww���E�v�o2�l	�z����$�ZL8�2�u�I�7�(�˔OQr�-K�卅�N������q�W���bv�Ǜ4b7����!�l�7
6�ц�u�A�P��N4=z�m�7�mq,'j��ܪ~�LZU1h�o�t�6���@�c��x�3�v9?�U���TM��w$K*g���MYXu���*�IaC�2�d�巢M��������?���j��3ڴ���}����m3q�yq#�GM��nȘ�ЙL�|��]�H��î�Yb5�h*:��-]�:y#���8����5��@S���1� �l����Y����f@!#�J� ���k���h.���f�q�<Wt�c�ݙ�ߊ�σ�����o����3�Zn]$�W�ƻA���)�`�I|�iX�.�W�Cuf[�[7P�=��"�2]�}h�gOTN�B����V���UHV&~�I5�
=���b�F���t�Y�ov|��"��,w�
�A쁌 �P��L�E��*�.��QDvr^^�̸��65�N�P��a6N� �/_�+CS�XS�!9-3�x�?b����p�̅�Sd�:4{~̉Ġc��P��䵡�����C�N��Yy���OՖ��pr��qaU�ef�� �_/����|u�#��e���ڭ`N�Z�r*3��8<a~�H�Q�^?�l���+	�2��zm�I>�b�6K�z�䬷4s������sc���m#w��e�mE�4��k�1���S>�C�t���Q}��֞� �q�Z�ɒ+�7G�	:P)�|��#}|��0��"<OWއ$�[s�<��Ў�����0���]\B�-���1u��WΎ��w<�l�>,�d@+�){]����O&��q󌶟�*Q4bUdq�������6��r��mXa.���)8T5x�F����LrVgf��e�&˽l|�y5|��,~�3⡴�AB,Q�p�:Q!�0�U�Z���&�~����5k��6���[��N��c��i9�O�r�@�*�{���n�.Y�ޑf5.&�=��L�)y�&j15��װ �Ŕ*6+pPG�l#~v�H}�2���:-�ҷe �L70�a��b60���ņ)߅�����R�co�CNփŴ�����a�(d����W_ce��i�����^BԦ���5G������eGL��<A7TrG�d�u���hʒ������Z�tE�9�8)��6��{$��n�Հ�؊n�_9��0�Ψ}_S�25vr}..7>���c�\U^a�]�A{��[}��2�}0�}X\ӝ)�A2�N�E����D�kR�/��9�c/�UL�0"�g�^�m��j���9�鯪��Bl��(�E��`ؒ|�6���_�c����2�c��p�lB�783oችMj�r��� QC{��C�3�C��<��:���{P���%~�)�>��Y�1,��8��02��.�V�/a��qՄ�[�Q��}Z���������zAB�?6�����v�H1�o�����}��}�)$X5�L�R�H�-����� ��ޖ�$K ߭ZZ��"�t���z)"��`��k��3_1�do�ǐ����CVU�<6@W*i�.-*��/佲����^�hgPT�q���1��G����.��;S%�7�+J���w ���H��tH<�����O�L,7�8��k�E��4��M_�yh1��R��k��� LI	�Q}G�����ө�<jEpϧ�#�α�"K����<��t��vb�����\�}�C��$I���1�r�o���~)&.�4afw�4!�ɔ /`����=��>x�A����p�)s�����Z�%�g�E�_
(��[�.�bk�x�t񎨝�ɤ��YV���W�z/oE��	��J��;���w2&���U�m�)��VI�M���F���+��$Q�_L��ޅ$6�%�ۣ��@�Z�RO�8q�����.�`&Tp4J�L�ַE߉�)9�����s�y'͗�l�썎��'�1*�S��JTZ�.�|$�)w箳O��g8�2#�ZRE
��~�]w���
l��)�F~<T��]�;�z[�AI)[-n�c5F��\@���ٯI��9q���]׋�V�_t���e)�>6��&J���*�]���ߚԝ���\ON�9
��o��O����/�]�ah$z,�e�1Y&���X lk�	�A��󓻹�"*mDh��Y�D���!��2vƫ�[�
�x����������ѻ�4mA&��J��X�D`�8�^}�C+(G��G��N����Ht�����w7ʾ����v��E�A����� ��l'��`�8Ss�"'�^I�Q�p�yN��ޠ���Fh��0� �I�w��?���0{Ȇ�Q��BZ���Ȱ�::q��Z����Z@���kH���Y�~X����L��8gŕӒ��ˎ��<Q��ϵ>� �[�3!���%Z� ���o(���qg��Lwh�N�DN�!���'��? �'J��&�\����{�C�	cMw��A�l�r������-PwKSP��;RiU�p2�ґ�,��a��K�Y�˨o��t؍v��CE[�WX�с�C&��p�[��t�k}�lP�!���(�}%��W�?{�KG�M��[,���ն$����n�V${r�c]��4���u�	�D��B;;pJ7a2Ay��[�A����F2	V�h;�fZ�>�I�R(���X-`�B�{���1��|뙹����d�m��n(y�=��=��iڌg�6&�$U��/��ʒ�՗��m�E?EN��*���||u6�|y���\;�v��47AR"+A��RkCwB��[6|���Q�ܸ$X�G������E�{��D�o���E��X��0q�# o�;�ޅc�֖Y��)�6��T�?��0��)I�s2��H��T-�R �٬��=nD"�Ҥ�	г����ֹu�ǉ/��6��ف��Apn��r:$��+Ysٞ��^����x�����1,���GEn˻o��:(�q���U&��+�!_���oi&�\�׸S�DI�/G�z��o�E<a�N5��e�x�;�I��J��-?,˪e1w ����#y�h��p��g��\�����=���~�"�DO�f\�3�Sl+/Z���𵺂@�jI*�1�J���T�n�j^��[��Y~��x �=�蕺�8�S�?��H���ýwI�!�%�����塞f;��!��Q��C�K��V��S�U9��<��g�4l��!ֆ��8�#v�L>�,��V���҂�)�[��ov��݀zq�5:1�7ZO'�tD���?�P���%<��c4d�}��#BXa���vk"$j��8bF�SJ��C�O��j�̸���ee�X��ES� ؠ`6�w|d|ռ�b��W���l��N���d�o�.�6e1���\l[<���e}��6�I%J�@xk���u�S��X���g��JS�Hy�_]p<Y{��\�����0�L���������-yO�9�|��V���@��0��U�}���mv�Z�!ʨ�Xh�*G�eqe����d$�\`��=�)I</�]�k&��S���ݍ��%��eBfQ�nu9OMy;��J����5�2e���Y����2ލ��G^&7w9?� �ւg�3��]A꒚hO�0?�D���{lT���A6�f����ud�8J�1������r�A�qF����|]E��y�|�QR+�ia�+������_��¤~݂��م��<�E�MvdP�8��}�d�;b&7��*q�~���	XI�S=$E'��Y�F��vuE��;��؎'l�>��KS����XqQ���z�ȷ�`E����kS�q!4�#M!��Q=V�2�\����OF�L鴺�d�����2�OYם�p\}pHq�(�%}Bi�&`���>h�Y^Ŭ�c/7x��4�P�s�!V	ey���ߟSN���>���H���'�5�����|�P=�9��Tk���:�;3a_c��d���ΐF
3��6�.D�Z�!���>��C�f.��l4Qs�Έ1$�b^�� Q���q4���y�`�0;=���rUx�7�%
VJC�H��|�O.+��C��D���vh�&�c���i�<E����[wkS��U��.X�ܼ�l�-⶯#����w�{0N��C���ˀ;�gG�7���	��T��M]��),�Ty6�q~���0�����D��[�V�7�Sz�.U����T�����2�v���W+�KZ4!ܶZq�ȼΒ�@���_
�+r{��i�gBJ�(���E��$J�^oea��7�4t���q[{�)�Nx����.H�������L���Ƣ�!�]v\��	1<4*_ �X���{�Dڦ
 ��ي����@
�X��iqW��z�h�gU!�>���b��L�"Wt݇k��-#;��RgT�bW�F@A<)��**]4�6b(�A��VvEeYkY��دe��Z��� ��yX���$�q
��O!,���ж,;*k
)�U���|g�����P�hL=�=�l�ٔ�
�&9f�Y���u�7k^��t~u��5�����|��i�����', �ٚ_j��pP�����Ɏ��On��e�ۑ_6[3I��8��3+�^֩�Թ��_[/4Z��1GqZ0��V�"]��;z�����.��U3��5���1ͽV��^���s:���1b����ȠN��@ qg�|vl��%��{�����J���.�ۜ�Ɠl��ߙ�b�OY���ә�O�;ܻ����vfH�Y��7e��}yz��d�@=$/��\��E��0�GP��"۰@�K��ws���Z��%�2������SM�qJ����A�)9�~�*H�-�����j1$Z&]�R(O���>_%Q�Ű�1c#�"�Ҝ��]v��uϙ�Ə+%Wgx�T�����N�U���/�d\��]gTV���&�ZkT�����7�x�f����jJ�T�"�l1T�4��-Y�ZT�"V��I���
2��ϝ炝
*�h��`\� |U,Q�a��:�-�Sv2�3Wwt������>�fP�C�垺/�#:Zn����0�t�W�Cɢ��Й@;W�?K�N"G4�J�l#	u$�[ʟ�� h�,����]��E��f�O�s)�����b�f��td����x>
��M54��A)��P���m	���R���a=���y�t�����$ T/M��ߜ8�|{�$)穉C!�����,���Լk�B-Ff�.�*9���Z�PK�9����ķt�����HQ�'d�� z�V��Ig�Y	�Q�����pPK�x��La�zP�/m咥(~���xf��"v[�d��G���P e�@?Y���t�Jĕ�H�[��)��|}�v��0��0�7n�'ý.�.3�ha�RUΘ5��_�¯�_�O�w$k�	�}Y(���I�Z�ɣ	���}���zU��L�*�/K�� *�gcg߹���e�pȨ����<��*C�:�u%�rJPLڧW3qG��/�uJC!��{�526�ʄ��Wv2�5y2d�4(*ˣ���}~��!�̪{��ʯ�_G���8n@�{�|���:W�m>DqX�3�]�M�(�w��/,׎��ܱ�iW ��A�)ѯ��%8�<=�CV�L]\�W�d�{������kI
��y?�d�`F%��f�_0�����p�8ÿ�j]E~<9	g���� �J9sy��L@rЊ�b�	١K���<�U��̝�Qcjl����/�s��D��C(�nA���hz�qĆ���6g�~!�oo����`m+'��
ٍ��q�K�%Q��`}���7m;�����6��P]�@@��!۵P{�2I�S,0<��"�����b�
�������k?�T?zwS%��D�Pшh���9H�:��C����D�����C�Y+
�C��r+�:�k�%��f~kz�F�C\Q��z"�h�8{���݌��''ю�PU�K��ǑH��B�vqO@"�n�j�/t|`���8$H��wr[�.�Dw!��r�ߖ�cM�
E�{��,?�[<�|�y��b���I�jZ��K��e����+ޓk�#&w�a�/k"���/���JB���O 0s~ݛo�K�Z�n�(�h�TI��g��S���U��F*�I�}�t��Hk����2تB�����/x�Ε�W���� $���7��~[႕.��m�(8��O��ÃA�,u���sԞ�	g��Z����J ���(���7��:Yd�8=�xz ��g>D�$
��7R7���v�.��H[�&dp��	�xr	���<�;҄��Tp�=��V���:���r��Y!fK�E�G�I���V�h�}�M�Y��H�_�Q|��k�B����bb}�=��Hֹ�}���3����{����B8��59�>f	�o�+�ӲW��D���C"�>�r���N�+�QD���USa0�>��_0r���U7�n�|oe���z�?L��K�'���OɌ%��Τ#�.���+|���e�a(�" ���P�u��_&�̟�A������%��A��L�u�׳�b9��Og�;�0���+�H!�����*iD��QfZ۾35�q^�m)��:��4\q߲jǔzlT��'�B�(ΐ��\���_�]���۱����M��K��sy��9��pa䉾"vt��:�U5��"^��W���,g��-h�p�nJ�z�¤�&�`^������&8�M��Ǜ����I5�:[�^��8�������x������I��C=����}�k愐�>KaAc��&��?mպs��ߎ���tV��1A�75����5�*d<Z)H1Wu�E�R&�N��f[��;f{8̻|�I���?r_A\���k0�T?������*�30�o�X��i�H馨�]��+Ѓ�A�����H�������r�WA�oo�����5��
�9�^0,~_n�9��� �������9�"��ݛ��s�غ0B��kR���lɒ��z*�$52����jr�2����M�	�<	g��6ıCs?�߱���;�&^�9i��Ase��q�����U&{J�&��\�"&�����E�?���c�j��Qf�8���(}Wq�Z{�K��`�/H�3� ��RT�WN �����dsШ����ْ��c�]���(�!
NTN"�Sa�mm�;���v��ȹ@7�lm@�t�Oe.��~�5�b��eT��g0��T������>���h>�������0��_aZ\�<`�[j�I=p� t�=���Ҿ��=
��O�R��/�jo�Ey���n�r띪��xj� 7/O�q�0I��<)%(�C6T��}E�*��)���������*��(�h�U��q�Y4�[u�t���\9f�i�d��^���4bM�?����h7�H�J
��}?-�� ��
���@Rj��7VB%��W�7e"2H��y14��|�@���p
 ��xzqV���f��.�E�y����rP�d����[�~��$ߤ!�6��AA�"rt8V���S"\nU�`��?�1��Ts0^D4kE*��L[@�Ӥ��#��_U�2����� {���8��w+"X	�_���MD�M�a�P���>�l~���$u�{��fo�ouv��c�������&�(@cm2M*����E4�՞\k���ob*���.L�[�A<��J�����H�"����R��N<n���9g.���Wg�dS�g�I\����0إ�}���8�<�]�l�	|�xWh���VeǔB��v@�����ٯ�Y3������y�
o��j��p�$*|q~�1����׀ŸZ�M?(;�k�wu��Y����>[zg xR�k'�h���-��A���׬g��9&�d�՝�@�x��q�\��.��ڸ߷r\|����ʔ+e�J��I�׭:IK�ar��w�PF0.A�KɅ
���ۦ*ceN���ءvUTw�N;C[������9;�A\�늮/ԕ �ά�;m�bn�9��s���6����^�'�Hi�7�ISݲ!�~<w����"�63jY3�)fTui� �>�n3}��#|\����'ux�b�E�ت�j+Կ�6%M�٤|��be4n�
�H#�����*������:MH �:ؚ<�TR���L�_%���`�K^A+.rCfe?����%��7.G�y�2w-ӡ&gn�ɋ���ݖ��XA�Ŕ�e���f�?�p����]���C���MB��UqT�^�ĴT�a0˓D�������Y6�d��2��ߞ:��O�Kߐw�9��Y���{k��7�C"[`�h�L�cM�d���w.h'd�����[��D�8�(8��C'�'��[���(lQ�r ���+����=����,�0��ih᷃����D��sې'�'ES�)Zd�����f닓`7�;����QЦB���)~ѕ��!���$����(5[jt�h��%xe-����Z���b>o�#�l'��Pb�B}����u����S��,�9FAJ�8N��;e)�S!	�t��[!t5�9���5�(?Z2�| b0��р���!q�qs�p H&I��{4ܾ����������X��
�zѯ�s�H��⢺�'"�����|��Dٚ�a��Li04*�q�`l����K�=��Z�j�Q�5��
������q�u���B��	���J/�;�LEI��R�� �_;V�y�EP��X�O).�O�%�A�,2������ƴo�!��	�"�^HVi�"�H��Xi��K$8+�8�M��k~#�mJ�����?��n:��z�_g����S��m�p��H��s�]�8�zk�Pe��䦈 �d4 �h���]<J��}:Im/���\x}�)�6�Cw	�Z�`M�\�g��.C�9�a�(Y�}��&9t�̈́ò@N�4V�X@5�vFuJ�I�*��@0t��cf�5k�h�<:��(]K��o
� k�K��Y�K���d��x/+�K�r$�F�� R�ѫb��f���s�lΊȗ��T�:�k���*�k�;�獗m��:�Y3��,��5p��,���tL3�l�:�t�;�n!N�[Y��D�ej&:��.�6�ɷ�X�I����n��+�Ȅ��M�c���Q��b�#�8��F� ����[y��kf����t�f�w �C�'
�U�[� ��KF���_ ��e����T+��ʧ�g&j�������%	NQ	�
	��xUh���)}J�.1�+����^[��l������?=Z'�.�Vu������/��i8��ǟ��p�n��6�Abam� j-��i�s�c�\��k�BbA[/4A�SР��j���d.`����"�O<?��"u�FZ!�u�����+RkV��UIk�E{��� =�So�%� �ݦj��ϩ��<ز���2F^���`���%h��o: 1f��3��L�qIM��������΍Y�	@TO��pG�;�
�s�ՀlK�?�6f2n��s:���z�)web~�������6�K\oD��z��w*�z_CJ�<���8Ok�V��V��u���h
���~F�Ri\�u��E�ř-�����@�9=�+F�)�ԡK���_�Um��1=���e<����͘�&�І�fSJ
{������Ҫv�*P�rs���I,Ǭ��)��ޫi8��jc��߉���,�Hx/���	<�p���g&��F=���&��0��]X�����ϪQԍ��<�]�	Q4I?F=(ɧ��X�O9=�3"��eG��Kb�;S]�Z<_�#X9�mh;�{���ڍZ��HXw�X@�tG�c'L�����E����5�y��~h��Y2
�45#V�u�P����<m�m�N�U �YH���/\���#|x�LMy3���#�FѬ�l@F�� ����
���
u*of�}�}U��%q⯹�9����@M�#6��B�o�Ӥ�����p.W
-񚹍2WE	~Ǿ�f�z.��h5ɞ�������KJ*F��R���s��7P�*�Āp����c����T��j8b��/%~a����HqJ�\�|1}hF,�Ҫ��w�&�˒����< nLe��ǘ���B�WG�Q��,��=�����g��K������x�.'e�-fP@�iT�/���� ���7B5�����y��wAD�L�!]B�sr�J4���J À ΢r���-@6/�f=��"��7�M����F��]�դ=)������=��ФĂ'{p� ^��?�Q�� S"������,,g�1�Hf���5=���7[2�ђ�S�ڣ�^�al��b��_G�TӰF��
��*$A�S}'8״�������$	a����y���)F�M
��uc)׊Ʈ��g�8'ŧ ��Ȏ٢W1p��[����,�.%��:�Py��vͩ�%�(��љ1���N�J��&޴�*Oб~H�!q���Y]�A�>�\�&_����r#M��m^;b��<,w����٧΋��D���
�������`����,�jn�:�HN>:�ζ!�U���Q�����<z"Q�� 2����w��:�N���`��N*����������1�)�� ��`R4x�"�Mq���G,`miߊ�H����	nQۗ1������&jD��}O�?�p9u}T>o������a�W�_��7;�R�J(x#�L��*�� �IR�j�L�J*@���S��<�W�����)�;�Lω�'�<r~ˏ��MWt�O4��)�;79*�V����ń%�����'(�>����x|���" <�׶�-0B��x��L�Mbn}HzI.��p1�������6~='����DhX�Sѷ"HH���p:wV.!z����2�cǭ���re�!ƑᘚG�O�H��Y/�Û�AKST�ơ�[�19��㿪���zL��M@�p�m�G�jA��Y��	��]���Б����.��SJ�j�=��*R�of�$p��q@�d��"�ӭH:��<�}�k��aX���N~e>6�~����v���4�PT���,-�X�r'�B��$d<�W���h�X2 �s��!�|:۬��`��+̔���iQ�X��e:���R*�Ɔ�����ϫ�! ���&�2s/���JU���t�pFIm0l�m³Ӝf@��
��-ߝ��n�o��c�ժ��n�Ӈ�o{�r~.���ݳE�$�g �,�x� {�G�U�-�ᒷ�R���MGx����������R�B�K������4����#�!�n+H��<IGQcAX�o��6�	�@�Q��l
�!�C)��k�ʒ[���Dc;��o� �MW��@���$ugEy��َ���?� ����&u��#;�y/N��N/���A��ޕh`"�L�b:T�����O��)ԋW��4��9��N���t@�pY��v0�*��@	ks5�%�>����i6�Pc푵Iz��m��R�5@P�[s�ۤLџP��D��������,V?0�_�$@��0;�澆��IO�2�8�f���;�n�b��]%Y�T�i1��^�k�,"h���`컩�w��L�����?|�ӥ��Q�Z�ۘl��)a�� �(�,��K�{��l�\�!ÇA��:����]O>�0��87d�U+__XnT��;C�*#�����>�W���6m�?�l�{JtT=Q�ʅ�[2L�ְS���x�H]���s�-❟)��Tt�b#��P�Sk�/�\n��9�N8��+d�?2�s�"n����Z���¾������E��Y>I�d\��_�v�ő�{)�)�.����P�#�x�/�5��,ij�ɯ-)�����v3w�1�M�i�� ����h����f��"���o���/<g������fb�[�!؀��ʶ��*�i��d�+��`K}��� ԃ��aqf�MY��"�]�Z��\�骭Ҋ]�r���x��B�����(��D��	�.���"үaD�E݈��t��IԖy%��N��o�C����ӡj�1�wf��SCQ�Qly��f���zr�7{cC�*�r��D�Lx�ʗ�Pu�?�[(n|`+&r�2d�����Ĉ-�n�����?k������me�s�X���Բ������,�8�o�ک
#���GoV(��*BFsLN��{>M���v_�E����.��K�@U1�e�C�&.UQ��β)-�~�ɾ��Jn�p�����flXp��4������ӌ� ��m�`�n��)��*���X���U�I��m������Q�i�r{՞�]Pp#9�(�w�*��g{����`�5\v�Z^�)��+@�:3eֈ����G����+OlBg�p����jPb2 ����Ha��2���9��П�J )�����C;"1QFY�����G�~��'���N�_�?i�Yza��1�P��H��']���@��u�%e�ˋn[� �ޖ�1݃�y9�]n��8%�ꈭt�gb6�7^��+
 ќ����V�3^J&���bV]�b�n�����Nz��c9�ji���v�f'����K�>m�]�g7�T�:�/	�"��aG�e��pD�h�!�8�!<~(�x�u!�*�W�=���cm��| ��0��ژ�7lQ�����stZ#�o�"R���y���.�ܡ�� �J*I�3��ᰳyk��R�Db�{dU�K����#D$�Q`�mK4$DG����9&Pc���}��`�P����D�������Ҩ:�X���u-<����R��
C�f�>(���k���?�i��Ø�Xշ�j��2�'m���8��(UH�=�Vm���pfܐ$����E7<������,L��J��t`g�9�|������`lZ�/^���->M`�X��Td��l��B�R��Q�l�#�� �$��^Ӳ�,n���X�岦g�:L{M$>��A����� [���@�<3�W�Z^�~R�|Ό�L�}۔,s�t���H��Q5��z�^���m@y�o��<V�!����d�	�*:jz�_n7>���8�q�L�y+{6"��Z�ϑOI���G�DPV�Hi�j���<�?k#��yov�W����&�Й(F��L��B2$�r­����j��B��i����{�諛�ßǑK��ҡq���V7�&�ι���ɾ�y�?�Ž��d4.b"��`�:E�޾�ed�5�M�0Reۅ�X��u��s�/?����GyV�jrDl�t1��s�:��������<Y�)e�W�Z$�NL�oj�0g#��%�V�4u��6e)6%z�	c�A!Rg�w��qJ11O)�����?ɇ�)�V�or��e��&'�(�=�_vc�W�8v[�7�C��E�����
�[�Su�Х��!I<��"� K�����ɱJ[�z�@R*(�7BYh¶������0a#�o�Oc��,hQT�����Z�ӓq�����9c�k�	���Ψv�/mwߺ���(�چ�q�ս����V��U�&ȁ=�V�:v��Pjl	SG�jD(�����v|7n�t?FN��ǔD~�,3KM�eHZhv�??&<H@�ʨ+��p�����?����H��?�H�I(��
/��J���<�N\>�40�WQ�E�#;+>UV����"�ų��}�Qu�\`�>���
�K�"c<�:�t�q�
-�a�3Av͚����>�oz/�ʹ�Nw2V�l���:����3i1�[�W2$�i ��_�����b)�U�K�J/�VT�)�p��qk��1���'��6����z�P�ȯ>R3E�*k5���e�>.\�!'�:mjD�}G��i@<��s�0�yWҿp���P�<��H�*�	�Ҹ�1n�3�G�|s�-/��[p���k�ӹ��Y\��t����x�{/�܆��Rd]RI?�[�0�R�a�Y�AW*k��8�jK��d,�A��+��3{(��@n���N�_�� =r|Y
 Lc �QB�?��Q� R���Y��*J�����_�L{j�l�J�4���̣@K{#adܑ3Q�Yo�Fm�o���#TD/'±�������#�P��T��*�v���	��鞂,]i����n,�P4�39��|�=���-7Cy�$VB10m-�i��j��v.�L�%�yW�̕iVTUR�(]�R`"ޑN9�L��fU���C�=I�<#�n�t����.(���>���RgQ�;eȈ�lx�7�(L5�����S%�W���Qk�.�a(&��Ԋ�s٩�Z�	u�c�TϺ����{|R�д���i���,����lesg���I�*�.�����i��EH�tg���T��|��jD��k�N���h�n$����@^W
�o�&����'z-�cT�k���p������w���m5�U�df���A8VF�I#�?J�����<,k?�6��������ő?a͛s��d>&���� �A��J'�K���o�іƭJ!e%3 �T���'Ah��3k�6$gL�1��Y9d�~����0�����Cf�kLß�D �t�2H�H)�BA�, �F�*��#K·�ko` Қ�;��^Y)d�_�2��$�s~�cj��
i�e�kE��ۿB�P��E&��Vx�թ9��&�h��s�����uLO��v������#��!�]�H�fy&���Mk9����覄��E+PQ� ��yi ��U���ܬ��SQ�q�QΤ���;|h�#���+_ר�^�z{5��M�]�<"P���R�N��p,��r|)ߪ���6�i��W�35�t�r�Nҭ	F�Q�|�299% ��֧��!§{O2�<;���<�����M�� v�Ɋ6l�eս*���p�����.Ǵ�kL�]�g?�D�����/�j=Ώ�c�O�'z�%�|O�o�i��$�er���7v��:��+D�,7O�����R���NL� <�����R&v�F���Mq&���l-�o9%6��Ŀ�%��
�ѱ`)n�E7��ST{���I��3�Եj7��S���W7J�w{L|�,m��X�w���o �Ԇ��=�.��٠���!�X&?���\gk�R��{�!T�g���f$����0o=1��3˲�ux�\�|�<�w�cC�A\��pk7��������2��N\{����f¡%7�5�7��?�6��
�ENӂā{�������M$koAb�ن�A	�D��B�T�������T�3l5]:Xk*z��E73�E�yck�5���g �����U�ǅ����2r�^�l��,ywve���2�O��� �s^h���5P�t�����K�В6������c�5�5z��K�b�X��2���H8S�с�7�է�8���{�e�&��&I����y��- ԯw�{�-��]�0�N�Y�5_R�!r�]}�1 ݅��Z�R��9E�/�g�^f%���� ��7�s����'�h %�����h����,�/�D�.��>J���X׳
��X�w�a�~040�6g-��}W܀�,h�'�wK&�/X��cAk̻� �	>��z��X��b��F*{	rC��k/R"�"��_9�j��ד_�?���``���x�_�kS�C&�����'e]־��Q?^-���N�E�Vi���8���O�!~��# n��r���6a�5��Z��#.�:����}�k�X*s�LcM�b�l�I����0{�9p*mmz�o��0A�	(QY���4I�9�� �ŵʩ�ij�.�|������Y������7�>qbd�?����&�����P�s�Q[91ܒ�?���r�;�i����ږ�����FKW�^�4����Bů_�N���Z)����V˽b��ٮ-8Q��q>4c ��G�n��h����4�5����1��a�s�i��-��f�>��#A��l�s�5���.ٲ.;Q9����1G�1�N�i��剀�<f���H(�	o�M����O�F�9�4������	�+���@��~�Zw}Y�Xg����;̏���g�h�q+z��H]g�9oZ�G?ì�=��'�FFx�*>�8�3�T�un���;����H�w��m��5����%'f��pɧ��8I�ŧe���/�n��Ԍ�T�I�����ةA�1��Jc�g7.ú�e�>�U��T��S�ab���#J�'�XmL��{�d�M?;4�;}�lQ�u?(-a9
M.��B�����8����6���>(�,�*|�0+��t��V�=��9W�T1+���t	[��h�0C����/go����3���k� ����V��"�k����!�;Uw�*"բ>�{_� n����K�ӛ]�kaZ�u�y�a����A���H��C	HO�Ny��Q���S���ԡ�bP�G�[�dx*d]�+ͥعhC���B��\ �/H �T�3���yꊔ:�&��Ow�#0�f�w[�W����
��5��=EyT#L��WL�`M}N�V�-�4P �9S��5n�;;ď�?�%?�0x�� h>�=��UpЕ�����ގ�S4M�*w�6 �����<a,���S3��&/4��T�I��,B�Z��	�q���3t'R	m��XsO{6��@�~�~%�?l�e����y���}�\�Fw����C�A�}�=������dl��7;WC�M ���O��u+�m��go�+W�}g�&��h��~��oDo��B��2���>����$�u���ִ�>��xݷ�/�)p��8p	!eG�Ĭ��[�&7$�N�Q�u�����Û�=?z��A:dNx$��eY�{�@
�0���p��yڴ<��ڕCw���q��A#p����N�yi��s�oPB��	S�K�:a����Q��j��26�6Ud�7��s��i�1c���Gà �p퀦]��5�{��΀�K�1V��ȣ��U4���#R��fTk0<�Ǔ�Vj�[5�;T��gگ�
����m�QrZ��Jq�3��p�Z�t�\�b���Q:;zx\Ȇbݚ��iD��u6��Sx�������g�e	m:�I6�;c7ʻܸn���s$�By[��7��Y�N��`�#�v¬��-���w?�� �Բ.ć;���lw#C�4��B�:d�}{Cҫ/�'�G��&ݗ��w�j�&��"�.���]��h���%u��w/�W��0�u^":"6�B����ȴ�Բ��)���T�LiAii��=_�-s?w�\a2�þQ����e�)��M_ �Zzs�Z�B�-�W�vc���WJ�p�&�+R+^���+R!�ͳ&!�<�7ۑ�V&�g���:i�A�K��G�����}���V]}�"2l�"Q$X5��[-����ikZҠ�=�w6��Is���P)c�j�l.�񥣰�k@P�w�O>ᾴ�-v+P�u5Ux.�D-�78<�9O���>������u���YV�t�FM�>��;�\�5�9�r���0��4�}�Z�5�Ad���O."�,R�t�� ��)�"8��u��c9�3��&pd6P�q�ߞ����N���o���;o` �F���
�ނ��bCElI:I5���b���5��*Λ���M(㝝;�Z��݀
�W�4O?7`L����M5��᛹�;���v�^��w�4�e����T9���՝�hQc�/�g�C���B��3��1��8�}3H���m!��R�#�p6�K���E_<�.�%�c�ZJ$�ck�({�#���Y�nt�u�Vl9.��&9�s/�k���;͈��1ă�:��Z/a��N�r���A�Bs���l��db��&�P ���%o����$8p��>��#=X�|W��+�=�oj Y�n�E4�!�'1=X�S�阑DO���Gk��w8��T~*l�U�ةp���\��mU)�n�%yQ ��	�����H��6��/"{���Gm�:�5v�L���,�S�W�b�o"��;!���=#>��\�giI&�>�̀��Is-�9$�1r���کC��աi���Y�yvhD���o���|��I�a8sV �K��jD���xM���ڨݧ���X �X�G�mm�i���_�q��6���Mkn�;n�����w\6HE:+3�}� ��x��g�R����╵��o��FM(~5ٽ��O܏o�� P��pڭF��N���
��X�_]���DԼgmjy�'#	�c��{ثA,thsҝ-���:��"�d)��A4vk�o⇹�ԺO8h���*���0_�rJ�� ^ki�z��LnEw�7�1|�o5e��c�ڍ��x�zH�ƑܭcD����d/WR�_�yBs��p(�
����.z���ylx��΀�vC��������'o��x����3��!4Min�_Bs���{x����C�+�hΓ��.���\?u�);�]�Y�� �j�� \�#CVǌ��P�F]bD%F�f�����0$��eKL��1�,�U���|�xH`ܻΌ��|-~�%��?W�(��k��*��>�<�e��W��.f����g�rN�V�Y.� ��m�`וq���ô�x�����cV �P#7�i�-K�7�  ��e����3�$��]�[a��	��r�L3��άf�E�5�=x���̨2�-�5��@��Y���,����r37�r���_�@�{��p��W�Q�J��?%���E(��k�M�d���- �>@!���#?}G��6PS�V��@��׿��@�I}�0p
�r��hJ���,11���֤o�D)�ȹ{8����$�X���Xq����I�}A1!bi����~��OS֬�x_�������RѢy���#j�Y&�e�qʂA�t�&����)����E(@.t�1�5�/��"Z���w��p���
���B�>���"f��)�
NM���U�O����"���nS��1}�8��|Ztb�v^�u �ϋ��r�٥�-�Q�Dn�&�| 2���Ȣ���=G�H��I����O ^��ͣ>���C�oP&���lv�|3� �.ɛˬ%����O��pWF�g}T<��� ��]�`�(��o�l�,�9��mV48�q��
����P	渞BlEw}���!��H߅	�>�BH�*���2zpZ�՟m��8��qC��CmwN�	��m���D�
.�?���5��	ÁE��Wi�$�s(�-Z�È_��s����Dz7)Λ'x�$nUHF�����,�뻇�֢]�����w)�GLg��@�����V���'0�b"ߘ7��P��N�s�E�u�lFʹl7Է漌���P�T��t���]n�5����f �L��<�/ƦD��%�׏3��Z��'�/�q���#�Ĩ�ֻHA��#Ka(�ͱ��g�?-�C�sv,@��11����A����^��9�Q��RF/�Y�ó��f�?N�-k
r��z4HCBNy(I />$��qMҰB7�GY��m&�(�׺�v.��*�yf��d��w����i�`]y��G��U�ZPjv��@ĺ�^��Z5������J�_�ȹot���S���K�,�i�,�r���+��P�k�?��*�@PF	^�S�V�_�<�	51��.`/����84�+l�P@� �JR1�� ���l̓�p8��a��I�*Z��]����o���J/M���X0Zu�������.�[���xB(=2�*,63����Lv�Vȳ\� H�Am��q�����~�5S������3��ȚU��ĿDjkK��F��wTOfx��+lf�/;�_.�OąO�kXg��3 ����_���$����C�\�+���O)��	�9}K%j�����|tK��C�T�%��z�"�n�l<e�@��HT�:���/�+J���Ŕ��k�"��qZ�ۏ6�j�����zW,8֞����t�_2��}���0q���:�	Um��X�@׋�/P	f�<��L��f�)[��ө��$2�����ަ����̂���^ׯ�r<'�F,����"�<��d랒�x�J�򧢳,F%�B2��� ��9]�8��J�2����~��pz�4(� �?���+[��#�W�a�*�2ڞ�i���
EH4���'���I����w�Q��V������.�I�S�b��#�Cl�k������Y7>Uw=�<�t9��??� Ӷ޶|Z��av$-LS�`4�%"aa9T�z�h��h��Oh���b?nL)v�F�"M�L�:%�z��m��<�[ }eV���]ԡѪ��bP�c~��|��֏8ݼb~A�DطPR���Zt���Tk��F�lѤnf\/B��t,=���a��q��q��?�]��ᰇFW�$�8ǔx�}���͈d_ér��>�x�\���٥�4~慾�4Jt���<���;Gsc٫G�?�zյ� ���\�UL5����Iwж��9R6]���>�ȏ���X��W�,��%3�LVB��H2!��Q�&�sUNH�J	gFz�\}�]�1���q��0�i�9�a
�]�R�dWr֕�f��1:_�p������l����m�%�O���Ec��CG! mq�H�3�yA
R�pbq+�c	�2!��I�F�uB�p���U4�u�4��-�QƤ�aZ�O��0��<��植N�qn�� ??B�!�~Q�7��Pw�F��F��5�6/�Mq-�`x�pǺ�ҧ0�U�̤�O�)I�H(Z4~�!�Kw^{�o��0{	�#�1�g�=�)P=?/P�*����	�_�-aʵf�(׷�˦��C.��KBӣ�;Q��p�d�(l-r�q	T�`�XN�%pn�P�2P˰�MQ�d��A7����Mi����]��:��w�k����Is��	ȴ*��}K����� ���#��T�\H85W�dA5�G�Ճڍ*I'<�ν�6��x��i}�Ҡ�����$�a͜2����q�O�J��POF,j����hf�HLL/t���_��R�$C��Aw�gi�������h��SFi&��XWN����(��%z�}��e��7��v�c�)�O�� [��;"'�ZK��+�ǘ0�m�a�����l����0۶w(�!�Q]����o�"���l<p��g�7��qƇ���7�fvZ/�l(�ݕ>��b��{Q6����ؿ�2���9r�X(b:##^D��g�����`y�����V�{���L>B��U�%��	yE�V��G�Xx ��0���T�����΄�tgJ����{N����A&:>��;y���WF��3���T�9�q�a��ė����/˶���&�.�݄�A�Z}p��e׉��"2��A�f�(��[%��W�h~<�qvρ�����z�=�c���~zy��~)�Y��w;���ؕEp0��"A�).�wZ�l�z�s$�6���n��^���Ē����՜"� o`'��M^z�%�Ӏ���AIso\���.Y�4as.�9��X������:Z������ϐ��'����7p4�[rZ�c	�d5'V��̮V`c� <���}�T'H$������s���Y��/�

�J �ㆽZ����U�Q��l�݃UR�+KTz�v��q���Q��:e���}T%��`��_L�"� 7ү6�'�Ȭ7���Plx�ނ4{�����a�w�����fNr��nkz�Ϳ�oJ_�kX�7�@������$�*�����5� 5����J��̻�j�h+��neW	��K���R�9<fK܂�uHK��i���@�mE�Ý�X}&��Y��֝�F~���R�׀�]���� �[-��X%_J��Ƹw鴅�Z�kN�kNҿ
��θ?%[�؍��f���hRsΫq������M(~��<+Ђj(�&����`e>�.��4��y�L��Zf)���$?�C�N	Un��w�;�}�L2(���N�]�N����g+O��>r������� ;&�]^��wݴ���"��3��A��3��!t�� �J�_���9��s-{�Sr
E���qȾ��o �S:4Q�q?��sg���|����_�����f���3TY+ʸ!��̉3����BK���8r��xѻ�}�x��'��)T�����햭U�^u����0O8�3o�q9�J��^�$�Ս��Ec"���z'��\Zh��]AX�RV�;�6D�)��`�|�F:��?k�p.Ұ,�>���"T�rq�^;�u"��d��Y��wX �LP�U��O����B�}'%��H8�u�x7�ۤ�F3,<s�쎱Pѵ�P�� X#�! ������e��������ɭ��&�3.7��1��h)ʟnd���~���Z�>`�k�A��|Q���������L�?(]��d�y#�z~db�����>���չ��`����2��D@ #�F��\~B˷߳���1�
nJ�D"?k��}�O��+wݚf��$e��`�3! �p��O^ReS&�e�5��)n��($�Z��A�T��܍fJ�f�
P<u�)#��]��
���rРS�c��d��M+��X�kU������ˣn4Է�z��_}�*�L�x�q<Ǹ�?+BV��� Ӎ����yg�m�'|��S�����k18���&��5�)�5A���"����ͦ'���褩�
u���W��	��O.q��
��.l�fO�Z���ՏTO�1�Ȣz�d""�oi�2�d��+�D���d]���4z�w(�A�ʫ�F�P��ń��r�x0Ӊ��5v��qe�<�`x�����J>��ku�wt["g�BQ
���;+�$Оii��Y ٍ|x$d4ۯpP҅�8ٴ�2:4�Q\����p���<��B�]-P� E�,��u���c����tÛW*	-��B��@�D�0y }t�K�;��7�V#��S��h��B_����F�u��R��чgw�_9�搉�,߷��l�G��T��q��N8��� "_m�ʺ�Xe�h�:��ھ����=j� ����H�떦o�-	��$�s�r���v9V��I~xc��X	�s&
��$a�:A!� plυ��e3�\���G��:��ppuEh��7n��ƔNV�OP��#���l�eE����F�e���e�j
	�$*
ҟR��9�ðR��T�h��A�YE��+����ޭ=��E{�F�Vѿ�O%J�񟉈{�)G�#I׀bEϗ�q�-�"��#Z�Q��RN�P�DFJV��z�.m �V`p~�I.Κ};���lt̻0�9��*?��I��"6�8g�8�\4���1@c�'	P�1{"J���N:��Ap������T뭡�5u�U��Qv�Z�W3
��Yg
�x�֥.�2j8;t����MtA������o�y����1�D48����'�zM��7ʄ�0*��� ��}����3�d�R�"�;�$�%ñ'�a���Ɂ�$ht���j�f^1��~����'�ԉ�h�խ�Ǥٽ�?	k�����Z֜ו�$�����p�-�O�;Ӄ�)c��O�q���ԱGX-$�!�u}"����+S�Av<��av%�o�4jC8 hZ�㶱>�p�L����f$>����P�d�vl0�p��d�	L��+�:� ���/�6� ���K9����,lA�0�ޔr�v\����D��x��ԟ�ZE�^�jZ��M��Le0��2��kLf�<gG�ex����Ǥ��p����JݜqQ�3�U�ҙ�L�]+�,�v>�#�vw�����\�U���y�hV��`W�{a�<*7�X�v��m=�<���<:B2O-��}�t�JE�E'���U��`+��%Lb��S����%ۜ���7�A�V�\�Ù��pmr#�oþ�4hqSX�=���ϴb����Qt�+'S"JH	��Y럭��$�?��(��'gf*�)�҂�냯����G�f"鍰!G�u*)F�;��p��1��0t��u����-��j_���{K>�c�ّ?8ZX����W_���l���2�t��q��T��6O��D8�u�.3�뛯��&�O�KX6�{����x&j����,nk�o*��%�=��@�8t>����W����� Nn���R�������+�١�?���Ⱥ�U��4ݤ�T��_��k�A���R���׀��I����,4��:��}�]d�,��H��k�����;Adr*e;O��_˓����ŧ�`Ǝ��Z�LO�
sJ�Z�ϖm�-��P�Mɶ�k����;ug�{T������6�&N���Ws���@
�mL�2���p�߶���xjd֐��zѕ�þٗV�,����ƨ�/�|ՅdK�,�]34�6^ex�R��E�,���"�:l��*�VL�.<ck��aA��e@��6�T�� +�:�yx�<�|��8C\����6�xr�x���_g�$	���3�2�Nr��C��I�º��ih����k�\����P/��	E���565��n�c]]��q�;�\��w'l𔶌x(��?���7c�;wi� ��93tߵӊ�e{*'	����7G����I��tzr�� ��Y.�K�/]�)��o���xW
�*c��f��`�-]WQ��T����tvΥ�4#	n
�(���dVO�b�wħo��T��@C���=����3�6XYH�f	O���e�1�t�#<@�����-Fä��"�L�h�Z6�1�Q �F� ,�$�M,���!��/�>�b�'��&�2�2� x
O=D�����+7������:ɒ@�L��~E8�a>��4ɻ�����C�W���9����v�|�Z���2!N�f��e�R�!Z��e��-#�UP�f�@$Q|�{�\D#Z�\k8�|�X(oi����NUG%���B��J�zI����
˦�T$Oi�ݖI?/�!�HX�V�%@y*�m �MrZ�|=�7$���@KtU�h����!���O�	�XԛA�pr�+��=i}�z�<��a�t��L�[52�u����Mva�URl�"�D+0 �k���X����aNM��@ߐ.N.1g�ϩ��O@l#ZWm^֢eo��M�T+8��n#���}��������C�E�v���rZ|�w]f��x��ËP���N:ɿy~���Ȃ���gc7[��r���h跢���{�*{W}�[�F�v�d����@T���m�]�2����<[U`�&��wbjk�5"=rŷ��Icϫz�NL=�fD��M��������G"��V�Ȣ)�m�}RM7۵���S� g�b���0�~Т$��6nD>l���O��S�����?B4�AT��׏E�nfg�+��t�T�������C�+װ�]�S�r���x�ώ����H��ע31j�
�Y��U$v��5،&k?W	F�R̵�^�V���!N��(IH8��������X�^��v��4L(AmR��؇���ѳ�����(�{9��S�}7FŻ�h��㱴VV��S��@/שL�6����Ӻ�Q��l�/��"���*����$�N�u�\�\�ޱ[J��FŰܠ�L	�L���Fn�h����#�B/��5D���[M��5���$0����^����(2??���YV�hO��z@�=�g�oS�I+G�{�V�$���Mz��1�M���q�u?n� �n"uR���9U(ٝ7�2���Zc_��i�nN��7*H�wI�/���_����h�H^�(�<J�����S�;�����қ��[$����P��#�L��wًD5v��N���K��W�����=h2<d�)�Wg��Ց�C$r����:�m���a@H�!�˿���|_ �&�~k�w' X5��	_�^��Ll뮙��/��s�"&n�ʩ/����.h MB�����ϩ&(�A?�8�r�a	*�[&���^�z2/+���6�gn�ʵ�n��3�ԥD���G���/�"lK��H�e�n�h���4j�6�U��e��;��Y���z�� ���?"��!D����Z�eA,�#M�ۗE&ү��i�� ^
���f��']�=p����oG���I�WҙR�b�m��H�X�G���iw�SR�Ni���V谂���@F�Xr��\{�"�vN/����G�'|�/����5����0t��Ux��PdV�;�-=�ӓ����t� }�kDe�N*��+ÓVEvb{�k#��	R��Vu��\������T�ѦR�rb�0�	�|���}ؕp�H�t�yw���؀�������ЅU�5�=h��zk-0杰Al��K?�Bd��n+��qfYP��r�kx�y+���u����j��?b��-�|��v��6'+-U)��d����F��q(<{��Aj�;�*��&t\g����(<	��jJ�(i��������%ٍfK4^�ӝ�cӲfb�XqU�o�����}3�[�H��/flcq�����C��o����Vc��� v�nfpp�aQ����sv���.�oJX�R^�����-�����
:8|�V�5\�ff. .=t���l�{*�B��
Ƽ���n",��<��į�u=�$��^����<�9O
&�@C"�)8��'�R���p��X�	�LpJ�9��䍊���������X��\���F�I%���?�-5�}L�$�,�����Q �:l��Mf�a9L�LK��(@p�"��.<�u]�u��\����_'9�n��S�-�&��Uf$�B�?�NË?�893�%s<��*!�P�I=� ,;%K��Ly�	�h
3�/�3��#�,��{�Z���'A}W�k8:Y�)1�-BY�ޭX��@)m�Tl�Wz�w���3;��}��~�)Hrf=�<h�#�V}P���e4Y�F�G�{��*W�w�F��M�rB:�E��N�̀IV�Z�>iJup3��'qYv���X�W���i?*��ݸ�JU��U�wB>t�>;YE�����5４K����d��(��7�^���F�j{Gz ��wy�PZ�az5|�	����
��/X��9���:N�,QC��7~�Z��9�o��NѬ��+�,�U�Qj[��A�u�*��+����|K2$��Z4��:b���-R��`(_��j��7?- ]��`�K<�Tl胑g���Ú�]���gݟ���i\2J��*��&��L	��|Umf��|Pb,�z�|�(��-�]���ex��%-
��sL�G�&���7���g�� ��F�k#uV���.�CK����h�W�T!���@~�VM�j��C�9s��߶���LR��]ar;3B��6�ו�ʩ� ����A�7,�T�˒6��.l�.E�U���۵���`[C�钮Sz�-]h�a$�w�>u?��7ۯ�Ꜩ���x=[��ll:���s]���hu��e�ςx�i�';w3[�;>w��h�j��Z��V��Nk�Z�Olŷy�ŀA�G��!�����t���MM�l�%�۬Ly����(l;���=��g¶��e2�ۇ���U�>AG�0u�����&ifm
o+h�������3֊�ן&L��U'so�ݿo�H��[���Z�[I>4p��'�9�c�ʿ������,�mr_F���qJ���$��g�m��h�޸!Z����
�r�T�)czT�Ԟ�#E����uh^}A�	<t��\S��6�R6}���f��.�����)��l<�O�?��L�ˤP��h*m Kظ���5�˧���/�܊�Bw�0w^������9�t���:�ߕiU�+P�����"3�A$̓�=��nX�n�^ �w�<Q��v���-�O�]|fs�r��pg�AW��x�tY&)�X���oEA	mj�CF�\���Y9���}"o��&Vé�@��K[<<� ���tps��������?�߇甃�h�ȱ�	�$��^�z�}��
(O��!���Ź#W����l%��� ���cZ�d+j�w�ɮW�̨��31�����|?(q���)�E{�K}�V����(�NZ0�H;��"񎍪p���w֠���\��F��޻F@���?�ᎁ��� ����;����)p�dJ�l�U�&r�q`�C(�j�Y�������ي�9��s�H������?�0M�����)~�̐��%�ћx�{�;Z|�T^��w*��=v�؋17�`
� gs�*Gp��m�cw~\n�%$�S���F��w�.�1�{V���i,�=�G�L�ff��A�b ��{6�� ��-��S�4�ʙ��tlOC  ��K�]�Yke���� 緲A���5 ���%
�=��?Σ�l��{w����=|��k�iy{3t��;����ו��A/$7��[ϳkR�"@���q�p1��W�Ɓ_q����M��.C�*�C���Xh�]FSi�sF�e(���k&�!KX3��pW�1�̴�p���k���$�%V�Va=Hle5o4�Q9X�P����V!w�5t�<�fgN���}-��W4��=|�Х�2s8,�Z�d�t�Q;�Ǭ_�b�~�%��j�z3Ϙ[t��z�?����B3(fŏ�G�_�;�c�f��e^��'=OY{�Nl<�2��n&t�#����ƚ�|\�`�ceWt�P+v)O����U��]�v���E�H����S��̶/aCzs�;kZ��Kg��B������s?u,@[��;�����t��<�T��0���d7NFdI�!�v-R�^A�(Iz��W0���7�B�1�g�1�-Ðf�$��T��2U��Ӕ�����E�w����&�)N ���3S�y�9�b����y79Mf�Nϸ}�"�1HЋx�:�	������6���?�C��`n���7eH!��[@�U���'\��UU'R��@-��7W1~9�q����?�qu�F$ʍ6�%����p��'��u�˿�x�̅�S��U�)�,��`�%��]ڧ2 ���>X���������>�}�
.hK"�x\v���c���	䴾{�D��v*í�C��L[�YKq�p��]!�z��yF��,	��Q�xo��������
���͆�e'|�e�:e�Ѫ��7��5s�5��o�Y�3I�~̰
.�T2�ZcԷ� ��G���﷝��^�
8��W} Ph����( 6$�	I&v	~�1q~>�%,��1M@9�.]��S�~�b� �u�À̱`t"� H�+F�6*��)>�2�����m�9D���;�4'��h��������5��2���C�I��că�sqy���L���y/sR��#�3j�1���Þ-� ��:��w������-���@J����#2��l�|���g�s����+��[��(�4��H�l}Y��Q���
�=t�;��� j,�\�ooy�?�s���~o�A���..��B�b�EC]sc��q&vf����
f�I����=u�����ns`[�
���Mg2�1R	ْ�Y�O� �o�S˼�����o ��|��.G�b�om��P��{2���n�(�%��6i�Cv���;������GN��簴L����F�4]��cJ!���
���W�ᾠm�xY�ѤN���;�5N�ѯ��1P�=�	w�|�Ю�܋�$ϖo�5��[��l�1�)w��I�\�c��D���7��s%%W� x	�~��
�ܘ���w�Jei���K'�q��6 (��۳�ow�u����A�ܨ~yL��?��p����s-�<��U���Z^�?S�k�ڒ�m�T q�ag�Ymok��6����卟�E=���psF��vu!�Ȼ�@Hզ�6C�O=x�ܱו:i�i]f&T]���0Y�ўx}�\.ѢX�Ls4����:��	fӽ���;!�M-x>L_Wà8f�m�I��x`MZ����i�m�Rz���f�4��9Go���ŧ��Q�+ |����?qXؒ��c\\��J�b^T&�!�8��K�<�0Sq=����7��O��S�K�:���a�=��ي� U�+��B����˫�.+�牮����yP��:˷���:(�_Ϩ�Q�q�|ｖ�Y��R��d��ײJ ���n�ٖ��(�+�;$���Uk�@�"R�z'��!.|g+�����65��U�>ޯ|��GAH���w_���.9�Io繋���"Y����]��g_�CU=n���(���.$�9v�$Dʥ�2L��K�@����
�KT$�^*q�[��B�'���D�K���"NCQ}���2�4������L{i���;�bLW��4�y�\!wx���¦�&р���]Β?���d�@�^/�k�_��Y?�ϬHВ.��~�SY�t��}�@��uΘ��<�u��Љ+�b|�+i�i�~��WH�3�ѓfR�l��@�t��F�?^�'�s���}��b&���o$9�+O��sVy���x�Mj�w��t!�`�iV1�胤S�lW]1W��GiB�?�b�o1X��0�P?��߃�5�
��9=*��d���='��t�a;f��*r#7��P�2���ߵb�������{�<ְ�:�u�#`G���P���pd�(�&OɭNby��Dcp,��W��n��iJ���H��7V�(��$k�}g�Ӯ�^�V.���^�,�a�j,�uR��~�V�,�]vp-6��i���mW�Yyʗ֚C�@�ǘ�N�P�K7v���D�F��� ۘ���uܵ-V�4K����X���ɂ/�gJD�>׵cU7��%���dzr3CE�X�m�f�8�S��1����� ��fU
���؏�Y�� ���ʔ�&֪��I�+�H��-P6��$W�OL1)����_^6hc��h�AP~n����>R�='�D
�Ն�Ny���$d��r&���8�����eo����r�����j��9l*��%c��9��|��e��"Oؔ]*Oݙ�PZd ��ߠ|��DI$sHI��j��P}Daל\W�M����ޜ?����ǅ�e��j��
8]]�(b
Q��Z�G{`�C2�'�"]�a�ʒ�,�)��5��Fpg�E/9�2s��y��;)d t����˟�M����D�~����i0�k4�o�ixo"��;��tS��l׮�&U��J�ǒ12u%��0Md��n8��y���A*������T퀯^��W�CI?˹Z�]3�Dƌ�:ͨ��'�E�Jk����]XP���Q촨�8�5�H�,p|���o��"a�d��A\���2ۮ�.ܞ�]H|]TG�^�mx7�����ҥhM'f��ݥzҁ,��ͦ��<*��͕��y���>`�� ��$�f7�R�֖�����o�0�v?4r3�h��GJ�hB'�@��
�XP9N �Z ����خxz���ۛ44����:�*��RӁ����3`(�~@A�����\P\)�w���
0���Qk:�ga[�������k��易q	o�?���tڥm���?�)�����$�y$Q���GB�B�;b�߿ӌ�g*<T�	ő��\}�pB���o���ի���~Dd>�B0���M����O���ū�#���*;v�p�1��%�v��ߤś��#���<�����.��MGT�l�Ƞ�d����}���tqَ����V�>ʳ,b�C����]�+�Z�~��`U޻ e�����<�a��B�r��YY[W���J9񵁌k��¦2�0ֱ �8M��ޕ9�i�!f���R�jdie�H��C�Ig�н!S^&�� �xJ��B"z��%0����q�e�v�#Ӄ��҈]2۠��P��S��9�">�b+ډ����l2!O6���0S
�D`e7�P4�ᒗ>����Z�_�g{{�S���T�^�o4Y�'����x��ih�Z�J��X�.EbK7�Z����y	eܫ�Ձ�ъB_+[:����R�'��C���**kՔ�J����C�'*��w�:{�D+��M?W��ݥ�
9iR0В� Y�qӕ��=.�����.>�ϙ������;X��uХ����u�e��W����.A�n*��R�Z%\�xO�G�4{����ټ���s,i
m��������� 6J��Q���:��yo�/������>7h*Ԍ;�pPy�<Nݯ�ׁ��b�$;=���1Js������-@�M��IGl5�w	�&8�.=GQ�=�
��hy����81#>���y��-���V|a�ܲ=�0��#:��,�`w>|�i����9@�%��y����a��b7Nd������.�c%�0�#`
�W��uK�/�*���S1E��t�ǘL��?�Ls]'�Ik|~������״(�,��˼��3�?m�M^�H�5E-0�B��z�y�-D���.�0���:���?��Q2=�{P���L�7���q�_���\t���V˒��)�)�#_�:�>�ƺ�Yڨ�ч�(Pe7�B�$DG~�f\�(�Q����*-Yo��]�J?6|���a��F-��;�a��gZ��q�	a��vg�Ċru�`	h`/��Ʌ�j.o�4�`�_�'�t:��Vv���
�p
Њ����m�d��uU���&�C�i�� pkv�Qi2V3S |����"d�J�`@�_����I��*�)��T[x#��{�@|T�ۿ�A'�ذ���ӱ�#�8Ɂ�a7᳄胸��*Uc������o��Gp;b�J(�x����"���xFb0�E����bb���6$�m���r˃[K�h��$����-���:* &/�[��}x��������F;�Z�6.0ӱ���#�ص�L�� U�����=�K�X��v�ҋ��7�P�}�}/kT�\fpPIYt�h'��B�u����&��k|�NM�sQ�:h�|�
��{�P�8ψy�;�1����4�J2�NLIlm1/L�j4����q�"�}�O�	���;���Rᬷ������6�iH��3�ff���T��d�";0m%wD7���_���Sj�O%ëjk�,R�"�f̫�deuT��܂�Vp���l#��vv��'�����ڝ	R�r�$���I��P�gt���9���%͡��ȫ�����CI�?�F��,*�
�{O���E�[��x��~O����6l���߲j4)2j�;��׭�9�����^�	}��#�#�A,3�0��Ī�yW��Q_��Y��Kh���T�-���xT�	�QC��sbwʃ�o�ŝ�)HH��ҡ|D��¯��ÑO.},W*�y������2q����eC��?�k�S��҅�����XKtޫ�ԏ�6��4u������6S�z�D~*�����(����#B�[&z
�O9�Mȴ�G�H'?�a�3�� ��k[^��u�����ǡ�w�]�_jwI�����B]��_�e&P������������v��P\����C�A]�0Gr:.y
!�h�I�B}�޸N~Sl����n�m�p4�����?�B��2Q�'���e@G^f��4�,��/]g�������u/7�����x����Z0�[b*1�WQ�(���x�V�w�uדhR�	��<�A$,�L�sY+vZ�>wcM�^O����K!��JG��k{|q�0$NWѺ@��]�j�o�(:��Q�gG*��.��Sz��>A�.+C����tk�H;��~�?陲>)%��e����� �G2��Yxeuy�j4����-�V^R���$�į!=�8���/5�|rK�?t�qP� o`�Q��_�x���+�HXa�T��pwʢ�7��(�jSM�����[��*f���ɋ/�?�~8�[!���~f�~�Vj�&��#?�q���p�6;�"��"����`�'8<Y0\}n|�p\��R-w�r�E�I��k���X��q䲪L\=�*�u ���5�G�4�'E5���cM�&�v߭�ä�+Z����P�PO=pךfӚ���p��uӃ�s�V�a�'�ޏ�΁�uS�\}>�{�:�`b,�pjm���������%	_Lq�a�Y��`?ty&;^qˊ:�-��e�i�N��`�N�E�$�)�{<գqPN"
^�<��l,���.3�h {��¢ǘbg�W�Xr�M]2I��̭�!1l���}��U�6���B7Hf��[�p`J(�j�[0�W�(��D��er���+�Nt������ɶv!��^�D+M�z�tE�Z���擂�|dn��i��#��.�1�b��Ҭ�f�dU��[p��v�k��)�@Ok'p܍�N��	I�V��(�u�Tǡz����w�L8�U⥕�o�%:�Q �%�t班��Xt��k�pH��^�]���g�+���	0
VI�M���6����N]T�T #����;7\������E��Į��3�O �����"�Pwe^���,%�!�p_r�'#�G�9��)�|�{t���eE|y�֮���:dF�' ��˔���'Y�g
+����n)�Ș�8�I�mw��!��SO���{ �T+��߉]v��`L�ؑ��(8
��J����ޟ�.y��Ԩbi��@�'7�	ܯ���U�ץ�mE�, �]�nF*<��TØ�P��4l�G��\a[�\�Q��>�熔=�u���KՌC��l/���Z��xø��#{������)�;@������b,�?�2'�h�^�,~���H�$��d551�9@;�����M���$c�Ehf��y兎�f���s�	�,���_�w�!:��Q��RG9�-�����R�$�ktrɫCZ>�?f�=�p�u�W9N��d�4���u���dM�_����|x�?���:�����Z���OK�\�y�{/�ѝ/Bf@S�20�g��[8��2q���u>J�>�	���'�ʐ���M���vGZ,y��%+����M��q��J�h�Z�+��;��3�tl��:;�ڷ���B�GA�M��z��9Ǫ;�o|U�oAm��:ɗ�����;7���`�r��E=�^�p+7H�{�����&8x�k�j��6~)0X�cnXJ�u�H����b/W�Z�I�1^��-�y0�rH2C��1}�8п}�酸���W{��C�v$u{:�PG4��ps�:��6�6f��t�*��\%�@Jr���&p�\Cb�rZ�s��1Za_ǫ�=o>��r2�pO�WuX2E�$�v��ϒ�d���@��ע��> ^���Fe�C�;0<��)��tS�Bt�k�O����d.<V<�вE�*�q��3��g��g@'m�`yp�O��2�V�yqI�?���zRw��?T)M�KuU�m��Қ��`)��K(����8i�{��8x(�N
"S���� ص>'f���\�}qW1���o��1��qLn��}�/z�e`����q�N�^�.�y��M�JY�0/�zd�FI����1��Y;��O����X��VV��|в�f��cyL��<�&�Y��:�R�l�-|յ�\��+���|	�_�D%D� "��7�}Ұ�����´�h���U����m��H�A{e����}J��igS�.$zx�;�r��4�nAϩ�Fb�9mӶ߽�}'B���ɒ�S��	ݛc���Z����|�<��0���mV	��q���_V��_չ��`Xn��vB�T���~`���
�tr3ZJyJ�~{*�݃ɛ�=c0Ka�1���ˮ�!�-��إ��0�e�nuI�a)�;� �v�B7r�Ϛ�
�+��7��+�  ��q���n2k!��D���N�Y��yi��,�6�H5HN�U7Q�40�>�8���>�sm���8u�-�<F��|~(U�\J�L�,�X�!��Z�����PT�A�!�3ΏBy(+�\��kCM,���@�ax��͵��euB�� ��!W��к�s��'^%�T��m�����w���
�.�`Z3hh7��#ɔ�ęqQB)a ���
���Rg<x��|�*�ȇl3��0M��>��X\�,�?��b�d9Q�teW�<C	��o�h��a��8)���Նj;�m�_KN)��x�M�G�y�7i��a��j��1�+1�?㷴<�ç��*��k�B��l����]��5��=P^�Y�[xT���'��)���t-�HI�~����scU}�cy_q�SPE��+VcaL%���+�q�������9�
*�`����
Pʤ��p�Q����J}������Q�T�=<\o#VDH�U�٬u�栋��7�d��2����tL�I�H����׀�lp�<^�h]�&
���P;�^����4Rh�4�:<1ט�����beA޽�a�LЕZ 3VP�p��U�ĨԪ�����h��AJL/�R�ݯV�������[Y�^־��_�*�
�]���s��u�I�3/�r��+�ڞ�>*�S������]	�"���`w�7i�7eY��k�s��r�Ĝv��|��gw9�"�g�_��N���K��÷�iJ��cD�	<���#"��ᇴ�T3�ݷz/1vy��N�ҊW��ܻj�ʪF��z���k����̑Ud�	� ����_�knJ�dj0����L���}sa�8�fp�ѓ�i�m����Z�`�S�z�ɷymR�8I �~�O�Ѯ$����Q�v����֐�B
�k?��e��*�z��T���S�=�mj^|nQwl�ܦuA
��$s���+�zD�H$ Q���'�����)lc�a5z�o��#��6TP0$��l����Ξ}x���r9D	����"6N1�� �sqv�R	�������?�;�{ˁ�D��q�pݍc���������;�v�{G�	�, L�R��3#��1Y12�=��	����Y�,l��CJǪ��ZZ�uO�u��(�RJ���V�����B��zB���h����c3.dn�c��M��I�b)��/ ކG��	���
�Qy\��ZV[L��<<ݼE�;ދ�j�H��6�s��T�<ݝB!��<9]���;s~>�iG2fz��dA�o��k/Z?M'��6d�^��j�G�L�..��	���|)���X�"��Hl-{�Y�j�
���:=z�V���G݀ўza��c�V��`�G�~7��-��k�q�Z�����LQC�ѡ�x,��ϋpi/|��f��2l�'��2u���IĂUO��:Բ)�7�^��)��KRˆ�o:��K4�-�������A�.ǥ�i�'V���ؼ�m�}[2�èW��nG��ﳳz~\M^辜}���Tpa� ygw�nW?�0�O�'͐d�)��Z<0�~B1/Pݩ�����$\�.%��3C�,:��\�^��^����L��l�(����l���^����!~�h��:�B{��_w豁�}M��y{�q���.~����LZC��|���V�*_��*�T�1�8U��[:z�UUaWM!���'��ZY��8�KQ�*�	����5�L\Q�k�x����٨��t�_�M���W����77<�O+sZw��51,�n�=�'ZH;�x�i�v���n���3Sp��n��:�֥��-�X��mV��uX�pX���S �J������!���B)��<�{
�T�1�o/g6�1�,��-ơ�ɮȇ2�S�`�/�-Ľ�x��	M��gP��K�\o�D�����L��KM�>��]��!�,�z��c��-�u���QSꞰ^��&S�@����SC܈ECZ�4]���8/J�۾��(Ϊ�?����t��>(I�;���y� 2Y��}*�m��[���)�ݿ(W���s��3���S^2���:+������i���x���r;�"�M��@���~�J�L��A>���ϔ	�1��Ү�U����.�KDb����x=��������8=��Xck����~|�C`u�tyЂ;�ǩ�t���|h.z�0r2�}�78w����5.  w�k��>��Ӷ�ᱍr��p{�k@���^6N�	[���t���(�x���(������*��n������um�H�f<kw@�>�6�^;�usW*��<�m�78�q�Xsϗk)���e�Ȏ���#���=w��:8�����8>��]���3`�3�^~ʱMgiyy�+�i5P~u�;ˏ��LK�4������jc�������B~�}H���
�I���E!���\MZ'�ge��񠼶���`{g Z1�ŵf��c�.ƣ�O��F �Uo:���߿��U��"����Z
��e�ETe��|Yƪ�X��촾��L�y5�����6F�Y�5�����Q-A���X�Ƣ��˧�/P����+�t�������5��@�sd�ۙ�½�Ԣ��Ws:ɚ��ؙ��,v^MCr�a�`f����b���?Eke��?p���k[ؿ`�6�;Nvޣ(w�oN�(�2��f� ���&ǎx�����T�;��Vwp��Eq�����1lԣ�{�eX���hy�P'ǔ��G��W�1^����u\�],�-����;1�?��n��x�k'�*��;�p%H�\��_؈dTL�
�(-��JR��!n뽥����
v�
Ǉ/O~�עJG��{���p�������_���	L���!�[C(�H�F#O�{�V;"�Κ^}s��5�E=��q�}���e���_�Tz�$ɵq�!�8u�48�9-��{�婃�fE@�p\8���ult�N%����O1��d�y5��K��њ�m1�v��re̘� ���-͍3kp,&H�u�4Rr�ni$�Y>��[��7�����& R�c��Q���_�x&�����vo�4�r��u��mwd�{�6Ҭ��[�.Dӝ�%D'������6S,�Ubl�e��J�B����S��4V��g��\��^A8Wօ�`h=sxg�s��n\*|������2#ON�#ݠ��]��G��x�'��f��Z|�/Iv��UrA� �V��^:��(ߚҏ���Mß���7�ڳ�	4)�y�����(K
���_ �2��vR�u�.ۑiu}D_�ƪIT��N����W\�kd2��y�i����Ff�J^�ML
fsjJˋ�TǱ���mպ5��#%��4�C�@zŸ�:�(m��u�M� ���]�p0Y@D�Id]zT�ѿ�W	�WI�+�Y^��_��+=K7�!����v�@�ros*wk�껡�42W�)�z�ҡ<z����$��+������
��?�?����S��I���5~�3�G���u�rM�������F���������|?E$�})Y=~5�)y7TO��6�
U��:�J��ǫH1�^�����oo[���^�>�
��
�]��K'���A^��@
�6��R��c�W��ܻl��Lp�h��e����\���n�&X�xAS}h� ūP�
{L;�\%������1�ӆx�����۫GQ��љ�U�m����}��/x0Å���`�F��w^N���X:���A�9�Y�I��R��=E���y@g̽��+O~v{j��G�Ä�MS��������'0^���+��S����H�e_��Z��o�����mּ�}���fYaݫ;���''I<ͶI�/������j���n�$îbsf��7]f�:�x (�/9�]~�t<��t�&Oy��5ʐ��*w~n�����6����t8�����8�r�T�o�X�5�Z�m���t�y�u{��s�Z[׿X�x����ʿ���q�v��D:lX!��%��5���o��᱄������)B�����q�;c��]�d���� �"$W�ĥ0|��8�������TAGb;Q��o8>����R�4,:��L�67�\�{��DѢ<U�{!��Lз����S��t�S=ǥ�7�|�7�����kzfʴ,�!GT6"n�ʶ���G2���	YV��):����X���i�R@�-Պ�2H��������ec�=-����ڝ�v��d򹻅�2��(P������F��&�ϼ�óf6z��@خ�6��<�z��|���!�]^o=��Ԝ�|�����n8G��,`��I���@���؛��Δ�B��J�o�i���CFW,8������wXv��Z�|/��/���#U�n&�~;�s�0Y� u�xMWiѿF�}c�3@%9L�/{��|�c����=}Xi�������0��_@o��"k�1��Bk��B֠��.4�rĶ�oBy��-$�h����x��׾F���g�:�a�$h�9O��ٳ�,ҡW����'5AB��>���K#'��1��i�n���E�A0�`ӊ��1���W0�0%��	����w�-f�[�Z��'��%���T>�,9pF	y�p;�D���ɓ0 �4�g�%~��O��@|��;�ֹ��B�@��J`�k1^��E@���1;ڀJ��h�b�?��#m{�-q�)�ä�鏉P�n���E����23�.'�9���e|��u��<8E��  �_x��Y�d�|���Pև���!|!qX$�5|j���҂��>�X�Wi��I�P�>"Lٞ�S ���U�la@$jR�B	�T������ɪ��`���~�5�N
��x�`����L�bAdS}zSCjQIh�p�p�'�{���j�,��{�$,$�X3$����ջM�:�� �}QaK��[�[�N��tl��<���`�b��+�۔���m���F�޷���:��6�$^ϏY ������O'��a�'H�y�,�|��zSҫ	,��h����@�X���p�wӵ]ѯ��Q�lr��2���?�?1^�"Ȟx]N��σ�8M*A^~\��T�="�޸|��vs�9N����N�/�/�W�+	��_L���hIy�_�JM��24�"�T;��G5���N�گSt��Ĝܦ��tQX/�;��c2���Oq����E���(L����#\l=��������^��}��ɞ>�}wc������?����x�j�TS6��(������U	���6$ej��Զy}��o�(������MOV3E�G����S��U�ԭ�V�f���_��r���A��צzp�T�QV -�l�(�̭�CW�XĬh�QO.E�2)^��ɿ���KH��_�|c1��}��c~-�Z����s����a���˪O�5p:�k�&d����kIN6,��%�:$V�k�t���}�/+5���o�S0+
�E��yEb�����Ś7��r�"����**�
��!S�R�`��Y%>��cE|�Y�/"��<�9{�T�9f�E>h����+��@�wZ��M���=ֆ���Sv>�D�A�V�����QU`}j�#_ ������	���}b薡*�{C#�f&�0�kg��v7�yY�E�8�3/Ec�}]�.c}	����n�*����ҽ���XT$ݲv%R$�ێYI�?�oG0�z$h�� ��n<���,`.�d�s�������W� >a��.$���j�Y^/M���1W����`<;J09W$�W�aix�O�W�+`�gbAOD���������5����~�+��K~�(o�3�!Do�:3|~��Q\�o�y|yaS㾋��E{���P�4���E�s�κ�q^K��]��&+���G����N���팢!^?����ٺ����W�%�=����0<��#�_���Fo� G}�3����j���ѫ���J<���U��3��ؘJ��i�Z������+�<��eU���U֗h7����#ɜ��X .�%��5�M[N�Hva��Eg)A_��폛j7|@S�{����	F7�M^m�g��ҋ`�_�aw��ҹ���!�c�C�."�����ǣ�Ϳ�h��(6HD��2�p�Ձ)�ұJ��$�$��܂_e�ߗ܁���V��G}ȶU����HЈa�eG�����k�?��u7�x�6
�x��g9�(5L��Df�����Y��x�'�~��A�D�nq7�b'j��T���>���.A�g9x������&7l��ӭ�p��L�I3�OکnX{)�j�H�����l�E,|���+��1���R>O�⎯�c���q�Y��`F��!���V�9���Ǯ@S-56�&#�W��16%yq��f,��U��tJLM(!�eέUC�^9��"+�0[>�
P�9�hi��-5#R�c���J��L9r��uJB��l��3V������Q���	fL���v �)����s�]���LM�b_��n-����c�1$���OQ�<Q��K�\�	�:��S����lz�51]��!{h�.�̫C�a��?pݴk��X��;�l�;^L�sB�.R�Z�����s͛�,7��і�1Nօ��n����r_N9B!U>��t����0�N���I���݁X�Q�x2�K79/�yv�\{�x�6aG�%@������J>%�-��P_{��0�ر!�a؂�ͱWo� g�� e�|w���W�sw]���8-_`2��r"u�E��Qh}ݣ���O����(��}�H�Y��֎�}J@���� �Z�Ҭ�t�j|蕪��%]�R�&(���IC|�^/_ym��y��ÏCH9�<<ULT��O�̦����G�=�yb�-˫N=���ҮM߅c�_�D.y��Ű�~	�I�s����Õ.U&:}f5�Zl�-纅������4׻�T��O�s�1��t��WN3��k��5�&��i�J6(°�~�'&�����!G*pj���L�ŵ7��~�B*��$x�Dh���l�ê�=FM��!;=���>��~�J�PB.bvp�pr�Ց��~�Iz.yF� 	y�Ց�3bJZg�h�A0�b��"EmQ��=�EJ����9�8�>���o���h���"S����u�X�9��)*$�X:���u�sU���^���WP�繘��a���c���%��.<�)o?8�0˾c-Y��z�+��8��������$ ��li���t��Ҝ��K��>�
����Ǘw�]��+�����n;m��52����i����}u{��~��Р����3�j��ջnI%�h���u<�i�z�ɟ�$A�y���S:���{���1,�� ��b�����	��S7)�1U�E��}�*�'Jc?�[Q+ ++|������#J.�����68��#{�����*6i[8ohc��l$��"y�l�j�x%���lu�6�����;)��
ۭ�`�Ҡ�
�!�P��u����B.L;|���x�(Z�\dѓ(��<��tRɛq�Ȍ��#'`!g�o�B����g"� $v�$9�9���0�%�_V��To�Ϝ�&��.
!��VU�2[(�	��̤L��Up��k�!���{���N
;u��	�
7��"�Ԅ�,wZ�mZ�m���a�Z�w&Q����yq�URdG�%}�'KSq^�&�xNÎ�@��1ۢ�K�/x���Ǐ�W�r6&˔��̫�.I�f��������F�V����b��t4�֯�jo���AN�zs��j��a	���C0y:�&X�j`Ig��`*��K��dvF[b@�g�bA8K�?ӗ74�er��q���[���09(Av�gH�t�C�F����u(
��H������S�C��Yf�Q՜�?���e�C��m�!��w�t/=0�ĖI)2_���\ΊW��.S����!��5�a����g�Ժ�� �-��/���V�8��L:�i/�.,��vm���:�3Ǭ6�O�Wvhj��_�
��
ksʯ�us{A�@ɫ)y+w8z�^;auzD�s�$qg���
HJW�9G��������i1���g�.Վy��;Q~SCxnh4[��7��c=��+kA�_�Z��#}�ij�q;�Q�/��wKu�Z��j��H��z�Dl�(b^Ni���h ��˻W;�w��i�� ؊Չ�`����]jt^iB��nr�٭^����F��h#�b2�"�4\,���udc�Ź�ڪ�o�`�^�}�{�e<��J��~
+9��O���\9�N�$�6<�2,�;�Rr1u]��A����Y�	s�W���������ik�~s��Z^�mY�z<s1��Q$�����:�
K�v>�d���ͱ`|Q�*��[P/kv�MH�&��h'� ��?n#2�pB��3�YZUV�Qe�$i��C,��6��-;a>[eG��~�$sob誧8�C�r�e{o���oٚ�اDo�Qe���
��{=к�*5GVm�]�e�4E��]���j�Vr=�,��i��q6���HuhM��*���}��!'=w&Zv����$G�G�b1_�=���q�	��������7#.�t����_S'K��s�y�󱲅T��-,u6]������������cJ6����Y$3����8����:�[�>�9q@)A_K$���U������
��=��ǅh*��}m���L��	����O�yo>�S�i��1հ+�x�2���������A:�G�A	s�hJ�=���zRi�o��j��L!/)#��h�\hi��)Õ��Ci�i(H�8���Qs�x�(�+d�q�;�s*��iOb�Ѓź	}�.#
��}�X�"(�IyN��Ү>�\�-���p�R̨�,�P�އ��t�44�m=����bqf{�zz���m(4w����]�m�Wݑ�{�W�}�J~v��v�`��sg�����+�.L�'��6�^�/�:�%��OP��i��y�ȁ���e�ŚX'tt]:�(�4i��C���"�nGy����B�K\���c���䅴&'��9�?Rt���-
0{��x�;�9v k�OIz|ƸZ�uR��5$�|�,>��-Ē~eڙ�R��+ٳ���8�?�-���͞�t��uR~�˵:��xL/n��aaA�z<�,��5b�e�SJ�����[ϵ��|�*5|新A.�پ�S �'����=:��^��&fy�r��@=Ò�D Ha�X�o����z\�3��V�2Q�d:C=�XiAn�|�?O_5�c�#��v��
��w�U��%pu���r� 페A��m��r!M1�* *�+��U<�R��g�
��3�,�M�ҽ�PO
�ś�'ڠ��#8�KD��2j�(��~�	��Ϊ��5d�O����}Y0\�茗̝v�,}� &�R6�y�!���<�����'��ƣu�����/���51���mZ*H��]'ޯ���ؕ�k�#rz�/��+:~G:}�<��=�����9�V�Z�x����l�#��Nriɾt'��pfeTr�@��M���n�I�K�p������e
���ג�mV���S8��μM����e� ������ס)�o����?�P��ui2U��2�h��5�
w�3��z9	�9c�$�3����Ү �n0
41�,F�VVV-�!����H���?����% /(-=��$�b,(v�JT?�����w����f�{�3��m=<ݏ'滌�_�+}ȕ�;Goe��V���.���e��%z��u������,��/?����(����|�$Ev����S����Oo��<܋Rt�`��D�h��Z�|c_��W���3,����^ye��=��7	��>�8T}�L�f�J i�'r��zV����]����پaLO@���@"׌g�Y ��j8���[�ZՆ�ZU��|�G�s�%��u�UT�k2TǾ�d����ȉ�P\ܒ>�`7~�z�K�b���Y.J|��ǆ�ٽ��]�$n��L��V;f�����C%�;�ze8���D'LL��.8�}�����b��,�ug�y̥3_0&�RP'��]�rC�
^��b��v��5ڪW�Mi2+C��N"��'����	�t����E�=���+�KA�Q��|ԧ�x�xxN����,X��ʱgNw�Ύ�8�����Ma[mQB�y6��ӗ��:�'S)�%Z~��BI�\(���� ��J�H:�_i90���:�L���8����=ǈ��V
��|�"�6���$5#k|ظ*�b47�![ƙ���چ�j�z�DLz��&s!o@)+Rf�k*��k����(���83`�eɂ�OR$(Ia�`�[���z��v�(����%af�!9+7�3�
t*�i�t�5��V��w��T��6�:Z��'���F��]L$� ��"3� FPW�{"��#Z]�6u���?� "����n|�
�a�q�}Q23��:v�4v�^�Yp�1�ކؕD�_�Ƚ�6(d2�r��̨�� �dK�B�i���&�"=^���x��$S�,1���_���H-�,a7�R*{:������F��U�ŕ��(*���z�5�
�*G��=w�H�g�\7��c8�&L�����;8���� Oh� G�x��n�jĴ^�P�e��B$��ߩ�\�M�o擎<M����e�(qWC*�,:a`���j�i��̈a���E�e�mѭXz?��2��'��Ukeœt�ɁeTV@�fy��r���˴�3Qi@m����4/a�v�C���`��w����`�s#����`\,�?�_�JG�>ׄ5���s�����\�}�KZ����fv0���
g~|_��q ��
a��-:J��?���ڽ�\3�,5�\8O�i�������2��ů�nOk�ϙH��}��|��[9Ea��l���|'_X����+������˱�D����+�И�m)��m-�/�k_o7�������1�5x��E�#��"G���ʎ~�����84#���%߈�4B.�X����S!��OR�$�Y�(�A�l��LW�|2��5hMԕ��p$H��QE����l =$ !��!(��9���RĻb3f���.;x�9:�8��ۨ�5s�X�
�ףa�u�UNJ5.%��b]�e\Y���"�/l�{���PR�Ƚ-Sr@�I�"��K�b�S:���Y �Ɂ�����Wo��ƫ���m%��t��ܒOt�����I��*9����ʡ����n��Exd�T�d��!߮�OǝΆ�5����׍�"ʮmI�������_|� `�!��ۃ�������U�P W����	L�F��<q���:��Et�ճ&�c��b���Ȕ}�@����R��O�-,Amt����}� Y�yVج�u
	d���ۅ��KʷN�8��[w&�1�O�טN�B�y1��:K򉔤���.0�\��V"P���q�bW�SސV}\u��2N�dl� ��V���W����鐼
��Nڭ����y�Uڏ�8Ġc��ya�xȆK�脵l��CI"�
�Y(�������M���L�k��)�93]�pwb9F'Z~��M؀�����g;�kXSHH�8	d5�]�_}�Ĺ�(e����u~��M��#�7��� ��c7�6p��cF�68�
&�"��J����@�y��U�y� V�Ԥ>)��I������ ���F~�f��ڣ�s�_!ه�`q:acz��Zͽ��}�ۘ3�z��g��)��ɒI��K~�b� ��ps�W\��< �H��B9`\7X����*ř=���tn��p��m�>ǧNf~L�-�E�E���[C��p�,��:�1(���0�T�f~��J��.I~ǼD������y��mC$�Peu�D}JH��E�=������()�	����.�ᗇ�6G>�����=ۛ���6�f��ǌT��[�r�+4�ԍ�G�GP�!���������M����u�����Bl6�x$���n��� ��ī 6�q�=�����ꡲ�@P�g�A����cdKB'���SU���M�*
'��L�;��w�,�p�������h\��R"�yg
^�Э����!p�	fQ�e=��*�����F� �^��]����o��8K�����w��󂡪�ź'"��M��D'Rb� (=���]��:<�n�1�M��zǑ"J�,��'��72��Q�l�'{*��/����ק\Yw�����-�_]�?���!}i�K�}�ύ���>�L>M�vh��D���u�\��M�u��T}j��A��	����	��d�Ό	�p_lmU��fm"�x2)�w̺Q���"!��>�!�����OD@��)+����l׉�!�S�4�S�P���
Ȭ�W#�?����K������
U�0k3߅�7�����9�$�S����jhޅ\(C��|1
T3iN!�o�CA����pQ��G�^�\?F��dH��'�9?�SMT&���}1-����µ� �K�d�9���󒼮����vsN�B�Ƭ5��3I�1��R%b�|���i>�ɢ�#Uz�㟬�{G���rw�}F��o��*�`��p���	`ݥ�8ƥx�a���0��c�l/�R=�U������7ŲCN��GUo�:��5}?���h�~�J�Ҿ���W�jIc����?�7�����������ڟ�(�	�H�$��M��<�KEi���y��!y��A�f�Ρ���*0T�t)����g�D#y]+��,�g�:g�9�����CsF��x�IM׭�G���M��4�)��px)��DH����� ~��`x~ϻ�����ո��\���|���0+���a��.g���͊�+�n|:�G('��߯�fj�-/$�IC���Խcq1 ��TT��#W,7>݋V6]+�P0�F4�cՈ��b���`*���BH#��\U��Y�>���z6������.m��RSVPcޡ��B��a��~J�#u9���)�P}�v�J*l���MN��$ �7��0��fv]by���6i@Rg�R5[~��i��+�j�tE�?`P���z*Al���?�M�CW}i��,�\�I���3d���b�f/������6=���q��uz��bY\'���g،��A�w�s�{���!�ߦ�*5�K
�����&�(A|S8�n����}@�-A�����w�{Y%PC�.�����E��Zg@�"���8"�r<�!����}1G"�aK�]{�T*]��ˢqy_�J0�o[�<�
�z�S}����ɕ��Uw�Ҫ-���*��G���&��2��Gp߶L�	O���u/��Q��-~/g�j�"4s�/5��g�7݋�T/��XH��;V���IA/h�O�7�&��a��*���E�E�UNk���1�K���v������	f��]?h�2&�( �܊:��Ћ�x˞�(G�,��G���],Ə4�I��N��Ɂ�o4`w���V.S�dn��
�3��h��>��ߘ3�_���x���ofJ��4L-�����(Η�G��f%C�f"-�@�|�5)jK��*�, d���/��0N�M``�"���,H\#/g9�.�j��>| Rd,�Ӟ
׉�X?v�����h5LoG=�E�![n�PI�#5b*EFu��c��%�g!y����W�q�� +�	��������`��q��X(H��O�F� "�3k~H �=?�>�m���Q',���K��&�{f��6M8/NC��d�!5䤿����?!rj�#?��� �< m���\��x�3>]�e����œ�, ��fK��qeӼUU �����J"'s%��ɯ+M$�}�%۵�0ȎJ˸�4{�s%jJ�Ћ��� �~�P'hu����c�s���I��t�7y��*n���N���&������WR���}Խ�ڡַ2�G��g S5
�{z6"]���O��G��d�~�<8��
w����F���#���ῠ߭���{A�rX�m�yp>��nnw�#,�����F�'݉H�\T`*�"��!T��R5�ؚ^�D �ω�b�7�L*AΛn9:��3a(���&���d�t5o��.Ց����U��{QWk5�'�߹�L�-�İ��+�,k`��6H@����*{�� ��F"��ØI�*��#g ��,���4߈~��.��[����I�XP���f7�U�<�媉K��m.LM�ڍ%T��4Vd]HA����p�U:�Ǣ��z����&s�o�4�s�ď\��XNؤ$�B���|���nRh7���T>���F�5ֱ�B���\4�%��TS5�ڪT,:r[z�(j d�Yd�;��"��a�[�Q����%(��v3xW��ZS֮0/�b�#�-��~t�F��gӹ��<`��r�
�Ə�1��a�7�7��	��e�1�����~����E]��V:I%�1j�e]�Ƥg]�ȝV����2�Q k%��k�؄��|ȼr>�L��0���@1d��.up�ğ�A�C{	=c3�>�����J�؃�ȝ#�h�wy��h�>Ђ������'"�r��A��]��T/8���_l�.��*�T�ŀ9��!!A��Y�;�q%|���
�g��6�e���0!Sl�ЍF0�G�ځp���)�p��/R6�*e^`�5u ��b2:3u��O��f�m�U�(��۾T6��>8ӎ�W�Ӎ���y�4f�s2����#T����=��=��˟�̟�R���Ǌ��_J��~�ω�ͭL
\����y�o����Ё�:��+�ƙ�p+-�/f`�%B�D4��4�\�
4d�U%+�Vi���Gv��tgp���_5FC��4�.���:\�݈s�NT�x���y����^���[�R���<N�Ŭkj�J��%�hH�z�\���d\���A�J�t���c8���Q�7�m�1�f�yi�S������R(s�fsRe*�2�y[�T&K���uU �O��f� ��*���[��~�k��uU`����M���C��\�������l�z�3���cF�7�"4��p���)7��뾬���ȇ\��(�.vL�A�Z[|r��PJ�q M�%�l����22��3OȌ\�I����1K��*t���8΃S"�`��z�yk&�����;������3]]�[�/������hM�'���zm�,`v@���}5�ݯk�k�o��>�A��D2|} �&���N�����*cR���le͕ҚR5�΁^��V��J��ۗ*��F�˱��7�Dߙ��b���~Ѩx�U�?�����W��}<�H�;\k|񁟪Gs����k�E�7l�Oʨ�H�᎛�*j����r�����}������ �4q��d�/c�赯r�IxSս�H�A�
<;IvW�q+�E�� �7��6O{��Y@o��r�e�<���r爎б��o]iXBA����|f7iȌ��9dg�������j���+;�e�f�g%�]�Ӽǈ���8�!��Lʢ���h=��c5ǜ�����
6�9X+Z_xS�������%έ���Q��I�@F��vR0qI��x2у���J���v��֣�cA���/�G�����R��ʿ/>��t��ڹ؅+�+F�1Z�ơhvf-�?���1�����Jᩌ��
MȯWF�?7&�q��]�a�)\����#D�1ء��j���̩�ZΧ�B��������56T�fP�׍�x� ��vnY���&��	׉T_̹O�~�5��R�R�����v�LD��ϔ����iP��-M�9#���l���t���m�ƹ@r)w�}t4��0>-��d	\�_�b�y���a��D���Ը�u��6t��n"��fӿJ�܍'?���\6� �{���l�1�ږ�������f���c��-�(��yoQ�$�`�B��'�WH�Aiċu`2��� �N���$=N������c]��)%�9��D�F{C��/N��Cx[.��4���,I=Ɯg8�P}��7��)g��a|�O,ӂz� ��NZj9vi���*�Q.�!J���A9��Oe]�D�u8��Ѓ����C��0F�5$�����
Q�'U��1?׼�u�"��z<PQ��S�فy�y0�ٰ$ *�@�c�4U`-Ku��y����:�-"%G�@L3֑Pl)����SZ�����_�p}�u|��(���[ OB���q@����-�au�[	�/��j�gX��OrGg_F���p$�G��'���lV��O�!��EN]86� ^�/�[�KMx��E����s�՝���}h��ߘ
r_��v��e��~�/��S��k.�Z�>�r��kE a�>�͹u}�J�b�$T/fL~MKF�5��� �K-pK_��9<%)�7V3W�]�P:�$�򆮹5���S2�=`�:����:���k�C}���YxH��n}ѵ���E�� �1^��dҗ?FX�A�y{�<
�Z�����?�䬨vM���0 i�z������\,,m���u5ϧUb����6T�#��j3�,+����j@{��~��q/����Nd�^��!'�閾zA�3{��e�bS����}�zO��<N'�);9g�(��7S�x�x����/��mW���+;��3�ۧ�]���Ym9)N�ogzVm�;]�8�]���o���y��Lk�꽨�R����iҩs���N���L\}�Ï�WR�pӆ�	,�0�e�G��T�&�oI��b/�F�zlU'a2w���ԱO��OB[�'�wc%�>V$I�K��<b�h7�VKJ�U۬(�*�i�_M X&�=���K ��Ҭã�x������KR��ΌSNNر(z�!�+H�Cz�@�UCo��Ϣ��Gem��0o �\�ua��A�2����!�qQ����cX�o`a�CJ?�P�&bYr6~@��4T��j�t�d!�"v䆽x&k�6ymV��UKʅ�G�R�-��/�ˑ�ـ���8��E��35?���i
4ǅ�&ôZ~o^P8�N{��J#I-�n ]��g�69�,9�<��j\�Y�$(���6����,أ��d��.O�D"M�ЋU��'w��P:틏���&�JI�����?a��q����2+��y6����f��q�����ag]*��^N�쥗u���²��<�[|�w�@��
���4��:��ド�V77dsZ��̳�ml�+��{kR�H���v���@��8��9��Ir�)�QN�q��퐱3wa�nY�Q�)Kk\����@�"3q���!}��qC,bD�͜K6�3��
	�G4e����؈b�pc��8�1Tmo.���H���8~88լ)��x�ѽ"W��a�ae�{�TLn�5)�{r�:��-��ɵ��[���@]߈��ZCA._
��^t�3�q�r��[�[[`>"�	�^mw��}�N�`��7�i���_bԕ����i�	���ڻ�䙋Y
���)���{��@�@���d 9N�̲c*�T��!��
�R�ژ
�j�Ǵ�t�0���s���ʎe�3����,QA�-"�i��Л�P��	�J^F�k������G���^9I����ʃ��Lט�����ﺠ�F� S�!��)HTV�B��J�u�k�;u�g��_�I!�|����S�ѻ^ϰ?6Y�g>|�ф_�h����1�W�*�M2�KOꀯ2Ιi�a+H�'��L�"�Q*D�<�K���x��>	����ܖ�6��H�!&-k����;	Q���H���Փ&��5�6��] }��8�HOQQ��S�C`���Bs�4��yq�r1a���A�B��0�zٌ��K�:5s~����D�ߢ*� W96q�W�2�������{�"Ws���O�����D$��� ��ҡ�*���M�{��� �w1�Yl��<�+{�G�������Um̡�#H� *y�����9&�Lѫ��B�%��+��4�Ҳ֥��Bf!L�����C9xQt��*��D_����j m���blRi?-P�-I m ���o]n�&,�'��\,bRQ<�z�m��E�~�T�=�׮�< ����cٹ���B_-��Ӧ	�ςs���/<��@o�`G�_�;'���0�I���/[�`p�e��N��xWޠ�ٱ�97����ş��On&ڡS6��T�k\3�L��f� �`���4K��)��{*Un#�I�X�\P����4����a��x�?_������da���B`�w���_vP2�+��}��|܌�!oV�cll�Sz�m�����,H&<1K�9�B����{��?�apF]�3����tw,�����ϛ���y8>/�O�k��?�V�D�1m�v/�FMڒw{��	�^�+]˜��B��sz���S"�*�%F��k1k������}R�=��G�\JC f�Eh'#�vӜۣ���b��V�u���Z�\�u�x������UxS2�i32���$��| n!CI����^��T�W���4'�)%ȯ[�}�C�Yk�$��6��t������*x����U�ɟn9^ͣE�>z*w�_̍�� ZZw��B�����tA��.E!&pyY�8��X��ycd�̼��À02���!s\T���A.{?����S�F�;M�&�/J�A*W�LCl��������j8�f�^�MZ���y���y�ؽ���F���\e��������v����G`����r5N����Xm���!3h��>�3�ٵZ7�{��!��_r��@|`d�ts�XX��YS5�iTʹ�۫G�z��%�=���7�94N+���>�ݷ��՝���@Q�o���b�ya/�Q���.P8�Jv��T�_gg��hF|�3)0�h��>Q��umn�l�RB�l��	��.5�+��o|�Qנ�N�kt�d
��;@ɬ��E�h�Z��5�s�Rz��g�:�d��������$�8>t	M%�7���7�ѽ�a78Qh67��@� ��;�"`����gS5�t_�=6�J��TgDK�tO��t�X~�;�Xɨ{�[��})#�S��)?��ͽ���fR[��'����)z���ԈA��(��١�O�n>ɡO�n������pz��Q�1�@��nzآ\��!٬>zq!��j@��o����<kfc�F��HR*QO	��(�e�̉��ؤ�|�X��>�S�J��(m�����&�m)��D+X�����܉���{�i�@�3D�mH��6��~���s�d$"]�����9G�@��u�4�a{IC_z��������Y��Q���g7�)�L�х���9`��_�;1�_���zߑc�U&g0���>�i�^+P�my��#ʍ]��_@泖��!!�g�h�|���x"Ԑ�vC��{����Oq<ț��]�;��hK�ɖ���bY�3F���E��#d����Mf��a��寒���*
����;��㭁����(�=��L��j��ߎ���q��H�fY��(u6�d?��EDή��(�&h��?���3<�"3|]���֦�͆�(�bߚ�4�Eڽ�]���{xk�7^�B��	m׫l��.h��;��@u���ݺ�3)9y�|c*�b٤��|��(��S�����7*m�~�o�̰qڭ��w�q�v��ˑE���X����q%�ҧ��Q3��!Z�|3XP@rbkV@_�m�=����Dy�Xm[`1�"x�43��X�ۮ�z���4T�>�~r�fn�������bWu4�N�`N�8L{��
4?1��n��󥒜���`�B����1�9 F�i���xT{�k�ř��όzBV4[�r"Q�u0��ۋ�r_����w�fSx��G�F��|��ȭ��/�A
�u\���H�\�	3���Z��Ka��7�F��5�Ax7|�_m8Ɩ�oې�Ԭ�3�ǐg+�l��%����)��#����*߾�.Q74�Ҫ��+�#�r�xG��=6�L���
���:�jφ_���b�f�Ϲ/���;�7	�Ո��Д�%�����yn�'_��]�?�����\!��*&�]��8���>)�v��q�]��
2�����$D�kҲ�٧������ݏ(����^��t�T%���{:bM��H�-��hC��%����#N�C	��QN �wKt 5	��V�ny!�?U��Ƶ���u���g��E�����D�iel�ԑ '5�,w��U�i!y!��'��y��JD3`B�ȴLD�pI�z��F����y�V����jA��oH����]|�B%��*Խ�&I@K>ƫ���+;:@��a%5BGv��c�zgB�)�D���#���󃞯���m����s��4�Fh�R�=���G�f�}p�t�CL.��L�J����������n�p�,N'F��P��]�ĕ�(�����E���o�rB���$*89c=�[������u{�� ���ѝ���\"��ሹ@=f��RA����h�r*&d��g�|��Vn�"�b$�_�(��76�
��ڠ�2�C�BO��j?����b�; ��Rey,k�p)�M�a��!���3�"E)h�w�O4�n�!��X�@��F>��λ��D|��ؘ��l,$	�$�Gh�#�-U�յ��	>������,ۈ>�RfZ��%V,�:wSɣg0QAR���Ƀ.�35�ͻ�ӳ���&f�U�v3`/5���xRA
��E��%M@����3g�u��gH�d)yc3����%��U��8�yu2���Y~]D��Wf.0�;5��rsߺ�'Tt�[�9dL�M��~[,G�7; ���A�{8.��S�^��e��h�Mt��T�e����oLzL��+&�WB�':�1����c�#�>��c1�ZV��"�kپ���#=w7Ct��Ȝ�{�m�2����Rw��e.�%Ҵ���v��!9w��l��5O�!j��1����gx��0�X\�2��ΐ���4�a�g�����W��4���R��6A"r����H��珞�����7j��<I�p,���e�l(LT��	5��݄���_7��y'��D������X��|�-�����R�2�5p�)i>O�)~���TZ݂C�j�yT�6���_h�%�#��Rq�@�,8_$�=�V�5��w���9D��W�d��:c=������"f�G$`�\$���V3�X	[A�$�������]��̓*.��C�07RO�f*��6�%������z����P
2_�xt�6
:���A��v�R��9����(df�n�[����)G��(�78�)%��Mt��{NæR6=��3�㥴�n=��B�N�kYc<"��4��Z5R�^��s�$���mo�	�x]<�)�N����L|>J�e����Ր��1$g�(�2Ul�Q���1K҆Qw��Q$,��u���S�
|297m�ŉ���+����@=a%�����9��뾛/�P�,M���N���o��uo#��o�ލ���j��N�y�ǥ�/<7{�קg�7�%�@����G�D���X=8�ԯ����|���[�����l�Y�Uh�$0�)�K\��)�mC�9#����LdKM�iA���N����v�p��§>3�Tnϲ��Ԁ�J�zn���v���݈5��*G+���<�ѡ?�>�~��P���pc����}Y,��Q$��-ל�y�=�e7���=�m�H�8�5�ޞ�u����2,<S����McYj{k��n!_h�f���%W�߉�u�y�A��6��$����)$��}�Ȋk$�r�8naw��Ga������!�hI~	-u�N����p��O!���[�jCF)o��vї�� ��� ��k֔_YIֹ�0y�.��E��}�<��=�l[���Y��E�}�gn�h�?�q��N��>��C�� �LCf��X�i��>@��|�:�w~����Ӿs6@ �dW;�K�u�.,O�8L�~Bd�-�azo䚂����[�|��6���[�l�=��W��c6������c��������*��� �������={A/y>�L��8�eyq?ǠM���xp���P7	�1�U�֍[N.C����BN:Y�hѨ�W�!or�"���$p��G�S&�l�`���&9ch٧�����U���{�C3�� <Ԉ=��G}�:֞��[!4oP;}��*!�{?Ј���?���xFe�^��*Bž2�"�hO�o�?7^��Nw�w�Z6h��Vu��@X�eO��A�Ş�X,o@	�]�WO��N�S_�B�
)"R���T8��E�{:@����p޲��"���z9��j�m�@^��5��t�g�]���m�ʥ'�T���1'bZ5!��3��ҙ�-��Zih��k�3��[�D#4/'�e/^R��*&�k|��㰰�����}����zn�J���*�n�����z>!��.G�W�Bw8�0N�F�l�����϶:�pJa� ��N����ra��)"����-������D-ej�K�o�g��/{�Q�(�&��g���g�kF����[jQs�����YtF�뻍Mؓ���#������=d�,9 (!+�K`3]N�[׃�����c��
��m �����4a��X0e̠%u�K�;2�X�]��"���!��	�)�&�v���EV�����Q��%:�3Y�s�U�l����I�����혦J�8�|^[�S�UY�Ky*�Bl?�˾ߴ�����wm�pf��.J�d��W�E��G�D	҂%��Gg�!L���E�H�E��Yn*�̂��<��fNx�/Q���2�)E���QBE�yk^\��5jĦ�#��A�&�(
D��{���n%��D'�X>��2���[<�M϶���>V�	�@�A|Bc��|��ݢ�@�\���J�~9Ճ���+���G���J���e����˩"���H���}�g�&�;�QTy�
�B�X�����w��@V�@(r�wJ��SC�#�oEf�ڷ�8�1��X8�~��C-B��}`H�_���D(���/"�~;UB~n z��DYИ�_e�1wh7�b�6�xJ�����*��T�Cs���Y5#E�/D�wf�1�nM�Pۿk*ɴ�7��d��FZ,�ڻ��ďJ(��ޑm�h��#��F��:\��T��	�Ê��b�k����O�Wͧ�,��4?�+z,���k�L^Z�2�cc��z��{5�����8�-�5k(�W��te�(}���(�[�����C�����ҷm���Ϋfv�u��G<��Z��C2�@ĸ_7���X�m��{�#��}�.��dIj4J����IQ �Ǖ�2�k��%����:������Þ�_eo	�t�����'���/3�1�������h�۲��;� �;b����v�/Hr�3�~j:f0�����,l��)��#zQ�� �"��%y����b��Z������AN�]���x:O�:\�b�Λ��8�G�n����u��B(�I�^�շ���WBãK"-��f�Oe�/����+&����9ӈ�Y�a��MK��NR�0�K�q�e���\��\��L�c� 8t��9�<�h�,/	���'~���{?I�r��B�U��1ɍ���$�ez��$F��ȉdx�Y�O�U��%���.;��\�����g��7�:��
�켮�H����O��ٕ�E�PC��u�no}�Z���ԡA����|͕�j�����O���;���Qjd^���肷aU�h��#r��H���k}�X)�9�'t�:��,Uh�o +_���ɥ�TZ����5�T�{S��p��$F:f�峊Ž�6���%G���U,MB��9ē���_{��I��0|Õ@�O�;?*P,g<���b��y�4�T���#WOQ�U����Ū�"s�B��
�L�eV���C���5�Vo�7�!��[�VՕn�xU����o�7�_�H�U���7�^&��G�8u��=��a�6�>9��"����~��S��h���O���??K�-Y�F��>O�^��w�Zѐ#?�O�
�{��W��.g^��#7; ���/��v��,�Ca	U����ȵb@!�r�y{�A�y��o�NT>���ϵ�i�JI�S0p��K%���u~���L�ҍ�T6v����EL�A��ΑRF4t�r7��N�g{5�*�	�N��5x �IU������}{J���8�DO	4��,+�!" ��AH-����ָ�Kod�Y�a��;��D݁���5)b�zMwA�)Jܡ�� _>[\�}���Um�<vIϱ�p��^�Y̙	l~59{�f���	�kZ>Bs�_gq RD͢�T_�]�L\�)C9e�:��
?��PP���VFPsP%�1 *�n�3͜���6��8�0l����tg
�� ����_E�:�\j]xi���L���<C6,��d�c�����/!IX�?/=<dRd����0Hl��P�%������pfP����J���Pɏ�E*�b6�X�yi3��;�yP�|�㻞j ��#S��}�gaT�ƭs�u`����c�(�v���sb_v�/��ou���];_����������C
����E�,C{p�1�&ܘ_��X>��f���A���I�j�N��Ͱ9�Lʡ��J�4-(��{ĈA��p���q���ՖE�ѣ�5&4��)��pU����*(e���	8
N�s�W��"'s~e�G|�6L�ʘa1r���/6�7��|�eN���,i%�ՓPc�e�.�5��(�U�~#6ɬ�Ɔ�KD?����QM�J2l�%	�@x���.�bO�Jv�P��*��z�*.}��1�07%b�5�h��C;�������]��xGm���aI�����p�rƪI��Q�}S/��I>ʵ����&�mQ!+u�kK}~I�R߭�(��G0%�>��',ԃ&���l�Z��9_���}VO�|���	���3U�`��aC��> �U��i�Գ�t�:qs|	���Ɂ^E/���~v�a�=�p����0�/4�=��m���(���/ ڈZ�+Q��&g�eT��+6Hb���zѥ?*\��
��x6D�b2w^֒]j��7��:�S���
`�ả�1�|�͘�������Kv ��;��o% ��p}��P�B��oq-�ń1y=�e�8�IpK���+����i�8�5�D�]����.�%t�Χ�@�n�G3�0ͥO^�a1F4�2w�"�>	���#Am����)�I���,�s �Ya9��͋�C(q&.�C�j��J�Ј�o�yT��r���9KD�WWȴ�9��	Sh���ڗ�QB��y�+72�e���I1��l:8���HH���Q��+�) ��ˏ��6���uI ἢ�ՓY�R��p����s��o�sk}���p7�$AަQ���>�J��鰲����mwqU��q�o� �0�9��NE��R�G_P.@�G_9%Tc̻�g�t�w6�娲`��L�$-?�B,��� ����`YM)���d]���x�p���$K�?�c���)`h-s�v1��8�.5ٌ�?�/��
��|��kW�4� �r q�'�l�������<�i�M{�bv[݋��6&��MC��$<_�w�>LNS�%�����2^�:pO��Cq����	����0��;�������~K���D��-P/1���g�ľ����c�1�e*g3�@krGe�,�g���M�E,��~��]����t�a��h��]N���m����qy�� g��QBv�=�
s�!��n*�u��e��G2E����l��_�V�}a:V|���#��J�$����o5�@/�*t5ڮ��y�VyM���0/Q��&�ʪ 2��ߎ���<�>��ώH{��!H���_��c��f��k0�<y�?�is�bF_��y(^3D��x]����&=�$���޼�j��L_��ݹG=�Yg��#7&r���1��Qz� iI�촷'���׳Dz(��}z��RTe����E������&��|�+��_�v�=�����{W��9:�����������"�nk"܀W�}^�t�������V�s�z�)۫���M�BU�9�i���	Vb��G:������V�*�N'��������hb������-�#�W�t����o�(N�˷Gc�z�����g2iW!���Y8	O҈[��=%E�M���am� �k�J=/����6����^F�.�ӊ���3��`�Pt��_킳 �$L��G�:�K�e����X�'��k+W�����s%	.������?��e*߇��m�;A)e'?�L��룫qT��)�zwvѻ(=��;8��HG��P�������<�z�K��x�g��,a
Y���V��,�z���=05�L�hV��Q���k�/'�����.�$�������~c�a�<ƿ�g�����7���ݸye85Kњ�r+���L��I��`ծ|8x���̫�2X�WБjc��:�f2���/�`�f��p���M6�
@mzMT���q��YS�r <� mW��_�4�����[ݭA����bF��Z�2}a����ҹ��"K}O'�:ۀ��,�E)��wp�0�o�9#l�[��B�o�l�/G+�=�$NǼ��ȏ�-���lPp���Q�)������b�����˜���ʌt'�9�k~�ȝ���NP"�y�k\4n\�N�s��{��B����� �=XF�15����DI�LO�15tc�y���Af:U�Gc }����N�$!�j�P��h�Jl�Ӻ���:�̕ܮ#��G�;��#<W�Qv$pD����1��	ji�e;��B7�O
Ծ����ѧ���ă2Qẓ��������0S��`�aC#L�GZ��R��3.�S���^�8���O�~AH����րV��ې�|ɰ�b��l֡M��∯�)��YM�<���Z'߹@µN��&(��I[8�[R���2`"`Q�|��7�+`�t������t$qK���A���ew�C'p����F��l��Cq#_�oUh���A�Q���}nJ>+)���R)���M�"�]�z�L1�6jқ�X7П/@��텱��4����h<դތ-)��1���f�a��a�"��Y,�
�L&�}�B��|[F|�o ��3��e�<B�n6lb���+���,���c~a*s��!b?��f1���H{<�ɿ~�$����Fy6�����������9���5K"�c���ز�R'�r)�ٱx�\<T��<<-]�o�,�E�2�����&��W�>52O�L`i ���x��79��S�a�ں�0�b b��vD�R-|���T
��{!��*o�d���z�c���1�����@��� 6e��=����"=�7��^��ko�T�����+ƚ�iY���%��׭	}7&|���ö|zY�7��L�R/�,����%D�G)���������Hf&3�w���"_@�x�`v�4�
\��$�.9��~N�0(�� c���r��8����8,����)�q����.=[n�t՚4�-c8���G��h�[roW�[C���#���;�a">2��ѲZ�J��s���A�$C��:�H1��]�:��q*�<��=�0ʰ]ԯ�I7�[�y52	���ಞ�����!Oܫ��''�q��W���(gxl�tc�x{�4�Ƅ�H��N��l�jiT��鍬���W�ԘT�]��͡��L��%�5����_�q�Bة�F;���+���;<WfG�j����+i�#kI���g���о���$��5��D�u+�P�'���M2�+�v{��	��;��eQ��ߛ�a6�^�_�C�K`v�*��0�]8�V��q~
o}�ȠF{S�B��$�Q���5��53����:#]�����\�q���[d���CFf��������]�E�
����*-�������΋1N_Uϣ_��Cߧ^A� ��t޸B���x���R�B|�`ސ교��/�?� 7�I���k^�(ӝO.��l���2-]%W�4�Eĥ��T+�����ݗú�"~�Rlا+��Β։�מ� -te@�n��Y�*Ads�%�n=����wZ�
�:
*����Ȓ�,���s�u��G=��P
���^ܩ�S������V#����ö?���.���F�5gІ�Z�r+\�P�3-E߉^b� �ǧP�nX�������E���fSĲ�R�a�������
��bJV��

�����xᛘ~�%2fV� �Q�o_�Sb:���L��n��m��U�7N�g�rК&:4K{ ����i�����cr��2�8��Nә�u�d��]�1~�PrGY�����^�s�ȾYC��� �_�	�t^���%�Lű��%w�,�?_w��eM�!,������nN}�e�ӌ�z�B	�	�Ԫ`]*��+��orf7��< ��=ٸ��J� km_�	�:����x�������Z�&��LI �f��Z��g&��e�Ga`@���Vtl_@���E#M���Mx�N�'����,��q>�C˾,*^N�#�Zp*�?�ܛ���gڪj�)<���Ck.��b�D�c���M�\�
ӯ�.��֤[夌�-�B�M�HV.�r�$A �=w����<D�Ѯ�F��Y������q��8]���/��7>>��3��1ފ
��cl��S���IfQ�L�A�HOū=��b�4�'H,N�l������_N�N�%�Y��<.6\��	8�+V����dP?�5����5A}i��O�q�ی G�����;�攝�4[�����3�T�U��i��v��h���Ͻ���F�D�;���t�Z�j�?�_��O���d�6JSN���\�B�O9�Zu��:��if0M��W=��|s�rV��Sc	�R,���g�����ܝ�QE�$�BY�DD�YH���4Z���&��.�|��<��%��s<�(�Խ�E��/5wۧQ�����2X�3mԖF&�x y�I��W�_�u��+�`�AM.���z᭷�7?:ԡ���3��j�ߋ��H �| �upCIH��^�/7�����7 ��E��1��2�ofE/ՃD�`����y+�Ӎ=ŷ�{����Κ�s�,�)�,�Ğ���%����	%�.��XMO(�:� �E�Z��e��_��D]����K_���Ϥ���W�v6�N��C�P@wZ�`�O���`�&���]/�
b�F-F���7�;?��p%��X�l���OZ F���DA�"Ԣ{��+ p��RP�$H#�U��,��o5<�Ô�G����w���d�R�-6,�.�`��0��DlQg�-�)iH��2[����7�C�l��T.��>�r	�=�y�.={:��CJ�i���:j����@���Ja.�1*|���HS �/p����(��-��})F�局�K��	�gM�W�b~�~&�/u,�	�b��uo�TPFv�6�KΗ9����~��"
���j�G4xٖ�'?J�11��`�G�q�@5�.~�*�飅:"�YG N�����+��?@O�a~;ϵXv�k��@_�)��q��YS���%�ɯŀ�o���n0\�.���i�AI�P�j\er��	����
Y�4�ݑЃ����Eȅ�"V�����f�Pr)&��E�]v+���T�}J��؞�{yZҡ�:��-�A��1��a	�6ٺ��F��\
Ej.rw��.��C��
=Q�r�mz���񮹸�B���OB`Z�ѫ h�ֶ�U�2e*�!y�u��Hh������McvP�5G�1�'�n�O��V���Q(<s�K�Rՙے/�o^,��'��/INi��8��c�\���[v�_8/�]���o{����X�v¸$�D�#+@!G��v�F�����V'Ղ��.3��5�U�� �קg
��!���ІN:K���JaI�/c��Ȏ�|y�p`
�*���;k9��#TƘ��M>��9b�o2�E���J|��h���f�.|ݲO��+���N3�fQ��VW�~�A����R%���M��[:�-�!WK"9���Ua��s�΢�2OS�N/%CO�*|�
2�T�u�Ģ��w|t� We�ߜ]Rm� *�i�帺����$��i�u�D�����wEˊڼ�Ե����-�2�����zSB>.�+�?d�|�63A%b!�i�"�\���Ti���ߣ3J���Wnj��}�4"���-���1p��һf�~f7��u�}�A�r������u���HH<�EV*;���N���}��ۆ�v2"�{%Cb����5v�����,����]_���Y�}��q�*�]S������Fa{��ߩ-�
P�7�~� 2x7����r���_&��jc���B)8�j�
�	�|���'���Ғe�0���L���Uُ�tU�|��-�ھ�vҹ�WV>��U�
y,�/F$-Q��%���s+/E��s����k�r���z�.D�?�.��:P;�J���E ��}ug���|�Iz>�W���M������6A~?՛������_"��.���Q�n|gW�jjy�Bn����D� @���n�O�WjߑO���פ���s����^�q�P�oߪV+7,޾؎קn� 4vK��ft_q9�6��4�zѪH���A�oy+�AS!� ����8���Mn��Տ�<��%&����WҌ�ף"��c��]��3��*�J�2�m�4;Y�~��M��z�'m�/Ap�k�a5�1��J>8�:ε���̛�����.��C���X�9���RW�)�#����F��i���m���r�q�R'?�4��+I�ws��&d��,�;�)zh���͜�M�q�n�xY@-$dw;��Ė��AJ��9\�ЅBz
��;9@����f�v9�iA�F�`���zA*XX���b����[.#��f�[�;s)`g� s�\Z��"X�x�Evy�}c�P�(�~gR�MKe,��%l6x;�Y�E7FY蕦<��x7�<�q�-��*w�� ÔRu�aa��[�ʐ��s����A��ڎ_P7�Do޳��4���2,wٿ���}��BM@{��=o!2��r��4����b(����%���-�7��	\;����"�ٔH���:���	�B� �C���k�u�ğ�+Ҫ��ԥQ�!��e���,�0��g�%���:߄3&�I���P[kq����x0��31���,XUӮ �L\�.+M�~r<M�kѲ�(8��ڈ͉��*�\����nRD�*��p��$"�D6�qzh�����0y�Y������r��/��-�f�5e	��;<�pM����]���.���@���4�1�1���+J�
���w�L�8���Y�eWZN
�o}��5Qq���B��+]�!ۢI%�g��m�+�8VB*�W��F;��xrW;��k��)Y��lŚk��!���P�4:n�6�ٱQ�
�{D[��j�2��� :=��̂�~Q�KD�g��T�'�x��O�=�O�,�d�o�@#8�&���J:�Ʈ����F���Y�)���Q4�%�L�A�V��R��EE���.������ԥ���旻TeI�ls�X����K��F$��)�q�xKgTn�	�W@@u�dWi���i���
����o�"VQ�45x|���(�<��/i�	�흳����G�ߧ{s�!�w	K�����s�eV���)c/�4y5�u�����u,��_	S��MB52��8y�E��&F�ބ	Nٗ�G�4��l�+�ҝU��+�������+��E��AB���+�Un	΃����J�-Ѷ�~���(&m�\��>$N@E��ն�^�N�������\�'4�I���=0����dV���^�y���|���?3ir���%az� I"%��6�v�>���T{�؄��<�xD:�hi����"$�t:�>�������ܿڌ��Z"]f��W |��9	#2����u.It�}�Nj���D�2���U�ϵ�������r�����كbb\�-[g5^��-���h#�8Vd2�Fd�)�G\D;'�tZ㤔����c;�{�][��c����(����[ ��9`�f�.��6��'��f8ί�EGǉ�-�=���R�%1�fC[J�E2��Sҵ�6�X��c�8[9�E�RD_`1�hn>78̂NhYb�F�O[�2��73��Y�=(��[���Z'څAU\Z�9=c��Q7캁P�-�]`*1,>P�M� ���MxǦِ��2����x+'�&nB�!����;��Nʏ(��3�����:�8�߽���!du;���.<�Nq��G1��`2+لSA�T~s�L���H�j�|;����������Dp�6������J��n��34�S��(W��6!n��A���#�¬�B���H��I*�=���u\R�:$���"��j�M�if���vD�N���ѸC�Z �Ձ9.�]�_���x�OO!����6O�4��⼏0�@���)�����3�ywmg}�'��궖F��N��<Su�}h]��2�-!�!����m��'���I�v����$�%95t� ���$ ��9����d^,�¦ij��ΌX�M���5��znI�q'�E�&���:1�
|iE���%�M lĉ���b�Ɋ�D�;�m|�~{hZ�O�dɬo�e���f�v��@�xk�V����B�>�}ϯ�4hɈ�^`�i^p��6<P�F|�{�;
�e��_Z9r/.����$������Rz뺇-k�HP�
�����^�8?6��(>6��u�6��tM���2�S��n@��FM�tȟ�5}�|+�O�{@��E��y�mÕ5�s���ܣ�e�Hj����2r8�-�pf�J��<�0lW }N��ֿ����L�\.��&e��h�igU>�|%�I�/^���g��L.O�<%�����Ea5�>Wey��
�;�#�0�uADiC��M�hC����r��oT0ӌδ�p��uJ�����VD�D:,	0$n�+��0�+۰��I�o�,�$C�s���S���{�Q8�#S��zf��K2ā9��#�V�@����e{��s#�������t3�ƞ�;�)+��ao�~�-(<��މ��ޤ<1�oK9&}���g����.h�(\a��^�ӒG�O�Ǚ�Jl�+���%Kw�:��sz��(��s8�dz��>����"��a�5v�]�'n^F�#2~s`%z[�������<�x'�%�9�	��j7J�:*�ӥK���Fo/÷=���l"�����\+�V�t_�����wP�OB�ն�E����03��9Xo��{ܟ��6
Lu�����o��Y���n����jc
����ejU�L,�J�_��Ct�m�L)a<�Y�^�!In)�]��=G�K�g�N;���dVב�R�`B���2Y�5$�"��p�1o�yr�,�<��{�lli���	�Z�U�i:�ފ����y��`�]�( ��	�5/Bq��N݋'P2��ɚqC��!�kH��YM�o�2�P8=�h����]�N��B�gE�XqEj�.��2�Z�x:4_S����ڊ�`a{+CA�z�1�J�Kh[sl}�5ߊ�/��d- �oF�#�P�q��%�������Ҥx��-�Ѣ���e|�M>9�v��Ƀ����3#k�~[V<#�����ߤ%֑�������eŚEW��z��i��4wzK�A
��ռ�����}NM����ɈM?�>�Ӹ�_��YF��s�$e��]��$aT-1ƪ�c�N��h�(����	�B�෭z���|ArU��Z��	_�_,�k�(���y��{~��n�P��Oē��뚣��x��~�?�yIrx�����Q��I�W�~@�[����������	B�$�"�Ͽ��]��jHڕ��Ӕ������������� ����Y�{՞�
���F�F'
(H*H5��G����}*S;-��2���D_���0gom3jN�(z�{�. Kr������t��K<�Z9�9�[�*l�!��ƅ[�T�%����e� �y���K�n��+_-���hU�4�/�3�P�ʑ	W�jyut�G5B4�4�)�b����TV���0q#s��/ܮ��MO. 7t,.��8Ɓ�{�����|wi�mY3��j��$����e`m�v� i����M�^�����F����|����I��Wy�>���M�v��ڔk��!�\����m|���u���C�̐�B��r���!*���Ꚋq;�T\g&��r�b�� *q�E�Z-���D��s��������_��ͳ
�0bHKͷF�	i�j����\��(�h�x�����zS���y�d-+�Y�z�sP�b�܄���2᭤�V���-ʡ^�f'8��n*V��Cά�PF��*���ޡ  ���s�iZu�_�%I�`?S���;�h�{oα<�rF-"Q0�@��NUQL}�3[e	���o1^���q[%��4z	l��������I���k\< ?��Tc2mt���7`�-���r�d��#�Z��!�?�B��4�����s��Ev`��:SBb�ux������l�"��)c���!�������?A����-9���W���I�pB*�4M>��Vr�� e?!��8�/����9��3���Q;Gh��MC��V"��"�50��`�#,
�/ ���JB��v��@Z�}���Yn7\c���9����j�bA�5� Ԫ�pMݖ��pg�����1vI�Y���+��^`��dT}�a�f�(o�I��p�hF��^^���r�mC&��Nƽ��¿c[�T���_���V��w���he�x��Sz���3���]�`1s/��'}�SL�-d�#�e�
3�^(�}������eV�I�>�U�
�5P�Y?���Ƙ��h�@؟�N��4�+��.�9�9(K�af�m�u�?[��=���Z�� Yi�zי��C�~���;r���(t�(.�o��"��H��v���I`6?����( L����D�*SV�`�m�zҸLpk�����#p���)/X)۬�t�Z�|����������>a�UK��C}C���J�L|�ϒO���s���fݴ�~��Σ�fi����u���y��S��C�;���+�}:;̂�Y�4�T����#����+�5ಇCʑ�}��W�\��@�<Y�+��dhe��s�#��b��h����͞��]`;�W����9��-->��U�v��n��#����|�9B��R�m��*Ζ��w��FQ�Vc���h�u6U~yxߪ7�7�i�8�t����Kd��Y&�Hs�6���_$��e�K�D(��க-݅�Jh��G��s큑��}�����_�P��8�7{��t �u�~it��L�-�q�W�הY!Qգ/"��A���ᙚ��jz�--y]+��(A��-h80$��Q�]�c��[,�:��xa���S�
�G�~8�w&����+F��g�y��Q�\�����l*;:�L�x��
�l����KX���O���h|�S��{	������ƉI�"I�`sŘx�}%�پq�{�֭Y�|��;0���ЇH<<�_�e��v�ր!�./��9�'��K�Kufo��~&(d ���U�87ML��_k���@��D�ˉ�v{�E1�<]/��/���zO�B93A�ޜ���S3��-�]��9�`OJe�;b�ٔ�����G�i$k���O����|�G���j��våOM���-��zn�d�g�!�Ӱ�}��p��x9�}{X�:K8^�:��*���.�ΰ��[x$##7YK���	I�
�=�W۹7�g�t���ݠ��Š������ h2��p�!�*X��)a�}��*yn�&�9���l�Ȫh�2�sJ���r`��s;�>�GOO�w�l�Xb�+h���GC��MV/��3o�sCOpl��9�e�]�B!�;�Ko�r��Q& D��R0C}zH�=Q�	�V�����\�I 
�n��`ϼT�F�Я�����2Y0�9כ��� 3��=��{r�"��	���v(�ih�7#z�E�H�{�m��aP�$'r̸�6�+ެ�v=��?�4�w�=J�F����"B�D���r��Š�0��(z�kT��-V�Ϙ��kV����|ɼ5黰Xl�a�~
�Ɉ("��m�!�]�͒����!c6�Lr���;T"�~Ѝ�u���
|�t��Y΁�۸S�%?ܩ�:���W��PK���3kVc����PYKVW���$o֣)���Ν�ux��+Z��{�Ak�\K8�-h�qF�B�'�/���/��>�N���"�2���(i�AW�[F�Q?u��U��D���eO����Sx�G�KR�$>���V�r����S1�+yO��O�6�g��6b���8���d���@/�"��o��h�B��#h�,���e%q���aze��&"j�H���D��4��y���rx#+>:n�i���h���Ef���y x�Dh�}�I�����4݌��L ��(Q��YT��-�/Z�[��&�ͦP��YꯄXB�l�/��
Y3#�V�Pm��P�q�*�o���}`6H�A1Ȋm%[�a��=T����s��)8	1r�!�
�B3t��d��}�M�Vl�:(�Uu��w��Ʀ���/p��2�����*ޢ��.�%b���u�\�w4QR�XxG�����u=W�DVj�h޴ʍ�+�qլ$_���#@T_�c1�)�S�x$����9Q��Yh��=����iZ�t������<7O��c-�M~zc�6/�Y���@G�3T�i�TH;��>���f��!�P�����غ����)X�28s����u���Θ��PȑA�h7Y��%����_����f�x�U�>�6g/�k )ů4<�W���JYW�mA�,���������G��p��f��E�ѩP��V�z��9 �����@{"GyE�YAtT�,)DSٲ�2!J+��@P!��o�X�u�y�*P�n��0�����3~�X�#�\��ʧ����D�m��_�K�`a�zܹ�����ʦ�xv"[���*��X��wg��U��-��ɋA ��g�,�F����\��e��x"�%ta�-͎�'��_� ��1��`W�.�����f�;�qk7��#�'\F�懻�d�w������0��(�P��֨p���&d-����~�,�T�b�sL���U�?/�;��>C�I��u�x�V��
��MS�zGG���58����QSv����{H�ƹ0?�3�b=~�hO��9�4$�m �j���`0�żߠw�.k�*�Hu1"L����0�(�ىB2k���YcMn�RS_VpO?0���|�d��K�_��h#��[	��1���'x8BH�� �8�~k<W��T�l RJ8���t�$O�8���]mV�EV!j�%�ub'�@�Q{�q���3�8a����ϣ���.�L.Zlc:�q��4��o�nN��	9�q��(Dm��z�.S�Q2�4��gK�r{��`oj�w��Ad�|˩�j����9���qиa� ����c���W�m][ع`��^����=R]��,�
������*}Ԧ�/ʱ�h_�j폀'#�7_Dw7��cg�p����9���,3�"�6:��g&W��<�)���nE��y�%�fv�*W��a���q�Zu�Do�J�1Q:=�>���!p�`�{�m�����>�+&3�<������\?\��0vA��E�&	EQx�p�0����B	� !!�tm�䬊d��]�L�$F]W2�Úf�t�E%z�������"x]
z�.��ܱ�,(��ҕW(9J'�]Q�(���f�SK�f})�l��h;4�\�Kܸ(�������8��97���kAۯT؎#A�ٴ_�j";/�0�[�i�J��H=���/�I�V`JW�m�Ua�
m��w�ip��Tp�Ä����$ǻ�?�� q�e_\v��#��>n�:�M^P��o������������+�S4`r� �33�Wԡe=Iu��~QEs�%}y2�j)fG�EE��-0�A�e�*�^�������͘���I���0r#��C?��9�62/���Y�g�â>*��~
v�U�.�h4��_u�c�y��Z��4O4��d (oy�"�x+d(E��+	H-�#���d�V���rhw$��[��t2����>3�2@K�0�eaq�G�jO����G�wV�/�)+w���b�gD�=xHTc�Q�/��w�ڤ���udz�*[�w��
>�
��G��h�����BKI2Z���7�J�&(1-�e=+:ݱ�}8Rݞbr|Qʁ}���m~Yo�}��D����C�q9�ܸ��Z�ܠI�<�.q�D�R�g
%�v�Ƨ6��4�$yL��$$�x�Π9T�\%;�V����A�I��iA��.qIH��{=="jA*^<���� X
����m���9�՟�D���ҽq9[�&��{���PZ���茟b�
��o^�A3z����_�(��G���o�ɝ�VKװ���t,;� ���\2��"I\2��1J��nz��c0�+�/&6	X�cΊ�+�6# �;-`��pÅ��A֖��ֱ�������ľ\Y��zgnИ@5:������[:��;���wݻ<,'���M8�yxtĒ�D�<�B�<����N9����Y?r��#���
�tѭf�Z��g��r��ܳ1�V���1��k�k7��F5翓g�p"ɍW.� >:o��D�eX����꩞�������"-'���I�w���?^��v3��B�a=�[�^��t��~Դ�F�}WI�ejb�/��x��?��XY��o];�������Y���;�pK�⏒�����P>���i^�$[O�h��9��G������9����0�v4 �G��*I@��@�I�rʑ{"����3��J����S����i�~,Ś��Rg�)�X~�6'�v����y���發���R(A?�8>�R���37�XD�FIS�?F��qkpB��r}��&ɰ�.�!�����2�T�d@+�iI�NTvS2��L�2�j�!��uh����R,�v�!�0,O��,~���D��-�![;ۇ�g�U����4�<e_!1OT<�eP㘠�����ޢ�P�t��M+�`�4�.ng���[hL��f�����
e([�Ň8t�O_H}�T�0?���eEW�å�n^�����4�����/^XvF�:����3�G!H�WL,q�g�]N*q��h|�]����?N�+����Go��� �D�J�Tm���p���])�Yjן�ZEG�Xp^A^�X�rԇ7Ǿ@�!�.;��2�0��k>�ƕOݠi+1����V��9���1h�x>Lhg��0�����a���7��`=���lH��׉���'(T�̤`�9�1k��&��,5�id�&�iq����Tn��}��]��2`;O)�˞>`�J��T���O0��Q_09��0>]}�=قM���H���8n���0���d.��ɡ�6���={c�X��i\���VNq[`�$&�7�v몺�����a���[T���������tJ�ĪZ��x���F�
 P���bo��O�-������t��;S��U5ͬ���4�y�	���i���v)x�˯�S��"@&��z��F�k/k��RN��w�O�M�9\�K�6�ۇ13�]kh�z;�M��}��]�$4�����eFf�!����Ϙ���=v�x��:�|̴§���D���}�ҹi����1��,~m6'ZQ>�bV�`Y'z'��?��'��ݍryն Vꡉ�E�f�Bl�g����-_e�BY��`Ѵծ�0n�B�(��X!�~�����f�س����&��
2������+�����V�
9���}BX=V�%���'ǁ6�
���� �Uo��3|el/XM5�X�.�`<=1];~����'{d])v-d��1�ܷ&����#�%	��.�P�DÒ-�x�YY?H��ȲY�M�L��(j2�����Q��ߑ���4�wB��t��ZWQ�ޔ���8K�|�q]&Pg����/�q&���om���d���*�	�L�1��ˀ��9�.<�����(3�c|InP��fu/K �E'�mn�Dy�Iu�"U;1d�f��l]�e	ԓ��*�ӅD:���ڍΏ�.M���b\�ws����N�2�M�)D(��|o��xM!e���g�ϕ�a�;�B��24�S�6��XK�unG7	rvg �?�^���)�-�;���_���ZA����&6Ӥ���7\lP���"� 1E�W�<c�$�"w��/�A��?y��|�<M�^}Ũ(�ʷU+㏔t���U9T���b�u�4�lPG���<X���&��d]���K��cafv��^��"���t�"�ۭ���t��	�џ��Ӂ1���������z��Wzr+�ۡD<S����������0V��V!ơv ��f��p�YX�V��`�Z���ޖ���"��%�!2D孔�1?J��O��-��fd�w.EdYa��e�VL�ƘWI��>�:X����W1�
��� �"�c��X�3�h�f5tz��R{�\w� �N�!�BQu{F�#lB:�Q�s��	�ܨL/��W<:g�}f.�HV*6��]��+p���i�4��ll�N��,��B?�;�	�w�s�!Tgf�B��K�!�cF�|�� 7��^���2��dn,S$��׮���ظ�*���ڣ	�ᠽ`W���XN��mL��T�����g�����A���������h]Sh���$0�o	{���PF��Bi������eD�]�Y��5LS��-�o;�V�՞᡿MI�5���74)EZ�5��<�0��\|�n���C�M��R�d�H@��ޥd@�k7f��<{��zL��8�H#��|�\���%;��qt��`T"�e���
��7 �����"�S�S�O
C���R^���i���͜;��ߔL��E�o�fW�~�·�W�0��C�o��ٔ����.5g�djG�y�̽L��aۆN�з(�����Ӿ��=��$�g(�
�7+,�Lz�t��3�˄�C ��4a���Ζ�����}�y�Ԥ}O�갹��>�T6]Mz��m������	(E2Qt�o��}��bI �O*%�n �-�E��0���H�_�feh7�)�~"wlQf��u�y_~w���	�^w�y�&�u�2�/�X�<֜r@�l��7$��M+m='��nA�A�@D��`	���� ���1��7q��B��{uA��%T����j�(�T����Ј�X�f��V=�[�}%�e�E�B�;�=l}هQ�6���x��=w����*=%����g��,s�SZ�#C�-��ٮ:y�^B7�آ�Qb$������9�FM��g?|�^�\b��=���P�ov�cg�Wd.F9_����'�O���Hq0���nS�-�r#FE����e&�Hީ���R����{���-e.��\±�V]�h6� K@����S�VOn����/\��U��L����s�w���Y�9fw��]���PD\HXC;-��A�Th�)�d�|��Nȫ�.3�NEM�z��3��Xɟ���U�Ȑ�D9�u�[�Ŗ�c��A��:��E��o��N���}8�������8.V��(qg:�%�~;r�r���Ӝ6;D�Q��<2T�����z�`FGմ!>��y6�m�P1�E��U��,�%,��V�m놱\��Z�o�?E(\ymա�͵W�� x��YBy��3�����t�*!�k��2?j����DIRF�pZ?�QU��O�n���"C���&W�	ɺ�Aⶏ淳X�>��	F"�޷u��u�tN?;7��eR�M	��|Bj�[� !�?`��(rg$Z�:���"D���M�*�>�|-����šD����s!E��v�e�>$��J �uPOP_�
F��6D2^�ff⯙
D�A��]���.i	��i�l�o��B�:��̦"5y{�2��q�Y�%z!6	��_S(����ƨ� Nd�.�(gT��t_�9���w'�8v}���pH��3�W���m��߮�������wD��0��7��BnOU�s������{�4
X:����z���]r�_3�pܩ��<zo�/��_:ک VE����p8�/������`��5@Z�	�K�{���
Ƶ�Xx�k�:[Y�n�y�@sfD������wd_���`�^}�
���~aȟ�W�xq�㵲YU��ω�p���z��<L�����y<ם��A5��^���ŸX��(��AJ���F~�\��봓��!<~;��:侪t�Mh��]�qX w+�q);z�O~�8îj��d�V�D�}�K�6�LR;$3��'�en�d�(dG�<Xug3��(�̝l-B�/�է�����q�� g�S��-�C�Æ.B+�
��������)F|�i)0�(+H�������r-\�C�pN�H�^��-���U�u��!Z6���ء�G�	4�����S����8%i��XOY����O|�g�=lV�2��˛�>��9�#5a��ᛎ�%����	䢓	~i����>�nɃ����kq��]�%9�x�B+c��=z�֝Q�7�)��E/�9�8}�H��aw����eZ���'R�Kh$͏�>�$�y~�QV�ڏ�{t"i�	)M+�.�Р�T�J��K�ځO�L6��A��_�~��w���֛-v"���$���D��0(~���W5���;��{(�3K���g���Q���#S���'&�qj � Ǧ������ߨ�#<#����e%9���xз�z��ňƯ��L��G6����E�t�;����Z���S�Ңg���!W�[Z#�3�F�yx'�:�����ǘP2�{�+�R1zq�P���Q勔j{���e�w���.���ћX�{?�-�]N�w8j��4�HY Ҵg��G����7c$�n��W7i�ܖ�!{F�G�/���t�1v��A�2s4���U6y�@j���--���5�����V���_�o4`7�/��D��N" ;7��Mק����=�6���e�*k�)��?����j�i?�#7V���D���q��ǋ�rȟ��5ؕ�tzQ�?i_�[5jxF����&3��#�F%����Ҁ�4�o��D�\�rB��Z���Siϟtm�_��O�[�+>	��M�>I!E�"�A�_;@��|e3�K¤��6��R?�ȧ�8e�Ծ���(���*�;�*�¢�?o���+�)MU��"���e {��Lj7S<-;�ߴF����e��R��\Z�>����>pu[p��5���y��?"H��m��#����裓��y�J�������!/�h��o[�����A��"��XU$b�h���˽���שT{L'2�e�ap��ަ�hhc���V��+�x�� '��� x�9���h�^`1A�j�v�G���ܝW9^�یȩ�w^��ǻW���
i#�2�	V5�A�
���l�d��Z�9/K��0-[t�FqA���佄S��`���r=K�mw8j�ۼ���N�E��]�kBO�փ�]�7.6��{T�L��Q�y�KCE�I���}o��mxP��hޢ�ׁ�'v�q���ޛ�փ�`�;R�hD[ʝ�#�����l������L��h`�2�[Ơ=QB��I��k�^��a]&���B�. ����6y�>ة[�y���i��},�vK��Q����I�.M���5��� Q�6h��1̀�(�O�i����%�� �g�K8�,��2����w旰C6�w�2�h���zdmS�J���m�ws��� �(\w'ڑ�>�Og��!�?xvv:�3��h*�~�}�,��S_jyԲ�հ����R
��h��4h�C�^4�c��`r��N�۽΅�*�����V�>��@f��Ѕ,�x���*�+:�������#=++�� D@�2��b���xM��X�)�M؊���
Hԙ���р�sF��[HA�=�C՞ɮ�=L�魮N��}��;4{������~�:FwifY޵�Sp奣�Ke�*ޒDKK�u��������i����{�����4#�S�h1��u�C,�L=�w���@�����ӽ�	��_SW����0P	�7�=��M�F��`�1rc�aI5=�[�aeN��IrsE�%g?�L�XJ㪶�0L��Ѻ�5�d����Oڒ��1Қf��V��n�� ]x�z���?�ޖ�CU�[7!��RI����G��G�bpS�f�Q%ng���aۿ�E�n�Y��P ��Zh��tA�z���z�1-����{��V�e�\�2gHP�>��v�t�>�<�{L�J��U%�o�����d����c+ �Y�}xŌ�A����/�_#�/��n�n�jU�\����L0�e������,��Od�c!����ve����:%;��td��5I�3��"��C�±��~6Cj�d-�/� �h[,#6�S
z�Ck�󧤵��z�B��q�&6Q���M���]#�pQc�o�$;,�t�yq W�H:`����+�{6�ei7�:�זo�TJu��ekB��x橯�y�3<�n�V�Oe)*��x���2���� zN�2�+b�=}��P�ut��&�A��j���Ynrı"��!!�owx�U�� ��߸xD��oA��el���n��?�><��,�&���j�ϡa��F<Uȸ)^�0���X��=0���������w>����T�I����3���/�]aW�+�L�/.�R�kbp���P�g���גQ���x�ۿ�C�,��6�������k@��M��p�����#q�9�-j|��ʆ|b�����ʤ�i��#�FV��St�Wd���]s��up۟��I��8k�����:P�h�6��p�%���X|��C���#�nJ�&ͫL��D���ii2Q�jn�kѢ�k�(A�*�w��F�2�"{3�ҶXG��}n�	���^F��N��i��w��2ص�R|��P��{^�vL�½U�CnS>V."k�5n"�Ou@n%���3�:�����5L������);�~�!�-4.;zO�N��3��Dxg�S@��*��
f�=�PS�C�_��� �b·_��� �N9�<Q���{Oc����^+[[^֯��zO,?�1�W��=��0��&��L�rlx�1믽)g y��u�kIňu�	�C��x��)s�4��S?XFv�[��r���=�&��ɓ��.J:*xg��g�l����qԔ&d����k��qhk��(�~Y��s���dWk�78�������?(��5�%����Pb]\��p	[���f��c��ݏ*�Uʪ�ޠ�d�AB��$&��K�2	N��z~�9Uc��l��\9�k(e�&��I��*[���b�A�%�jZ��Gl)�|]f�}��)��<��|ĥ�&+������#L�OO�^g�Ռ��n-q�@$)񀃂BL ��}�n�1.VZ���ޱFC��̠RO����/B�Is��U^�}0�0h͹�W���O04T�<���Q���	��;�Y���ᤉ��n�nI4u�.�AU���m<�X��}�v�W�Ge3{��8���=���1᧨�ٶ5���/*���Iw�����V��T "�k1�V���~����Mn��m��������DL�;m������0`7�������4��D��k�p˜�e4Bjd$ �]sՂN������q���承�hF}W�(sy������f�����jy�ɴ����3��W��M����"D� (E�����٠K�,�=#�6~��{Znn�~���T�
�综9'�{�S�|q�[$����*���H��x��h��{�6�:�^��Nڟ7bsD�$'9�����@N%��tb�	"Vۡ��u�	�|�S��P���(Q2�~d���B����� �=U�� Y� �A���5����w�,� �uF������5��@#8��E]�����\������#�K��XH!K���v��!��r����{i(��A�kgb;h�==u����L|gg=\�� w�#��}�E�C�z�;����H�Y��!9��0E1천���=X�б��ܨ,p�����9a�vI�t�/T5::�dS�۟,$��ͧ3a�]��Zxy�31�$��=ǸM�iUGt8�
�!����sn���qF�֛����(%7�����K������R�n6'$��Q���LLĞK�z�	�H�
H3<��̮gw'��+�o����ܱ\�<�1E�uh����;��S���R��t�la�J��m�	Ͳ����\99&�C�9ƌ�Y�%3�'�[�UN(�Dh��?p@�'�
��������(kf� �`0�ܐ��>�2���*QAW_.�A��X���S�k��+xn1sa /	�j.*!�<���=\�(\������n�)	� W-/(04�i�Ib����<��~�q5�L��H#f��0�#0zo6 �56�g;�.X��e��ˬ��h�M�YlNx�C�����X�.A�9��q���(xM�Op�O`fx��7�2A_�wҚ���zk���}�uV���ۃ����`��]f���X��1�<�p�����n8ĵ6;�s����������B��8B�����TL	w	�{����\��
�Q[� �G�hCEWAH�T���67���r5"�~f�-b�M��87oД�Q��܅�@;�J��fS&.���D��ā~�[����#g�Ŏr��@1��7WUL#��y(��D�$����T�HR>��"�g��n*�HV�8w�A=���A�{�`��[�Z9�����P��{�n}e�
X�殳*�A�e�82_i��5?�QW��5�~핥W�&�bը������9ʰ�@�� �o����`�p?�<��q ��q��ʹG�{��N���C<�!k��/$����~�L�N�)��K>o���@�/N����L 5�<o��d�`�MF�����.�Hh6���=!]����i��>�Ē��?b�ț-���J�/!��2�{��ԍCJ5=~r��'�U���\����)OZo�F�*�R���SAL]���3Ѻ�~�l^�;�nh�1|g�g�n��tРf\<�}S�5߷��J��VV�b��<�1��)�l>1쪲f��7h�5��.`��5�b���u�o(τz:(�.��6�{?�;�$\u}
��� �LcA��o~Ɠ��E7�ض�AD��w%,�E!������'y:,�9�ۉ��6�Bb1�/�v�Ch֋52�����<�^m��=p"h�l��܃�ү>&ɾFm�O>?�oJ �xa��՗2ʠ8�)�v��^7�v�\�ZAg��*�r� ������v��/������u|/qǐ� �$F�����"���$:�ܳmM�?Նe�P}���oА=A$L��k����YBܮT���ՙ{����w>Xw�s~����v�p
#�;V���k3�	���|6��r�-��V)kNQ��I���J)٨�vO ;���
�D���E֞�l '�oT���Hw�	���K���$�u��-U�z�)!𡍶���j��8�T���?(�XP����"�
���P�TS��e���`٤t%���AS#�er��gE�+s9�j�(ه������1_)9�IR�����I�d �~�c2�4e!4��,v󖹄���c���"R����*?�w�6Ab�6��?(�b·���� ������(lD^ߡ��p�C�Ƥ�t�ի�!ү
ʈZ������5�c�+[�n��%��R�4��w���������]�3��|���S oW����Y�������_���e.��|��rpI{a�J�(U��t�N$d�E�ύj�t��e�Gt6"Z�f�W� ���j�]�tj����(�d�\�]x6����@�	�޳���W!�3�Сv�F�B���w���y�����SfA��}
�L�5�Nu~l<tC�m�mwX�� Q����*=T��
���t.c�&����|�ϗ���?v�jҝE�i ���6�Ј�YT-�a%�rLO*��g�����g*S���"�	'�W�����Vۉ�(�8P�������c*w�����w�%y�NS~(/�}W�܈��<_U(�L뼀�1W�mf��t��XV����ٜ.xa�Y(��^�:�f�u�y�f(�{�Α��)ߎ؟Vkr�X �kMQdIOK	<���1k����D�-�Of�l�z�5�c��:���_T��!/�uZs@�h��Cp�X{r�v���*��gU�x�R,��&D�9\��)w{Y6E�r �����FI'�s<�G�4��M�p|���U�� @i�Oen��w`K��@��.�����rh�͛[R����۝�,�'���!`&����L��ȴ�c��,{�k��?��LC��]���SP�e�K?S]�|�_��ӆ;��Gn�����3q
G�$�`��cwpl)e���17� e?�~;��]��97�%��h�r�-���b�Y���f��QbC����QwG��t��٧ʁ_���P�� �z���Z��Rhj���N�w���lH�v6�]�`��s�Z�(��+BM�8�&\*�`f��_Wk3��VT.�|����:��b��|E��u������F��@M?qaCl��~ ��������Ⱦ�[�=�U�������y���~/�[�be[�)���'���MlRK��Z�8R��1_i��<���T`D�㟇��V��o�]e(�=�j�Wa���8%8b�G5D���qo�d@ [���/*.p��%a�?�	�t�l�4�ųCB�/����U
1��0�� g��X.|m��$]���ݗp�)� f5����v,��;\�Vm���18B+U!���}e$��A�Q���OP՟J�񼼇�G�AM��MRT���^��q�&b�m� )Q��7C����\��M�3�6K��bڇf{�� ҃!{b�ey�Vg��;����?�Q3��\��vb2<Lѕ3�!�J�v�ذD/�I~V�/�me��3��k�S�3�)>����[������aD��n���R&CP���B�Ad� )�=�LV��J�h	�@\.�s||C�wz#�����[��kYG�Ԍ��K���x��� �r�����c���6H��I�ew%�L�aA�?"�K�
��7���x֝U�!=������b���"��a�P��t�D���ϥc�`���W��GεK�s�$�i��PD1���W��4�>8.�cc�񋲇�X��D��s=�ip�dAg��:��;�#�b��g�Ĵ� �뉤	�vs[T,���6M�W���t�Bj��
�(v��'v��̠c��������閎ϼ1� �.�%z�瑡�:���%l�D;6{��Ta�{��u�	���P<�t�׷�<β���?OI�+=k1�LF^�����B��ϙހפ���6�r���!C䚯T0�'E��.3H�Wv51���w[Pg���ڕ~�ܴ����G�8��krӹ�_��$��xxQI���~��HI�<w��@y�S�V@�P�p�D�i�����^P����g�3+�Lp��h���O��_O���e��յ�����(]:f � ��F+4�d4��uz O�&g�ߑ� 9�etY�M�x�y`8��%,����V�^nK��#Ws�61��̵"M_I�)��YT�=xS�`D����#��LC&V�t��Պ�>�y��N�nOS��=��A�1HR�h�Z�t�g!n.8�2`�%�y3 (�w?���� �~���j��Ǝ��� 'ԅ�[[���6����{��&$=w��xV� ���ܐ�*�ē��`����+G�Y>���*��~E�/}���C=��0R�h���~����-�y�_�Y{�e����J��H ���Q%>ڟ8AP�[��z�%���K9�>�~���J�u��*Z>T��ש�W��q���������K��*w]|ss�"�,:�I�P���ڗ�c�As}��%��ü��rS�.�Om��u���������֞D�e�Ӣ�V�W'���
��C��p���V�v�Y�=���=��\�{7�@����Dy�Ɗ�h�,4xA!���	O�S�LN���c�t�ُ�Ǝ�D�K��_rʇ�GDK�I���ծP/��4�ͺ�ldeO�T�q7 gIZ�՝*�s�.Y؏h�p$�����I���b&�`�}z����WJ^f��is��[ I�#C����^zO��)�h�E���@|ѯ��rS(�8��A���O�G~x���#L6כ�5R�аC�_�
��C�V�T��Y���0�F��X��Pwt<�n�T�_	g������>�8D5쳥JB5؎��.� ���u܁���IR��!IP䩉gQ#�o��aX�3���E��gr����(O!ū��Ҡ4iH�a��M���8>�Ұdy��a���v��N��Y.(s���e�j�;{+LUoπ�o���veM�@]���VcS>�O��ͳ��'C�){�P0����+���L\�I�(�g?�����f[�#+��*6�&�>��5

�xʮ�������3�Hx�9pP}Jo!z�j����J����Z�`v��S���L�+.iVU���4�����C�3��Tzf���>���E���EC󵡹?[&#\�>O�l���e�`��?"������T���V�oI^�D�ar|u�>��x�A�?������i����4��%L���9!w�?��d�X�rU;�����;��	J�������'�qJ��$��\t$��݀Y�Ћ�W$n�w6V��R�ئA�S��8�X�.&�B��I��P�[��Ȣ=o�$�*-3��"�j�a���b9�;��Gmk�g?��*q��}����`ђAN@i����1�v��hwq�,96+��:�~�O�V�1��w���a�B`,��בݎ��qk��������U*��]U	�yҶ��e!3���B�Q,G z)�\+��D�#�  N}�<��Y�|��sa���>���R� �����3�3=Nj���y����	�����!.x�ɻj�\�<���pZ����p�xU�������yg����i��mP�X�?�;�S&8�Q�A����*'`�^Y��2;���0A�S��J���0�'��tLֽUh'|�8/���¯<eV2�v�)b�yE:�*xje#����2����*�؂����#��'�F���L~���o01EK5��f�֐��͒��U�H-�-U������B��_~���i@�24Q5c���r���w���81m�9�P�n�5�Rdrg�M�/-ȉl"0]]!Њ���y�;��	��Hg�]��a8����<R��]Ph��+�k��`��5�Lq��(�x���r�/5e@�����
��0�$!|��{�q�:-�q/c�@�&��j�58��.�QD��1>��w��≽,k�qkhl�O��"�h|d�eB���b�<���ĸ{5�^�jED?�E��	�ל[,t���E��Nyb2�Ĕ�y���'��/�����Z#��E�~_g���]?_�����j�V@��bYB쇓�Tg�c��C ��T}RI�y���Ev�.XC�/r�,�n4�w�I�%!��1���I^��SF�Y��f�;���a�d�d$B�a�'���+�����b����F�]c�#Լ�d�h� j`��v�?�N��"�N��
��#H�F��Z�t�'�;5t2�M��L��̷�OD��f%�>�*����b'�̞2�)�B0=_8C� ](���Q���V�qfI�`�Dw��n�C&��9G=_�6N8�c�y�t��F�H�8�����د�V%�󞯘�[ފ��2.��/�	B;Ҍ�02$�מ�����h~��$��D�Ͱ-3���HSy�ŻMrFfuח(lX�8�-!��l�|���v��M����N��[�o"dh���^^3�Yz�(h�U���;ȃwTYa����b�G`$^h"�H��6[���w�=��������:6<�t�R?p1�6\�Emy�������.�U�3g��}=׃z�]��m0���`��1���Y�AikA#\H�EY�"��L�ǻ��_���s�jQ́,ټA$z!�;� �~�}��n8���pV�ј�4�h����,�<��b�� ^H�\������5����QNU
x��{�J�O��	+d[�+�]G���|e=]�@�^#
�I��Vt[���,�������_� ��w���}=�= �[�(7�;�(�����L�r �X���M}�=O:�����H���|
�w�$�N*�i�� �?"hasD�.��.(�Dj�Q8���B��v%�*�P 21n�:^���y0[B\�����ʚܭ!X�3�Q7Y5���b2���~���[Jx�[�Z$hJP��Ӯ,���R�;�2�E��=$�7�����Y��j��N��K��b��
�E�_��K��9��&Y%���-a����]3��j�9���#z60��D�#�Y$X�A?�j��W��_zk��RD���Z�g�m�y+�ߩ-�k7؞������
�n@|r����&V�&jE]�#�P��ػ��?TSL�n1 ��@]�]ͷP�Di�v������[!���)����m��ԡSn�0!�-)� ��-���S��3�{u���\�ױD�-�w��7���xz�5=`��@�hYz,_D&�����ɢzLLO�~���)${E9������^��ih$Z/�~��A�ە�[�@�P#��z��0�'���y��C�z6�E��O�Ҳ`z��V��ⷍ��.�����(�4E�-��tO��6OHR�JX���:3����q�0�V˧�_Q���H�Z0B_�Xy������v��iM*���� +*�|�"ʬ�tK���an���n�D;NP,U\f��mc7��n❴i���g���Ms�gE��J�f=���&5�=�kQ-g����_����%}�.BMQ^ş�*Ѡ0�#G.�~�oD�r�	�֙Ň���[��$��`���c<�9�M�`t���%�t����_�F�$�?�	Ǩ����&k�|����b��)Q��ŖXI-u�2��:!(��*@�Q�$�8rQ��܅`�_�!����A�Vܲ�US�R�!���*tr�puZ�GX7�G�~�4f�{9��>���A��e��i۰�H���Q���R�B9d���7�42���+y�Έ'P�O2��c��ӍR�����d࢜�v���#ae /q̈́���^�R-w���K��q���3+x���
��K�և��gjg<�Hh��-+UƯ(�9ԾѰ�Iy$���2��6��M��-�A���"���씯�.���F��?@�px���J�#(g�ӣ(���͢�!���E2�������1�k_��-�:����b-J��&����YH�t㸒�����m8���<1%�Ӵ�����1�y<Tg�l�s��2qF�NgRc\T�!�_��_ؾ��L���|(��4%*R��^f��Wl>Kvax�e=���.�Ih!��	I4�Z1�M�y���8�������K�x��������!4r���Ka���U�o�%�NM� �LC �	�K.�H5���xxJi �)�4��x��|EP9ڿ�nK��*��s�x7���{���FD�'��!uaz;�Gt�eB�1��H�	��f�>s0;fQ���JʯV����H����$���Q�*�v
��B��mn	�`�A18]Κ�9QB�7�7e�e�H'���(�_Ԅ�^�t�Y����~,D=�#C���Ԫ.?��D�����7�J����@@]⬖*?����g�3���!�H5�Ŝ�X0�>$MeCK�8�O����V�u���Vӡ�U����>,�8��l�7>ޢ�ܴ��hX��Y���������r�4�3R­��2
�i	2�B�� ��7V�K�$>)\E.���U���$�v��C)w�p ���[V}�8��)16�{���_�i��������RGڴ#D��h�U^���Gun�i�����ˎ%'J���A�z��ķ����Ƚ6sޫ.�A�  �t��:�� �"�ޟp����(�	���������H�'%a�W�Ma�N_�Ԡ̓TfE1����B��!nk�^�{x���G����X돱�7���2I��,9?�~;K�h:��k�8 B���o;�k�uf/��$ʦP��,���z��YS�޾�}x�$�ƚ�D���o9�2�H
R��i���v���ոx�MI�n��r��Q�6�X���Ƌ:=Z4�=; pg`�1zܨ(��}���˒�X��!��Ĩ�Pv�h�F�`��`7ی!�����%%����;K��#�r@�gs���f�ػ��R��g��f�@���;�\20�'���Ţ�!Fu��w1���
	���J�^�j�����6x��b�?%��x_����,���ؘ:R��)��$#R�[�J�l �"3��'�yx�$%�:�f�2��9�*6'&X{j�`t�TBY��b����a�k]t� �ػ��(�>j����>=�Tk/݅��2�:$�k9�&�j����}s�^���ު<���5�/y'"o`%�T@�AZ<�ܢ�ݮ��}�J�O*��Gh�X9�y�ޗE�~&��o:��3�i|i�e��,����7&�P����E��#��Y/�f�7E$���v&f��S�"a{�_�+y	�x��g�W�g8
���e[�qsK�|�"��E�C�d��yB��Vt>��K��&�'���eq�8�b��J��j���y�;����0`��!gp���D�'��������|u������K&M:Ԁ#<lQT���JGGxܰ#v�VȨ��*����j��	m�î#�@�C� r�C�~Z~��B��c�l���з���驴q<w�%T���g��y٨���R�T�\oN���8�vw��
+��F��h� VNY��LO�U�d1V�G���(�����P��zNG���MӨ����	��;7}��SHf�cw�2�ᗙ��0'��
���Xq�zӯ8gl:�y���TP��P�о>�Ŀ�D�rϒq�F��N+�u.o�q���TuX)v���F��m�&QGq�t}��xX�]�L���zɿ�6�b!vC)��ntM��?�~
��6`��p�GsF��l�1��DH;`���ț�~���/��=ޞܸHD�\.$3E���o�Z�K��܍a�G����5�xkmo�ڮCUn��l �ޠ���ɭ��VU����B f��ptڛ9�?�b�>���+]ډ/8W1ҨC����X�V�a�?�i��5�3(	�M��᪈��m!>�O�Q��HBO���X��;|����d���0؜�Sע�cP�H�H����F��*Vl��aآ3��$�`ՉA�(EVK@W/��KP���v���x�)t6��}�B����Y��������¿�Vd}�>�8�ח�e�O3]~��z@���W�D}W㩜U�R����p:����e�Z� b���ב~�I���'3�I�<��$�ϴ@]e4FR\2$��o�������D��F:�RG�,�I�d�r�~�t���Va� f�8�T�^w�QM2m/��Ԡg~˝��P~�p���� �Ks+��ռ<�,���>��۷+�o +�)����`if����z��=`�� ]:�t�;�U9=��ŭ&�e0�1E9j���U��j�G�S��NE����E��pɺ{4؄�~��E�w�B�ʋ��SH4a�H��P^$��Q�Uh	���_�?��j#��c� �Δ+�ӈ���L�4-\W�13�2��B+z�3e$l�*7�s���'�r�J��[��~�{�ˣ�Um��$����*~��9t���ͫ1�8s�B�$��7h\k�K1.�؃����~�yMƘ%�8�B?+��C��i&"e	��w1�m\�r�-�~EE����g��#�_�$���N�H��%ẉe�X������Ҙ��#X-(+��!@s�2�k�|�g���x��ᕸQ.^{e!w���D?R��w1?��rw����>q��������0p��O�&Y�X�N/��Y	�T���"�m��ۈ#O�SN�UR�hs�ʊ��7��/,hP�y�oUx�d4g$� �n��в�����FY�x�,|T��C�F�<Q���%�D�nӚs�M	!�"�Z�]�*
�9�L��N��1�Ir-a?'Qy�m�}ƽ��")U�P]���R��i�ۄus�l��a��u��Y��uQẖ���V��v�O�x��W����!�<2�����O������|�{Yr���g���-x\����٫�*Mr�K��Y�������e�+٫����@Lj�+v?�VӪ���*d�<1��vc�k���U����c��-M)�l�����M���KQ!Q/x٭�<�����w~��e���3=�>(��Y�n8��9�&���������߉���t
w���@(�u[�4c�N�Tq�]p�{��-�2b+t�x&����k|�V�g9z*I#��qv�>&��T��ߒ�_�Epw�z����?\�׶4��ƣ�h\#L2s���Us��֯ ��X���:�S���	�m�U4���k�S����V�b��Y/ڋ$�9�1�sXU�P W5���[7^���`l�4�m�[\�k����v~"ɹ��m�6 00��>?F�h����m(�aZ��뾋r@N�wd��L��\��f�D��G�b��[,jO�BG%LYq�jAC�偦��smM~�1;H�kR���41N�n�kU*,͛�[FH�."~HgK�ep	��+� p�1d鞴3!q�E��:���q\�KWl�g	����,(�.<�:���9�O�zs��L������h�G8��M����E��)X��a��z	ڸ$�҂���2��xZ�r�\7~�:�0{ׅ{ʑ���]��z���Y
=�.5ueI�`幵}]0�%?�%�8ĩ��U6�č��ݧ@��#��8�\���� �/e�S�@����8Ú���P*-}>�3sF��D�������e8��ӗ��G�ܦ<��S�Q��9���4�e;"r��_��`�m!���d]�U"�5��������݉�V��3����,���gܠZMڅܫȡN���}�{]�O0�V���ı���1;�����âfS�,nw��VDc�6�Лܲ��{/�pƕ����l���qJ����0����O ���������x�ۋ 'M��������e,d,`Q���H[��W߿	Ivl�3�rk�p�P;�%0_ySZ7��i�{*�S��7GN��'yGu +��;$�c��3�������\L�T/�U��Ϙ�9��xnM ˍ�+[^��H�,��{����.����N/��m󑁮�)�����7۱��r/�-rڜ�?�N�����[� id(�������/u�ӲB!iC�I���kx��eT��u �w��-0��f��5���b���eM>�p!F0�jn?a�L�d���n�&&��3���R���O�]��E_>��ZI�.��Ā\�<h�#�a�1���h��\T�j�CE���U��2va��|�!����vـ�{l�
��z���nF�)�,K�ARW�&���2'톁$W�4⳵���mR���܋����R��iE���{p'��b�g�g.ݶ���<�����\r���yuH�9��������V��"��
SV��I�,�XM{5�;�:��Wv���SGSm�|=^?2f�a�C
��NԽ�p�s��-�[�J�
&Z!2���Q�m�� ��Q���/
�N�̀6'Iec�>V���d�ZoY!��bp�p�A�!�����;�r�ADE�ڊ���b�_y1 о1Z���'����3 ��,�к��=�$�"ex���Qs��z�(�.1]���iW0��3��5�� $��C;�u,�"*\���˂A�F|;��g��ߌ�c{��"� �Br%Z*���ړ���U�i6ю_�&�6�ȹ��e´Z��C_u�b�}���r�
 �~4���d�?�P9�c�q�W�'߽��?}Ų R@	p����sj�zm$�V����0���ž.��B/�@���*��CB?:�9>0��frdY�[D��fzB�F��Rj��Gx�����4�,D�ީ�"�޺&�`�ރB�J���gA����W�쉯��˲y��ވE��ĩ�o��Je�yj@�u��S�T��LŐ�i���Y<�.�]a�X�J�;!�k�W�-�w��/Nz��������K���DM��,2U������Uc2�J;�x8�����m*$����<K�R�D��L"�J����ƨN���-�+ՙa}��ÿ��XA'|��W��iDv���(ݝ\��=L�PKfyl�ܓ�#��s��C0>{��\��?S�D�F[���4�"�^����{�C���cC�����i�t �Цj-m��k��`ꢧ���*�����R4괬�l=0 x�렒[8{���7)��ɵu�Ż�B�/�]D�����6O�y�܀���l�����:"P�'|��ќ���Y
Wvl�
rđ�c���'�KƢ0�?���a�Q��oГ櫠Ne�G��c�g*� 26ʩ��&���+�ʫz��8 ����U�{{9:����d�-�R�;GdZ�2��v�Ò/���>Ҍ-x�����Ӣ���G�8'�B��;x^�~i Uf4-�p.wŘ�((���t��=��CLvS�j�uI�v@@�H.��L��vд�b�:*<��Ԃ�/��l��l��M����Gb��������@�B�r��9-n\l@�p��j��9g���k������uhF-Y��k��lL����Uv��$�\�P�'l�X5Y@@��9�O�juP�bY+�L;do�|ߤ��(�9�Y=�>�#�u����yG�b��ݛλk�=ň,. �������W�c�� ��rNM���g܂j,NF�Z��
^{L�'�k���ペl�2pZ���E�ę��#c�H'a�}Ε$�$(V��U΀�g�-��x�m�6��^�񵌺�¯-;8�� %��6Ԓ�������x��T�� 0]��H�if�}p�$˖*�y9�a!���ܲx�Ј�H�-�Cu�[@"�tOh������㳭����r�.����
�m��AE" ��$�� �\�%d�K�&QVc�kK�mWL1ɺj�뼕e�6c�h;����w�8�-�U���F��(	؟&�Gm����Ŋ,����%�]kyk!�)��m�*;'^	��k�乩��M�ybo.���{�%,e`�+Z�L�u����XZ���wg�K�M�A|���K�����m1���!�g��m�t�}o�d�j��t^�O����u��&�F��f��2�s�o�ۿ�A����Ŷ��������ن�;����6�j3E(��"Z ?�ͥ_P�M��zd��4�b��$B<(+x�L�������wE���1��e�����el��t������=�7�����:�ppɟZ�U�":��]	��r�����"�	��U�~J�Oklr���u�l�
,��2�+�z��'m~����g�������Ն��l`�Yg�=��d�m�B'�� V�I�r̜�K޲3��*�5(�#�P��}F&u�Z
�� ������+� ���k$�_ʝ��� 5�f*&p@�ϸ�g�~A�k����n�}9�ߴk4�� �WZXwo�[��1`�lw�b����y`E�fk�����X��M,�&�AM`M�r��e�Z6v5L�����NzB�CS �@)��J����u+���̡����Uc'e���m"J�_�Zf�	�"�U�F���a���I,#�,��֬0a�E�-��,Z����,E7���twSLCD߁g��*��9��t�����y�-�%�ĺ���ID���̓ v2 �	>�Cl����pk�k�>T;�XU5�$'V�zbu?R<�+�C\m�N�R��qT�=�d�`������L-c>�a?�{�A��������i�:�����l��W $U���`��F����w�n�|�S�V���6$��3�\�T������]�\�bXI�x�ĵ�]�)ֵ�~��r� � v|T��^a���Y��~XB�/�#�)��>�~{�~�Do�Y��p�9$��aև2�P�����w3�o�v�(��Ux�n��d���~�-iI������ l�"����3Īo��B�O# ��;��P�N�y��*��F�w�,i3��{�Ӽ:���fm�7OYg @}�A��S�5'"�LP�ϱL�͒����>�ʰ׶�a׊ƭ�I���ɫW���/����2�#�|Qz���uJͯ/�ʴ�Zǡ�Di׮稁S���bu��h��.m�,�j�y@�@X��V����(�����U��X�m��9�V�r�	�lZ�|�*?��2Չ�����xA�Ǭb�n]�`P��$��w����Iޕ�,vO�	8�|�B�첹>ؘz��X��y"N��&�(9�,a��x�'vT�qy/Ahi3:^c��Ǎ9�ri@�eK�1����8pX6ͽԖe,�<F�S�w�myIQH�h�T�.��M	�WyX%�����^��@f�Ù�^�+ Gj�đ��WM}z�����jk�@���|��1)	����?��e7���G�z���N]�}��?&�6�d3>���7�Lm��[�g�|�#�h6�R���I��8.�ߡ�!���m<h]�i!Nb�;r_�&�I���sA١C�y�O4���#���T�H"�Kx�S�t�ݖ���Z]�6#V�G��`	ԑ�$�|#������ ���kK��yv��b���Ƃ�����&�j	@�R��i=G[����I�QT�W�� ���&�������5���-���q\I:�t���aT4�p���]��$H'�z��#�S�*�v!�}���%��	�@h�6�3���o>f+�	/����1 �/����u��CRl�z]�
�_%�:@[���
��UA�=%�,�`�]��R�]��r����{�8>՜~��RNԮ�B�������������s���&j�=>��\F����'t?��ZU�Kd	琻D�l�5���W���9+x�a��)%\
Z-�dˣ�x(2��� �e� 9�����m�}rN���\�l6s�mS)�m ��r%G��c��s#�ZG�Z���.v��ԟ��D"hF~�i!�Z	DMo	��mp�t�%l���j��_$ΒyP��BR���3C����4�A�xL'�A>��'@HR!���d|�E��-%9�1��/$��0>�$��Yڙ��O&���mK�$�m4]��}�=���&T���).V�D�u=�a�t��b�鶽�_�'.b�C�9DPn��Z��={P_>Nj�i$�Ģ�C7n<{4Y\�W��D, sL+<r�[�jA��A� m��{��6�.7�'(=:nY�L5�BN�����S��&�L	)��L����`��,�(��M����(U ��2���} ����Dʺn:��}Ŭ��;���9��:z����pC�X�����oR�_�KA���h`���+�?��P�e!@��A��;J�;�w)Ry���a�9a� Yx�]�1b�Q� �~�B��Zv�8s����J���(��yQ�'���d݌c�V&/��5�=Y���]���L?�[ }�= 5Ѝ�����d!��!�N���k&'�3����te��	�°;jm�AAZC��������$f�b��cQ�b�Fw;NJ�ח�2��n�T�� `�%��_GDʳDiG��b;�6�|��H���Բ�+T�����$*h��Z^���'%��xT~UW|܊���!�'��R�؈��|��}�%uk�<ߕ��P�ա!Z,�m����B��А_x3eYз�; /�=i���J�����KD{��1oƠ`ե�P ��˼���X�}7	yHJ6~��"�)�I�t*��+ &�v��f:﬷k�����7	nM�q�e�8��� Nqd�ǋc�%'�
K���{?t�m ����2v�$���8}ʂs!��^�o����u��w�3u�^q�	:_�+�GT�v�l��q){��u�U|c콃���]�h)늃u)�[o�������A:�8e3=s�(¨�X��
z��Id�6�����G�r���N����g�>�b�>�ad��?O��[������Jp 6���`0Fd'�Qɂl�5� ��P�����4��_�(R�'���@�_���#	��w;Jg�
�I��& `�ԅ؞.�����m�a���*��UJ�0�%	(���Z�;�i&�}B��hߢW�{�E���ہ���e�2ҏx:$��]�2
����-�&E��n�V2�v�;�G1u�����*�����7f��+�j�E�}�Ғ�U(z���4{=�Zm&��	R��p�J���M��.b�hQ�t��6�;(���l�U���_�O'_CI�/�.�(m��!,9��W?�#	���������@A�Au@�Җpb�<��C�G�37��@��m)�8R�ŏ��!e���Ȏ�3�
�K`]�Va��E�{A�`�
UXz�({R��G�f�y�2�=U̏��M]^�?�J�=<� Ȅ쟞^a �DB��7ߟ�ư�ِR�3��N�>�y��׏��؅̉R$M��{ܛ����C��a�gi_�c"��*eo@�rX3 /ӵ��k�?�j�,�L�9��j�!�ˆؒZ����o�g��O��ePD.7M�m2|�h�����4�)�6@ NH�Nɹ`���"�u����@-&���	4]wJO�mI�����TG���Ȼ�����[���S"�i�ҨE�W��^�)'����`�����]=�c�Ӈ�<�%�#/�RZj�S�`���"d��o��A|D��7}_�D�:p��B���t:(	�QB.�%��:,�[�F�k�aV����+�S�3VK�'X�h+�s�&^i`$D9�&A]�_��_(r�)*��!�`vn�`���":�T��>���R%��&�����ˑnxS:�-�i	ԕM�;�O�m�b��+�A*��PU���58�<�&�jjb��c��q����Κ�>�ڠE|�D.�3��=kӿ"�s��:L�㬛�CI,@���q�3�jNJ�QZ�h���E�hRu�2:	�������k?����f��qE��H3	W՗	(��/aEb�	�Ǘ�2d'�$�Tw����=�!՗,�w��P$��	Q�������������{�HMT �52�+�o`%��MG��I���u 1�8���W]�o%p~ �;��_z����}�倗+�e�0ui���x�\��s���U�au��4��_�E;�c�:��I+Xā��NA��ڶv:����妗��4
�T
r^����$oh*,	�͉!�Σ�aE��dD�B��SP�B�Cfj�P�_�(}��Q4�$�`yT9O��im�+rk���i6�NU�������~�ř���T�Ů���#
�B�lJ2!6~��t��he=_�I8v�כ��ĺ�4���w��Ȏ6�w�����"ļ�oL�\µ��a0��~�����z�Q��:������h��VzN3�h���R�]<��c��kʪR�`Π�QO��J�����E�)Os�]��=�4�,|(�ɔ�_ܟI�ز�4@��N1������ǂ��C+�y��
�e���5��y���\[���~���*>��Q�_���c�ǰ�	��H<Z��v�)�fn��/,�y���\RzZ���6�ҵM	z���:��i�ҍ����+��H���d�7�V0e�׈j�и�@QN *V b�gr�h�6�sc\�:�׃��'1���r
p��������R��5�!uH����iu/{�f�A-��L�~<xn��,��"��1-���/�ބ4�2��W�f@}�
te��:�x�g�aV=�<e2̦�,9�?�Iۃ�P�m}小�6b@]K��X�R�at,ZSжJ�c�G�]�g*�ב��/2���ķ&��P6p.o �o�T��ޯ��*d�
��(�]�<��z-�Ջ�ߠ�#�	o��ZH�*Ei����k����Qx����1�ė��5�氟Υ��2�9��٠[5i����+1/�~��o@��CgUW�A�_�u�{�~E����	X0E���z���Ξ�4���.��A��Q�"�5�;mX\��ƕ��o+��_�Ln���ge��pf�U1?�8��~V\e#y)�
9�!e������֌U�B� ���lvq)�}�K���_�!]q�s]!K�L�M�^y�:�+ӎr8&�$Ҋњ� ����� �4�;��#��YgWC!~_<�!j2Z��1/��4ԋzr܎�c�Ѳ�T
��&�
Zݔ�?©���9��Mp%u/Q~_�s3�����Zhh�KPӍ�i��5�����A�[[�YM��*a��b�����&W�r�:�0���W.��ɵ}_'�X��SX�lQ�y>���mF���~�'[��h���ނ+�*A��\��e1Eb�������������g�����쟨��T�~�8��?@Œe.����d�����0-�UP3��rmC��0 �h�
۞��F�;p5�C���W������8�cϰ���۷ ��{�Hi^D)�����t������><��P�V�6��\�����V��$����%ٝ��C�4~3ػa׺V��m��b)I���9%�� .�Qx}G"[�gv�ٶ�k��0M�V�&�81�T#��Y���A\Kv���w�I���3t�u�����F=#��~�u@CPaZ�l>�E<b��nx�m���ݕ	=�:�߿��>t7���_H�W6+q[�Gě����A7�v���P41*��4i�n$5c���_:H�Nۖ���E�}�)c+�Y�f	?nc�|v���qc��VO<P3��� d�a�.�	u��<�Z��ᅀaN�����+옃�#n�_����u�L�� ��'���2d\��ε�K�e�w�J;�*��MAp�Q�p]�	8��k�C����L�g���]��W�cFN���Cq;�t�h�R6py�{B�>��4\�e��B�;��R��J�Om��%�)@�y{�f�&������%�o�R���<�'VQH�m47[Kpjd��
lC&ր�W��/B���mg3��{v+"l���p�M`��zF@8P%2
���+���L������)�2'Rvq��#����`z�XB�UeRr�P1j�\kv$B����.�N��׷4S��q���~�8.����x��!!$L~\8��R\-���7�I�Jz��Ч�hV���
��j���
��r���{��d��7����곯�c���0J�&Z )P����.~?"�����Q�X�k-Re�5�@jf6`�b��G����t$�iO��A���f���!�9� k��Bk�?�l!@��ɮn~���S�S����}�\a�f���'#���k.(��TE��y�k������:+(�g�	4Ϫ���Q���aZ��Q��8'_0=�����f"8+��rK�_��z ��4���Mx�wƆ�����aj��3�ςߒ�NU�lXq�~��?-
U[kv*��ؿ��nz��캶q|�޹���Q��	� (��>���z��/B�ֲJm�gE������M��k���{�Ax.��ɑ1|Bߎ�Ƣ��/c� f8���m8Y#��m��|C���]>Q�X 8j�my�ҟ���e����c4�N���(�����D����27�7=!�x�������T��T�3�!�H����'nE�߄�RJmb$�Ҿ_|��q��*�e���Cr�8#�޹-7���Z��b�����E��O��h����.�	���(y6��U�+ $#(КA�0�o�nk�>��|3��8L��!X��Ft��n���B��k`�Ug宖�����U�Z�IP�Ǐ�ߑ�&�q�2h�'�p{��C�ݼ������x�L�cj� �U<I}D��U��z�-n�즍B�s���Z<�Vt=T`���`B�s�:��Hnʦ�E/���`���g��Z��{���aG�g8��Z�ke�7��B�~u����ݡ��rKw���K̅�qi�O�c����m!q�� Dz�U��}	�L�zz,e2��ޚ� �j`�����&3�u��^�k	3��>ѿdp7�����
�O��Lz�|����CK�0t�6�A�H�8��!l�����Cy��0~J8��)$��Yt�C('M��[U�H(oz��wx�9b9��.��u5��"�}Ƨ�U��0ӎ���3����C���ce��УV1[�7��3������� ]{����
�Qq%��s����[SȊ��>��?��~����Jƪ�pF���Mp�N��G�١i����5��_	�ߛc�s�w냒��
I�+����X8!J�43����x�Sd+e��t���v��Yi��	_�vϤY�c{��
����d��*U�6���V�a���Z]3�0�k'&�2U���Ƙ��G����ec�#N�_�4��.t��T�}L�X)�zèx�t�Lm.Qk��^֡���'HO�#��WE󟆷!~�nR��m��U������!�g�ο�Yo�y�ӈH����h(�}�I��<�Í��3�fȺO��f����/�� �����ǁ&�-�&�~�.��߻��I���%Bـ�{�&�4�?����Y���N�,G��|�F�7 !�\ڽ8U�vV���x��b�5��7����J�r�^P^�I���4��d�L�ͽq���#��&�
���J5�}��b6��|MX�0{���[Uw_/��)r폎�7�.�����ܠ4�ַ�����I���S.#�݈8.�fj�m;'_81Gy!ht��sA���m�ĭ�d(�G�c�&
b&��^�s���i�w����7I(��0Hg�4�V(0�]#�2���h��C=*GY�Kw��/���*����$��3�,��;x!����B�Q#��߳����wV_��}mTR�>������D�n\��$ �lnλ�埰i�&������(�E�臛���s������^����̛ T��o�=O"t�ƈ+�L�X���B��Q� >����vm�g\�A![��Mw0�6}kf9L`�`�d�},���
�**!�4�*k2��5�`��^�V�xdcMw�A�N�B�u{�>���%�����nZ�|�6ǏP�s�g�ءe�sn.�g�۟�P�D	7h��MO�,z�V���fF�T�ek��'�6�7:�b�&I�<� ޫ�z�,��fOw�J@r�.�d!�G5�ud�y+����@%(9{�i�,C��Vu��������ݦ���W|L	2��k�T�����w�d
ɣT�p����F��)%�_X!m:B��8*�E��?iKHd�����_�S�����*�����LH1�U˸�k���
�p~��6i�QrlvJ��)Ji�������NU��$���zgi�2���)�	[HI��xR����ًs�� ��j���{"&d�ˏ 	_�e��pYn��ӛoZ�on�~4�'3�Q��e�-�ւ��uǛ�)Ɩցf��f.�3P�JT�6��2ք�
��0*vY��qV�!@t͝�ڨ�kW�;��+F]w����Ym�^��w�uX[W���`r�������k�Ti�_��Jx����n�=k��C�M����r�U��Sd�L�m�y&�܌�憀'j[?�P���8�s�|��BT��E
!�>)�2�֠3ء��m�%�-.��0ir}��Q�I���:Q���m�.{�(�)��^�a�y)g~�~�ϓ��:$�49��O젓\���쑚 ���H)�a���]�ZN�,��Ph�=�jQD�<���<�����z�"���.����?�A:jKE	TV5'�w*j�x�5�;I��f�Ha ����f��&�?�7�Y��-�i+�;�-*��˽9�N;�mXr��;��p�������7p6
���b�J�&.&�B�ޙ|�����j�Y4��,��WA���2��q�Η����	'ל�S�9ݻQ�H��
2��}i�b��g���/�����?�A�������m�����~������7Z�i�k֬��^����5�����^W���,��q&d��n�O#��oL5��aO����Va��W��c�I��j��kP�ij�pO������=�[��W ψ�����M"�t��6V/9��v�"�iwdzk�:��֨������A��;�B�r@q�4�X��Y��Q���~�x?gvo����)�L�E�=��	
�t�㪸�Z��K����%0�B<�R�܃�L���٥�cas�l��I�cY�49ڡ�q23�g��{s��^���$���/t%��h��Y�!V��0��^���]����O�>���&�o�q��m�s���	�|��;�j�4�������ԑ�U�-]��am��O�g�t�T,�mms��!'�to~}�K(zf���̰D/,���C��/��㥫�0��)z��hKo}�j�0#�������d����6�E�
��X�yp�)�`t��z���I�������|cnM��)���U}�/����bA����f��$!�eUgt'�Q?ooĉ�4z�#�*6ϴ�����>�.�\TL�����"�g�#~M�<^T)�C���pC�W^�6�5hrQ��6�(��wM��/J��X��UT�`��?۳��N�S�sΞ"�@�LW�_l���Cl?����{�R��έ�˼����f.RӃ�ӟf'pWX�w��5L�ST�f('C�y�J{�,��"7���{x������:k̯������?��8����B1�
t�n;��*T����3@�)$A.GY8�{nv/I��{��J;Ѐ�j��p��2�T��ю��?.��`��^����ǌ�LjIn��g9rbs�ѭ2sz�n���hX�e�\�b�ˮ�ld�V�\I-6�)QL]&�̧�B�u�d|�h����~�=\I������>OD�sB��Ȇ��R�ƹ'Z7�}�R�>�'���ِ�>�:l��S ]��H�]�<�E�\��,m�Wqzx��
�\v�ߡU��托��J���&�)�i�>5��ҁ�H�W�l������m�6%'3qϭbF��m@��d�nA4��\�CD|P���V���H�DԼ�3.�OL�gفd���.����c��w��Z�B5��ݚ���Y�B�㏉v��ߒz�Ҩ�:Yk�N'��U4m�f��Ji�yݔ�D��Fz��m^m0��zbQ~p/�lӰ��wz��2���믷Wl�h����8ϋ:J�'�\��s����9D\oۃ��{�YDRV�Z�2�ϲ^⡜i@=dׅ�7N"�n0'
m3�4������/��iU|[��-�k�u�`�k\�m)���� �eTMqEg#<�'9pyvo�ͽkL4�[�Sf���)f~���*��Y%>�+jѦk.�������ht��[�x�/��I��Vjה��] z�V�ex
�)U��;gh�o�(���,m?�S1���E��?�eH-��o�u�g��	t�bg¨��S�j6�_�/ϸ�_��
6���Ư�d-u��7�\U;,��="�mgCy��Q�Y��o跔�eG�{=�g�m��㏻Ixu�l�%�mt�ы�I=��qT��W�2�*
�!��F-�w�{��u�V����J�;�u0|�����I��{�� `2-�9���b �8�}�1K�(=O�Y�V�0�-K�u��L���'t�i��9�H}@U��V,wM���6�i�p�J�Z�a�� ���523���䌇X�Q�[#}�G>ol|j2�HGf�QѐQ����L�70,"10��}?{�����e=��,o�:d���Z·�¤p�yN����mR�$i�P���
�E��J'��޻C����X�q&ڒ�t��z��kVP�1X����aĮ��&2�4�l��;s08�H��<�;���&�(��`~��Y�X��Ґ剁�>'���Y�lb��h
h47����g�����9P�,�����k��J�r�_����p��=B��d�Y�U�s�?��6�$@�}A���S3�K�Fk�>�����jfu٤C��r�sG��Z��N& ����*#G�I�7K�?�����r�Cri�c.R��{jd��r��zj`��%t��S�5y˖"
�s{[T&7��c� wk|O�]��Y�,��h�Q��H*���Ѭݙo�s0��8��2f�`�T�_!H+�(	#���5o�Ԯ�,���wӦl����P˄ �x��Oi�R�V�Ր��qۻy�d
����`���x��qj�HH9�w�(��x�^]���:T����ehw�Ф(�'{2|g5*iG�Wں��'r�##k4mcc�?R�h21b ��!��P���бGBA�Rb`>��'���L ���]Z1-HK6�&�_PO�ȕ�n@^��G�Ll��?�.K�;�
o��S|a 1Uٟ��n���L�r�?�臑 ��Q�b�@͚�W��<۳��t������l}���%L׶�U[[X"��Sh�ЭpL&��
��W���6��]�.�FR57%�O�������O��*��;�u*;�@)b��e�*$ I��1k9L����G)��N�O��6�IN&�� ����a�k~K��KP/f�������*���R����ꇩ3b�`@�
�n�!�	�n忞��"b�o���A���94��k����	��w�1�fݷ�i�}�v�b�nT�
�.���]��o���<q:D蘘�*B��R"hB,�*3�0�rߢLMr��|���D%Opd���2����#���ʩQ7 )��* �7-�i���w�S���M�~6$^4�R�·��RB]P�۱��0"u�zӫ~�`��W-UU�'���W9��=��e्�^s�s��4�N&J�0d<3,YvӨⲚM��HN1�D��(�}P�L)T�#{�б@�t5b�JG��]��"����%��|���`���/���7���/
�o*T}m�-��%l��1�V�I!KR[��D8�֬�E�N�<�3����j⮓4�� �A�Ů�O̊58�r/�'~�D:��'Bo9��PdD��H�T&w����ҋVwDɤJ�p�HMqW$��;uTc��� ^��e�]a� ��P��ǽ>p^��?m0��m_2O��x(�ͮ[Bx� �[�"����v@V���mr�-��̯�!WZ���ʓχ��>~�Z��J9[�7�ڦ����<Q�+��R�l��T�iw2��h�^��t,�ie2���?��	�]v#t��A_��?]�V|���Z���Colue?�}hm6�4'ʼ��&��&����^��y=E�9�ɟ�������hJp�+s�� �F���3ۂ��ߥ8���xwN��S&'�K��E}��^������2/�z4�ݺ��eZI)���-&�de�v&*sܱ�!�=������/��d�As�ތ�鐏[�#�����!�̓�
���]b,��T��Iw�1�;[=�wV�����8f�|����i�y�+�ײd<Ű�6�2*7�\(�������L-�;����")D>ۚ���qa�!\թ��%��b�f "���MF�Y1�i"H��`2�0T��R�/F/lQ��>*���bK��%�Hu�rC-���p���O c�KJ�My%G��v^D�v����!���N������?d��}D����F��
�_P�2�%�pV�9t�[�C�
%���L^\g��u 5�EB��F�*�}��O(�y�4\M盼n�wRBJ�	T9�,��m�n>�ɛd2̎N�-ī��:�tݎg1���,�	m]a�'���c�%�)�O�:�S��?)���|���We��T�?sf���~�Ĩ�j�����%VJ��W
���h�\\���MB�?ީ*w ��5�7��h��2��XwW�:ąz��Z7�J 2�]*�$*�2������U��n(����,���"�G�{�JPQ��#����� �)qb�2��~�h:���{#�� ��q��9�����F���:_��6�HgGp�Ļ�6WwZj�)/N�)Ő�;_Iv��|�ڔ!��`I�"�P���&�s����ҡ�����{�j�ˈ�"Q���=,�7o��p��5PDD5�����ꇞ]̚pT{�4YB��b;�>!^�xB��᫚ѰYtsSGW X�Γ��<��j*4�!<���Y6�!��z��h�#�_Zf��	��䟇�S�4��I&J�!*x��Ԗ�+9@L���x�O���S������-N�7��e���[��OuM�	S9��e��@$���>�7d��g���_������kf��A}�>q[��3���'���"�1���f�����V0�vZ��U�
�^��v:P5���eI+��H�?��s��[�����.3�;7})�=��8d�����8��3y�Oq��x�>WY�"Y� e�4�դ���ɶ�H�r��qc�S�M$���5����{	Ly�uc�u��_(�Μ��O=�4E�~�vWZ�j['Yx�G������0�ŦAL6_6��LL���O���3��d�t�V32��b���Mv#�F����Ʊ�*��g[��mg��)�N9���L;j��s7�D���\
0b�D?0��L��G�#r"�DSsj�(%T�0M7����s��� ɄU&Q��S��?�>_I�eG������������M�^g��������Z	����F����+��"�8M����F��qV���e�3y������E�^6��d��9�g@��M��䰳��g�B�&��0^	v{���p4���/�%}�_����5�*Mx�j#��?n�!�R�LJ��,Xڙ��Z��
Wz\/%��̨S�zb^.'2��e�c�(�T�S�m�_�G���c��z� lj���~�~TG��Jm�K�57�3���j��(�owQݿ�� h�Ib�H�ѭp�D���:�{��+�{/���/,r�M'䬛�F9Jݣ�sA�Wl��T�6-�%�}x���u0BT9L�J3����ĭM��P$�ͯ��os��B�2͋*Voo�w�̿G��9�7ϡ=Ah^�y�0�/����h;EX�%�T{!����M��Z�~{N�!g�����P��ݴ��X�]c��P6V�H� ~qcMa�AW��a�v�x������l��j�BCJ�E\� ��s��[LS�����#B�m�(�!zފ��gf���1p�Z��E2$菢ԉ�0����S��:�X*o�yJ���M,�����)�'���٥�ĭU�.��
D���}�Tj�p`T�wZ�c������ #�3��6Hv�ŕ9�6��_��)|��ONƤL�RnUTҏ"��"&w ��	UZ��F����We���3"`���q)��q����>�}�^�	����U's��L�,�����s���1�ְ��5փ�Ja\������	5ːn��dџ��6�da��1I�����J��?Me���չ���e���(�j�(�YTߦ� �&��q��@���>��-.*p���"�	�����mPPPؐyc�P�U�����U>������cOB&���*t����U����~�]�d���$M�j�,Z��m�����|,��2�sm½�
Æ�2~#`�i���<��X��P�
/*M!ՇS�v
<��s�F:8����/�;�Xm��R=Ow]�#���'I��jmxݡ�MnN�`��M����9��DmH꡼7�ӧ&_x�a<#�c�\VVkR�V�
�k�bO��O6_V]>�n���Z�eͼ�9�����p`�;��N*�&� �W7�2ͯ�  ���ǨoN��_	������=9�wy�䦂-1�sf�3Q=P����aLye}g�|��B��)�"�/�'r�\ȚJM��r!$f>ǋӲR��`9inF3P�)����Z�����*��:-�{�~�	Y> �fv�M��x���[�e�iA�2�p�x�V���(U��m/���1BJG[�����k3�2mLm�a����J�,�
s��X6�U��S1��o�ao�DC�T9�<��6c�fw����r	+�m(��@����������������i{�{��͢���q]�~�'����L�4qDo�Z�t��16e�aS��$-�VQg���*B�Z�70�~�fK�q�1K��S�����$��wI�~ۈ����o8��ԗ�9��W�A������X]�"�#~���s����ة9��AU�����"ơ�3�2eA��T��U�{�.�(j�&x�=w���ۦ��p�+��>�>��X�7�=�G���N#	��<����{��^e�#�lǰ�{X�Kc��\�b�s����S�f�_68xjè+�P�����D�I�Hc����{2`9�r�X���oi��w�?1�@��,��|1$.����8���b�jI�Ŏ!�w荶K5O(ܒ~�)P@��)}�喝`�T�y��s��,{X@� ���(��	7?�}�Zd��↩맙���'��	���o�S�����q-N�{rta'Z�}z�nk�r�@y�����I�?�NX�J��k.3��x091>/�b��Ї>-��q��^���Ղ���[�n�JS����ż�K�$+'SJ��c�w)ЊEO�����p�/^��<��{Y	�5j��K ��KŦ�+v�;L���������1�%3P�6)E��	N�Q���]��j��^1����5_�KV��%�ť+��h&���c���̝�q�p AkK$Jui"���-A���]�;�6Ga_F��g�9͆�"�A��)L�s�Q�h����w�'ǋ8Y�N)�]A�I���N����d�`N5pٱ�s�Xzm��!��Qn�7}���jJ���I{+!���5ة������|�V���g��P���c��^o�]��T�G�Ճ�'vݑ��Y,�< g�+�|{p���*��v�p~��Va^ΆDn"X�)9s��o�/Q
�x���҇��xt�pR�-�s�B.C��Ec��W����7<��棑��l�6Ѵ���y��5s��k�- �(X�,7d9�g��+	�'��Sb-�?�����7���J�O�v/�K�2E��k9�N���O�ڿ��w$���:!�r,a1h�~�i�U[��PaBB7�-����ϒ��V3��i�r��T-:94x|q��-��x@7�]��ns<��ou{����`�u���N�%����{�:��m�.�_6V�4���t1�S"r�O���Jo�����]Bi�A.`��jqҩ�5���;�B��b��l>��_M�_$��\�=�� ���%�{�yR��Q���f���}�:�Hc����.�M������� D�Rbq��Z��� �+�K��O���`�b�pWyD�0��.E�t��(.׆4��a%��{7$J��=L*x ��1��_K� �*-��'Mt�P�{�-e�M�W։D�X�=.v�To���;c���]A�f6Z�}��L���rP_�Ҙ�3Xd��k����~4#
22et��лJ�d�9�p�	�	�k�ޟ��3yvQ�3�Fn+CgI18w���63>�=u%.��t�w7�K�{���PSr��W���H<�
bT��2�p�;,z�����
��5�O����CC~�x:R��B���q�d�)��Y�<��o�X)���.���n�4P����&?=��E�$}�ң"J�-��
�a���U�n&��(i�\�Q��U�B�)��G�	w�����s�JA}��q���b�⋴�E�/m�?���| d������ʈ�	�քU��
D�'�ݹ_)C�MR?��`c���Q��e��x���2p5�,�@�%guEE����B� Pk,��sQ�R���젅|i����as'��R�>�B��V�: 2��I�0>p�����r
�/���`�h�Պ)��3�8���ƊVe�5��RM��:��!���'Ӯ^��l��5�I��ة4ԝQ#l3�؏Y<{X%g�A�s�߶���"Gf�I�����[����\�(��4͓"*,?_ƨ!��V�C�������>"��G��,����2�:���z+��.+QסF�5M&Gi���9�N �]l�p��?A�����P(�yI@��1O�"�G�֣E�oy��E^�y[�:34��Q�^
?V��5�oï�j��X�8`��|J�����suP�!(Ɔ)g�t����d^��A|_�aA5њ�]0��^]g1�!�V���Y��j�!)E}�g]��Z4P� ��R�j2�l��ԗ�TT����2���(��)x��2X����y���������.��9�a)ƹ��"�ݶ��CF��|k��k��t9���oī�e���}�݂C ��k6Q����]�f(M$�o}̗/�t���p�95�I�DQ�J�D,�BF��fPwPA��Y�r�XL�C BnE!�d0,���V��x�ژî�quF�]sԪ�cc�B�:�+g�+)�@4�"���#��nOV9gʨ�T�/�ɬ��f�V��I1�Y��!3Cq��9�L��=�� �*����6ɪ��g��P#L���V���W���Ƙ�1�~}�'F��w$zL���1ќH���!S9�\z��6�:L��SL#��&!f���Z�S�\�[^L�^��������d�U|N�N���R��Ō�}B��-�I껡K�E���4L��3�mvV��p#�X�u�{�
n(�͔��P�'r$�+����	����O���P�xD�S�_�T᫶�]�4�]4��y�D�FY��\���lt8�M���������+�Zj/r�F���e�6�@�FMK�n	̀^h\N���s�PCrm�f���!
�Ȝ�o�H^C�y��-�=��^��k�#��t;�/�~�Y><F��q���]�]xNk����u<y֋�fm�@t��6��3�����`Ĕ�5�rMtc*�cd cN�@CZ�u�$��X��^�/����m6�c��@���2�Y{�ST�ߣ�Pc�������<�u�/���l��~K�#"�zp`~v8^wn�'	��XР.�:��ei�)�D"�4���3��2����ŋ6b	��k$rj5er�(�)c\b��*:7�([`q;�Ew��0"�,���q��=�c��&e�TPC׎R3�}=KK�΅�2�1��v�'���-�Q�rz���|��i�' ��/�HSޣ�;�*n�3_$*��G���h�Q�S���#X����a���e�9��!|�_{�C���5݈�K�:�t��r���n�M�*@��CV�.q��׬FC9�v�F���u-�#T�6�����;/�!#mhtqsY���¯��w�05�Q[�9�㦌t]���j�}��0���쪮��Y�#��W��C*��>�'��w֛�T��z�����H=����ow�eOlB�2-�Ց�5u�C𼶚Ք�u�?7P��]�
��5E�L�Cєl�t�團z�C^t"��:�����ܢ~S��ԇ/�S>����6����y�eeI�B ό6�M}������ĻW�ƚNT F��_�['g���V��{��u{$胦)��=IQ�NK�S�.�5��Q)U�j�߅h�ï��"L����\�/���R�|S��$g��3��S�����v���Y)������R;D����m��2J�ɻ)�Nk�	%�G��F�1'��G'���5�,(��HXlr=g Ȧ��L�YwpN֏#���`t�6s}��]�*K���+vzbhM=a���� ������%**!Bh?��ϧ��S�DO |b�ת��:�=Wƌ�8]  33�Qo����zˌ�r����<�u���[�i��t�?zJң�d��p��d���H�]�|�`H߼~/D�^B�xP]��72���4@� ��sm�6"���]�@���Ƴ-�l����ؾSG`�x��u-�"�6�X^��s� ��!Y$�����@�.�TQ��I)*ܺ]F��Hq��� 3�^�N���[��4��e����r}"�>�1L^�[�$��t��o���ı��TD��B�Uu"�\��qJT��k�C�4UE�/pa��#�%����C���;S�M�Gl3��_�J4S�4GrZ(����hw�<��V%ØC��M��)�(�ek�JA0�r]
�,E8��)L�Qqխ- E!p��t�G�*(L���Ku?���(u�Pȋ-^�5|z��N��ީsM��mq�I�=P�a�I�G� N��p.�!�z��ϦWW>�A R�R�n��`�H���H�V�97|�3�#� �0��LC ݒ?o����Eaa�p��`{�ou5�u�~���r��f�,C��?�Ç��{ԏ!�U��!M�]�$S��q+�|������N�1�,��È��I�
��J�f�]Y:c�a*E������X�jqPzQʫ������ݎ���زدMh,t1!�<�K�tfXͨU����TbQڼ�S��Rx�n�?�W(gC�T+��P��s-��'ܾ�%���w�:F�	T'�84P�%�]|��v�;Ar�N�/��>y�-9i*��˚��ܑ\kj*O"A+;ەX��(�q� ��x>����|04���;�~���A��=>�`��^��X��
]�����~�^5��\hjv*�����!(�!Z���.�7<Ƿj�X�e}�|��6;�u�sH�nx��)������f~���>b1��e˺6i<$�F�a�G�K�Z�<g�$�l����(�~`����kq�ٍF�
�Vb_��&;��4���#q:�?���R�[�#D: s�E�Z��4D
	c��*c����3�;O�����	S��]�����5�B=�kM>3�7(�%*���.$B��x�`���OI�J�q�R����`G�Y�7��}T��
�����U<�Y��ɒ�+� Ȗଆ}-�*��V�4�(Sf��a}���e�$9a0r	��ɼ�>�e~��HR��0��R/�}foiV��H'p/��|�MP�*fe�(j���pԄ5t(%s�u�,�?y�E�ۀ����O���F����mh�Q���(���%�9xш�.�Q }��ljh�L�ֻ�A/�._�Ä�\_$�G]����+�nf�)N��*�e��8�9D3" �(\�B�}��,oQ�z�]HZ�U;V��$U"�#N�yB�s���K��Wٜ��ϭ{�\$��<��"$�;��c&$�q�@՛�I�{įm���;G@w|^h�_4,z?�kﳸ&�� ܫ�/|P�\�\1x�p,1������� �#dgj�/����R�)/��,���b6!N/z\l^�r��S�X���%���:�(΋sɅ04��UCᯙ�����7��������F��}pL�����Dk�V-h�	:t���!ʙf��&���B=4� �ol}�D9��W�5�΅�m�*��3���Y���ل���EoB%�\?�NJ���[f�����G���1���@�qc!I��4}�ڀ�)��u/u�L0�Qʜ�}	�Ϟi�C=	]����s�qkNCK����q��� �@��n�7z�&�[���s�PP�W02_n��\0&�����&�!O��h˦�)��F��e�u��3�����4��UKI�6y2�@���J���CݙNK�W�L��Ln0F�����Wfv�����OMVD���K��|7^�-��,�tv�E�"��Y��F��$�s��e�ˉ�o]_����s>/H�� ��t�~�)7B	�F��@��ƍΟW�hlV^���_0�Q�> H;VH$�r��(ʸh
��I,�0wܣYՓ�xb�yP��+F�Y�� gO�CļR�:���W�:{gs���D���9�������M��A�ԟDȖ�cizAҤ������-���'\�+^i��	˷�IJ�_&���u����$��#�1���p�k�Ъ9��	
� ������FS�c{������{.裓��� ͂�_�����ex��\�V?���*[�r؄�ZStc�W~4�9�����]#غG��M�x�_9 �N�CP����< �����3���'�>�gwTA���qX��J�햠v�iC5�u�Ubu#\���A=+���E	q��2ve�Iq��IZ�*��	��@�5���IEكS=�Ko��:��tb��u��O,"��k��U�r'�y��^��e�߫�.3����/o��Q�|_П��Q�#����^H�*q	�ǇDB�(Y��n�_jH���r�&N�aNH	@��=^h����������Yo ��`T��$��c����L�N�����"8��N��u*a��2�增�Q�m�ߪ�Xr}\�n�%��cC�_��<�Ǩv@����ɐ������U�KH��\d;)EA���ȂE��W~�Yrc��6���::�nO��;,��6�?���P�1*j����<n+��+:@{��5?�l�v�v^�|ǘ̄.�XJ��W0N1h6㥾�TȆ��D�UQp���|��
�l�s��ϸc6�����'��UF�q�����~���D�z=����ξ��
J�o�Q$�*������M������`��ϸ�H�C�wI{06���ɾ��_�Qm$��7�)��ɗ+Nj��5�1�2 �;AJ��6P�sx�X9U'�;���I��/T��*��;�y�J�J��maf*���<�G�G���`?�uf�S��'p�ٕL �$��eEh�ܧF*�8�C����^d`"y���F���[5?�nm��
0F�)T�r��K�έFl�ps=����ز��ZQ���X�l�y�`O����d���.GT��<|�Mn?��_��%?����%���+�j|vjp�U|H��&Ņ�e�9��&�	/*~��ރiADIz˚X�L��J�U����I��p���?Z9�X�xQ� #�7w���Q��U����boۻ��v�
 �u�ռ�I_U([�ib�n6�����R�ocM �dza�SB��o�~L�A�����ra�l��ݶ#.J�) łȼ�F�K���ݝ�{#��ñ���EǄTl�Wc~�?�c�BCm-C�.��N���\��)�;��	g݅l�?#Δi�=I��]V���S�.-Z�샞��tq���	�q����$v:Uh�����R����P�饛�
���r,����`�K��#��,�Rp�����/TN��u��!�iHw��8������@j�\��GBe4]#P0OV�/ß,Q��^�<����xD���Yc�`OĤ)�!�^7�e�8<����;��#+��*�[klH�
=�n�MX�� x����
mj�ktvW�ea���;M⟓[5�K�(_x21!�����	D�W�é�9: ��GXr�����i�_!��uK4�c!H5���ܤ4#?�Q�&�}�.z����۔X����*�G<������V�k;�L�r ���ٵ� ی�	�fG��T�N���|��F��֑���sR���ȷ���`x�
��xG����/db��ڬ��+l�%
In<#��H Wq�M����+���_J�(7�u]��^J=E��R&o*��B����P.W��D��|ʖ2f� Ľ1��MNk�C����>�F��O�y�ׅ�PV3���ҥ�Kn��ɵ�RxJXd����34,	M����{�9��v�e��jH����9�u�]J�� J{����Nd���p׿k\��_�~,�;��}h��t1�y��|��nT�\���2
�
O~��e�M��M��sX�87nD�+@6���_��&��#a�����ꋐ���I�4T��}���n�ƍYg��bF	$�_�l��nI��n��le�&�u��$?�^b��,�~.F��!��N��P�=ĳ'���5���f�lk�¬K�5D�+�p�r3ED0ݒn �k�"�|Ȳ�P�����H����\�6��>��-�(V�I�P�JX�2�Y?� �?�ڦ-rV�	�a�����mW�O=[�H��w����4
�F�-��1
Mwrѻe?�`����Ґգ.\�i'2�-ȴ���I�6ȥ�VI����C�U���Vh���ٜft�} ?fG6]A=�G�aL���4�e8�]��� a{�i[U���:�<�.a����	x���یtNS��U� �L����c��
��t�p`V|��f�m��7j����%������ׇ���O8"����v����	��W�U2���V^��osnO3�p��M z�1_A���
�P�	ś�ޛ�Č=�?ud�e�UݿM^@�K&R"w�w��2��i����o3�3\�]�נ�qq^���A;�� V.9g>a��i e�r�9�h�+e�"	x���ލ�m�f�%��$��D��qE��Ьg���Y�E�n��ʹfّ�HM<�l�L}Ǵ�I�Kȭ��0Q����]g^����3���H��s�N��i��
ei�[����%O{����m23T�Lj��}\�gч˩��A��z⼽[�/y	MA��a�����pmu!����􌥽~`��&%�<df;!���q�K���H�f�Y�0d�
j];
m�J�K>�8�����pw����N}x+��qvN���h��a�!��8�JA�����wpԦ�vJ���jR�����b�K��j�TE��M_m�����J2�o�S�{}�e?q�f�)^���宺�X����!з��yXE�9.y8�u�&�9n��2�3ƀ S�Uyc�iR��V������S��K�6�0��2��9X��!y�Y��KP�Xg���9�n�������:��-� U9�V�A�|�f{τ�EC���O���f�O� �V��TN1�{�N�x�-  V����x���n��T�_,K��~�+�Z�ȦҨ�n����ɮw�Ξ����Ol?k�*��A�l������u;��)������*l+�I�Il�#	pGS�H�?�:�s����G|�fo�Hcd1��y����o%.�E0��<+O�⠎�� ����=�D��${���˕�ǩ�#TĬ��� ;}p�� �^���R䔀�u�oHr�X/�$�o��tt�q���R�ڣ/�~n@�~�y�m��{%vZ6lo'Z�tg���8�~l�D�SNx|ڃ��b��Qj�Z�@��N�`}s2+π9�x�r��ɮa�FX@���,VLD���-���%8�k��Dfx��L�ڴ���.Oj�Q�WK6�����j����o�s���O�Դ�����>��<l���X$y��A�Z݇9=���@�a�8r�G&��j��{W����-���J�m��n9?p/��� x�)FL�ܼ#A�O�_��2K����訢[��V+��6jԂ=`�xΰ"$_��#��G��I��cR��Y妴�6 ���-Pq��s�˛��^=�!�w\yHq����~zIb�ܡ�4a�W<��R���3�s����}��k�f��"BA�O�=D�qTUE�9���H%����S�^.J�[/�3CYd6�Z�~�L�@��V^U�
P&MU�m��V:ܤ�b�(Zk�-���Ɖ�{�G�ݎ�h�ݏ<z���c����E�Z X�GH�_/��ha?��������!^(�k[n³�ҝ����2x�+)P<?m��QR�Tn��*���5���9�;���^�5)��������32��{�?�X�Q1��OՑ�.g*:#�Y���6�8�5i7�P��,���"�����!6���!������},��󰨹גN�
p�>�,��rq>�?�����O�Y�ݗ�y4�������TSq��W��v��&h�w�D�a�?�����7�SW�j�_n�{�z������<��]�J쮮)���(i��"�o�L�=5(N~��r�4�t�'7��Ɉ.U�*�o�;��M,oxB;4���{,K���Ϝ�v�X�{9�Kc�����}�x������IH�Z�(;Qo�&2�|�
m6�r�rp���ٗ\�.�o�\�&����������0���������-<����xۍ�|ME-,�ԛ�F9��@v��h�6.v,����*-�L�Qbo��_���3t��ureۂST�1�Þ�uCh�gP���0\��-�hڌ~����x��;��UܣEG�S$��\��q#���ΰ	Qʹ�ZYB��M8e[���d�)������q�5}����lZH�]�}�iCK}^��\�*��6��'Rsh\f*V�:�8b���!R�'l����q
U	+^^Q'՘�9�{�b��+S2�����(K�!t�nX����$�T3ghm~�������l��C�OR���70�	��OM@��źq�t���F��M�����u����.��U�(�y{ݸ��kP̘s�wW�%_p�Ϯ$�`n_#K�(#��lT�4���Z�&P䥃�sy�L-5��y��@�ۅ�A-��  _B^�%�h��j7����BNB����	MP�y���  ��#Z�Ջ�jժ/�pʙ��jCǨ��+�'�8�ɧ����@�)l�
�.��~��YIp�PXw�J�͢��v0X�@�ɛ6��W��pT���:-BG� H���d�����E��q�U܀. ǀ�ɬk�Z�d��Ĉ��pI:��~J �Y��~�+��;y[����}M�do��\�;l��:���9)�d)8c��-`jۏFvU{�RAJ�4HW�!�hW�N�����@�m-R�(�i)f]<5���ѹ���a��=�l���D�+��Aw4WƗeUH�ia�@X ��ޠk4'ris/�خ�h`|��lA�*��%�۰�M��&����ӫ�M�+�{eBđa��Wp�3��%
%)r��ګ0$۠�l>�G��|v�B�ި�uk�{I�f�f80mR4��\H�~��M�2�rV���sK�x)����1k�'�b�˛��iU�|+)���NH�~,�G����3R3뱺p��B(Hl�;��iʊ７���P��NHr�%�u�! }w��քy�I�I/Ũ���
">�:��g��L�gŧ3P!�^K���i����0�̭��F�\un��*�	m�eE>���#T���JP~}���=��}D@��K����.����B�#m�}�����6��o���"��'�������_��I�\0���8¬���ގ�}���>+ǆE�E�wOt�*x$l;NNz����7Њ�	[{��tr�)�nі�4�95��ӳ7�m��*�zN���@U�����������#��o��;=^��YsS#{ɭg�ݸu� ��p��xG�y��4/c��C�M[��hCR�|�P��0����SĈh���q�����K��w��g/"m>ZJ��<��q�o^m�k�JLٱB�=����s�v2�,Mc�й��Q���9�3�/dҙ���g�E��, @�$YI*��07�qIy�3��Q�bđ��:�'Gd��dJ9	8�r��4F�sL��J�`���2̠	���j`��bi��P/�*K�V����9�n�����ڭ$��F��e*�_oF�7CWHFo`���[]�(o�#=�A����\XuP�<gL�X(�;ي��v�4(&�xG�߮�d��[�:�Q��l��c���T����g�n�3� |9\/KW���q��ȗ�L�ۜ���[k��(���$
1Q��*a=e�X\:ì2�lb]�p�k��w�L��I�u����������[Z��lq�_ٯ%a�	�NA, ��_�(��s	��⮑��F�F_R�ɝ��¿Ȧ#"	�q�"rk>�h<Bu�Z�ݾӫU��[��SFȻG��t�ܴ�����jB�>�Nԗ ��S*�+O0�1�@#꠮��t����IY5.�w�Y�侳N��;��1�1+�@�N�ӌ��X��n]�Wµ���c�Ik!
�րD@d N5����.Uѧ�r7Rj�
�m+Mt�'��>; c)�.=M?����!�r��A]O��L�*���稤%P�-{f$�,fg�7~;>fϚA��Z�3[�[yO1�p?����\���2�U*_#�P.r���S�i"��~� $��d.��o�D�����!!�3�}Ӷ���*����Okj@(�A�IJE�n==��*��wfy���)/��(t��U�~?�щ+�_�[�6˄Oʧ�>��S�����ۉ����A��m��� ����!�dZ�q��C� ���uM0��]�׃t}�*t�����~����k�GxY�IW�)O
���$� �vI�/��4r�3�b���e�N�H�J`e�ef��w�~Fnd���&i�2R;iz��>�j�g���"��=f����$��k�3<�x����Њ7�@���A�F+yQ���z�~T��;#q��V,0n���P'�����h/�R�/#++�v�I�>�1��U�3�K�f��)|���vj`Z') B�[����=���b�'�QC���.VEx�pC%T�pb���5ܑ���B˱ |A�IoWz����5�!�V3W�(�b\I %
�=�Qe��^Q
�����Z��&pU� ��2I��&�җ|=[��}9Nt-�O}V�M&���q''"���.N�G�	��Љr����˓Od�p�٢�3�y����i��쟬WE�H@�ꖱ�My5X��J���D��S���i�&_�;pP`��/�HV/�wJ2Q�/A<�H��	jRl��#s1�C&^@Yd�]T�S������7��;]?��&�����T��L�j��.u:?�ue��{yyU���l�׶fx��ck�ƾF��'	o���_B������2��ȭ;2�����~�,y�T���d_�nrsХ��A�p���{v���v����j�3t�����r`��+ɛO�SL}��!`9Jrf�|�%���5:^���'�L�{\���Ztek+'6 K8�`Z�P�T �s"=�G���e�3������C.��{7: ��>�O���8R)��8��z����T"&Q��tN��>y��H�T"9>�����0'啭Ӳ�����ߒ�QT�K�&QI���G��ˁpZ�6+R/B�r��v
��O�hLQx�'&��AيxS�h��l��e�6�����	���=��R�Q�~�i�̦��Ζ"���R�SY�Myx�,�˕���J���L�����E~�b�$0����$g�V��)G�"k���"�6�y�l�Q�3���'Q*��|ʣ�RXb�JbE����^[Ȳ�4�_���Nvr���d��Z���R��	�_��-_�b�N��x�3�k����6����3H^*f���N�[&����_!�$\'1��'X��:�wT�Ȝ�������q�#�`>+��=�H�Y�,Z)����.��'�l������A�]�u��1����L����ywH0jx�>�9��Ry�1]1x��<@u5d=�;㱬�9^8���R�����D�b*R�<|45�ڠ{2��xa�yw��sV��~f�H��tU}9�MbsnL�s�|S�&�b@�H�9k�e�9�ΥJ-������A�&��?����=��݆��M��y�֮�Q`�a��.)ag��� a�YѕL�y�:(<�ƌ�-�{ʞ	�遝�20�]�rρ5@x��E���ǫ�.��WY��9��RK�B�u,���\�¼K����L2K��S�� "/�ޯ�
*Nђ�;��2]�x��qb9^a���𡅄[N�٬��n�Q��i�*�P�Ysʉi	�_��|�G"�q!�������lr��k cٕm꺨��<�H�C������V���]�o�=[|\V��5T"��R�.zk���	ݓ����O�gI��.|r�h6=������xuc�'�Ͱta"�OMO��b +��ō��|D�?�yBڎ8r��%���7ԢC�	���$��\�cQP©��M2d"R ZRƵr�.�l�0��?W���O���i��"���B�nG�Cz�{J����c&����I�x	�j��I�pW;�6�@��gH����>^L�~Bk�J�[\k7�Ye�i32I4��X{7�N9��A�Tg����P��8�
�%���Q?#�84f<�$ޛ�6��T�� ��^�;]W 曍�:����m-�T��^_��sw\!e���@7��G{ X����
f>�������k�J��2�p���$.9S�T�fQ
���.>b.8��A��ɕf��p�Ex�����mq:���?s=�X�Z��Z����Ȼ+~:�L�"ƍ��'c|{fO5��]�pz%��\�V`�Jԕs[�y�v>��ߥP�z�/!)��C�L�/�nܦT{I�@nұ�f�H?�#\����H
	�y��L�B��ӜQ����heQ�e����-��N����i������;p}�am@�˅K�7��8������'7��;������3�:cq��9���!��zE�h����FI��5����`� J�/�U�������t�_���BIN3J�L�8ꪜ[S�P���>�����~~�O�7Q����3�Ч�y��Be�������G����p�i[�� ұ�F�w�Ӑ��<pSv�Tk�^�js�K��<�'ƑNH���?��3�ԅ
`��<�=_���RU��J����Ġ� nb����iO��JF�|>��p�M��&�nnW=�˺�Lڄ�ױo![���ò�L���WQZ���fv�B/z��o�m!��aw����`m�23���~\9~5�hszH�AH�tx�Ŗ?3s�L�h�YD�2���-N��2\����ڟw����"6(��y��4|�}�>��,�?Y��w-�%x�"X����d�K�]�۝���;`X���pm�P#�\�l!K8,����+�o������k�&����$�j�vn�:�ʖ�m��t����1lwȼ#Öa��מ���P�JLg�q\O��,C��(�8mwc�C3�
ȡ��|�]��ݎ��į1�!�c"lu2j�2fR�4U������(���j�Ts����<T�N��&�$���^��m�ǟ�1�f�\V��ۿ�|���z��Q���#R��y��a�Гo_�����O��r
o!�;A��ua�M���513� G��-�~�zE�A�uR�S�˕M�A4�i����)\���l��]���8�tZP��,��=B$/iF�׸��&
�@iv)[�2�cA�����"iHZ��a.߀��e4��oB�+��M�����,5�-���K��i"a���ѡ#�D�ڬ\��cQ=��Z�
B
�Z�U�dn�(���J1���^�i�Mn���b8x�u=1fyʔ2�l��E�@��{sv2�4b݈1����%�c	nУ6ֻ(�q/z���{ 0u���(���\�����.�aB���� x�L)��U]��r
����=WQ��HsN��!͹T�L�]�.��6��^E�'��	���Q�_֤LB��#�1��/E�?��Sl;2�	÷�r�$��dbDh˒�֕ⓝ6�!��Df���YV�Z�ώ�ʼ;]F��t����934��f�<��]H<#�Q�R�4�T|sz�ZŒ����;�rGqO�M�{����I���}KL�T�1�#c�Yt�.�,��@m�xF���/���*0�m72mo�ŞX�/ �+�ٔ�.8���G2[��}c�ne> n� ��rS���)<J��^�@��&|���lQ�)$������R�d~0R��9M��z����]�R��,֍3�H0���� �ʹϮV r�>�0y�>|�5Ub+���a��w4ǘn~�M�9K��������^��_�����x�#]�	--�=��r�]\X���ɠ�oM���0m~%У��j������&ާ+� �:�׵��@]���O��E
ޞ��3ixjI��	�� ���3.����f��$����t꾩�D�<ۣ�2���gSX��
�A�,�6���Ŧ��R�A6≵�\���$�&������ ď ��Lo@G��qǙI�/#�v����42�����=
�]N;��-��M��ِ���B��J/	@���{�ҦZ�~�m���߼'>ς̫c���Ĕ�u�Б�����m?���������ę�ߣ�~V��տ���޽\�o�rh�`��-��8��B��֚S�~;@֠���d���2ͤ��UI����˳�W�AS�y/��{N�e���������r�ݾY}F��������#�tWE_����"g�fi�F�b��TϷS�:9*���PO71�����0���e�)/����P.WTo��pP/wt�#ÑpԸ�����%��v���O��N�9�Z��n$�F���c(r9�s���x�/WR�pv��[����p����WGF�d(�������;��(�4$���
Y�˱�n��V��x���'��ys�F������ڛO��.�@"ʩ�_7\z�	�n-�������nBċ���/��	i��)�C�M[�Q���܄��l�\�ٙ�瑒�!���T��F���QR@hH6x�K
����k�FyG��K=3�l��L�|�NsTz8�ky�a�~�kʡ
�X���b�/uf���_>o�_hȭ0���H@�|��.�P݃˚-FW�t����c��A]l�^���(��zl�y2�����Ī��<5pN?i�8H{Z���}���D1��}M��lʷ�D����+�'ǹ>AM���n�'/�z��O;�z6@&����X�Ev+w$m4(���X�a	�*�jB��# ����ВL}����g�h9\c5<��
���nO�v�[2�]�ܧ�"�ɧe���E�\g�1ŚTc���W��؞O�Ӝ���ܛ?���d��:r�&+��l��a��ػ<v�_EmjH =�����>���B�D��s������"�a_~JO�������-~�@]؀��V���������R��V&�t"]�T�Bꏚ�~f2e����IB(sy��:�w��tC�Ӗ�B�#�@J� ��L����"S@�7(6!���i��v4|"!P��Fr��p�⛹��c����!�K������.&�y��(u8|��MC�w�,�[�2 �:e��Z�I�q8�?�r���7cn��l��ه-i�մ92��ص�����
4_fg��O�����" �M� \��M��뷦�c���۳��2zHim�{�?�--��d�����4s�sK)UpU,<Sz�s鬔g��=�\ўo�l�\�8���X�/J�oq�Z ���"L��ϫ������C��Clp�)1w{%�`�C1�FWv#���MTV<��ZHD�>�5j-�/�uL��o˳����g��(a2��Q�T���Yʴ���d�NW�b���F����u ǧ���0��������R�ږ��LQ��-��}Z;X)���^�?�2,�srea�ln�T�ⱁp}��c�X$����uL��Ե����;K~����{$��bI2�`��/�(B�G�<�ƫ�Fj�h��Zw�G/p��S6w�o{��R=�_�u�Q���qd<��#�ϽB�|�-D��e��+�²i�O��3�-$�(
���:�����4�+�X��bq�T���F)�_}���נi;Ԡ��Fz �����3n�.��Ӈ�ŀ��g��:Z	���)����&&Y�W�}=@?5��*g[�a�iq���4��B�v���_[�]�O�:�ދ%VO��d㿙DS�劲lY-�z@F��6a��Nk"R�@~,���E��8��,>89���3Y�g�ȏ�}31����=��Z�}���m)�(���sβ�%�%�U+�L%�2;�e �L�*���N��ұ@b�ߜ�6������DpW���Qu��ǔ��z��I�ĲZڰ��2J
>�2- �l2R�t�+�砭�G���R�F*)d��SKx���[j�5h���
z�5��!�j��<�G��	�錰+i�Y���)�L<7o+�`����{�������:��Py}[�-�|��t+��Ou/��"2�m�bS��:�:}x/��N��|�{8����O���on-_2��Rs�g�h3�y}
n��?»f"��~92V�_"�o����`��Z����Y�U�X��0��&�kIU2Y�����@����h{R��_�����\z�I�FCL=( �,�euK���ا�p$k�oc,DnP!c�b�dkP �)y���4�F׫r����ޤ���m'���(݃`�y��A*j��_d9��Nꦮ�[�[���Ͻ��|��
�z�o^g�������W����+W�2wʌ{%
���1�z"\�!t��@h�����z�W�Bn+�4�s[�)Z��$��GR2r?�$�� �ɺ�`��ߠ	� r��=N^���)�
H��	��6��y.�L�����a��@����k�2(��&�%M"��6��k�C���A[����
���ܯ��C&$#\�=�6� ��^A+I����3�i<9h����6t�����R�85�А׏ٕ�i�땺��s�KY��%q�_�V:��&u�+>Z�*l"�i�m\�]ڿ߲��tI�sA)/�z�PsJdA.���$(BACY�_�S]�-W<�<m�~]:El��PW�Y��"������ڲ9߇zԑ.�����6�l ��@Z���H����z`�FMX���<ګ�]voT�'�5Hm�֊<�~�ZJ��]k�>�X"_9��� ���r��/S����3Jv�f*n��	���	/�yW6.�z�m��,r�#�Y��1�|�n�2~�!~�2�
cE�(�x�b��G&U)�[��g̋?����lg��"3�|�r�l���92���ۯ�1D��}jR�i�� ��;��	�$����=�u���������	N�_�����<7ƞtN��z6ر�G�5	y�\�@��]����Ge�M�/M�`��ƨ���v�PCa�,���ayy:�n��0�Ý��-5s|�k?c��c���u"�ី�Mu�?e	����� ,�ܶ��̍P^e°�} ҤmRqN�oRٶ���WL�Ǽ^<����Ծ�xL�'	(<�j�����1��8��+�y�5��y�x *�q�f����E�;g۲���TCj��I��ք��y�͵������u#C��2#=���Uz�]�7�W)���e@_���(7´#�G6�C6_9z�qw����ʟ��t8�#���{���U����*�ڢ�x[<]������&<HZ|Pq���@�>��!��w�jR*r�>�$�C�3@�C�.D^|��1�*�����.M�y �	ۦ�$���+���wp<߱X����eO�oT$��A�82���|�ר��i;�ܙ��z�2��4��6��
z�{��h�1e)ad��V����ϯO��5���V6 �F�˜�q�v�&�L\���*����
 :�OJ�D�8��lh����(g��˕�E3�O��R�	0�^���Zyʟ�
N^�\ G*b��|07��t�݉�?ӭ/��q)f�8&�=��r�g��:}jx�3���T� ́�|�Y<����� ���5|����d��j�k[�џAy��~҉k�&`���� zF���I������T^��i�I�E�SF�>�����K���_�Mi%�c�����`�T�s_�|Q!(�wy �t�ת4i�aM\��m�F����E�u���wZ�",;��Bb�U���_	�U9�M�S][�{������%Vv����h4I��~{[����D H�'d��@�z�:���EηT���J��v\����J��z��MW]:�8[1��KƬ����!�$gD���M��l��2֑�>P�ä/�A�� �[2E�����2�x�����	h�����Qm��IB �fpa�V�JK�kkG��~hb�Zmdcs��r4w�|�&�I}���H�l���F�g0�ѻo\���x�\�s��2��߅}.�����Eф�ꒀ�q�]��{7l���z�i�\S:�k�%6!���m��5������]�)5�
����5�j�P�����;�z��\F8����p�MJS8]{%C �Y0���tBͿ��?���+����o|�<�yhE��uT���c������kq�b4鐮���e�ַU\�c�c��˪��:�� �κ$��Ŝ�gY�'=A��I���^:�-7H%#`�8_7���Tl�P��>����h���w4^��č�ٝ�-KGɹ�q�MȾ9I�����ʘp)���._�M�1�jn2�6�tBJ�x"��@	%B!J��aY�����p?f0zL؇E�u�Q��;G�"��8�?����g�	;S��K���˻�XJI��9G%�����X�v�^Y�l!D<��mL�cTm޸�|y����j���bI^[��g�M�C����m����&J�#�����AM2ڻ���J�?	%�����vh柡t|�	HM]|7�K�JS�3bft��7J|D���l���m���_.P�*[���7s.�:b��̉r`A�f̲�T}$�۶+�l��l���ҫ���}j"z�Fc���A��N=1=������JX�����r�At�r�w���؝�&� 9;�"^���1�'��[�7�x�0}M0���V���!�N1V���=Oci�̚dC(V(nJlc���3W���-�#�e�����H��ۑ��2�h�pw}�d2�U��D�H��H�Z��ui`!�.[l����'�\Y��f�n�^���bͶqNZ���_5ĝ���2��ڐ��h�,"���|53����t��Jo�0�!K LIϒ�كe�#�k���`�����r^�ԏ�&H�H��Ļڒ�G��)2��Ӭ������#�t�y%��8�S�9w�۬U���v���/�RS�Ų���.�e<H^R�wT7�4����_�����BAO��Q��b��"��@���Fܨ����&1�������^�N]�d�iE�ַ���MeI�J�(��u��P�����7 ��u⦼A��^��S[y�+W������I?iKi.Px6��V,��V���.�oQC�`�J�y�H"ע������ZV4�s�)�Jh���r�()����-���;ʁq��Q��Nɟ�<�SA]�ޓ8���"��~�~�'��&Ͷ��Q�j¨��x��Y2�M)$�B�5���������H5]ZH�qQϲ��ֺVFR�[��S�t�A�k}�:&Q��@�{!�Z��P���x��7)1E��:��l8�K��
r�IFG�-�]�78W�P��1|�hd8�T ��򄒽D���x|y�j���&��}N^���H��p��䴷��S�D���]�[�ȅ��6��mMY�>f׆�o3+����M��60B{Z�њ�'X��v��R�&���2�h����w��I��i�=|��0>.�Xc��7r�wTq!�
����.8l�EjH�ѷk};�%zA�Z�rS�i�'&�N��m����P�ꃌ�έ�^Pܼɒ<�l������j8h�hy����ʯ�xC��Q��mO�W������<�� Y� ��,��
dRj�˖�`_/��c�$��ՂY���tG�S>1N��</�9�����1���y�i���G�f���G��_W��H���Y>����\����5Y�A��5�t��!�ʙ�\}�_<�חa»�M;�	d�Z���hC/^��N�)筚�f*�lI��B��{z"�^�Xsr��F`-LY����y�nbW�,�P��f:G��g�{�b����(��G�>��Wш�-S�Ġ�K����!��I�$��X��v4ṿ�="�t���Zx�,eȊ��];ka�,�1Ɣ����a9v�w�}�	y�̉�������!2j˫܉�9�����^Q�?�k�D�~�2���FŰh�.�y�����i9������?3�A`�^����������_,X��+:���������/��s��KG��dvg��%E-bGu3�'�ь�ifv�W�H2�0P���R[����[M<ӈ��#D��l��~._kFx��D��9�D�x�HD�q:��(��5p�_͏��p�+u]�{F�����68Ef�!+��_�(����ɿY5hR��c�!���o���v���`�8yY����t��2��#r���[]��k}rə�E��"���4{��!D=e�D�tc~�;��+����t�x����2c��Se'�Bw����o�/dX� Z�����Ġ,���~P+������>�fY�m��gWZ�fHn��Mz�ٮ��<O���[p�[�`�! K�q���� �W��$�����ӗ�jޣ�
�Q��z��6ǈ�)V���I���'��v�P�Y���s,WdvR�����:�O�0�i���f��L��f�$���ϧ���Lኆ�`��v'0PeӀ�Ǽ@(�ڎb�E!g��J�o�?|V������ީ�Ĺ��
��J<*��Ïb�Q!��e��
�*�WI��0,x�x�Щ����I�571�Ѕ����z�O�"���H�� N7p�^�=>F��-"���	v��~>���1nt�N�	A)��ޮ��������z�QD!O�����@W�K�qp�P����`ZUbvמG����Ɲ�����uzl[2�3�C�{I�}�'v Vb��֎y���
�lj�:Yk!�4�8���]����j�P���"�Mp�n����ҡ,���,����X��!�$�G�ޙKzR�������Jk@@��=o��3���?I���E㸝IvB�m�׋c��r����Z	DϚЂ�R�K�f�Ϣ|"�!��Mإ��XO:Yn�ܣ��ѷD����5^N,�~���^e��Z��5bX����5���MƝ�`-$b��	��q9�YbC�@ *��A��wl0�|�D�,U�T��[���fa!`m������|Nv�v�wNi<�ؘ�!�wd��H<�i��$�k6�[-�J�ks��H��u�M:�x�ঐ���<խ�0S5n>U���2X�-���������Y����� S����!&��^�;ԃ����l+?&�N��jR��0�j*��<xMx�!��?�;�����������;ل�ŏ�����Ι=�P�.,��1��Oj^�` O��欴�W�(��|E�X���X=��3ȝ\�����N� �T-�#�_� Y&�iP�HP��A~~3�z�avz�T�j�D�~��m�O!AA�uڻkTO3a_�A�WF(�h�$=��bv����)
o���TV�e���L7Ts�g�L��8���<�|@
D8ԁ6m�.l����#�1ބ�M�.�R�@�1��)h,C�p!�`V�?�qN�W���8��mrZ�u�� ���dH�}�5��Hf���dr���u-Ա�޳z4(˦�][���s$��F�e�Y|;ܲb����buƀy��)&�1l����N]1�W��D��C{"�_��!�/2�,��˨Ӱs���?w�?z�t�C�.�='�iY*K��ԛ����rU0����%7�l���w���}Vze��n{����l�*����E��ۇ�N1W�K��cv�r��>�f��� e"���x������$�Kk dK	��V���A�4����]Nă��G-$�������i�x�c��0R�Q�w��XT�͉����8��]k��)�l�8Ҫ�(0�����&�`Tb����S�{'�#S���WZ�v�K�d���X��:�lm�����-�������@ćܥ�M�������蚆
oE�)�A��.�Kl��PKt~���\���(���)��ܺh@,UP�J����*�Q���?w�c];��O��J��.��,�G�l�)ِ>�WT�3ԍ��8o��؛��kٔ����E��U��q 6������I�Kk+���ܞ�'�q��Qz�jd�O[ۤ:&z+q��8RX0L��������e�ć��ۏm��0�����<M�q,�E �aA]���Ǆ��L����Tx�uH����b]�b����B�[�8 :�\y0���"BϿ�p������y�9�t]G���K�#z�����2é`�h�u-r}��g��p�
�3Hܶ�0���%{&
�P�`���Z�)(-|+�̅�&��kc۠�;�����w#���y�����y���v�`V�WC܂-�b96E���z�60$]�/3W�]�C��l��^-�NB�?����C��i�B#V\��k�3(Ő�u�l�ԭ�B�
��x�
"�@�UA����[q��VE�>���u&�t�|imD�TUs�Sڻ����s~:A���B0���b�U��40=h��,>��pdLx��� ���2aNV�uM}9/>`���Z2�T"�h+d\7�޻&���mc��F?�	JAܖ���z����h\3���/0b�9��Z͘<^홈5 ~9�Ls3`V�x03Ka��U$]�޻���0�gAQ*赲���y4QR�L��@&pCC�&���%�����Z^��~w�A��S��A�@���N�M�����k�XnG�+=lF�&=2ƊO�7��=��Yz���ό��L世�葖B,L�?[��JD��<Q���0Hf�$.e�C�����
,�CT_��h�~a���6G�d��|w̢�J1d�!���)1��$y쫱�o�_Z��6-c*��KUg@t� �_���CT�}N2�(�8�Tw�N�}$�搩�ĕg�h�9�����	Ѹr�HQ�"�륏00��K��vI��`���:�ܗ��}/?��w��K�%p-�Z�N �N��8H5Y���Hq֭���p蕜~��wG��x�+�'��!%y�Q~|C������\k��a_�����H7��^޷�{p@��P-��f�R���m�C�ċ��r�m����2*��'�����bC���ɥe��7]���~���mvɭ��C�H���\!䓗���:"��(G���ӟ�"�)pk�r�Z1v���+��n�m�x��A�wE�FLV�V��y@.6Pl�霑}�m�����tm�;N����jcg�}��me���~~>�c�=E.�y����]i7i;�I@A�M_9����Yl��'���j� �H��=��[`L^�fF��/�^Y��y)
���	��k��>�#���b|㯣���(H�ސ��S����0�K�C�z7�.!d/�Zh�y��Ŷ*H
>j~�V����p�I��+�h�ʈ���'¥گ��M5p7�b��j������!\Wh��o���ѵ?���4�1{�'�9��H�9�+�:��|x�tT�X��^�Id��=��]�+8��Vv�-�h�Oץ��|,o��n��^T�0y�"���/�f���Qջ}���U�&{�A�Q�0Z�q������C�%M�~�W��5ǘ�|�Y������x./�}+r��!�O<��v�F��Hc�:��0-z/�_ʹN�G�AI4�_��܁V�n��W|q{�x�L��e�b�[yx'��$���!�Π��y��`��F<���1��'�5��ѭ^r�������Q&�j/�4��5�P"��>B��&��a�Ծ�"N�0䰋�����ɨ8��Ɖ&e㖚}Ff���Ν	��� �J�(�ϯ����!d�#V�3<r���0��?�>�q������/���b�7q�ک�fK���&�ִ��;�z�̠���!䙿g܋���O>��f���w�au�W/Rc�#&߱+�6:�v3�uն�$+��	A�3���v����ՀxFEeȞ͘�Ʊڄ׎,K;~(,u��#�M"*n�L�0hW�������1>	`�M���#x��~�^w\���O��<r�-��
��Yg�?|ƀn���v����]��B�䆺��C@��p^������W�c�Rh�Mxj�9���[�����ڮ����<�Z}q�8;�5	�V�@%����Jk4A�q:�����Y�r�e	4}�2�R��D����N�%�ReNEI]���6�w��0:�Ȱ?����v_�\��·1����[�Ʀ����3��Y����d��n�`�UA�v��J�]�U����I  ���~��RYט���[d�3H�\���6.P���8��#�7��0�����Ajv6���(+���q���/����B��a-������1"��ׯ@{��O��^"d%��� s�#uM�r+��Xpm�%h�����\�'��� ,Y���rl���U�z�(�Yd+�b�ԭV��2�(m1�$���as(.���=��m8����k'0�����ՠ�j��34c��� 2��f ,u0��oq&�n]�
��R�J`?��0=׽ǘ��Ϸ�9�X�G�m�0�Ug�`��9՚�w�l��'�tj���+S��ɇľ"e�%�hAE3-���`SW��<T:�p�u�����~k]���y�PkJ��+P�Z�B��.��Tā���l�r��{��f �����E���Lf�b����'z��no��qCA@���|a�o�̱��Y���t�&C׵��@T�O=P��h�ش6K�����mh�ے���$c3+��S眹4��`zs��+��2�������DI�Ϟv���QX"N��Bˑ)����Cf���=Z�m�Ң^_�ڏ�@_�pb��u�1'H���Ү1�N7K�l��w�2�hW@�)e���\0�0��3�o��0�j���_�`�8̓-/4�����jF7�xvqA�M�5I���s��Ȥs�\�s�GY�O�B������:~����Z��!΃L�5�'���E�i��[go��VE��!�	�Ob����%�^�QTf����+��^p��s��g��1w��{���q76�nt��:Yߧ �:��Gcȧ~�,5*��p�Ht��_��Ǜ�$ P�/�F
�\z�2�#2�K�
$�G��Mh�k���m`n�Sv�o=w*���tv��ȵ�9�̿a���(�᪖�Z�M<�A��W��ֶ�pk�ÙjK�H�Õ,����\`�z�KV��A~��,6w�M�RS�A'���w�)j�Y}�Y�Ί�܉�I�  =]�Z�z�G�.V[y�.���t�M��l#'��wXI.W�e�����q}��N�p�Z�~ϲ�����8XD��0�]E����ӱTw�G�7�	D2�7���sg����~[mue����������qpnX���V:� �[���͋GVm���UH�}��*d�~��<�dc:ȫ+�E�3�g��5�����zΔ�Ava���#$M.�e���k�w�[H��_�D�3
R�^��D�h��4G���~zI��Z����+��[%�'��F|��Y4ܻ;�`��r��T�u֪�s5�vom:N=� �X����䫓�C�#���7ʜ	���� �&�U~��TD�ݣ�����>��K7p��FQT�@����;�q�xH?�|Eo�i<�����N�^��=��a/j}���^�;w|�nM΃)��dRSN���IﴙO�n��E�����X�ik�y�$3�x�:|����T����V"��,�;�/��Yn��ת ���&��%��,�h�V�'֧�s-�:oЋVN�F݀��t����b�k��f�����li1)�5t�K!]Y"��E��[�J�kh��KY��]���-ϐ��x��E��`?I��W���x�)�8���4M���l��MhSLI��"�=����ɠ�I����P8�x������ȴ�)4�0�����z��>���1����e*��;������Pc�>���>��]G�8щ��{LV�m��R3��^1Z���1֪��c�ҩ�"��:�O�TS�Fu	����>�x'��-T��~�}jF~<z�*Y��IpJ.h�0	��uV��٫��x�OIj|#����	��#߸���r'�L1�����Ļε�_�v{O&F�si�DH�	�u�&��}k�TM�`(h�K/A�K<�bQ�x`�o7B�,]*ǉ��� L��7Ǳ��@J��轤��������<l˖����q�K�oǏ[kaI����et0���o�S��j�L�f�1U��;-�f����*� �:��o�Irǣ(�Zl�<��gbԇ��?d!���B�{��6S�9��z��ᅔ�Լ��2�}�0x��!���"�KN9]���`y@OG�@K��� ���׳���Y��,p r��� ����jJ��l59K�\�D�bqsݨV�w�ˆȟ���,Y�����|ǝb�%#�$V��I*]ٍ�� ������q�F��	��0�q��
JTcqb��|��Ԭ>����C��S����\ӜkN�9��S�g1�v��!�|��鼫�4��pv
^Һ��PSN��"?T��ոi�ʍl��rңL�����MrHA
���"����Ԩu\��>>y����(B��g}\�!��z��@��V��شx�a'�T���$��c��3e�Y��\��eT@#h�-:�Ρ�^HƈP���n'��?��$��2��xqI�P׮^̝�H��{I���Q-5�tQ�t�RMrی�o"; 5��|�[�.����%ЧA���	R��\O�(fk�mL�r&jշ� j+�6'J� ��3"�1P*�y��;ͥ�3���l����7�805�` ,E�3��A�-؉ �����JYy�&7y5��v6EQ�5�7�ܷ:@���I�~���ǖ���S��0U	,АP�K����l�`��-s�S�]pA~�[Ā�9��$(;�]�b�	��@%=��J�/:*
W�\-'tN��4�܇�OEr+i���$$8��	��8}�Ԑ�Z�i�c�O�pO��ٷ����&M�N\G�'G<��[��ӪX�l?���9f�\�?P�G��_8�����5fe��s��!d(�v���ܤ(0��qJ5C���븴I:�-��<��D9:�g��-�Vz�ό�;[(�_+\�YV�Q��Q`�v���CTW�Eg**����p��u��ΰ�
�q���X)�gz�"�+	��v�jLM��!��֙�]O^N[L�H�¬�n�4�-��f�Xg�M���o/����S7��kn�j�I+GL�@�?�M��֙��K@qT����Au��m%S�&3h������q��q�lA�د�(*�k<J�+�0^�6JW�BU�높V�P4�5���)�j��v�'��[.��rd`C�F��#�qE�wg�f�k� ���x�6�<�" ������9<��>�C\��j�M�\P�V��ȝ�oz!��N��5�=��uL��Ρ�IG�Xk;)�᝵�V�����dT6+�p�=�u'$��!I�~aE��P���_��v�L��)�c��~�����R1�U�C��?g8I���K��ν[�x:������fKi���B�on����7���Ɩ������U�� �Il�
_���������g��yl�����uZ-:{ҩ+� D�-<��$��!E"��qG���0����uȥ�y���l�8���A(*�6XEܻ�9��AV����;��^�Ի��� ڜPJN�qU븽�F��ܮ@��:b҇����YIUT���P�}����'�z"�ݠ;�(>{f\$s��\�h���U�l��]�\�z�ۇ�����Bt���!,.���e�-�/
x_��bXĤ�@�&8E;�"�W$���9������ڒ�J��FHo�sS�V����_y�@����2�߮6����.�yS�%�Tw�<���5��#�.&:m*��ʨ0�#���#�Tg�n���ܣ�+2�u�E��o�3)?����M=Z֧�G~��Q�_A/����G����!��<E�L;��=e�X��kӲ^l��`��V�/��%��t!_�,����z�,b:8
�1��-
�޳���|%y����4����FD^����aM>Q8��!�mȉ�$9��椛'JKZ)IԅyO�S��O������L[P��Ђ���ܫaK�o��7v��K�����b-��i��樘����[]=����A����d�YwڏsULa%��טb�㸔^q,i!�=�����DpE7	���E��ɋ��/��bJ�υ��k��0�
��?�v{�:�ɮ����{"�[ J<�nJ�2V�����|����?�`ʏL-����q��U�5�CU=.�9hE��Hw*T�3g��.%ò?'�&�=���V��m�Y�9��u����(c����Ea
c毢(.Us���������sT͇��6/DF�ڏ���t��:����J�hE6ʍK��N߼�+fo�Aٕ1R��r�D��|S6l�$�:6-�Uć؈���E�$&G��U���=���(#yވS���˨��ɧ��DY���"9� 0Up��'N������XS��jC�������[�gR�O�6>�krw�~�'R f�D-}�1��B>��V7�ө����;�7UYu��/`�㟣Ĉ�A	�?�K{���G��}�m�ˬH��c*�!�;�Z��`��n|��!�x	���w�P�n6����JO��(�M����O�<�]�Y����6l�o�!�>��\��t���01@�LTΝv��-afNi� 
q�h�V�p��\�T&�K0�(���Jp�ؔ[��K73�^p�r���vѮp�+�^_l�&p�hc0RV-���yRz��Tl"����܁�8>��R%�z���VGt���R���`��xi�́a44���q�rr:������j���O�0��O4����͞f�����J�q�Whزx@���I��y��`�Ot9ٕJ���Z�i���g�����ˍ옱������"oٛ�j�S3��q��]��VD�!�%D����P�d�:��R��0)tg��������3y!SjK#zw�����Լ� �$Q���+K��& I�I�0q�ѼK�a�Aܾ��X���.�0#X���i��g���սb\L���ʕ���Zw*�WS�V���wW<s((��2 �\�m9a_�p�D����%�N^HBywM�S"D��byX�ph9<���3���-�.F���=�������7=���k�X���L~�uB2b+��F?������?t2dՇ�(&��PxmL G-dN�yo��]�a��1���D�kI��h��C0`5���:Ǉ׵���Q����_�$	�$q�~5N���t��j��C��0 /v?����j	��
0���1z0�U��J�B ��<��J�P�U�M��CJt����I�m/����k5zAQ��M��$�?D�ܤ.�Q�N�0c�4�Ѫ�c�E��+�;Vqj#!�+�]a$���R�F��Z��4�R�����{������\�����"`B?��'O叽|�_�����8�M*wO�/��Q�J��d�W}'aԳ?c~'��LM ���a{8� 5'���(�~�y��.���&�[�3!��T�d5��C�1�a�q����85����B���v6��6�%�c���5x��K�ÿ�N��Џ�ai���' �3ˊc��Y���b��M����A��"2K�B�X�}/�R�LG�����.������9���N�y�i��B��`M~
+:�e��/0N�6\������d/r�7IY�8ԁ	OF��R��� ��,�Y(��G���B��&C�\�k��f�Ũlc#;P��L]��S�8�H���-cP��. Hy �3d�<Z37
˚Z 3��m���J}��+	���q�D{���i�;�L��Ԏ��b��ƿ	8�]�sS^i�V�TG'9ZM��S!f��U�]�����%֏�
C�[Rrq?�$�r:�C�,�c�� ��q�op/�3 �^S������6��?��(4���4���d����LX�AP�b���4c��G�*�u�5K;˫���.XDk6?&�bA\�$
H3[2�;���xF��+.����6��KZ���0ή����q�	�µQh�`�0�4p���x �|)�cG	��ZR����ZY��pn���ٝϰt�96��{-Q��ꂫ�l�a����G��^z�b�5j����e���I8Yۙ��|��'%��Qxض��K�Ǒ�l�c�s.���x��m�3�L}
��ϼ��503q(�1�P�ƹ����d�0�2-{��e����L }�<����ێ.ޒ��� �y�b"�`B���ọA=�0�#p*����NAI$���=�<,�q��t#�d �1��yAip�׵P{�n���#)�j~��Dޒ:G('Q��|S|7sC�:�}j1luUR�0�t(�-�pe=��G���V1J�bB}��\,���meN	m9E��I�UEbCs���h���`�s��n��%2�G���O#�V�XĐ� ��ݕg����}���^[�;1�eI�A?Ւ8��d�X�y�f����U����{|F�qf>/Jj9�Is$�9)��v�5�Zre�Fmo���q:AFs(�7�T�Vy������かR_�Gu��ʳ�J-�p^v׽�(�NC8�āQڕ�,�v���2����T]/�~�e�2�"�E+�%�*ƣ�U��V: [C��n�
쥕��3?};�����-�z�A�R�����A�?ӞM.��u��X��t2Ԥ�)EO �&S�i��V�n��NU���3��>�]���5щ�5Jz�㢒����p@H@�'�Tɷ9��u����~yɶq��Bcy	"yX��*�6f�~,'0�#�G�����HF�����2`sQ����Hm|t��ė�{� ���r>�x-���;{��H��ֲ�eMPa�6Q.���gd3v9�/�d�3�[U�eC$췎q�3��u��*2�O80���C/mdɛ�ᰂϢc��I�t���Qg���X#m�$����_��%M� �V��dۣ�j���R�N�$OĚ��^1_/��OfK�_��X�0>sz08�M�X��W�|h�D�-+%O5"�E��`��]*�T���{�ŕi�=7>�a_���(>z�_��p�@��v���O�9Z�w%����ފ���-J�|��s�a��ƃp~�ȱ�L���`/}hџ�K3��0��_���ޯ?��?�I�eL��{
�ᣬ�X�b�
����r�~�cI��>4Kq��!�*�47O"+aZ��S�2���U)��
�7wv}OT7n�� ��dX:��Y���#�+��^�S��͡�@�eƛl�|��O�c$�z���+	�����ʚUƚ`�A�X�e�&�א�w�����h7(��q�&�=;�Vµ5h��nɭQ��hDq�z@�.S��g�I�,ޝ�'cJ�b_p��t�l)���|�u����N�ȗ����b�g�q�&±<�w��v=�ՠF���t�����З�թI&�ќ!��\GT�_Ĺq>d�Hu������v��rj�q0k�&S���v���1��|6|��P�MJP�_����a1��"��K1:-[ϣ�ꍙ���r	�[ő�/����13�L�Q/W�c�ĳ �彬�(�`�e���4,z���q����[����V푶Ĭ*W>Ø��ukO'���f(Y��Օt�����lm|����TYHҎ��nbٟC�\�����*},v84 �G��4IA����
�$u�`s��Ԟb!ۭ�z�T4��� ��u����l!%�璮�2���-��n����]],��(�|qG�a��N��+}<�ƹ�R= ̑�'�>�����a�5��ЏZ�N��%s]֌=̃؊UHl�[�C��7�?�;:� O�k���+,���K"o�?u��n�����o�H��Mt�{.�aO	E�u�Uk�X>��JMc��!x�@fZF;/RD�<?��˃Yhp�~u���_,� �*�Lx��:�!���u~T�&7�X>߆+;L�WUJg+T�&��t�&~���m� �4R����8I�-^��R���	�q�-�/z���iU�g���L�3�c��3��)�Px^�8�
{��B}�����ԴQ�D����o�k-���#�WrN�hz�a!k����G�^	k��1�לý�)�_':dF*�|�� �9����k*�#7:i����WEʔ�/�+�ͳV��I��oi��2���,��%}�D�2ѐn��J�~y�1F6N�-[��d/��~�j2����ܰʃz���qV�;UB�C�]KQ�C��a/�(U*�"���z�3�;��}v�"�B6!Y�\����l���
�������ߟ�F�����1�F~&ˊ�h5Ф ����B���
t����r���<��k$�(�1xޖ�[[��/�ȣ�*�d�Y�mU����m�w|<��9U����%H��ٱ�Hw
���)X�`y&��̣;�x�.]��I
u��+cI��@C�s�b�oGԤ�१?��C~vC�n1��Ss7�n=Ϥ�B]���/Hć��sr�����b?����P{=�U|k��������y��ǫ9�6 �E�oݷn��k��t�y������d�;�[�?p]J���2;[$7��Y��/���ZǠ�\����d;=���;(��ݦV�k�τ|�ǽd�^^�r��q�M��irM�*�-V���'�+�'�l97-�q�qy�{����&��X ۫�g�
��5�d8P�g&ק*r�n<�0s-":�0���gZ��7�)���� j/2���In��t�'?�QQQW8�/]*t�I�������*���nY�S��q���\��0�7�cP��֚:��O�(h��x��7�S;\0�=o�.��ݜbj��ō퉥YwK&�=�WqP�;h���-�M��Ǉ��tt�R(�8d����BJ��!E��mJo��vK�W�](��-z��NC�k�y#57MU���a����� }:�&s>��}�"&�_�%��	�R�j�گ>�#��V�"3�����Vg����5a���z��+7|�SG&�hc9n!u�A�L|�#���S��q�3��A�Q�{���G�~��:��¢�
�x�j��7�a��阥��R��Co׸��Re�MN�/�<t�H�޶�� >�&W	_�'�%�y282�'��z��E���v�Y������D%b!�t+�_m��D2�YX�yu%���3+��g�u�*���a�4����(`�h��=�1�XK}X��VK��o��]k �ఉ�C(�Zż�_n\-�@,ЩbAn�u1*�IxD�E����T��ӆv1Yb{�=�v��e�~��k�&t����dg-O1A�^o��/��i��/�<�0���t:8���jϝ�e)0�')Z�Ө9M�p�����$(��:^��6vCI]�����%�zċ�C�uG6�CSdN��n�VCj��~���32!.�R�\/��~�d�M�����P;W�Ve�����?LS���^���(�M�Y��Ivq�/��eC�;� ���m���L����6��Rob(����\8���N�ք��,� �I���*�/C�Z:-K�
֦��0"�XM"I� �L�m�+*/�$C[��B�B���2������G0�v� s�v�v���r��EF!a��_�>�X�sb� LB-WθPo��w�!�e��Uk�߭�<�@���!)����a��C[h�T�w�{�q��>{�?��0Y��4�@�[} �Cx���̯��w��O̮J��'�mI��C��gk�m\C�
��Lw�֕�,{�]�B�8��^��DE��lt�W��%�V� ��ͣ���̪��X�э9�Ns<~&�!��,�y�ᷪ'���ѧ�@ O��'��s ��Xd�H,�\{~������O��Q>}���=ִ7<;��7jP���we�ꢤ��~�@ǌ��b���"�6������Ql�!$wGߨ��@�w��x�C#����]5Hz�<88$"���Vd8S 9aY��"�B��b��w�m�U��"�CC�}s"ѻ,>2�9ԑ���)v���U�_'�!���^��dB��+�qfe�;�����c"W�{`dp�&�$��8��3�t�|.���:h�@�)`D�S�7�o2�m�a7�$b1�1��D�m��3�7���nZ��yLͷ�x,��M_ͯr��Ss��?�6;���R
�Đ���.�PuX���&a~}A ��όY"J9p8n��1Y����NZ��=��7#u������Ho=���@V��]"�r�*ǥ.�s֪Y���~�)���=G:�o�E�&T��w� /~�Dc����-%ib�l*4eU_�|i���eFl*�V�:�(H^F@(TQ�}�W^��P]�x�Ɲ�ԇ:�=�7"��h�IQ��@B8$j?wh|��Y'b_�����,4<��ߖ�W&��/��]	-�i8M�P�j!w�hg^�i��������I�l�Z�m<�K���#آE<�B9�&qa$n����A�hu��zl�����TB���
MKFC�36��#������H, ���#_^-XK���ۮ��oR_�z����P �[c����|�K�a�z�'_�ZW:hғ-�3@X���0�p�r�$s͞��=]a�^w\�S���D�Kȯ�R����
����Tv]�6]�&�\� �]�t��`!f��3N�rC��s��]$͕��]$�na�,�������,=���`�Q�j��u��8���g1���
��Z^1R�I�x������H�$���_ ����'�!�٨�hW���?�����*Ĵ&�ذ;�\�,���\BPn�X?��cd���<4�/HM�F���O��#��k�-e�t�o�Z�3������a,�G���8F�7@�,q_��i�8��{ͱ���Ƃ�ـ��o�K ��J�[���T��R��޽�a�7��x6v���gT��BD(�l�%y�C�9e�uǊ�?���������-��/æ_�#��F7�Ҟl����$qD�2�`�����/�
+�6iE ���x�N�B���S��c%�A���¥�V�=��lGRaU ב�;<����NE��b{��oF�U���N�R��ιY�:r$!TP����3;���8����T۸τ�1G���c�e�,����~2z����� ���-����\~>g����h���N̏9Nj �s�^��u�V�[/�̴��O��̨��_���۳/ZHr;ǘQS�
8�i���z&1�Y�~@�20%��kYudp��*��AcQ��4]ʔ�V�{!�1uӬ:�����>sn��Ie7�� ��f�Σ�F^LJ!� m��Q����/X�'�L �ԫ���I�⧲ؽ�&ܤ=	��Wi��p6ڪ/5 ��f$
Xa�f�f��[��=}�E�S���uܬ^?�W{�梹�E�d���j�J3�G��%�R�[]���l����~V}�r-�L���Z��5�0�Փ#�Zv��QP���@�>XĔ��x�:3<?^�i��0oC�]i0�ƭ<7��t=��0�^��Щ��Yma�t��
��G6��yb��P�[C�G�e�"��ʼL�������#��K\��H���%f�KCm[��L�P �XO�W��$��Xxr��6r^>���0L�m��ͅ�C��`=À>���jα��Ũl�!7����5i����v�Q����=�-��u�.��M��&fՔ>�

�n���m˳��u?fG�_u˽o�����@�d��	�S�m1�q:ҡ���]7�� G�
Pi�<�y��qY�6��p襏 U}=j������ȥ#�԰Wت���5UO�Y��,>!�-�?���ăHf��	Da��Y_F�B��	�1�����t��$��;L}~^�kѰ�ß|��
�H��I��4�g]ʂ��V�8�N$& S�~h򹮭D�Z��@L��=j3Y��a4y2�9��xH����"xÍ�1e�ŭĉ'(l\M EDlL�Jn��5?v�-����v��h��{�Q�W���1cx�Xx`a�l�.]R�.q�B�!DkO��G�~#sFZ�u�h*�|���[� �iQu��Q��\�	��Yρ�-xu��[���^:\�"�6��ڂ2-��4��g����l4U����MgGM�Cb|�����S���z<�g܉M󽋍���E��}x��Wuǿ����)���1q��M��hc�˵~��� aq�������8����eF~Z�UP�Ķ1�^�:��� � A���Ej�i��3���ٷXTq�}S���ZV+[��}!x����Km�4���`�؅�Y�1&��(�i�9:#��.��Uә9��>����i�O!6U���C­�[�r�ӯ����e7�g>��ӑؒ�Q$�C����8ZH�T+$�j~'�� �Qsj4�>����b�3�^���c�x�8�Z�dȾؕZ_Vf�8 s$�F]���P9D�����DC9(D���Z�����m�c�]u�vF~UN���^5��,"��l��9������Z�?Q�y�ٸ�D���s�-Ļrʮ2��r��Śi�j��9�-d�ۗP
0{ξ7��{a�Y�k���҅�ެ=I7�3�<�BO�����qtu�1���O9w��#J\�|lS��E:�!��FC�5��֪޴4._J��,#�Lt��.��F��Mk��R<�������������_4�����x�P��J�����P�z0�H��u˥�ތ�ח����6��>�l7�.��Z�j�����*��5C�$h+�A�+���Q���6n�S����{�̳[���Q�
F� ��`Pi���h)8��8�D����=��3�z�E� 0��ʖ,g ^�ˆw�LS�eW��H�R������w\�Afi!��]k����Ҽ٭Gs,Ґg�	��LO�Ba"��J�����r�j�j�w�GL#k(���e[�0}������~{PQ'���MN���>~V��s`��Rfv�6��K���p9� ƽ^��8��ػ={���iyp���S_�k|@
�@0G�ҍ����W����� ���-6Q�e|��F"�Uڼ���wV���X�_�B�
ڹ���
P��ry%��Z֦e2e��� ٮbA�w~!-DW�b��wG��5ӥ�D�m����2����{��x�����|���6�.��Kф̭���ǚq��/K��Ƚ�B�E5��]�-�I�p��R��1�n)��u"Rz%�(]�!&hx0p#�wNӈ��pF�[ӈ�ƕı��o/�!��(�RLr�)D#aC�m{_m�N��ٻ�ҁx���_r������(p'V/�;d��?���]��~`sd������O�S���nP���y���D�&�1�E_�#�M[���c8|aX�g>�?�U�Q��L|;�eZ���:.K�r��J�U��1m*��Z��<�`X�4���]\p!i�~6b7��?�o1��4���#�ܥ��g�̈���n� �?���ŅP��kLw��v�oB(.!���Z<
J�����0y��� % <a��r�;o��p<8�u�����(G� �hRP��);qZ�3�ͭs�j`C�J��@r�JA����w��� ��d���LM�[R��"��49W���NŦ��������<zOć��.������5T�����TY�?��N�&���x�Kt7��ӥ:��/]��)��8��>�*1nD-����׹�e5K�yG��H����J�LE�z���ۖ&��~�>m�8���K�If���)�����ٍ�N��L��h�7��i�32Gc1��g��+�A{���ձ��e�FÏ�� �	*�1)HMt0E���������+6b۟[��on���Q	�hW��6?��j� ag��jF:�����9������>s7�Ч�nL?��C��̀�14�z��m<ie�=���3���t%��*�h33(R��n=��ߖ��2�7��t~��3�%���.7��=A�DI^u�dM��aF"Z�W��6�oA�x3y?�O/Q�3����Ņ!�b$�uo�w��:��l�5f���7���ƎZ�vH�f#�7�M/P��'5f/ft
�<ΌH��5��=�=�W�n�9���.��l:T6���ڭ0�T�!�&���x'D�>$�;>]a�U�WD%!q8G��wX
iWn���擙˞��䢬s��?�c�Ky�Mu��l7�a���y,�z�z��2��1���H�A`�f'r'���N�Fw} �W���7�O��5�Ĥ�����vQ��i}WǴ�'ޚ�����eX��	D�ݟJ��J�0t��3�J"�hY�a��2��$$���n�N� �1bC���J�a�z�����,ݔ��a�,� Nq0����,�3Ň�����P��a
Į�7SX�bޞ�l#Л��4��IV"���c%�x뚒� Xd��"��8d��P��6|��xca�ֽ�R»� ��Ky�N$z7_N�V��HZ�x[_��z��-��w{*gf��:,��BY>S�˖���V�aB�l-q���\D������:6�˞�2�C�����ۚ�j)H�[�r�N����[Pp��rDu�fQx1�Ҭ�g���|*�K*�O|�.������Az�y�k6Z���.�o��3Bh�ќ����I�]譐�t ��{O����D��n�z����ֻ2��i���LͅdX,�f�V߈�|�p)WPhz`�$*�h�J[0���N��k�Fj��	�)p�EcD@%�tw�T!����N:�\�o\ۮ�d��|�FG >v���;�!p]���w���O�jжâ�"� �,��9�p������$_CW�>�����;S���)5��=*s+�]߿A��<Zvܚ8<@���]�P�j���7%����e���:��i�����q�6&�ǘ�[a�EY�ᾇ��*�&�Z��9�sfR��V���TD���_��o�e������n�\kO^LC&~�JO_T@�(��σ��݂�z$�r���#�����k�}x2P'����ҧ�x�)�$~v2$���Ô�����,Q�^j�6��-���2Z��A>ߝӱ˜;@e�#Z"��L3`,zVF��D�����+�\V�i$8
l�K���˾�o0<����P��c6�W7;I��I)�����?�|Ɣ��3g5�{�i`$g�}W�R�E`,��u�,F�ͮ_�֍ꖡ�c��Yo��Jb�n+��Nnpt2.��rt� K"w�H�
��ݹ��y���f�o���(U����,|P>���.h4F�>��Δ�4��u��O?��FU�`����O-#s�I=��B�m�nHu(~�K7��+�E5=�L)���#��܀�]���j�q*4��B��g�k����#g�B�/{x�o���0~hB��w��'}#��O����]��~�w�A���\���n�7�_��\[���J"a#���v.(=��X���O���L�(뿷4
�O�����_�9>.1���7_Eo���(@�3��-McJ��|����$ ��;c\LfY�o��� I�,�1G�IE·Fl��n����{��jd��D��	>�Q�)m����1."ۏ���z^9-���Eۄ�KҔ7u�D�,C"�H�z����)Ud���^
�L�-���tf��@�W$t�	V�Z�l*�)X�sR���d�2����Fnml�	�W��l��<�8�R��Z�;�/"�V�}�to3c����#UG,�~s�2�c�̚\���Crd&�Ę��I���N�}�ߝd?�y�4� �!]��%�	7�?g#��W4(�2�?���Ka��f�E�^�.(m�۝��|����`�ltK�,�(�����7�N��Ή��|�:�f�pvB~i��'H����+��|4�~��m����;0���� ����Ȫ��T���`�J#��[�J���=w�
�u�>����]��m��@��R�"$4��w&�?�P�`v��.
nn��:�Դ�F�s�]�$K5�'�x���X�	&�f�F+�����ϟ�^ҽZ!�<�l[H#��Y��#$�}J0E��}���6o��w�٨�&-��IX)e7G���������3�Sڃ/!���j�9 �H�76�V��E�w\7i��7Kdf��۷1��8������W�Aޛ�GA��P� nª|:�8���Y*r"��|��C�z4(���,&'��nG�{�]*��X8���nQ�D�T㾼�>B��@T�<�Pdw�ȿ։P'S�E��l@����tFE)=�M�7�^���R�u���7��Nn>&X蓹�}�@̥�H��6#\N�쓴 ���Oُ�g�8�����[v��� ��}����C=m77a�Tܞ5��Z	�Q��&����k�$"����8��0<o�Qxxލ�/��'����[v2	�_n�z��<��Ҏ�1�E9��G�Q9��%� �F�;J�������ͭ�~�%бH/�WC��Nk+᭬��F��%<�5�1�,���-��G�O䴓c;�Ѻ����ȝq�'+
�
�d߰t��.����p�� ��-t�C��@T��rH������j9�*��~K/=�\	f`���'��B
���UHrc�g��b祲:}��td���-�C�����_/J&L+U����P��g�0�0Eo�k{L:N��o>������A�jN}��5{�`�Mt%3�~�$��O>+Gٜd�C�����\Vɝ)�	�b��xZ��IV?����R�L]���#^ɻ%��$�Lz�6���Q���%�fW.�Ʌ@�5��\>1���z,��`���]ǀ��>}5�q:�ߚ�ŗ�e���Ψ�+?�@"�A��u�'w��^Aw��tb?Yށ�.t-�z�ܒ���E�\�u�Z�IG>��'�-����;���г8��Е�J��[�=����$�H�V��gAZ��/��`�z~���v��Hih>e��Ή��zu��������Xmv0-��	Qs��(��v���k�(��%�f�C��'[o"z%i�)�kL����(@���ZS�&��k��F���l�ElT�!��<�-��b<m�����_0�;;K�"���D��l�!<#���d�Չ��*h��_krҴ|	�'ܳ��?�%��S���Tp��Q��䂩�ZlË~��NC"�&?7�j�M^��U�����Z�f��G��d�z\6L����o|g6����&~2=�}QO���X���ߓ�ξ��#��3<[��KP��mn����䆳�}��&���U���u�Ě��e>V]-�h[�爺;2�0�2P���~��r������N�'9<̗Fc��bg�����,-A���HM�5��Ё������|誨x����T�\�#&rt+C�v�����lk�j:����~����4r����9�e���F��3Ҳ��:c��P��`f��+_ja�
�$�f��H�Y	�K�q&��y�.*�+�>��4�Ҩ'���Ł����3�2���a汤	��ɶT�Iٍ8c��S
Y,u�N��N�� !���ָV�WC�"�K��v��>�
�u���H=y�$�z}Dbߍė��v+�;�A�5������L�?9) k�1ʈ&���^�E1���қU�y�8!cJǍ�a7�i�8
�>���G��M��AV��x-u0�l��E��z$'k�ۊu�z�c��&���g$�'�>f��'��A
�g��(�<ܓ�{="o���7ƹQb��b��u4T�c���Y�O�"��>��;�AgN��=���&=���$|����<��%3X�V��v^�͕!��*-��\�I�B6fg���[bR=���(Q�J��b��o@�h�<u�P�r��ϳ�8�&!�g\�i�.��.���j���2��
F"�=���PI�W/]
�a�a/���0�M^���tO�f��۩�o�5��ū���"�@�	�9�X����F/��E����Ϲ� h��Z�	����N�Y�nӨ���D5�����̗Q��>|y@1�ɢ�u���V��<s479��U-��9f�'�E�Qm[h�������w�BA�[-�(
����Ab��FЧy�2g6bV�����wΥ�ߛ�>�rdR��O-���#�i9��]�M)s�Csl@l��&�����_?IR;�tX�X'WI�G�n���˄6�o�nùn��;���%˙��o�'�Î��\�WZǱ|ތ�����^��%2�ƕ�w��G���q=�p謼��������0�(�WA�dE����l(z����Z��$̱��B郑
����;=1�N�)��Y�#�z7��}��;g;����qm�Xc���~$����W2W�bR����D\Et]Uc	���ag�1`[xm�F�E�::d
k?sМE��}�pF7�� ,o�)�����C�ZN������ �x�����t
>� m+4s�\J�l�C*
8󹱑�>��A�1�4L�yBgw0�XiĦ���[�[kr�{�2y粩��R�+yk���a�?Ɵ3/6��q=[GZ�ԁE?!�1~��?���qvtE�q��o ��I�O��3�k�P�~qI�����2pno�9�ߌ�~�`~ 8w���9�d,�N��עN�ǖ��"�b�o��t*������a�G +�V}"��1xV5�D�.��t�#<�}��&(����s����۟V���b�$������[^LI�*+Stm�鼋��_�߄=���Or��m_�����[a�
��$�@D���.H:�*�?�]����A���/�]����&���U;��e���=��N��tet��Eٵ������7�1d�+�'z+�aZ�����K���Bz��8(l<*7{6��10s* ����hh:�ib���VF��_�����Hcy��#��70j���3�B�R[!����;�J�N]G��yC��ٺ#uVz�)^daU�1�C����y�/��5���$�o�}^�^�v�Ȓ��������<�=C|��6˭IK�iw\.q���M�BTFGa�I�ԃ��w�o�U�DM|7]C�q�AX!���U�)�� Gʎ��@��c���|�+a�u=�_��[״m�
�{GEd]�i���b���f���z�&'ڂ�L`�:g@}-�Q��?(�M���-׿~�1>�S��'�b0p*S��!I�C����_�U�Z�'d���GD�`��0��P11�+�)�G�2VZ�D'͛��i�W���j�����Β�?�3�29cS�"�,�0[z�=B{����T:�5j6H>���+d9��nT$Fm��T��=\�~PDPUFn�M��U����/��î���!EO���ӵ�ķ�%��`I<�:�f�˲N�5	�C��v2��\��<a\q�3	HT�BԨ֣� ����5x�&/i�(�+�r T�'H�:!:9n���f�@d�<��G��;�S�3oR�5J���K���bĬzD����R��qzF��7��$�rt|�,�%<�er���<�!��i���u���:�rxa�m�Ӫ춅��\���;�7����J����fwU�uH/��L&| �a!��݃{`�͂��oy
{���Ug�<N7�%�`���[ߏ4G�D￳�����$�T˘֗	�=ٮ@�+��[9ě/`�	a[V��h{ȭD�"$P�����;0a?t�Wj�5޴�"�8�80���lΈ-�Ҕ�wufh5�G�,H�^�ll�`������;�I�ۻ��O��OgY���7�"Q5M�7x�s�)(	�����H��^����g.K�=㻘��q1aZYƳ?��,꬐��2�a�Si�9�z��/��U���~Ȅ*���Qŉlsc���ɶU6�`���0�����c��%�%^��w���5�T]87��)vu@�:3�B��[,��+�����dė�I_G[�Ӷ~A���:'~��V���%p�����T+�	`�s;��I(e�b[�a�d�y�
�N��\��Se��"RM�@��s:Ed'a�� ��� I�G� ��mr t�q�<�`���DM3,�P�ȼFX��ߤϘ��^�?��d�Df.������֢!�)���������t���_��ǭmz��΂�崟�j��6���� |��Nj�X�|E%��<1��*�
zP�c#�c����Utt��VLI���Q��_�^�'-ݾd���H�� 2>�$��]�*���.�טH2,n���{!?��
 �.`�����a���н��^� ��X��'�y/R�)w۟�ir3:�N3j0�"Gs��UA�غh
D��¹��03Z�=��=R��bc^�H��fh� �Xr�VP��/������q����f��uڎ��r�2V)DHIAv,٤�EBMe=�0�n����H���:�N$�~���SÇ�i^�#��"�1~B 7ݿ����1ShD�C� ��p�����6"^�����D��@9������#y?u�T�Z�6+�M��������mB�8�X4����i����/�-�Y乽�a�IL?�&�V I7��4i��� Ӥ� %�ڈL(�1{� �h_,�G5�h�y�ԊV�rH7�m�]��<�U�r�م$��{/���4��~�eI�����Nq#�0��O��u0�B�*d4��:e�\��*f���~��'�r��Q�t�tͅ��p���KO��ԥ��C,��5���O,90�Tn3נ��e)^�M{�_'g�w�a�AUaUK߄�D�F/`U�Q�,���b}�g���܋{y��b'�����n�z^��^�L:�9�_lޤ��{���)���������Ѯ�f`-�6��ݕ=}_�zk:�q�9ﴊ�e2����Ή4U9k��+�0Vڄp����5����?AjQ�amz�2����,|��p�cf�Ft1=Rڃ}%`Ѧ�r<aT�EK��ʂ�;�X�f(������T�n,�u+��$�Z/�~)h�Xr��g黧�]�7�G&�t�[¨��'�G��5�x6��!h�/Y�q��簰� �1�����r���9���S��wh	xL[ ��֎�V_p	��RnQ�����Ғ���3_e��	��Yw�GN5
F߯\�3�j�8/��ݰ�=�]�Aͺ�B�X��\��I*x�[�ѹ෼LZ��ʆ��3zX��{�Ql�4��%̬V`�����đ>�zʆ��m�y�W�ei6Ot;
�G���ٓ�(`�R
t�bO��}�q��!�^�Qq}���(g4�D����i�U��jq�s�A��0��G��DE3}��Jr�嘞\��#�)Y#m�Vؗ(�ݔ�������#���0U��'���r7eG�Y3��1�"Lp���Z����*욋��]*�k<z����,��z̸��x.)JǦ�Jam��7D�	�b=u#�b�����^�˃��J��x�U���W�3��4<����s3V�͆N�O&	��,��sJ�*_>)���`6K�6��A�ً,vX�n@��	�����(��ԃz�8|��"g�"8���ϖ/D\m��Ǽ�/�̆LO�q
�o�˔l#�����y�F���z� �>�=�<�5���Qn���<%M�+����������*j��� ��ay�ѿDw�z!�q�O�J��� �d���ŷǑ>�Z��S�#�m��D����big�/:�FOz44�r�����O)�4��9�/ �*<W�s�c�H0�}����g�D��:���Ѱ����5�%��� �R%}�����RM�и7���¹H��A���?K�n#�AF/gB�=T��ç��h0{`]H��Ȏ�ӲQ>=��K<����۝�D�o�P,��X�� �r�}����/]
5_�����lF����O�d�sp�az�m\�<�ȭ�Q<۾�e@ґ��e�/U���p��~5Im|���:�;�Sb]Jo�m!�4�>��Q����=��ܪ\���~Qx>�mĈ[�]�����|v������,5�Υ�B��]������~u(�=�fk�y2��љ��$�N�$��.��6�g��zo��\�܋&љN�s��lt�{Z1�E�/"��}�Ǵx�t Vj8����s��1LmЧ�����N�ގ�ō �!
�o�s#��ʏ%l�5ߺ�ߔ`N/�g)�1d'�CN砖l�JW�U[7'>�)��;�GJ]���[��i<��M:cu���42�u�.����;k�;���,mPX-	���3`��X�c7�WZ�G�D��>s�����"0���H�I���x[�$��YW���A��/�\�=���9���M�qJ���vƥ �ߣ�Rn��N�-@�CC�k��zf�O�-�O����U=�ٞ ��5�<`��7�Qz��簕 �"��oаܦ�*���ﶈ��#�xp�ǵ���P��t�1�K�D��X{T�:pE�ʋ�qɒ:vX*e�~[�զgԠ�l��Iy�ߦ�	��o<g��m}�a���5yPr�m
�V�����^�&^� �Zؗ%znK�ƹkv��/q�A��xɰ���W�S|b��Z�u�	.Z��Y�8�vm|�GPhH���M�6��-�c�|�"������r�D٬�}&�&>��)a��]�(�S��<�����{bݔ�F	B��d ���
���Ś�crG+�X1nH�|�4t��k`� V��S����\��cѻ�즶<V��R}[׵W�~a�,�2�5��gҪ1�I��1*Ɲbk	~�ǆ��}FI���;�99��4�v��� �}!���a'�>�J����o�t�_TŰ�H3�1Ql
���[�qs޺)O$��6����S�Y'�Lb��a��v�P-Q0�]���]���+?����8�L"R`G��E��\����&�C�\u0�|a˻~��6��T�;�_@c�@�-m�� �|F�;���Mh����ܹ���r	���t��[��9͉���ᭆ��4]��%-�17�����ꥻ*���٨?��iHad��[O`�ve>Ӛt�$a�A�i>Jy� B�T˫*\��6���.˂W;�R�$XW���y�	�;��\M$���r���R��x���&�廾l�n3�A��~��+G
Έ�$��9kʷ��zؽ��d�����%�ŉB���.Βw�z#K5�4�>r�> ���Й�kԴ���wS/��5�]���Zk�ɉ���N��Ծ	�v�Xs���I�/�I�9	!�A�$N�x�Ix��S��MgJ�mc�h!�s���C�����3	iB2�гI�|�W:��$KD߬Җ0I��t����O�)�Jd�Ky?I��H �o�}�f��U�"��ơ:i�y�74-�TE_7��X[�9|ug�i�G��ó�S3�y/=��x�Vt�!�Hi��X�Y�e��]���WW1�0����hx�3�W���y�ЄhX�~y����V]�uJ�s6��R�#���-�������3R��l�e�(R��P�æ��yʘ9!G*�?���[ �ʕF-���IM/��P����Ө!�^�!)8��;�|���R��V�c�A�F������I�GL�x�r��,w��f��cC)�͈ɛ�_�l�^�x�7^��㵟%[84꒖�q
�M�"�%��4Ԛʏ�u��	.��h<�t0w�e��U��Ft�Q�o�p����
g����N���rr�U�5����k久|�[B;����*���!�=������	���`d�t�*-H(�
�N�OH$���sxZ��H�ǲ�ظj@h�IL�U����y��h���ⓣ&�r�Y1�l�4��\�������$�W(���D�4].9�����W�w݀��0̔l���@�H W�m�����n��l��8�Oj�Z)�I���!��x��,�2�ʾtJA��ϊR;��"�Ϳ�V!��;�^}w�m/�� ����R��q�+}|w�c�c�|Ҵ�7�x�=-,��k�qU,���k!�,�s7�޶�TD��X�?8�Yb���4�T�`@K·u4׍h��Q�ma ����g��'Y�����Y��麟L�]�l�wu�uN�o��ѵ�.�)_��tB�>.]����/��S~Ņ�H����DD��@c�+��s�^�-g�@�d9i��
� ��78�\��/R�O�� ���  `;ꥈV��Q�*���<���vC�������F+S	ܪ�7�H=����co�U[S���i��O�}li���O�K�i\�+���ϟJ3�Yv�]�<�bNG�%=S�\���uj��L���/�Vn��ܑ��W��]Z+~�sR�������6A�>���2�4��<�q���A��.�N����G�ʨ���E��*��w�OJA��y�۳0C�0j�nT�Svn7�p�y�8�}�Ґ��/��Dn3J'�c��y+Ya��q���:{�%d��_���kϦ��kUR"2�Nb��7���˥yff�l>9���1w��XWl�zv
��KD�������S��An*���ą�g��[v�l�NӉ��C�*��ز�)ߒ���} L'+��W�����jw��D ڞA{�l�'�Lg�3z&v=��_
�g�7:�(�>}`�U��x~
���?x�Z(uY���7$>�]����#z6.��fӧ}=�㢴Kxo��,J-\H�vy����l+ơ���d*�W/�m���]<� �"�`L^3V���0zb����]�a�bO�q��܇zY4��]< �?�wN��D<D�Z��K:wS�n o̼")���@��K^+Pq��~��x�E��ԅ_��.��O�`�F���w���M�gI��U[�R	P�f�DL3�K�~�	I���PѼ/��($��e��Ч���ܨD��N�+݀�X��Ў��>k��:�����!�}a*��i�Xn�V%������?%�J/Q�M����( w�XC�٧�3oe�7�6	�&M�E�͕z��b�������6�����]�bn�=���aF���C=��C����i:�
n�A���f�W��n<�W����@,�N@��q�
��y��
T�&[�Lg�ӰD��ԝ2��*�X���x�)�.*
OX��$v,�xE��:�1����ǣ-�M�r�0�ug�[m�i�3mo�v:��'iG�,�J��G�L���;~X���s�l|
y|b�
8'���_H�5�>��	�)D�a��j�}�*׮j��$�^e�Hu��{��ҟO�HvD��_S�ˊ�P���]7��� ��o�l��_#R38��ΙPl�^��ܔ��0�Nz0񊆣㭰B�U�X��w1%���1�Q��J�����I0��>�G���aM���}�S�����]�t�c2�C��:�hzs�[b"�3�D�Ȟ^_�Rx���^cC�iy�s֨f,���H��U���;����[�$u>̈́�\S���+=�����e"̄X��-0������B3���y��<��-%�"� ��HpN��B�6=���N�\b���#t׋OYk���e�w<t���D���j�T%Dg3X �Њ!W�H(����3C�9��� �K�'���<�N�n<�5k���<$dT��?58��Y�����E��@hv �IT�=B�B#��'�iV�k
��na;~���m��d����df:�z��L��8��jR�qS�l1�����a��Gi����[i}�z �xoA�Ֆgj�\XW���5�*.fZ�
(��}}�i/�)���v��;�	?�kal�$�9j-oj��i��+7�]R2�|?d�����ao�0�mpE�����5D �����ɜ08T��L�&e��X���,.K���;��'�T��륍7�|���9ir��Y�3�N
ق�L�EV��T�7xH4Z|d��={z�/�`wlq ��,_^���3��J+T���s.cg���P�iV�����w�0���f���R!,qЏ�d�$�Qw���V�V��B�o��$h�(4�J'�����Y�"XܑG��˒5�V�@o�q~������:n�m�����0SP�a)��`��*�X�rNn[�A�/���TE�³����z�qD�t�s ����VA3��l[<�Id�s�N;���%�N�d��J�[U�M�m�6�>�w��Z\T� �}�{إ�2+�vݴ��>�FԩNy�V�r�1B�!ɩB1~� O�c�^���M o4��4�W^�� ńT�+�W���L�-�9[�,�&���#��<7��B8��\�̟�I�G�3(=��
ASᒫ7B�#i+�/a�|��l@ y�U����7��G�Ǧ�"���{�I����e�$���O������u��:�����N��U�%|���w���f�T��������؃����Ka��P���V<��R_�b|���8(��y���S4Gl�=��� !��̑rD.��P���"����>���qn���26ر����d�Q�#pq�wM�f.e=���:�m����xXm�=-���J+vD@ע�e<�{��R��_#�L���>�,C��I�-�$C��Ǜ���B#����_I�Z��oC_���)k�?�f�'�c$)���#"S�+���H���%�X,U䟶�	���Y��:i��J|yB�`�D�%���I��.C�Ș�"���+5'@ٸ���"�	�6ň)���*��b1��hImW0���u�_�C�)R�.�ÑA`��^[b�JN�8����Wc��ۭx3>(��]]�<K��`%޻?���]\����b�#a����;��M��bJT{�4<'F u��s���B�k۪χ�q�a�q1��@[����K#��: 3����9�9��rmsZN�i�R�,���S/���̔F5��Vo�m2���[Q�_O��wC��J0P�+'q`���5�/@���**���Np� rC�j��/r�ME�K:�GRfU�)#������_��A8��s����ꕋs.�����Q&��5D�z�)��>���%���&�z��v�L��(�\ǆ����h�99"![k��a7_9؟1��A;1�y ������b(����3����m��u�{����l k7;�9��A���7�+ '&������DIŏ�d��ӥ:�r|��@_G�����q)�\�������V�I:�$٩*�V0��ʔ�!�x"��q�|K��sԕ9d��z0U��/�kk�?S�"��8M^	iZ�*f��/`g�೯"�Ar-�g�ͩ�ANϏ�6׼(�ܥ~����kU���2C
.�&�{�F�'�����MW
�f7��X@�Onn״�ׄ��Z��o�t`��֒ �����@M���]�#�+`�[��*s�E��0��JN�49�A�>z'y���qG��Bޕ�aid }��{˚r���.K�|m(=E��*�E ��V@�aAO�R (���]-!�1�ڱ�>��.��J�CK�5�߽0)ty���2��-���Z����Ǧ���vxְ�T��n �RPeiS\�}���d�n��Q�Ye������G�ću{N,L��p�vFZ~Y�]V��ur�[��wU��U��U��rmH�S��52�������<@�!���_��p���'����Wa����=���h=z��V��8/�����a�خFh�I�+n�P��l���*.J�ɞ���'{̚|F�~�@m���|�Ĭ��V�:-.�Ѡ��#�.S����eNM��D+:����H�Z�����t�}v|��]L�i3���F�����[�a٤έ*u�{��o��P4�Cl$ �O/<���g`f?��I�ǎ����.D�e���Y���1��G�\8��&ط��Q��=p�K�-������Y&Q��s�ٚF�,&�
%oS˫&�_�"��w(��i�?�㖉�$À���g�]�������I��~ʍ�LYG�тU+��z&vM�.��d�|;qǵ��UJ��q
8��0Z�!tB����I*kv�S��Z�;�j�[ӐB�B�����Rӂ[S�	�ﰍYh���6���R�w�sCk4�^%��)�9�{ib�Ԏ�P�\�	��j.��2p^���vv�����\v�Vl�R���(��*S��k�<p��3��B��m��ZF�����/���r��^@�||�Z�D��Vnυ֌9����Y���>I)`A0�'-6��FZ6v�c�Yq7����S����Ȝ��wW�lʰ'~ܫ�.<��f�cIhwYA9�v��ClBі!�[����Q8���Pe��ʳ=�%P�n��*�K��ʙܞN��Xb�E��=�8-�MdW���}�83I�u�v]��*n|���Q��R��Yg80�y;���0i�}.#����J|̤5�h�t���7-Y�	ֱî���OU?��VU�T�%����(a�зz9�*��V݅�>w���sZ�N�<ٸ���<����dTޚ��>�gԡ5��xzq$�|�&�9C��[n|��_оp�h%�e���9�����^j��q�s�ø�k��М����j9 wS7���U���(HS�fJ���!Ȋ��Х��&�$�,a���F|��Wy�7��Ic'�ſY��Q-�M���D]�tiҀ�,�q���뤃X�B�'{�m�݁�������9�d�����Ny�Lq-�[����U����9�ƶ�X'���k4(���}�y/��c�T_Us�*�p�r��nFD�a���ٱ�_B�q�T/�}� �1:^���	ΑP7�l�#�Ñ6�'��؁L3Q4��]����E�B�Kl��E�$��X{h�~�WVOk���qn���OB�quh��T����ӌM62�@���2��z������ֆj�U�(΅Y���|�8��o^u�bW)�&��_���p|>,C!�/�;&h[z?�%A�ܾ'q�[�_�%i-�|A~�oT��-I���_8�PS�k���I��3���Yj[���1y �u(-��Ż|���XXz��_v�iJȔ���q8�,��w�̎ه|D|������Q�6A�������ԤL\��M�K0Nj�>��|�ɺ���;�!�ZQ�Ey[uؠG�2�����61�*~��r �;#�ܭA�-�oh'b�ƅ|�<��@?��s�̦I���ed���ă*�?J��qI��=���vY��b�1�}5��T�_�W��\�\0�^���`	&�T5�������%��!�s�'B*�+;�#!%�U��ǃR�YMR5��+�K���sTw���#T�!z���!�B�n��ns̜Z��֮1�`�Q��-�س���G��F�~���4n�77Qd�й��t���mK��]Hp��Ʌ��a0T1� uP�|���o|��^��F�� ��t4�%
�F_�:��a�)���g1e̒HMyrxA�1��f����;p����pK`����$�*���&0��N����12��#`�J��c,�۰IL��փ�s�h�|$��y�Ck΍
�Ǒ�, �UE�}:�B|̊��2u�U�89��n�^��n��-ǃ%{�S�;S)���H��R��}����1�xWu�0 fV�|R-}>�|����xA�"�~�H ����n^��D`��2��ꩼ�v�?�m!l�M�X��5}1��n��?�-�}p/�������A�1;��LY;���D6��K6��O9�j<.qH�%��[��:�j���~�k�̈�9�Fg���H�R�ri�'�(H��<�X-G�:Jy"�f�-�9֤��$�H�-�;<�`s����Z�s1�#I+�½w��C���^;FJ��_���p�5m�S�̌`fb��b�C�$#��T����n�ܗ����1 �qw&��+�Q�m�w�u;w\��i���R˒�QZ<����H�CKԭU>득<&�\��Cm�_�d��H_]S��5���nR'C���.3ο�O��Һ���%���Q1��ڊ$Ѿ����� ᶼk"�8׏���ey`a��ƛ ��*�$����Gr?��-f3z]#�尜gZ�π��(9�0}t�����w$o����Pi�a�ͼ�ΨJ��[��Ʒ�ȹ�%q6a��ș�S�@&.�ñ�V�,��g�#@����_e��ñ���kg�X�	�o�*k�
ػfZ2�{��	�nB���@J�|ѫ�p���ݒ�;�2��w*�g��0�Ts�-S�ح�KyUsyۚB��P8������7 �Zj�{�Fr�*_��mh�#�Aۏ#�e�.sĔ�ii͵�¥�7��1�����n�yD�ɪ�DG�S�������{�^�(��t�a���w5r&@�Zӝ���a��/RP��U�(��
tj�=[��&A)���0�c��Z�x�!ީJ�۴��%_Jb��2� ܝ�-V���?���*g��F#EM�m��s�6�>�w.�g5����*�
�,�o�3tF��+]��~e�=�>�� ���lt��{以���'���`�(�CŐ'�t������t>����aR2Q�����<6���#�ZE� ����[8�ƅ��:�(���l����[���ݾ�TV�Lz��*񪭖Loa�H�$�#}����c���X��:�|l�{Wt���E?2&�
�Nfi�/��>�ӝ#6:w�b	#�1�q��(��'���w�)�-U���7|�q<�����'\=s9N���E�Db�XƧ�e�G�E���Yk\׏4�v�h�-�̓�O1�L����2i���a0Z���A�}U(���v�(C�K�ǈ<Y��'�>�l��?]�6��a���J*���N��>}�XV�����z�٫6�N�-͡nC4V0�˲����l�!�8�S:|�S�`V����v֖�n�p�Ryk���~�<e�C�u��Ԩʕ�|���C7��nY�����0@�H!�k����>�l9���Pb���Hp_m x�M���WI�_=q�O)ut��G�+���3)׎s���͐�ۊ��U�2�}+��stIЍ��D<�c�^C�l�t��+��QNG������X%�J.����M).�p��۱<Ll�ߌ�~�$ ��+pQ���\4s�����2���U}����%���Eb�+���N��K�B}�\��XN�=��C4�3��rSL�(Nh>VW���� �BJ5V\�[���؋�%p�r�v�\���x���?��N�`	������~���Yo��/�q;
��
�aǟ�:��F��� l�������V<TP�/�oi����?��ߪ����4��A����fj |��Q�Mg�\��*M2����?���$i@2�����pt����벧�.� `�c�ץOI��篰��׼�'H�x
9X��x��R�n�έ��E\��̾/�fdJ/̝_I����c����_1>џr���31n12�a�GT`���A���%}��2Y�{�m�d��ɼp��?������[|I�n/3���$�(փTPpUo6	k�A���yM��>�����P��4��T�R�����x(�5*N����*>���!)���#x��!0ȨH�50$�~ӗ1໯�u�u��ޘ�#�dl�Z��b���E�_����
���HҒ���|��� �d���2���Ka>'k�.��� i?;�gv�/h39V��Kҳ���Di����~-Y���浺,���Y�6�@�.D"����� �g\��w���D���=�J��L@ U�ߏ3�O�8�ҹ� ����Y'\�m\Su��H迺��M�Ӕ�'�+�1W� �,���I݅����WO?������TGn̢wg�onG�f�
�&�T���p)�E�#\5ڊ������G~�u�/Қȳ8������Zl��)�.�;I�¨���=�H��l�gv �w�� ��tFՠ�0[.ٔQHzo;K����{l���<w֕'*�\ �lSy ������7f��#I��b��Ƈ�� #pZ�����B`R�C~�;5`��Uc�x�V?nx�߶��v�mπ-�{����P��of�@|M<x4�:	�ӗ(U�,����������K{�Xs>9<�A>�㳩e��w��/x�_A��+���]N��hF'=6��,�!�J�P����S(x RB�Ыv�d۠���K��;y߶E�\�0㫓V%��Æ��#*ej�I��`�t�o���}��*c���������C8���Q���A��Q8�����������sd$�"h��a��{pu��Y�j�hF3��8�*�
����nOZLP�X�u�,㽥�=�#j�1ݫ̀�d�����h�~q�����w��p����1��'�M\��(���ɶk4�b1����g���3��쏑�8��\Dk�P����E?z��*��R`�d��Z,Q�WmV9k�>���+e9~)�u}�g. �/�-�����s�_�$hT�;h̦���Zb�����sc�Ͽ�BNo�m�ы5��G�=���d�[��&����K��^"�6��?���@�1���i &?�����8��^ɍ��}y@u�ѝ��u�K�h���IU�*svg6��Mԫ���&*=U��B��
ᗸ�F7Fq���M�W���G������t�II\�d����Ǖ�B���$.���
{=�z�H+O�1tu��,|]����s����hu��g� wF�u@�,t|��*��Գ�����
k�'TG!>�/�i��Rnv����سd_�i*�v,Y����@ٲ_a��{Z�`���T��o�¨�8�Mr�lNI/�"N�(��/��������jE�]��k���$R�;��T!��n����bTY�&u�%�rX
"^�P�M��J<
2��I�\p�� �;��]K#����f\@����^�T�9��ۙjh"v�F�t!)�:+�l�>����cD~�1�EuR����=��O;�L�����L���GK���=0+�J���ǒ\~�(��A�mP�`>����:��6љ�?i�Q�]�8f(_Qi�ѧE��nEI�)P=4�c�u�߸t+��0��@b�(�Æ��nIa��v�-�~.U�b��}
^�6-��[&l�8�������
��J�7���Ae�^�W�՜�;�����)5'��Q|�&���+��LygW�Hi6�1V%��o����g�?�2�i_����'8��	'��y@t�������0����Xļ 1�U�cL��u�R[�$�m��P����&S�t�%�%�l������w�w���*���X��z��3�u��^����>��\�����8�c�ڦ���F��1�	4����U��-h��'��J#b\�^����Ԓ:�뱌�s�{��~m���f�Q�Jag�l�p8$�c�-ks�KӞDek~u5&�����fg��
�0��U�ow�`�&�!��@��~�����R�H�6Q������(BH���g�u��gz�q���J���;->�׍J��I[D���*�|p=3�ڸE�7ߣ&�f0|:y,����WׅE�7�V�6�~�m���`gO�.�c_{�6��U��;��O�蕘r�=b��G�1�;3.��7�k�@��"���?��q������q����HW�7%m�o�H��h���9���NJ��T*]L���(G�Bj�FX���N�)z�/nly/���쇆�N�{�s�2�=T��t&Oq�2^)G�7�H��D���0ϡ:�8�(VU�[�=�ȹ��#�)$�ח�|���Ga�]dئ�.q�<�|kQɹ}�[�����o����t�q�$ q��MJ��3cG��@�q�{[�P駅����Owk�ջ)�m蘇�siۜ��ˊ\j�K�����=�����lE` �!C�jƽ�#(�b�+`@뚬�,I�a;;������B�ш�sb�a.F�6�����A]6�:��7��=��\��Y{�a2d �v�#�s��ߋ�!�R�N��ru�����oe���e���pBѳ�Y��D��ȸ^��TYɛ��fegJ�Z���B�@�h��;�gQs�׸Kf%��~�DG+ڰ���W )��D3���c�C��g���-�����W(�����U�!�kaU�0����w��} J��4�F�Q
"L�d�CŶ��������!Ҵ`��
��9���/�aX�[j�Cj���K����F[)�A�9������Ż ^+2�B@�ةE����=������N�+?��6�R��]�ۮ����|�Eۇ��wn%�o���A�5��@+d�Ԭ�ib*�B�y���YE��"s�/"�ة��L@Y��>:��Q���@�Ֆ��u���xt1*��j+�����%/3��ݸ�#��L�,vS�xV6��D�]��z�f�&�;��"ɓ}��6���Q�s�^ę�=�u�a�v֜U`�`3ֱTq�?�"%��Sc�|�׉q:]�dć��ϡ�V^XP��8tʬ%��P�'yH�"���q){�&��k�b���|�C�,�y"�GoSaq�-o�|~o��?��@9�e
T�G�͕��e�d�K	�c��n��te8.k�ܩ�5�/����;�#d���"cm�zT�\�n�������e��@t8R8�����������\�֢%��Nl�k��v�A�?r�S�
���.��iU��1mf��ax�D�B��)w�6��spsW5B��NW3�Bo	�Қ�u�Rc�cN?��ds��YV�4U70GN�b}�����M���� �K�[s}uSE�X�}p{];�����4��#��e��L��4m&�lV��|�p9��5T�_�y	f{��nA�U�g|!�)6�-4���[��<�v��URtKH�tkR���<�J��/n�5���a7�O�<�4��i�W.s������,�M��SeV8Xu��*��{--;�������r���]�#o4J�m�x��b��|��S/ %�m�)�r�ڙ4�,!�>��_�kH�ڽ6d���$<�d��׭i8�fZ��?8f��<��D��E��͉�E��K�^�ґ0�_��(#�0�
��6�FEZ	��w��v�xCs������p���I�̪��Ӓ]Z�1�嘌LNc	�v��������� �ZoHr��40I��k����v*NB+��)l:�����A�S*�c����

j�﵆ �53�MS�9�;j�m#��;���˫�� 8~X��Zۋ�b^f���tƌ�ˣ�^�Jp���1��}���Pk�Ţ����\��d�ݳ=A�3��z���YW4'�;@I3�Y1���!���eW��ն�D� �;���٭���I�b%H��ϻ�C�����!yuھ�B��%w�~6��o�t�7�5� ��w��X��g;����%+Qg��<��!r�I�aJc�:z}�G�w�Jp3����*�����R��+)d�o\ou�
�+��B�6�-�t�4v���ᄑo?$G�C���1��cmcr{� �=r(<ԼhMb�eeU5 �=�>5���?�z)����ܜW���k�.�ND�	�`�W���C��4���65m�E/��x�+��'���9\�Ĵ�Q���a��
}
��v�����}�Oc����cɖ��t����hO~�n�X�?\~�R�CL�&�N���1j��:D���3<M�[p����t*s����!-!!%F+�r3�{rrK+� L�W�brn�kQ��oaU�
r\��q��.u������y�L~}���3��x��&���e��@��n���0ZC\�{��zτ�f��J����;��L}&�O���mZ�_��s)aq�YN�}7&�G��v��C~Jt#G������zs?=Sa�����(���_-����
_��n>d��R5:ښe����� �Ъ��S�)w
s�A����IE>V0��JG�[��ڡ�Js����Հ��M��s3X₺��HM��f*�{d�v4qG��1n�?��;�L��c��+�
}����'�}��F�Kf4�}~-�� Ui��%�~��J#bw��N>ͱd�)�Y`�?~�i�<an=a�"o�Cs��
X�	�t�y��^<l�3�/��_B+S�/�n,�O��<�qT�r���"IY^J�BZ7�uʈ;�+`G�	%��[�=4��A�@��R��m�1J������ ꪢ �{�����e �@����ڸ���2�{>;��<|�ɴ��i���6'�#��ۍ�� ��W�נs�yG$����&�\������V) BN�{.��V���2�ܩʫ�
Js����)�5b�sͿp�ɲT+��F�����o��cͧ��X�P~	h�M�/��YK�s���(1�ĝ���-H�P^�H�gv�Gӫ5u�|v��HT(��dĞ=Y�A?d�c����|��W-���5�_Jo�
��;p�R�+�:�/c�m��/D����V����VJH�p��$ ��o��y��!�?�{u��n�W��:����(�Pi�0��l) B������QD~�1�8+,qov�C�e�<���\٘��t�+>�m����N�6���<K��ϱc��!�@얀�.#o��8w��­��47s��[Nwo!A(�ݬ��H��%i�Q�>������C!�l��"�H�A�3G/Ӹ.P��Z56>�(����^�`ױ.�M��5��G�K��95�X\�3����mNg�i��ͅ]bs�q7ګ���t���������}�<I�\� ���9�#���'�|.b�E��k���D�0���QRC����VѰ=I��\��r����R��b��p�fƚ�r�{���[�|j2���e��R�/�=P�&'�&ٜA�c� Ԡn�V�~�׮l+u�J&n@�Nc�wF�a2?�E�f`��"�`$�2�b@�(���)��ר�AY�]�}�i)�Ym/�E��Yf>�
B�/~�3W��Dt+�)�Z
�����~-��� �*�u3(���(2CԔ�tC���cs�,�<NyVV�
�m�R6~1݀�b�M�H�Ga�Д���v�*�ͬ��u�xuVz��ʆy�[�;t�~Ǆ�[����\w��J�q��� �Z�크�O��[N��љJ�Z"��]�`LU�JV-ʮ9}�n)Mz���kf�@E�)��8�L["�@jV���j��GeH�y<DU)�$rk�)�����4����\V��?bA��xV/:۹*@��Hk��HCv�����D���j�v-p�T����_&!Ӄbۡ��>/`�%���:�IU|C�T�
t0�k�n�㶪򣨙:�]� �`sD^%a.�� �P+8Sj,M�w(/
V!��H�z�v�w����
�5 ��+g�BWp�et#��b�8p�Ow�����I�E?R��@J���H��mj�(xI�<�<�V��ё6h(��!�&�d�& m7 
���L�4S��&�NT�R;���w��.���?YA2��s@�z��qL�.�5�y!ɵY����;�y���|R"j��j�#�����	�b+J�`�x��1vO��8H��#Q��AK�f켧@^��l�o��x��Hw*��D�h��ŝ�H~8<����]��s��/֡�)�^���i)gxq�xQڤ�w��Y_�~�_�
������>�E	}�d�q�#���.��1|C�g���n�m�ݞ�5��@�t��l�^t�ަ�8��8 ����ߟ'y4�A��O��@˰���kF2�I4�Ր�� ��>�o_�D��ae8W�"�v�f�#٬9������(� �se�\@�Q�$I���]��{�W��g�k2�/���^�:��x��s���9�:�ץ��_W�#&IVh���E�E+:�6#7).���1	�D���# ��'�f�3Ξɗ[� ���S~�B���h��;T�!|3�X^ w�V7���j(r��q/��c�׈o�1u��K?a_r%�=ڬ~~�J�K�|:���4�D�q='��?��2F��$Ƌ����Qꗍ�e��0ђ������F�\�S�;���2�]?�/��=�k�>j��a��1�t��NQ��XZ�0>o����ĐiC�s9wx���Њˌ��Q���qd�����?9
�y=_�/EuE���Z�Ҥ�ԑ����y��n�\2e2�Uq�T�y �&a���U���b�2��]h3���mM^��+��M�4�b�g�GLQx��Q�t#��:UgEҎμ�k�h/k��UvܕV����2�m!e4Z�C3���R[Do8���?��N���� ˽�����Ib���VF��_�\�����e��Ѿ��d����
�(�C ^��5�S��O��뚠{R9)�X�fҮ��SF�X.��$�?��R�y�2`��u���((�u��G�����<�����?�9��\˥�p��~�@�c�4�4��������i<E�1�C���Y��)[��b����a����)UԆ�Β����2�Je�A?z�Q�7����}��@�<�0:	���KD�{Mg.�#�}��X,0�WW��ʉ:Z.����w��d���&�y�b��}�� ��/��۽��(ێ���ܹ�@�_��3�e^�4�+ �j}�r�PR6L�E��T5j=k8�<��ãX�0�*Jbd�+в���o�YG�ʳV7���
��e���Dh�c�#�>8\��r��a	V��D뱻��>߳w>T߷�x���5J|填α���[���NĖ�G�� ��by
r��yD�>�v�6Y�Fd>�gD�H0����&^J쐄�b�Z���r�|yT���b\��:%s�� �$�'ݘ�կ���8����(݁41,�Z����G����K��TZ򩹣$�d\P�xu�8�T���a�> ��+҅r|�DK��a���m�w珞��ԦU�SѽzM�F޸�����@�2*�#r ��$��[�m��W��~��"��bK���H��i;m��#\6#��N�LO�M�j'嫉�e����
���-�9�m����yf�%��[!lP_��/�;�N)�Z���vd�+N��h�賏w�!�%����#�W~��ʀef��v��9YjC���	�*+߸�:)((G����L�ᄢ"�/Q���B�;2��uBbI�����1���V�E/���u �������c�QD�#���P�N�7x��*���R�����֨�(t��9	�w}?Fxy�d�k�X9]yKǳ'����7�PGE�N�*D�RD�9ш`J~�!\��#��#��1�s=����x�����+���\Gy5F���`JN|Z�^�ȹg� �*�h��,��۾�Xo����zS�<%}KB#�%��h�a���<6�و��)�]�>\�-����<아��=g$����G4�W�%L���y��֯?=�{p�>�-8g�6@U�����5��}(B�ȓ
�Q��_�2&���@���F\쿇�	!3�RA��ԕTc�X��ql�"�I����A$s����������G��4Җm�̢R}XJ�ƾ��J���?W�9�Hna�'3�X��б�q�9�dk-��h�e(���J~��C���rI�N��C��\������Yu{���H�7�I����Z�I�Ma�~;��O��w������.2$����b�AtX�K�کLLzw�4�ZڈJ�p�o�V~rD���:��Ж�+�Ѿ�6(� �R~e�u+m�$]'N����uj6BoQ�yj���ꃇa�VP�����)��Qg=�CN
���fte�`�����Q0%��Ȕq�J�^�GӼ�W׋&>Y�U�Q˕�$�Y�;��u�ac��$�Ѫ(��d��F��a���H��W: g�[�������<M�<k6��5��z\\�'Nx8�>��^��a�U�p��Ӷ�x��\�l�2;�9W�����2m��fS�$>+�wb���- �IU��w����i�����Xo~��W*��)fi08gX��"�Y�ߗ�u�d�J���H����3[e����=�.��L�o�[��O�����n��G�����Mc���u�?��p��&Y�iZ��"�|���V.pd?�Z�K?�R��c�ɛ^?��Ra.��rC��<����ЩC)#���5P}ވ(���dZf���gp��h��Cv���g>�Y�U�<x����i����x�)��<ٰ��݃�~\��;�-J7��_
Ga'�(Ռ�I�X��C�i����A\\g���uy'�@ 	��]Ɯ$�5��������|&x��1:�Ch�Ł?N	ϱ��Z�i6hͻ��l�F����f�*+pq������a��[qP���!r?��΅�{��"�VEգx�c�տ_"O�s�z�����g�+E��3�%<�q�����'m�5��+r�x����#���/$�����5h!�e1��h(�^��J��^fBj8��m��	�)��4ܡ�h���_�y^L�'�O�]��m�"5�f�ٓ<~����jd�D�g��)JW���2��A�����&�^�OI5��w��w��h�V�Ü��&CY�j��9g���JK���ɜ�7��ezߍ�D����t o����@'x�H�Et���LZ�����m���Ō���#��� �:�������O��V��x�[�<tu0Y�\q��6���,�g�x�A�F赋�5�J4�%��PQ�������O�ĕjg��_�?��|E��N櫋�F�o�:�S�BF�3��j��Sn0�\����<¤�:MwZ��w������yn?���lZ��>���:fkJu����5]'�3-��(��v݇��H���]�-��@Ʈ�l�h���8H-h�����EPP_c��N���!�<@�~Zꆈ/] ��;��r�A.b�W��@�v�����9&d9�?�ơ��b��8��I�Zj?b��e�R|�H��v��=e�IH8.>�'I*	�y�������vD�8WQ!'t�be6��U�P�+�������s���Q�Hg�So\�D4V�(�X�B� �_�.��w�,�Տ�4���Z �R��y��z�U��=�l��u�R_�r��-�7J��,���E��0����5|��ܗ�ky�V5#�k���3/ݧl��f`����a[���^�&qH`Ә�Dfm��Z��E�*1�"�K��y	���]9���	Ƒ��UW�����0�/�8��H�h-�m	��3�%+�<�Ji����Ga�*�}��7���me���e?C�Y@g��J�� ��M_�)#��/,)1͖r��Us����n��r����]y��9�u� \ґ.�Z"o�Fs�)C���Z����\�Zk��>e�H����u���	:e�v"$d��̘���Qq��qZ����<�kڦ�k�9�N���c���y�H�lKqn�`�Kh3�n�M��7��ǁC+�I�wup.��(V�o{�3�<�
����:�e�4���ЛV�S�.��9
��J���O.��-��k˞���@dؘ�w�78A0���_>��S��1�� ��<A��>�z��w���ҧ�����	G0	�h�NaR�j@Y�����.s��x�C�c{gAB~�����aN_���H02��֏���٧�{t�7}XMWQ��Y�=�����T�d0�ӥ1ȩ�ҧ,Rg�(�fO;E ���U��4}9�75��%�-�F�g�z򥳎8�m��
�8`������	��v�\o���)'�g ��2~��*��?ࣗݍ#rX�0p��ߨ� ���0�R��<��3�P��ǰsH�<xaH��y�z:����a�Ц4�<���|K4+W�*ڴ���bH,ŵ/�Ƿ.> �g�`�dgc���[�6�]����ۃS�:�i�O08�K���D@z]�e4�jFFY��l����[�)H�������۟ic�B��[F9��yYE�3^|���~��[C�GM�*��_m�'�Ԗ��A�r�?1˽ƃR��?TV�Tn|�;�/!yϕ��^#�'�)��nΊ�x��w����lU�����ϑ���c4��L��	�(D*l��I'�HG6C�]6
]󀍾L)%g�06#�#����ѵ�  �qʎd��DX�V0���p:;3>O��}/�`��:��𖻄����AYS=#�R�����X
��x^�?w����pPF�YCdL>"��Zк����R��U�y��\�f�Q�"�5r�ׂ\�� �/���w	�he��Ʋ��B�o����}��&�
����Nd3�A5��e��E*�� )�/ c���i��}��:��-��x`qb6����`�\���ACS�;Kv#��0;��T	>k�����E��-еs}��Q �A�tKulY�^�h�H9�E6]���HTB���o7A�v!��|����^�$zo���q�]:u��.�~hF�"��F3ԁtxF��O������J�p�!���Y��/� ｅ�D�^.��K\v����-\6U퓵��652D"�uv`.��|ޙ� %_uZ�����o;��!��ūe�ҌԖK�z��t�a&��(�`Nlh�4Ac���u9U��q� ��/�ED�9-��}z���g�Ûc.Cި}S'n�W��=��������o��O���e�m(|��_50A�6<���lrr���v��P2��;fA����S��;I%��D�:�!(�|2[@�F\C���1�{ Y&I�ʓcq��ׁ�y��T��p��;e�~@
�K�o��})ӅB�[!<�0Y��ğ�x��:�p� �e�Ro��\2��I2!K!�Uy b��_&_Z"��I�(��#��0�4mҮK.�cy.�Ig<���w�����W{������M�S}aԭc��tLh�h��cp>I ���>1D���d��1��2�}�t�ߞחx<}fV�y#fAp�(8y��LO� ���0�^$��D[�Cf�o�ъ��@�`K �f8���4,%�q	*؎�D�x�${=˭D�k���ҍ�	�zG���������öE���C9r��Rܔ���?69tZuK�̽��B?CXt�c/ۋ1�s;o���po��ނ*E| ~�C��s��D.Z͔�%1�>���mEE��P'ⳬˎAG�U~�5)�\r-ς�Z׿J0���hmTb��a��<J��%̼d{�;8',RW�P��� �V�-3`cR-57�?Vp��oj$CO�1i��r<|��nfղ!�%� O������H�͹Z��Ԇ�o����C#�Ϛ\xb*��*�eVTC����o��x=�晎GQ�k�`�*�,P�Ce�G���n��p.��+�s��mm��̥-�U&�C���*];���હG���?���ܹ	0LE�� ;�5,�C�y�=�����s�9�R�0�Ϭ��,��G���ձY
c��3W�&bF��5cU����<�����J�pA�Sc"O��6�f��蟜朖�8KrYg^��=�����'S�3�%���⑮�2��0gbu0�y�B &E���qˏX�N�-7[R%�WP6�6�}�On�*+[5��3�{�s�o�@F��*3/���K�>��xI�����,i��Q�1d7{p�����Dw���g�Z�����]����رj���
kj�g�2Y��z\_��E����`�m����x<?�|��F��8�ke�����"�9�8Y*��.�-�$�t7�?�r�H����ɕ@�W�Ʒæ�յZy�����SO�_of,��:��iO�����!\�Y{_�l�Ӄ�z�)~���3���K�Ǚ�����&􁤳��6䎝�T����E��g�Av�O��@m�bFЇ!P�>7[%��,]�ǌ��i�[��ݳ	9�'fv#�}\�^u��{q9���_'��������Ϩ��Te3L��N�h��f��{���m���Y�-nކ�XUԉ��a�h��5b�]4�q��Z��Hb��	 
��y����i���}y���|:(�c�O����*
b�BhDk���I�\Jŋd@�L-e�������YM�k�q��Z5�#W
Aڌ���6�oyћ�2����Zl緙��1�#,39@��iA6Cӵ��A�����Ե��9(���5D�o-��0�{��V��2�'���K��8@_y����on���'�ιqx�c��p�1�ڵMrQ�([ 7:���,u�ʎ�p=�M\�'�"Ǉ^Bd�m��F��T>h��m�[O�>"�\�ӼKKc�\3dԝ��H�-S�,�4����g��tK����4X:��V��(��D�>A�d�\��rsݏ2|�]�<7:�O�Eh��p7��>6@\�}�����e��pr~�Ġ�}��E��'=q����Û��~DB�[���Y�^���4�{���Q��u���	r,'[��m��.�Y�1��|=a�RS��CI���_�dX8=I�ݎ��l2�;��w��‿�P-��;�L���'�/�ά0PA*	�T]S`�.A�9�hGٌ�q��j x9#�?���4����#�b�u����Ռ�4��27�5sL�rط[�C
�1���x]`a���$O����G����O�b|��rB��9�Zd3�����9m2��18u��-+�9�΍b�d�d��[{d7\[��1�\��U�8��ӧ�1�>��0� gѸ�K0�O��W������1Љ�b��PV2��%*�Fs���d�݊��~D2��@��η�D��C����J��dr�WlR���9���k��?6ئ�ʀ�����Sρ���F6f�� ��)V��5J�}��o3ݣ��V�$�w`�'?��9 %����p�7$�\�[�U��$KI�0��Fm�����cl��Ѷ����� �V�Wr< ��E �4�b�o�l���:�$�9���yB(9��R�H���RR���p_M*������ �����+Ll�NG7�aQ�#dx��� F}�ۑ��dhh�1,}��z)+O,� ׈z�P-A���S+}�gn��e��|9�K��5z5�Η;��2%X���Lͭ��*D�K�n��ߛ`�Iɔ�H��O��t��\E��M�F~<K�,��0��	�N�]=����^x��z�����GT��X� C�s�1#�����a�i
�\���ڌ�4�ܾ�ȏ�7Kd��N�}`�<����C�?"�"��5�@+Gw��FJ-�7��W���=B2����G�3�+������v[�r����e&�}�Z�����=ٝ�,B�f[�7k���,�d=r��W�l�o�
Oi ������Gϸ��;d�G���<��m4&7A����xg��/�@M�l��G��dp	ՙa֏�Q��C�U�1�B-?��E^�pAI�ɓ���>J{Iq���򍭺����E؆p@(=�(��x�7mlN9��7�RI��*�*P_�>O��QP�M�3A.^��Y(��yb�|���)��?d����%�Ax*VH��e'C���Ϗ�њt|[�K��>,zt��Yъ���a��wDa�����D��w�)�W��b���`!����Uzj�B9���A�,g$�m�;��4O�� ֖0r���R�i)3riC(m����^O9*w��c̍k�UXu	�I=p
�����$�,�����"�x��1��Bt�s�k?��G~�M�VR���{k���U[�'\�<J.O��F��� �2�5�������l�Mv�(���6G0���/�c�㞚t(��$\��MS�St�Eٔ���a ��<@@��wK�䤪�:$[�rs�
�HL�^���b|�]�~2gj6ڟ�%��xlgY���������zY�>�Z�������{"p�5�����>��?J?�γ9����Tņ� -�s2��i���=��},�T�0��U���`�Lze @0,��R0X ���5.eyӷ�ҹ�O�-�#{���ÙI*��_�.�f|_�������ykp�.�.q-Y�� ��z�>����ߊ�uq���\u�b��O���_��峁&�Z`2��uN�Bw(�"�)�Z����A�6��ֻg�'�a��d+�t�^���Lъ����|���:	/�e��-ۈ��5���H ��0*WM_|�[Zh#l ��ߐ��/�I9#��8�et�=8�(��a���Z-_°9����:��t�{��/
����-�)/��)����4+.C`���^ӎۨ����v#��.um�B�{@��Iz�ȿs�G����6�B�h��#u#��@�9��:���.Ψ(&T�N�v�/�8����c0U��p�Ncf�M�|�=��h�E*u��
��ܳR_�3^�g�J����oH�VkDG��%�7`�.�Y���A�����XH1��6R��P�rY��5��'�F_J;�.KN/O6� {���D؇Q�t���He����;x#�y/?kh�j�������0�![�Ҧ>��.������0���D�)��9(�D�� �W�����c�����T��M2W�G@�G���9���Ύ�H�2f"& l��O$ǭs�;H�������ĜK `R�uI�1"#���S
�ؗ�7(%8v{�$p��a���|�n��-���B��5u����=5ʤ�5���@�Q	<_r]�m7h�ԱVW��;���aE��W��L!%q��2o����)�!�&[��?J!���w<I���8��*:�y�Iӧ���xQ��ƍi��q�W�[�(f�w�p,l��\��<�C�T�L�m�Yx)֑�@W/J<n�E�*�t��UAv�Uj�p�Nv*���/ ���XTj �
��|1�}V+ж@]�j���Y2M�i�P�T~0m�}�p���� _��n{��Ws�
<Hn���d����P>��<�L�xҜ>\Z�.��US�������v5േ�c�^��"Y�a����#��*:��MA�Wy(�1�Ш%�/u��>�'l*���[V�uuț��-�����F�ѭ FG�dP�q�:RG[�Y�H�Q�e�մ��>v,��j/U����1�aFWБ'� �`/���&g�Gh��p)]:���U�>���_�<׺��ղn���q�(l�/;��fb���.�ϸp���� ���<A͐Aa�03��5vB�&��i��RB��0_"_�B�EW��i]j���N���G-Y,<�b���t9B�:x�i���oy�FI��C�P�3TS�`Iz\��¦��/a�H��@�>�K&P��a$F��_pH6P�E��ٴt���%jŕ�@���%�9����rc���IÅ4/�{��Q>9�^\� ��E�M�/�HX!A����8���3�y�[�,}Υ�l�U�W��~�)�e�o��t��}�pn���vߔ�|_Ԁ�=B�)Ǉ+�5�v`��Mv������'�F�`��w��T#���D����qu�0��򦥾S�Ъ=Z�2���D�s[��&�@�ې���u��?i��#�V�%MŇ��~���I������!�\!f�E����s����*�N�⛟��x.$~,T������� f��ξ��ҳ����'���X�>Ҩ`�5h4n�<H��U?8
Y��^��Ă���0��h�����@��8yd�`X�헝�$}���%�:N��E�L0��)-8�o��
�YyY��%���z,rL/kܹǄ*�Jʘ���\J@��z+ 905�/��R=�n��f&:^(���r��,k��5�f|=�����]�"s�K��l� �y��W�/�P�F4��Ht3��m�I���z�n�dO:���_eW12��oY$��,x�87u=���<��J�B!6F<|vʄ)�,v3֗��J��r+|1�I��J�f����|'�0H_n�,��ݩi�vua��l�\�8���1�ۈ#@��ڿ��'��ÿ�Vgz�"4����i���a�����W��"���R&�^E3e��������b��Pe������v��$��QB�L)���ĞA��خ��b�>]-�]����ɯe�d��	N�����BI�O��s��r��/�pծ��)>O,��=��5X����Qg
	#_)�Z��P[Em�G��FL<�, ݛgv����<�+�Ȭ<�4��]�zɖ�S�w���Ls/���\:^i�*GQ��Ne ��ζlgmS��}<�Z�+�-�fa�e�5-�u�F3pLlO�_�8��z9}�%�P��gVp\;
�kSk���c��Q֗oPr��8o�0�eږ������
�zŅNV�ºo3���y�m�y��c�����1��4��c�g��İ���.�c��>�OcP�9p�/8���5���I���a���������3<���D�V�/f]Z�iQJ���<���"��ZWY�ޯ��C6�4	j��ش����#��ư���|�0�5�@m�*�ό�������ޏW\�)7��.|nLq�������}%�ݒ��_���H�?o{��Y�=��N	��J�3�P��}t��E�t8f����E�Fi6ʲ�R3t��ʥ���k��\?�3i�AQM�o!YW?X�/��}�=�oG���.�QZ�KLT����6���k���2�G+y�����Z�3���;U��{��$���O�к�Rp=�Ŧ����it���$��[+��BʶW���"�ad���	H���I��Y$$K�
��O]�*�y�T��.�������B�v2����ŀ0<����^Q9�7�c�s�FB"�@}���l�K˘L�/B�7�AK�-!W80|�r�1����������w愀�G���
��?��x�I���+����P3����R~.�N¥��9��"B��xX7��Q=�\�&� e�r��li.K�)ko p�{�bҳ��ƻ����^��g$^GNg��,�|�^N�5Y�xL�[yQbg7W��g�t֡-D��@E���J�:w�J�@r�-`ug��}Gu[M���3~��1.�mT|N�6򬎰�0��p{rI׻��[Cb5��>+��g� l:ec���x�jQ�eH�����4�U���H�Ѕ�$�0�<��4W&�Q�D���!�Y�D�1��H�8�`��$�ڟ��a*�A��Y�.jxr-X��0O9g��X�'`%d�Z��0����,p2w +����g7���2���3�����Ur6��	\���D�N[[^9�R�ZI�����		n5 Q1*���y ���������+c4��Pho��21𼗺`6-�Z7�QU�n u���} ��M m��y��� �l�$K����_7hP,��@��z顰����ř��6'ž��Ǭ�~ ��;��k+M��x���]�'�,��	�t0~�iI�
��z���U7 0_�Z�jb!��:A�{�Ҕz�M��NZH*������1�)��E���d���[�6��� )C���݋���e�L:H��b}cwuZ����p�&}e�yb�[�G��&��[e�)��N����~y#Io�U}�8#��wʁ��t�ς�ɯ"��#R�@R�{%�#����	��UaB�u]MT^�y��w;:�Ϸ
�"�S������,��?%GJ;�'�:�dnǎ�,��G��G*�yE���N��\�~w8��P���*A�t��h��/E�q�ʅ�緯0/�4�������[}�Ӿ{y�o�lG�P�C�YV��%5�ĉ���0O	�����-���Ldp��%9�5]�@χow5@��3ĉ����m@�p�Z��a�\���������h��j���][�]�]��G���:B��������?��>ߜ�	M"����ZS"U8���U�d�p<�	1�w�����E��k����y0�%8�<K�-؃�o�WL^p�ܕ��V�q����:T�|�8�hDC����)Է�C�c�����tN��u�1H��e��%?8O�;,v3
`�E�(6�0�7B\�����s]o� ��J�&3����W��+�n�Rq�6��[�;U?�wt�
��6{�m�jJ�H�-7���5>�N+�?��t��o��I[c�&6Z�h�cӎ�>����;�R�v����Pq7'�c�d�YG�Be�Q��Q��u7�)6�>s� ��H��H�;ՕJ��g��/��
|�~c���`��|�Wf����L��Jj�j�-5�^S
!v��rϮ۔�=�MU������&�aFJt{�F��q��W@�ͯ�-��l�	��~?�0�ʬ����k�~��K�X��6xkB��K0%�� �$�Ͼ�u��d�����0��G%���0�R�SUy��`�j��Yg�j4`�v��?�AB�b*�w�rTsH�8��Y�-qS^�q��&%�; J�@���/X��������Q��9>~�m�ǤȚn!��O�Yr�s��c���euu�e|_+���V����i]Ѷ k\��a2�n�gKl�;���k��\gL�Yհ�(kᆵ��D��oĦ%K���B���?�m9���n��v�AGq1���G`�R ��c�w�L�2�O��3@�IǐGx�+���~z��M��)�B�	���O!�L�'�x����Ʈ d��=���j!H���H��Z��8�2��b8��B)��Z'�D��:���I�S�o��~%Y�Y�^������# o:[|�l͙jxܼ���qZ�'ʹ��|6������PXC�dvb�H�]�|�v>�c����XwN��ŖE-c��6.�=_F\$�:
5�z�ƚ�v������I����誋mC�bR�G*�_��c"��M׳ů�����<%��N4�v\���?�/���bô�0��	���]ɜ�W��D�Ö.t�����F큤��j����r�a����ġ��sV���^4}�F�u���f���V�Oz�
MM5� (�.*u}8�0�l��N/�u'N[K�~\j`��SW	���j4�����Ե]ΥD;OSq�4� a��Z�)��t%s�Bh�EM&���a@�d1�]�M'�pV�:87��Q}7����|�sDc�܅ ��$S���i�5�-��V,�Իb��h�HCı�s��I���o_az���ǎܛ{'�8���t����\[�Ig��}�����;��^�}R:�Y�t�.��{���ڳ�xRg��jÍ�&�B&o�pk�+���e�a�tϒ�jT��]�tD�h:;)��t� �n�S�5�\L��kV�-?���c7[��b��V_`�����ȃ�(/}&�āD.0:0�-���6��`��l |v(�6�w	6ו�~++I��ޕ��5�
������2/��ծ��vM*��g��!u��C<݀3��>���BD��7Dꃘ*:�H�yt�G9��g"�ga[�# 4�F��1W�C�\�=Ź� �XXĆ1����f�":��Է�'�Y,��E6�vA|��{ |�exi"����~F�!�M}�f�~�BL���w#mk��+���[q���ޠX���>��.�A,�g����.�&�Mާ\('���;}�)KB�$�C��Ќ��@%l�#@߯y�`���eS�-�i�,~��(`����$˵0���g��4Y1Զ�e��<�>N2c��
N�o�i페ؗ��.�7�F�� O𕓯�!VdP�s���[4��jS��l�q������RO�݋��f�Z�k�v��;���j&?��@�y&g�qJ��`� sȌ���D�<v��
�AK,6����,���M4���5�<@D���{s�p���Ht�Q�ꐔ]�Q���}���b�T���g���x"E�_��3AwG��(�f|��;ʌ�c�l-$Y/������'�P�Rh�PT���v{��,E+�z���w@~c��s.����`q[pn�s�~���m�`D�.���`~�,}	҇)X��Դ';�$m���g[��{�؃��!��}r�GU���Y�^O���<�vuM(;�k4�|���E��jz�+<6(�2��k�R2[��=˰�=ob������7�`��qc�:B7f�@����������l�~eCH����v٤_���<���Q�I�̻b���,c���kU���͚�.IZ�o���y/޽�P����aͰg�����n�\Q/B:�6�.��4k�fK.�J9qM�D�J�g o���9�Le�Ӷ?!<����|g���[���#���k*�'wO�s(5
��{Cg�c;~g��mL�V�l pg�s":`����R�D|����W}�;g��b��pE�F~���Sp�ֈ�d" �1��ܕ�c�ɸ�:��D �0��0��`����܀��T�e����^Td��Fz���JA��?ʧɤ�,$y!<_|qD����v�����G/;T��C�ȸkav2r#�$��+E�ծĤb���x���G�?�A�oW�iʫ��c�@]�YessoN��~�SYę�&�O*j4n���Mt3��|��؈�e;>?dx��)���/i'um#�:�YH[�_E���Q�>R����8��VOV������E?ل��}Ӻ=��5T�S��]L`�;R�q[�`ٶ�%Kl��C�ɍX�M{��4)���d��w'�2������Z̐��&oJfNyѠ˜��D���]jQ�����j6jL�ۨ�QFSxc�B[�aF<�I��3����V�,�<�Ren�b�\`U�wn'����5�ꖆʩ�^��پ���O@e(
�!�0�Q�c}BJ>�� �ﭾ���u 	��\�[���G}X�R�`���2.�}��_ۙI��L!<W����p�y�,8��"9a�(҆чX��zsۏ�>��/C�P(�U/��`�<?	�\Y=��%	j��=6!�������ėvG������dN����0*#�6'�ڧ5W����3�M-��-W�[��!��?��rx��>RB^���[��$XH������f鋣����Ɨ�n�=1B�nKi��zKG��_L�X�V�/�28*:z�Xq��)a�㪊"#c���2�	H�B����S�.\"������t�U1M�@XԵY}f|���08�z����a�y�c0&*����ؐ�)�$�&��i�igػݧѾ�{8V��VJۈ*�Z�t"�q38a�.�^>���&/�y�"��F����e��犺00sB��g��Q9���,J��,��%���F���i�m2=���	+_:c
������*��@!�js�g���[e~]-PZ'6��tV���^ s��z6��G��A]�7�CP�Y`�����7+�����ۓ�5��TA���32w��g5�i�����2R�p-
�hl�2�m0�:�w)��e�j
�{9E�)w!��Hz��-�����(����$��`��B��z��w������ŷ%�(�H�F�l��e��3�����K��rk0;��'bl��	KYդ���1d�9"����K�<��ss��h��TF�=յe1o��F,j_��9W����]L\�ѱm7d�2�v�{]�-�˨�u�N��㜽pp��gb>��������\J��p�ˌ�-�� ��^Zwi2�e6j�Ve~�<���]A�G��x��`��W�<8`����(��`�t��J�Ql�
�@G�Y�)��ʩR(�a+ɨOB�+�����y�cP���&��҂�(����IXG��;*Y�|�pX(��A!���E��Wy��n����^�Xo�|G��)IR�a
�ɑ�:@�N�!%�J�_�2��S�<����mXVa,�����Etp�[�����>�{��R��*�?ܴݠu^�'T�;[4F7��Ƴv��֣������;����A8����	��jyJ�k!-h���t�BV�C�W�KJ������K�W5 9�D4[k|�)�������� ���W%�x�ii��k�#�<G�R��pd��`�YD�l�����&|��ٯU�|��*���)]��q�%��[m��#.J����/�1�L����;Q�P��pl;�jm\��}{�݀ԧM�`�\&z�T���J �+=�I��:�Ȟig>�>��7���W�Y���9�Z�;������k
h
�G�ʶl�-�#� Ub�N4�c��\�:{w�����������c�7�-8��%\�A��~S���M�ǒ�W;M��VU��)��K�I�6����j�Ňp�A�V�:�Կ�Z�%?�1��C�d��=+ 	��S0�[��Rt�	c���؀쎁<xT��e���ճ<���J}>��Y,HF��y58��JAZ���d��4��%>잾�� ��Y��Ȭ���7i�5x'�$���뾜 rc�wgB����ɠC�"�E�%�m�	3Fu�E�q������M�p�$�q	��;�"h�.�m���a��c������#氮���0���2`�[��ctX9&��ſ�7���f��^��tHD��<��Бِ�ì2r��y��������2=��!��.\��f�L�nn?�Fu�<y�������q��`7?4��5F�Ǭ���M�Wu���Q�u��vpL	����Z���Q�{O@dF!<&��y��
4�`��v�8�tJ�й�Þ�I�fa+�?f�I��sW�G�C|�7��}li��X{�7��&�VJ�_s l�t��X��V�N��Er#g2��v�o4�n:�;���x\<pa<���ugnўf�
�+����U�iF|3�A��E�~��f�� ��1v`��
�5H�I[�M!A/ċ��Ջr͛n������]!����#D-rA.�;�����p.��App� ��ö��Bn���
Ϣ����GUQ�bk�N}�z.]�
�����?��T��P�
V�~Q>\���dlv̳U��2۝jEVZ�h}X�b�S}E�홧R,�=ݛd���[5��8`S�L��c9��p��: ��E������5�p����)+n�����?���4�|��<*��Gr�,�2VƸ���R���2l��&�֒�߮�#XD80����W�M���x�N�i5q�� �h��I��#���C�`�
����(ѣV����ґ�Z'�ym�+̈�2ETͶ��x�.�|OewS�U����p���-���4�#�4�#�c�e��	T�%-iĈ@x+K��57���n"��Ѵ��Bt�9V�nV��n�)HDv��_�F"'���{M��E��
�?��{<cf����M
e���8fc��e��Dь��h�P?����l*��˅�)x�E\�����99�(��-T��8�����������g�V�S�| ��3h�!L7�ZH��q�EJ��:�198i�r.��T�]�A�U���Ix 6��<;L���^�J�V����z��HJ-�҉�����/�����H�ꀄ�-0�".�?��<�ҊAIbY�tE�D�}�F!��ȼ�Ȫ�_+T����dW������zI7���Ν�X��tOz�q�����:��*���$CG٭P �K��si��r�c�m;N����2��v�	Rq�hx`��<c>q3s�w���<�ɴ�?/c8�Y�Ev�q�\���Ȍ���嚫4E��2�ς���̩**��/����GĘ'�(�3p,�K��C#�C�/j�]c~W�غ�;��Ρ�Mb�nH�m���y��q?9��Uť����������l�Ӂ�.Z�@��ug!���}Bd.$!�3�I欮��f9G>����xZW���r{��`%�	�#��7�q��e8��a[��*O�?`��D0�":�i�6�9�@U%�+���>�Y?��(��|.%�v�Um�	,<�W��OD_���Pn�B,@7����d'\W�`����;��LڸF�C�@Ϫ+-���7���(s �wED�U4���;�@��^�tܹ���L��n��A`'/�d���9��Q�{�6�-��J�lv"�^+G�����/@u�շ��~��g���t�
8�@��C��]}Ǆ��)��F:��z���FYB��l�@V��唙L��J��R���QL��t�dnM�Jtœ
�ڔ��\�A."���g �⵾��;�����cu�w�>T�*7F܁m\�}�q��8�#����Gՙ�D�P�r�ʹ��h7�_�Dl܋=[�f<�p�)�O/��:[�dE��EY��b�1q��e��r�^����X��
5^�Ft&�7"��I��� �ɾ�̌�)�=��츜��N̜��	�� ������߸��������l<�žNq&���jm���&�u��|����#Ԅ�a�6�lW�IwR�̲�x�|�20�"��,4��Y-��8��b���~�G�̜a׀æ+X��<%�RIǴ�({����̘AŬ��	��YÓ�E���yqcΔ��� b
Sv��ZdbI�[)G��@ʩ��vRp��-��-�B٩v�X�%�U������:ˌ��E����jl?�B�d����S�j����.#0D�bA��+_�u�K�AOlo=�Ni޲�*���,!�D����0�]rG3����Z�_".B�S�K�*��=�5r��{�&�A�E��Q�;Y���)*1wj�@�&ρGv��+}r~���eu�ڇ�f�)���S�~zp��I`g�e�@�	BF��̀pz���E��z_ֲϢ~b���- 
0nD0O��_ǋ��z�v���2��FC�AԲE�2�.�Y~��z�l���;�5՚���S)C7�<%���@BA�ث2gd⍣��:� ����2^�V�U��%��s�t���39�b|T���J�/s`�6��2�4���h0�T����"M�a�AUڜ��;*M�(�%����$�u(�ȱ?2��y�����.�}�i�ρǆo�9^
Y����x�;$�x�9&��x��~X��KTmZ�%��')��V�!�U�gd1����X�B�����״�6=��'���>�P�K�����'7���1)#PP��*1Ъ�d$z"�]��}�Q2��GMìpD�ǁ�^LHo�V��&��t�!h#�r
Ӌ��WA
�HݮXC[	��d@��9��bIW}q)�|ÑE���s���` �d֋P�:����٦峩ܟ�6��~�;x�1����'�-�,ˢ/��LD@���$}c���@u�d���d��wu�L��F�:�8�_6_���%<�E�}��L����|d��n��?8\��K�p1/����OH��R�7��	���(�k�������9�蝳YGWN�|0@�K}ˏw�ʓ\��̨�����/�˖��_b��/7 ٩`��v�5�8`��VG�,VhN��f����e�h��}�� B�H��sD�|1{�E]�jS�P���? �+bQL��u��m�*��);F��rQv�z_c���r�I���8/^!�C��Q�����Qsd�R��)�<q�N�a9����$8D�`�������Kid �7#�MoZ�jZ�
�9���>u���v�GQ�5�~����і�xș���DS9N�#{�Q�����;Ky��A�>A�[����{�>͛1H�1�� S�Q�&���/x��Z��@�	J�,c�nyhI�k� ��O|�<����Ӡ��6ѯ�}|��y�8E���s������Vx >�f�/e�$�HB���v����:@�/�)�l�?�����!D݀���o�]�(G��B�(��;@����a��8q����L^������Ϫ�)-^8S��Pq��1Y��*_ѷ��ħ�9��4&���8�G<t!Q��,��:%^ɺ�:�M�X�b�M
�#�v�>�GS�1{`�:hY���B�����,nښx��-�/�r���z��e����Z���D����b�VL8���c�:���dTp��GkF�vD1t���_Pv�?�[%�1�R(�H�Y �lv�퇈�C���	�І=Q��R�_�0���`�cs�.������7���`�2Ԫ��)��,�����F�OPm��O(�����0�'=�N����K�j�h���eo�:�;-�XP�e��G��`�)Z5�EC/�+��&;ҜC���KJ�'��'�,F�G��t���y��VxmL&yetm��T��1��+˒M9k���hԫ:|Sx;ˇ���uAQ"��w�2���0�$
Ɯe1�s������8C5Q�a0$Xw!�H�a��0��Dk�^Y��&��r����ϝ9�2��1U��Ј�����ߤf�2�Y�9+�ihu�c���{ F��7tfN3FZ,=FQ�5X0{'��zNȝ�G.�n٧�F��:̓7�c�0�ZcC�����xrZH����O]f	]T�{�C~��˖לP^&�0��띨�-����BX�IU�@�3�bf���t� ,�pK�D&?�̋���x8lܥ�n��h�����ޗ�@6�HkPC98	f���U3��Qs��'-K��N�_��u~�H=�9��!%���d%�\=r�Q�|�(�����&���' ���
�#�ڸ\�(�}g��e�����b~	Y��m-�Bz�D� "
�����5~��+�ƨP��޼��F���H�P{`��dL�6�5� ���7�����X�ʦ;a^����4�8�7��[�`�{���A�W���QǪ5x��,�&������i����y�i�F���y�u/����oj����M����\���?���f��"�7b�Ͳ���0T]�sf�GoOZ��lWk����_�G�S�v�t����V�����!������*l�X�5ʙ��-�k�̘���L*[&�&^��y�3�_i�P���MȠ�����TsR��M�@fXR�98P�B�<5)O@)r�B���<������o�O4c��NƯ�����q�єm���H\c�4_�*���R�[��D�=u9DW��Yh���!�㛐��1�B�k{�Ӿ3�T��Z3�7AKO�G�d�v��> ^y���b����^���ҙz���A�����rF�y��������c<Q�6g�z�d7RK��02ؕy#�m#&�M/�&F�BO�Q����Ӭg�v��|ˑp�Xuylf���7r:���5�ނ�*���ʷ�5�xdb�(8�����-�)ܯ:��������X0#ڛ�۫u�kS�K'IF�/����]���4k��%�����.����2<�5@aD�C��7Mȁ%^���.��^�2wٗ����٘�9(��1��'�	�wkk�%ԣ1���FSN��(����d��X��f���d̺��wV!*:�����{[�d�K'�k U�v7_k�%��rv�խ��ZQO�V�{��B��˳�K��K�4�0��Rї�"����n2x��������w%Z�K�(�)���������C:�����VR��d\c?�x7ly�Q�Id�k%��=ǘ5�v�%���F������Q���%4:LA�]*�==�C��T�K	����E���H&�rti��5�n����cZW<wٲDN��D���$JP��K�Y4��T=���?�:Zʷj�R~Hg�����Ua�F��2���9��
�3 oR�n��q�
;���o�u3F΁J����Y��$������V�ԏ]w��>�J�s��҂i���A�w�ls�kwR��s�E�'��E��N�+����-\ޏ�o��aYl�;z�5Mw:�ۢ+�g�;�"_�J98a�]�&��1�V.��E��Ղ$FD��5(Be�l�O��UW��A$o�A�F_��?	L��x&��v�>̷B��AR���Ύjݼc��ŀ<�v��I��ETg��o�I�yVKb���b���8}��`���^��h1{p�	B�Ԯ�g�<�:Η���.�
��,�ۣ��T=~���+X�A����!,F f�W��A�j;��86��ni��P��C"��<ؔ�\#䉥����P�+$�7'��,kf$� ���\VLqQ�pT��?sS�k�
ա�MW���s�Z��ժg�d��'����l�'�[�G����W{��P�G��[��}u'��#����ji�����+։W;��݌�E��}4�������F�,� �N	%����A�Z�D�������Y��~4�ix3�lG!�^�%1D��S�g��XB9 )Xl_ @������#�2U΁ZPe�u�UE�k6�+	�y[lH�4��zE��2!J�N�e�[��Ti�	�V6��u�-��G�������䚿��73t�@���X��q�tF��몜���TsD�+\�O5jn�U1���Lر75���4*yyrA�@��;��m�9��9H��X���j|��{]
:T4��b��}J�Ĭ�z����ꋌ{�l���4Pn���*�:��}�$�	AH�ˈ�;�/7��+�}4�S\8������y�Y�}>�o R����?�����r֋O���X�z5@	(4�FR�b��ڧ�Ӛ�FN1�4�NC��ܻ����6�8�_HZI-��8�Q���rY`�O�kn�TZS/�ew��f\�ϖg�U穿Zf�惶*Yl$�~b:m�9��O��6?��Rq�H� �F����$e#< ��Y1�ӆ�W7�pPo�dJ�<�\V :�s�9��ei�w���XړFv�_�h1���GzxP\� S �ER��d%�7�mO��V��eAA������L�H��e��_W�,��Hq>�����H"NY�'݂A���s���G��VJ��@����"��d�������		,ΰ��b�d��Yp��O.�}p?�P�zJ�GY-r��T�o%�,�`���(l6*j���Il˷��ȝXx#���ub^�?�>ɒ����		�`�uD�����2Y�{^�l}�x�22��l)Q>����D��!}!�_�-�8ĠY7uQM_>�$��g;�H��<Q�VM!��W��̀T�X�ܭ��D?Iy�t|pyX"�3T������W�f��&Mh<��b���X>��V*dS[�HT��2S�ݳ���������y �d3;� a��i: �4�yK
r���0i)M�{v̉$5[6��y(iy����a�%�g`��~vߐp�[�O`d��	U^h��%�|=��[]�&�GXr��
� ��Lga_����hn�����Ԟ>�4m1�pxi���AÃ���6��B0�'0|Sy���Z:����xňc���R��T�1o��9�6d�3H$u~��_����2/5��灾����9�X�8��:��9y"Y�jɝ�/D@G	�0@�j����8�m&�u�)C������1��@���	��ށ�O)�ybf��b�5�Dp���H�4�R��ѵpw����i��CւZr�k,����|(��7�Rzay��X�����$FNIݹ��k|̋?m2��.R�������	�\4NZ�v�f�Sڰ�ɔ���U*oHUL��x��K�`�>�]n��B�����a6�ʱ�<Z��ը+��_��8�ƺ�E�3�0�q�+��|T���_rV���]���tl9Y� ��$f��Z<�iOBP�0�i��e���f��.u&�ML�;�-���:;�h�kY�,]���$lH�����πO�}��*�;:�ms�,L,V�̆�R�R��Y��"��v�!��t���My8�2x�(2�o3�-��Þ���{Z����>"��@����ya�d?{�9gZ-#�i#��Z���"������'��@Zْ!S�_F5��
&��b|�e�\%�떧�G����Eފ��m㔩bv��9��=�ϐռ�o��D�Ros��g�͟C���������$2��sE"��i$?��E׆]�Գ�xk�̉>"b�G醝y7`4�����]EO8��I@�`� +�̔�1p<v��{��'N�P��ǀ-��
z����s���1+�T�-�pR�t�m�_3���5��Z���̥،��^9�`�I���k��8�#�핶n�|�8��M���r_��u��:��X�l�&�3�iPEh����a����T�~�0<��ұx�c��
�,T���.�&�����ޗ���4��{�?sUXR� �_�Q�;VѴV`�:}P��z�L9=li�c�!沁��&Y�1�h�z�kJѵT�3ih����Q��<�,��`�:|k��9���%�o��� �DmՎ��t#�f�&��6�S�)<?�S�=�T��2<ҟ7T|Q��΍8X�ȑ�K���v�;��e��h� �����1_��25����;�kjXL<�SlQ��$�N�v�� R	��Ch�T<�t�8i�/S0��W�oؚ�9M���n�Ѳ[��N��Hg��D�b1N-��;��.@����H�;y����@*Td�
�v���0R�,�<v-��<a��u�uJ5��\����7�0B_�/�$��y0^\�Ym�ە��_M��v��*�\]=\��,S���4Eӥ,�������i8��v���WՋ�QF�b�GC�5�*ܾ��b��һ&!�o�c[hC[4���ϔ�K�/Un�����S���8z�:��̷Wv��m⹊D�ܲ,�����6(�>c4�@o�b��
�2��b|�X�/%�l���,��Ƽw�䱎;>�
��yk��&�S��G�Pw��=�Gti���J�.F�@�J�mH:�M�d�����m9�� VW�Jh�Pm��p	��0U*�;uP�l�se��/��A��ǐ��"��T獶����㾈�n�}H!�"�X[��yVђ2������>P]m���%T{�����^7�x]@��#8�K~��h9��],]2Z^3�m��sB[)���Ą�|fB�$߰sA���k#�&�z0���c�B��xn�V/,"���{�wf�)�v�d�I��L��+br��/@)8�f����w��5�z̀;{�� 	�l^(��z����mU�/<9c�6W��C(a(.?L��/����F�C��UK)8� �O��s0;G�c�H(}���#��V]"
$?�MM �m���u��ś��U�mq��hN���%0���O)n����E�Li�-��*<�4��������:5N���iK_���1T-�丮�<ޖR VD	j8fik
%fA�T�h"s�C�|�y���nURwe�tc׈���@�;�W��o�7�V;Є���j�fA�!F9�`���:�S�s(t��Ȁ��5A͑��k�P��0M��/a��5ݗD���o@�z�B��JZ��풔���*�eZ�Ԭǧ�B��do��w�c���E��G!V�;I����O�))W��;A��)�d�?{\{�%����&�"�z��<����3���x�tU9����&�����;N\��eG�&�ݳ���(f~a�u���U���A_?v��HDJ��{ϧ�EOWX�gb�)���{�����2e#	�n�g��Ś��Ɣ�{qZ;%y�wa�H�|��7��'C�2�ߤ�:�2�m=������uIfGT^H`��6����@t��U���=HX~�k�_H ���%X@`���YNR+�G�I�S?J;@>*:�YKG�T�����C�/.�r>	�T;\f�1��<a�;�mԘ�Sֹ���o��wz��x6�}11�-#Y|:�».U�]o䣭��Q�J[ �z�?K�M��ިw4S�H� �\���
��d�����e~(��������rD�+�H��}mE�K���"��&E��ƕ�{�HP;s-�#`:�	�qq��/\�'`୿�ٖ˫��S�5�N���=M�-�g��Qz���� ��k#��L�1����ie����[����l�����]C,�FL��(=5>�鵨�y�77�z�C�a_�:��s�
��G�V��J�?X��<�?�!盻^��ŸB�x��h�D�xf-z��\�uO��'xx����S�3 �4�3Uѵbz�j �C)6�[�j����wv��%�`��U7][��j�+���ڷ��j(,=j�݁����ya���0�)86s9��d�׃�C�rO\m:y���R����SU��r3���1��|�D~�;�wp��;����Os4���Sq�v/�UpEɐ�
gd =L� |x�bF����k���frK
����F��83�����3*^_WyKs*�K���f�ɮ�!٩�1�T��i�g]�%�2�� z�o:���|�w���fe|��m�׀}�,��Q"m]����f\L@��O�T��N�Y����;��
�<y�`/�M���� �� T���й�,��s��3�2���<��j|&C7�4yQ�����X��״?�D<�-���>����h�	�ʨ����k�>���Rzד�dIb� ��������?I��ڸ�,Oف���"w���(��CÐ�g��Z��D�c�ϰ>�A����*X2ͅ^�Ʉ�[R��ϧ|M|������!E�o4������*>I@�2��-ʿ��V��� �?� ���W����(�	�8Y�������z?Fמ�lB���ReO�W1=G��Õ��F�VV������x|�E7o��Ǆ���>4��uiu�'�u���->W�� ������ �JK��Gv��v��'X��I�W`���2�E]��.�̼6B$eBޝa ��.X$�G�/�D�|�T?i�QN�y�h`Q�X��A�e �R�s\��?�5W;~;i��v�>�x�w����-<�Pt�BWzʊ��W|s�էZ��|ޒ�ʑ��1^fA��U>�D����"Y%z�*Po}�`"x�K���������	@�D�~w��j�? �Mf�̣�R�y��Iέ�%k�a����b��}cL��n2S�Ɵ掽"QtICZB�l���a�1�r­�P���J�Xo�z�vb�ta��u��G~�­���煭�`@��LM���>!Hu
���ʂC�ol)����j�!���^}�^�Cl�˽���I�&o��X8��y��ְt���A���k�l6�)��s6�_�0Yо�����R_�g]���̘�1c'����Z��,R8�����b�i�\�νWA�'>�6 ��h2G�����EG�P0�������(�X筨'WJ�+��ܭ,X���Ƕ`�<����U�r8F�l���G�$L�d���=ΣR�a����� �6�t��5Ү�UhqWyI�i���fp4�DƏi�����j(�b���J�h�g�&�BL��z�11�*���U%pO�BHo���[�}rB��G�5Wy&�!:
��$�yc;���(P*P��[��	��~�]=�V�Q��Ss�A#WƤ��%�#l�2�<�J�`oA�S��tQ�0鶬<H��Btů:����8,/Zw��W׊�*���#Hǩ�~2�ŀ�K�Gq��9�p�>��00K�q�W����E�d˭�|�zLOX¢O�ǧ�R�3���r���V��?e�55q����ݨ4R�7�9�qp�W�|�f��5��\Fe����� ��ǭcn�b5�BP�oc<e�������:YC��h�j{f,<�;��\8I���:��=Zy�}�Z�_D���(Q��MҊ�Yw�9!������V���C�A稕��3Ҕ%�$�%IX�L|`�QO6���� �B?IZ���ޕũ?�>�+Гe�T�Os8�"h�Y|H�<�P_UE���=����m:
O�A��P�D�M���y(�K��������&��ݙ����2�|.2Eo�TU�R ���o����rֳ�	cIC�PX;�C�9�m�8��5B���^L-Jپ�1?A��O����7��*b0y@��t���!����iF���a�>�6t���'\SJ�O��DuН�+�r�	:�. ��b�I���B����u#���^�$�%o+
�ً ~k���s^,`Q4�^���j�����6������0����x���I�����c��;2X�~�����I��+ b�JѾ��,q"aњM#��᮲��MŶ����2��6E���4k�5�szE/ijLtʶ����4�U$���:�{Г8���ud�E�P�Q�v��v�;6K/ف�0���4�'��I"ya
��*��9��eK*]���5­���F��=�j�J.@]Hk
G@�A�9�¥2��[$�V<Fw+�s�e'���M�iق������줺P?{ryD�}(�-�n91N��>�_c�Z޼�l����au!�Y�����qr�H��Ø^�h�qOJ8�[�s�@p�L���l��0+�7{��VRf���ᬍ����H��%�{:m~�1�ɉe�'��c���N-����]� 𔑅���a�y��|�n�0�+9�t�FB�c�}������S�O҅�]�"=��uˌM&�Qs=N����0��Mx�%C�4�U��0��)s����yÙ�-�K�O?)ܻ���R�ugCm�aE�2l��~H���O�hX�fHW��F��M��z\�ݑ�c(�FK�D����L3x��ϻk����&
�X����������Թ���K@���Cz�ə�(�ɗ�9�Pͯ�} �S>TҠZ�YM o����f]Mғ}/i~����qyB�X!kN~����pr?�_O	���xB����;V??�u���=�����%�ۯ��{�^Zj���_+{�[]�}԰�ʰF|�VҨ>��Í�j@0�[x�eI�O)n���c�0�s
�9ԙ~�rZ��$J䫅5b*U�:�BD'��f�o	���ǤyDh$<v퀢ǕԽw�%0�G΁iD9a;���^Y�����ϖ��k������S����#D�.�8bLk�5�?�*=�)�@�B4<%�Y54S�_����=�)w�B�mW�h2��wh�8ju��{^��2���k�q.��\�4�=x�G�	:��	��Y!�Y�P����Az!��:V�K�1�����A�[r�+���T�k��kM���T��R���6�;mC��}�}T��ǟ CϮ�|*&a��A����z��P��S���p��]7
�Ոw:��˱��f�X��K�����K� 7��#�@�0$TyNu���"���g=��˶�w��o����IVݗBe��6��麰�~��*2��K������l�Њ��_�yV��@��$g�>0�l']����m���fK��<���L�L���>��3c��nv�+L
����٥l��8ٽ>�5.߲$h�J�LׅɳўP������qG�Pn<����`+!���2Z�d�)����𣮔���>´�T�T�e/���N��-�M�\v���-t�1�/�����j��±!L�&ACU�$�bR��#X��-:]rt���}�8/Pja�E[ql8�O��_�~d�N�8��Ξ �n��h�1�t
h�3��O�@h5��X�Y���sĊ�<4��/۰ü�vϝ���yfb	q!�'2A5p�>�Ș� �OϜ��P��2�d,�����dn>X�qA�	�8������Gu
.������8"����V!{z�jlZ�`���v���FH�4nJU(�A��d��(��?��.������9�~�Z���c�%�D��-��Z���I�\���+C�q�����Qˤ�ۖ��ICQ����5N(e-���5l��R���j_M;��)��WO��O���H�s4�xHP����]��z��5�m�5�#p�@�VN"�3��)�D��W2��yv��ap�t�<�v�/�BI����JqN�f/�Ю�K�^w�4/a�[�	M�!HG�Az|��%�md�qZ[Y>LX�崙&!9 �0 ōC��0��]|�Z�5SG�Q�d��v_�3a���t����1jv����=�I�"���~S&?�J���R�Q��9�av�w#�����Ո����L����Bzi4eQſE�~�E<�,/�!r���+���a؎eSj�y�r����I�� ��[G�L@�;�䆮O�.&�m�uuA��NJ��N6�E �һ��AzMp��
+}N??��-�7X~��:���Uh`�nĿ�O���+9l��l��_��E{1�%G	�65R�
ДẀj-�	�)C��v;�:�L�47ݷ��^ �?�lMz�n���=z�P��0���8�o��!1� �G�d���&�/�q&?=���?c�y���Cڸ^��2��w�ѣ7�Fo ����ӛyrBcJ�Ux�Qp��t=N��ϼ��;�Υ���C�Q��0�D��v�7:(�� m��D���A
�DZC���U�.8AE}���H� mC��;��J8�!�6>�5���њQ�XZ�{\6#�wr���N���<�����FCZ:��,B�?5�"�2�$�;^T�<�A�F=s-b��n^�\{��d"Koa�"���������=�o�tF�dkŹ;�@�y��6�^u�Z�faB�;a�.0��Mת�lΆ�#�t�;�������U���$�>I��3� "g��u��zӟ�T��QCjJ�>RC��.�G��Ȃ����!��'u��7u�H��vUl�eD� ��˩�G��@��8"<�#��^S����#�����Ƴ�V�s�>�%��W�~����nc����pZ���hW�UJ��T�M>^���W�����J�8�M�����B�]�YB����!��~�AW<��yS�Kš���IB��>���!2�T.�\)�p�'���&:�%_Ȟ��#�Y2���"� �\�O�`�[�A�	�>�k>��)\i9Ҵ�B��H�<�ö^�5��m8���ue��ڭ~{!�Y��g�4GdAV�?c��,,�7S��b�QB�b�Ý�WX��]�%�y�� 2I�)�e����MU�M�[�F���i����t�9�y�C.�����/��z�����hB�A�=ЋI!̀�/��y;&�R�w�6����B�*��ii�Xu.M����O�הaP����1�Z��g�`&@X�dp-�8-��}Rę��פQ�����cq�J�\O���L���ˋ9�J$�)ǻҎZ $`J�hۊ;�jQP�,nÓ���Q�4�n�a;+��:�f⬽�����@�/�"i�ڣ=�0���9�kö��Ҡ�5̲Φ���R�$ {�Ȑљ5�i�U� ��8�Ѣ�7O5�G`[�^��*I��K�˧\�ْ;de)b����B��N�����.��|=:j}p�q)vp-G֓K�u,�}Z6"�q��S�rT��_SW��v���~'�G�?l<K�
����^�)�5���&u�%�U�k�H6Ē�CՄ�����GR��j\1���I���c��]��c(ctc��}�ɭ�r�,�?<6�Xq%e?y׋wmaίI����&��0��f4�cS�[;�<�Ԥ�H�S��M��o������HT�ǂ}����"s�-aųCb�q��?YUU,�L�Y�Z�[=T��^�v�e+;�Hd)�F�.Zi:2�i�7��ߒ�lEE�l�
J��zFI!PKV_0���c۽yH�a�u�̟�\ىf8oV�QiߗA����<TMI	Bh��?��[O�J�J���γ%�8a~K�����V� >?�;�&Q�.�u�4w�3����N��Oj[g ݫ�y��E9�����0���5���椮�??�䝺uʦ���;�N*t!z�\��˄$_�z��s	H���X|+��^�4Qpe�75u�yg鏐O����|/�F��>��V�+(�oĻ����_5�t��R��s
�����
�B�@�C(�"��H+ާ�x��%o�'�Ӳ\vZ��9�PouT���dF��|?�Wͼ��沷�����/v�0"N��fs��G�\e� ��ҭ��/֔Њ������U�5���' �vҋ]G�L/�Ki�/@G��$��ē<w����G���0�̛*�L)Q�b�K�"8+7B�U=a�_g�4����+	�;���p��1�.QH��o����e�2���ӛ{�ϣ�Á��FhW�y�U(c��x)cC.`��↠��i�t ���Q���檂LA�ϵSPw���%��qxK�%p�}�c%�cB��B��A�vT؞���~$ݓn��$�t�z��|qnSU�z�2��^:���! 	P�)��=7�����kcE��T��U�>&���*��6�g����:��:'!/�H΍FX�̌�\L��zf��4�+*�~�QAj����B��[��	����/*��̿L��,�V���$v.�"c���.��_��������F��BT߅��Y��
qӝ��Vǰ��Xv*M�u�� ^�퐴�Tl��\���h�S���"vOȿ7������6�Ő7��`�m�U/�% ��-E1m�[��jO��\��	�Z(l4�i{��7�Ɗ0N������-H'^�k`?L ��ə�V5u�$)Ct[N�m�ğ�++�#0� w`g	xb��6j�h|�>��lm};r)B}�o���T�PJ�����1��aR�+x��k<�Ϋ�}��'�-.`�ʮ���6EͺU���jh�!V�1/�_X�����w��U�H��ib�8�J���ی3-�0���ܖ|���+LEcWE��"m�Е�[{4�5��y���j�e\~S��$���9oq���ҳf_�?�6�|2��/��]N`H��/�PL'���(��I�e��,m�}��&z6���l�j�-��$4���;����'�"Vex�s����^αT0��=�s��Ø��Î�4g:�/�r4H��a:�&Z�G��z��K��O�7Ip�忪X����'�i��Z(:�n�ge]�6̨�Qd���k�0���`B�CƾoNi/���t�&�mk���)��qq�|��x=�pP�{(��$2w ?3\����@o	��.�PM��$Ƃd�����6���������Rm\����W���#���Vi��HZgL���${#Y 1��:g��z:�kj����Sk�_9XN��K]H����*_��7͖r���lobj���6C�,�IK��@�*h�����,2UP�,-�g���}�,�kޔ����W�5�p"/ǵx1fe�-��#6��pb��ιx ����|�O���4�ٮ��>_��Rr�B�`��:��A<<���
��3 �-��	[��G��ߢ�ދ�>�0�r:��u~�WR�/�Ul5@���s�-c`�f��]ZJ�`M�!@Y@���;�&�	?ڦJ�E,�Y �F�j{ �ۋ���"|�Lq��h@W�6�m��Bn��[ASd��;%&�4l+8ۮ�����R�A������â���D���E:��Jf%iM�yL�x;Ő*#[d�`���)����FS�U�����M@�
�.���7;�������/��������3#��hդ'�2j��j>�Д�XN�bI3�6Xi�qy�9�Q�0��Oh��xڼ`#�Z�s�}�}�����쓟O�r E}>}��� IO0�Ĉ̔ �h�v�6�
�L-���[��{m����~��4�C���}jMDt[�2���<ԉ�h�n����x��	˃���~yEx/������zO��&�SC�o�W4��"���
�$Λ�w�JI�z*B}��	1M��Ma��DaOkQ�S�Xc0�����0+��d��E�tÄ}V�H���g���Qm^PR��5�v��5U�{�7?���o�?�g�xJr  8�T�dԛ���"ZV����Iֽ��`(%^p�e�>w���-�5�0jp����.��k�J��DNp`������rB~,�WT�����!��>#�l�r�����x���>�SAt��d�G9:���c��#y?� ө� ֩!2����<D7;��X�m8��l�p��]c�����veG��G��2|@`^�Ge�7���	��iܒ��KR����n�k�.�獑8 �Ԧ%lM�=�S��hu,>�������l�~��+ =ȗH=Զ�F{�
�BA'n�	һ��8�7fA��s!�8�}����#7x��H�ǣ�M�͞���,	�~�Ř��ٝ�J�~��0��`��#��mB  #4-�˶�!z�v�{l���D�vC:��K=��b�T��\�$q��w+1�nS���U�7��`���3���s����φ
�^]�)h�Rk����T���d�Fi�B�Lٱ�|QSJ���PAAe�ck~6��vwV,��S�i.%�8�i�뾒�T�5�K]�Yf���U��l�h�?	6�w^Ap^��_w���-n�HQE�M-"�=&([�3fLM&��a?VH��հ�Y�r2�y3I�}ط�H X��͑UB֖�CWimp���
�pB�� �\��n�2g���em�O� W�E����@����Ur�w����ȸ*�?Ab,��U�#ʷ�Hp�f���������Vc ͻ>�zS(�\6���.�{( #�0`}S�:h.����<�C}�c��I���3G1x3.6���;�y�ϗ�D����q�
L[O��	�d��d˭Sb��S�G��o%�"��g��@�|��T�*U��_�Ԋ��hey�U�R�m��I��C�ȋ�
c�˓2�I��S1q�Z)ZF���.�%j.F.lm[/+V�}�ѹ��Y&9�V���EN���Ֆ�am�ϗɀ";�A�H�ߙ��t�:U��67����'�^+(�.�v�6b@�	���(�TY��&�H�]7�ub�7�2�0�2v��u80ϣ�R-�>�?ʮ�ݼ�눚���F�a����	
��0ľ�c�,��˭��QBut�t&{�>�"�xlk�	MU^��� ����e�M;�v瑖��������y�u���j*MTCo~���Ql g��:dݟ�3]ю�{��E��L��2��ˇ��X�K\76U=�m��>��D��+��~�!�8.���]�0��i�y
#�A�HE�D^Z�)P��/2�KVh$zZ�DB`ݒd?�1B���dB�@<��eD��enƟw2
�D�(>�T��H�`���� -}�(�� �NvU��	1]B����"�4C����r����9��_��-3W�VX&a�>:��h$#9��a0E��,��7'B����b��v������u�S0j��,zҵB/��rG�q[�|t1��2MSO�F"{R�n̳��R�ۑ.S�d��іNm�3����fNb�Z֥�(B�-H^s)-��w�ʆ ��iV���=���K��@����fx��y.��!�;q�'�X�U�=����8	�r�IcW[���3A6='�[���A6X�F��H���z�;�4��Y�%������'�-xT�%}�->�Ǡ��;��NMg�h����Y�c�\�W,y�L�X�M5���԰1^Gp����QDԇ�o�Z.�&�Dd��^%Y��,犟6�Y�Fc�ϑOaV���=��@�@���5s`w7��7�t��D� 'a�1���-���{P�K�P�<c��&�aS�
�Pm��_1h����t�O�@�h��D!�����|�����!��ƈ��U� �[`q4rq	!�ח1j�&��Ò�nW_ݗ	��X������e�����C�T�O�jM�~�X�����k�u����]���N'�koJw
�Uf����|�]�寐4��Kh���~���za���@_�<���<�"C��"��x ��)�,����|�N����w�d<�����J��B �o�(C���?_$$%K���+��SUD����D��|A�@I�x4��9��oZ��	7����@l=��-�}3�'�|����D��h��ng_�K���V��_�#%�zS��xƂA߀f	
?���_��s7���k�ƨ$���yj#�y����ldI� ��P�~��`�v�=�q����dW�,�|��u��;m�~)��e���⚃l���c-��Е���ܳuemW<��w��h���H�&e�i�G��i���k������F��suZ�:&�����R��w��[�����߱�]`�Rj���j&�ܘ���K ��x��<w&⌽�5�9n]2#ޝxaQ��Pr.A���0�C=�Q =a�/��ޛ9���a���}�]�3MF
�?��XÖE�N��(����I�FI#�R��� �W: j�K��H<�HR��KJ̀�`���AE�F�z�ɱ";J�-��o�=��N�����N�����2�f���ܐ�Rr6
n���zt��/m<��~�ಀtw�'��y�aZ��>g��M��
|{��o�E�T��!	M�� ��_�UX�+3��sR��la�)e8*q�����F�����*�kҏ���)�0��+�x$J9�{��t����k��n��o�9���e�H*{#���j����|զ�ԏ+��Tvs ��c]��ZY�)��DP7ԇ�fpѩ�r��f�`�!�a�c5�4+�{,w�� �aY�D�on[~ن
P�r��Q���j$sM��%���f��������?�D�"F���[>zjuN+a,�+���Cj��8����_�i`bapE"����U�Ӥ�;�� J	���y���S��Z��� �б�������j�;u�ş���k\LG���rB��Xy�WhUp մ͞0\X뛣P^Q���d�>�Ų����AƎ|+�>�tv�PJ�Z�ie��P�WBa�b���Mߋ�꠴��8�C)�
�E�r�Lş����̍�m+�$=9��Y��U%����W����\�̶{�+w�#�b��v�DF��Z��vO9>���繲	No\X��hO�[KsX��������g-f�,Ѻ���QP5�9�k���RV�����b&.�ݤ G�Vρ7;I��3!O���G�ă�S�i�j�L�SE��ݘ`�I�� S~�>��_�����n;`m2*�;Ah���6��՚��(٥Iu��ڽ�%��f�R��52v��y�4|x��s�(C�U���^Q_H�vaL�<j�`D}l��N2-���:�!B�H˥Bڒ-I,k�`�XuJ�N� s[o�O��B�(�7v���{L�#�L�EOH�F��Z��?����e;��g;�.�A�W��`9�н7%l���<1����������ۉ�v��7�>%��p�Ar��xp���˄1�:������y�\É��E��O�L�����Ac$��w=4���9�S�a�`Y��|D��|���ND�dob�F�ZةSl>?ۄ��
�5�r
�rx�a�#�6���+O�&T���q�pش�^�6�*�Xt�E�(�3M7��� ��{�|d�w��с��⓳-�8�(��\��վ�y����M[�7���_k�W�����'ⶢF�&VۭAlUO*{u��X��h1�|//mC8�c ����]�ER�٘����(]˲sy&o^��q�H�+����@�
2!!��!(HN�M�C=OEle��X>D�)ci%��G�G�'����\���hS���& {�vC�����`� ���O�{��=�LE 87���Ď�LFe_Gb�:���g��*�N�BpQ����_��#j�t� �Xq�I�~{��<ݗ��Lb��ۅ�N�TH�8z��skQr�4�F�OCq��B[J����H�)�����w^��"�x��1�ЍL;��%�R�@JW�,�h��5��@%��X �C�����vK^8��������&�_c��[�cl�3�@R1�d���1����wsل�gC�%ܼG��El">r7_Zd���k4�У[	�|mf���Au�Nu�����f���hh���H0�я\��1p����祿A@�������]�+�b�95=S
��i`4
� V����H���G�A��J�TLp*��s��:�M*������j�ɷ󕕵�$c_��N��h|P[2E���i���i�?�gˁ,K͑EC���IB+�յ�}<�j"> p ��1qB;l������O8���vj�ˌ��Y���bZc�C��w��o�� 
�4��T5�~I��n��ӝp�i�S���sn��S��/?�AO�"S�s�ڣ����Z�7�^, ��i�t����W8�ܽ��U�!�'�p�X��A�C��v)fs\Z��|4��%����8�Cl���&:���#�tn��O�\�s;Up�gyEp1	�C�F,c� ��Ѩ%���}�B.
�S|ⵀ8����� ����nͨ8�������.�?-��Ձ��pPM�O�=� q~�znN'�6��j<c!���N�l�߬n���-3�Ɲ/��Zj񚆩�󅘈#
�NF�c}���0�Lb/~4�q����o�M�<ſzX�)�nm{�in���C;��a��.���p�-�A��Wqb�ƚڬ'��8`�9�
[��h�\��~ŠOT�����&������~����2�@A�^V�Cm.3)��8ZE�������]�s'����>z]�nn��^$���m`���y��F��I\\-e�a�g!P�������M��n3Ėo���^htJ8���׮������'F�v�?��c蛋(Z%V���fY�A<LB�~��F0ix5Z��hLm2���Vm�п��w!���8mb�4q�5V�N�j�؛���!����(�)%@A}E�4f�W��=�q�>��f,�<8,�$�.}��g�3ŷ�S^P�	�>��8o���̕����i���}	�)8�����*wqy#��0������Պ9��{�,���B�sJr��*���S���ۘ.���[5^Rg>`	��ʆN��Nyf�Ge��lvǉ*	�8�{̸��WP+��m��w�*�N[�Fyb"��Ȕ��\_Re%oR��h��SU[�o�=�h�k%�
c��ى�$.R�#�FNɗ���W�K0\�xl�c^g}����:s���?>�Q�������w5� ��K���u?��-jWI%��:�o�Lq4Yr<����m	��aQ+��M2?>�٧u���i��!��+N_p�����[���ص;|�~{kQ���.�u ŋV�� �U��J�<e+K5���כ���vu�·A":GW��Ɛ�n�v�qU?���L��k�jK����?'���l����x|�X �[��,�B�Ǫh�s�^�	J�����ޅ6V���-�;u�-H�[�d#3F����h��a��@��<K�#<P�'�+.�0��/��ŵ�3�z��������G��_!#���s���x��Z���;&�~��#D�ҶS�
k��x\0 L5����H��"��"|��T8�O���j�MnG�L�9% �TR�("�)$/qĲ���MH��R�pd&�Q�r���Ξ',b�V��hL,� |��f�T�HP��߭Mc��YMG�,OC�k���*]Ϣ���mPl[�#*u���!ȭib�%Gf(��|��_�r|<�R2f�uI��m�h���W�t����V�炾U[��xsN8zM���#R�8[v*�B'MQ�Y&d�l]�߸�IT+[�ɇSϏ�PS�׼�><杣EA���^'}������"�o�H�&8���k�����-�Ҍ��s�*,�0y�O�(�[c=�
\��������*�y��ߛ�qG�3o�%;H��N>ы ���������*�I�VFZ,�f�T���m1��f�	��sE�`�E�~�����񦮩\2��Զ])Z�_�m��� �#��kqL�|#�����K�ѡ�� ���R?ɦ�d�Mz-��+�5������u��MĖ�^�Ϛ?�N[k��-��U����qHп�$�hg	E#�G/`��z솀n��2��ʳ��_�<��MyFx3�k��E�����oOm��a~h�X?N���u�P�P��`�������� ��dps���D��ԖNK�>� v�)2Y��� ᖬ�gt�
X������ws�}H�÷���&P�6w�yj[�R�㚊����������B�s�R(ԍ�}
��;��X_��x5�q��cE��y&�&��l7��tzç��\Ĭr%�)�E WI���(f���X�}���ɶl�Vݡ���x�Xkʐ]��KɲNy��e�=�Z�0K����#��(?7�5fo�%J�:o-�x�=�I�F�^��<!�'�1�}R���U+Jkv<$�/����t���g]r�6�unH.|R)��� �5W~!͈�Į�0R�mSX��ŋ�:�V�1��L�$�(�$���m�f���ڬm�~�87�a�~]`������x�U����s����d��G5WE�B�)1���m�.��DTJϵ�O?�r���dO]1��!Ϲ�w��t����&q1�/T!�j��a�/a�)"�{���p�4�W�W��d���"xn�=��4�"P�a��Β��$�ho���F`�O����#u��zUb�ԇ�������W鋪�S�<	u����ԕR�E��[�}}ʨ����(E\e;�����b��
��v8�J��4�4w�Sj�Zrұ�_3�]V��Č����=�Q��9"�3/����;6�)� �"���{��^"
~.ZܝR��S�y.4�䐁Ut�����x�����2�!>?���B ��dᴐ~5S�#��u1[W�b^<6R��mt��=�73��<���3��ˣ����kJ�w%>3��Ek��x��]�M}v�G���C��Zk�y�m����&��clf+];
���(����#�g<�����o��Bz���u���Hd
u�x�����@��r�"�T�"�"�D�|�����6R��L��++����6�^b	X�n�*,)-���)�csqV�_R&��;c��j�!��p {Y���)�̵��e�;ݼs�r�h���X��L.I�����g�6[*J@��>��2���'*�y�@Z�����|�z�G�H'��&z*_�n�e��y���;�Z�Y�|����I^�Nq�)U�4,���/;���gyq���`O�Lc��ۚ$��	h�ܹw ����9�erS�+�!���S�I���=\�<�+tg�0����T�,ٿ���$�٭��I�z�Ј)j�4�(˟'�s52!�O���Ie�����[)��"/��� ]m������YfР[Ъ����`�ֳ���|
V[䇿�$ǃ��1#sO��i�7������1�������)��v��#���;cY��Im�����9���5ɞ`d�pN��"����}�o+�
NG�5H0�	(-��_'v�O�bi��v�������j�C�W�+�gCA?�s�V�f�#>�Fȍw* u���p�^���A%�  ��͂�P��W����]��tS�����^ 0�\�<OўCrA�_��A\��+a�����`n9�-~Ƣ��ܚ�d�	#o���8���߽T���3s 0��l�K2��J�×�&H�J�7�PgȚt픭,�M2{fݞ��uZ�Y���.�(�
X�U�{CI�@b��~�\v��APz����)��@�H[Ŀt��ԧ
y� �ԯΩOj'��$E�����Ϭ�(
7���ǂ*j�K3&�B�����H�wM �[�c�2z��:�������^�d�ah|[*�W�;p���A�����nu(�z� ;����e�>�ӔS��H��Q�\fx{>�*�p�L����G���ƽH��Ju/مJ�l�;2���d=��7�cbnǴ�I��Ɏ��a\I
׫��M1���Q0i���e�5�19uOo��7u=�کO�L�^�0�-n�ޅ椔;�VF3�Ⱥ��|vfT��1��'�����P����	i��Kq�{OE�b+���:�i5n�n�)D��c�+� �X���	7Y�D!�� f���K'����Ԥ��x�g8�Y���x���a@J���T��s&Ν�LT���r�������j�uE݉���W�)?RVM�
�s��V*�;�TmIP��Y�Ҧ�Yj�'
 ���&�߄]�7[�
f��X��R��h��<Z,��ڗ�Т35J��'�&x�I�0(_ �WR:c��Yit�LU*��'�O�c�m����f-�Ǜn�w���Æ*f��@���|~^��I��-Ey�,Ϳ�*�&�6�r�1>3�)�ż�<��9b�6Zh)
�dV��GI�����ˏ��8�m�x�����q,�� �J[��3Vq�C�`���4o��m��Yx/���%v���և;F�1���5�h�d�T��pw�H2��٪���@�3��z�	*��Jz�k��8ҏ	�tE�L%�@c���*x�E�M=r�k�=V>3��tJG��w��2�.��9����|�>�N�a�k?ír�qr��o�UsK t��ˊWR��d�4��.��@���fw�O�P!x-w�EٲƬ;�*"ș���O�6:6���WNZ!ng����4v���H6q j�����m�,;���hQ����� �V�Q�0�y���C�!�i�g��EU%ƪ��� {�ɽ+�5wp��e�=}f^��UL��N�|Q��Cwg"�Q՞Hܫ$Y��iQ��k�GN�DGo{.L��Õ�J��ì8���	��|G��l34y&�5�˸7�4����V�5�kCS�� I�6�15�c�@-�pe���v��RSz,D�۫?�j#y=�=��@���/������"� Xx�+��B������� ���263��J�o�|O�h�ĪC�uM��"�E����\pY��� {ݏғ%��׆|���vt3�уd����dQc�? է�%���t��CY)������~��I�z냮���^!�.��$��XU�Iz���e�U�I�ue�'���ay��ά��F���S��{���e]��O�a�υ(�,��-�����>KW���M�D���<���S��jF�
����k�8�;��U�_�M��ٶ��M}���m��@k�:ӗν��| �y6��oT�8I�L�?T�3	�y�8-Ϣ���y݅�gs�Q@�'���פ��C�$։��m���#�&� �C�������4З��Ξ��������/�� +g�����ԚQ����3�͛���,���+��ut�!z�w e�l�����x��@k��m֤�EDI����/��1�:���t�MGzu�Z�������a���rii�'�J�}q<4"�0䛮N��;(J}{�#J9�'���䘎����_�(�:�]
w�����ń}X�L��Rx^�r�t^_�K�&�����C�u��v�W��7�����H���HŘ�{p������UazB'}�'
�le��4(�L���(L�u�Ӈi�}2��v:m��M8w�HS����t] �]=�������TF��~"� �(V��L����r�c>w��u_bҁ%I{���8
�'�TMs��yỄry��w���B����4ͦZ���C(R7�!�d��=�y��
]L^�����n��#�������
R�����3&ć�+e CM�t��h۶�t�&��)l�f�߶�;z�����8dφ!Y/h���b����h�pD��#��NO��Q�EЍ���s�,�>
��;x�-���b�4���ZW��;�P�#��:lpiGAG���sj���c�����E� AG���S�w$o�x����h���_�"gZ�K��ܖ-���ʮ��$�<��'.���;� ��~��nU��.�q˿.͢����帿��^�(����S���ђi'��@����J�D0=K
�8���I[���@E3	�������`H�P��������c��Ji�㹢�r"e�5���л��<�N��|�����_WU�h"H���{�0�5HU�3t�ې�O�l����ј�,5uL.�;Ǻ�G,�%v�q��G��g;ҳ��$a�,)!1���y����t?�PND�o{ˎaw\�ܡ�@mg(Tx����j0��^�6�a�z�2e�0$��H��"�o��F!��?S����{�hf�*3�̬�b/��ú-��s4?����Yh�T��6,���S�<���'�ΚpOdMT���Y����(�x^�/EYT�xZ�r6&�r��[3��LpJ�=�UX�f
(��սdJ�n���&���t�P�(;g�\�9`�@Jg�9��&��#P�=�o�{!��*D��.v1���n�"���(�H�"�W�L7\�fE���ִ��i3!E�ݱ5ko�>T�[��.���:KbV�toh|�3��";q`�A~3_�Cr�.v��r�=*	�ރr7�Ӊ�B�6A��]~pr�ϼG���eh��f�{�L�߽�	�~��P�@ՙ��8p,�^�Y�}Y��qW4���#�@�4�4%j��c��!8)l��A����:X�lb��k�vR�l���&F|����;���y!�����������1q�ԧe��jY_���M�P�ΕZ}�,<���^���h�nY<�����G L�����H.*�X��z=��|�>��/<`	����`q�l���W��ʙW����$:��t����*E�h.����M�뾆�|�9[~ρ���d<��X6�j~8�S��%�%�<0g~oc[x��W׳�_�m�vH,O���8��F�Ӫ"f���aQ��B�ZPAka}cGS���
�o�6�B�ى����M,}���X�v>����1��>U��cnt� .��S�k_�jD��i��KX�` =HF�i�`���[X�eOp%=ؐ��Ҵs�at?oZ7 Y�hH�,����+�����Sr���b��]��B������
|���/��x{�0�I*T���1��� f��y����"��6���y�& �JT��#��2��X��n��+�0;��.��r������-���!�H�Wy&i��ѝbFr[��U�#�>���Y���?l�.���^<p�"����0KZ��>���Ow�(�WW�wG輀��?�����h-3HZ�&�y��4�^2�J���<%�yg2:�iP�tny����S�).��O@�sk��z�������=\��б�njIʾ	���L��
��L���8w`�D����I)_L��C�-i�_�н]�� w7j[5;��N����ף�9��i�|mu�|:��·��~N��M�������VzY����㢭\t�*˂���Oo�Kyf�cjM�e��|��
di���u��V��h�ˎ!�K���-$��k���t�l�ο��ʕ��O}Z����!����}i�3���D��o�[�_]F.������EE�(9�ce�^&��m˩�Vf;d�͝��*rr�b~��y���-�p�*E����7��Z��g�7f�0Sƈ~������o�ܮh��P'k����g����>pEl"Ev_t�1��y��;���^��Iu4*������yX��7���3z�����ɯ��[�~��l/?��N��NJ�6&`+3�6x���q������� X�ׅ�c��(��۞�b@��,9Z�H@�����|$6��G	j����N�'f���q)���B ��.��GÅ#���O<K�mQ��-Ϻ�*�IN4H !�5������$!�(8�U̫j�����gc�"ĥ�D.�R��R#_a�[}���w:Cpzo���
"��_$w�4�`�<A]9{�L$��B-�ÞD"���B��<i)�=Z�+FzT+m�����#1�(� B�I��r;_��8X��x��
����l%�z��1�⼛�t6ߓ��V}������E�5c;?i�M21��a�w��;`Œ�-u�� c.p,Bz��>s������aŚ��e7I��u�:����7�� �y��FE�H1qފ�k{�~���nDc��� �3�����M�Cj�p�'��+A�V~^`,c��Y�w�?A�Ng-qj*����k����ԯ�����aIF5�<�}WkP��ߦ����k�_"�����-v��cB�g�qւ��=Y7A��ğ.�E@��np쭃lK�MT�\��@~��(Nmg荨���[Ӷ~
6>��h��X���@.&W��3u"�ՖQ`՛߹H��k��3:���`uԤr���4���6���9gE��:5�z�B�:*>&�GثRס g�z�x0�N\��U��s&�$E�ǾX���"�Ԣ3�!�X�����v�X�t (���8|,�t�����z��lZ��&����Y����r\��>�?[O�1Yܯ������d�-�{�t��F�,R�����x�[�'�đ���[�"�*�2�Q�)M �/Pg���EN�#V���W=�ˮ'=����㲯nV|1�S���p>3>�P��P~{�;��&?�փTCX^8�H Jǒuˡ����틣�C���y�Ȇޛ .dʅ� f^��
N��d���ĚWC�73��.�-����wx"���ﴡc�ʠk.���X'4�>[5֍Ϭg���Z��忺�E��������HѺQ��2/�����?}��	�0y���-������|�6�I��K_���FY"%�𔡶��OP2�搶�X�qmѮM�͍ �5a\�[V���Z�&,��)C>���H��A�9�	�\�׍y[�����l�o�1��,�d��,�����u6q}�7�wA�oh��? *$�_炤��pvC�â<�3�,2n���ӪZ(�>FWx��M%Q��6�
�rT�Zy���nf�/���T;��9f��퓵���āro)
����3�r��O�l���qwJt���5Ͼ���}�WT��ڋ�R2/�1��ꊇv�G3�wX� �R��s�6bn�
ʾ�gr�ǭORVN ��	��9v庂�>�:v�^�2�(Vi6�i �Ǟ����$�qAƼ��:��`�4�q��6`��5��^��`j������m~_V=S�4v"����'ϡ�&��H�&���Z���]�l��Tj�=�oS�PD�+�ݼ!z��*Oe�i��
�	i�`,����A���|~A"���P�ٴ�'C�@j��Z#p-7��M{ �Ѷ��;_�B����6rd��ه'�"�Ü�5e���X(�nY�F��D��g����C��4��0�w��^Ğr�-1#��y�Yk�b�j�/Ԙ�/��%�v2µ�؝��{_�r�TS��z��0&�a}	�h 1l�I�gx�:�����ӔZ��~h&q��˻n��Q�?W�Z�3�`���nl�Z���^��}`��a�X*c�Ш��PQ�O�A�������.tTs�Pɸ���Έ���w��� ��tsBi��S�0X3q��d��|�N�IWu1v�\+��#� �-w.d�2�����($3Z�%�I���OcmI�ڑr��YDIKwA[h�B�~ۈ��W^�w�^b�9:�L�.�QuZ����lL���rb7?iC�~��N��)W�}0��W2�>5I׬���hx��ź�(�J�q")�>ՙ�0�L�Z7��.~�l~����,�����ԋ�Ane%�Tx���[�y7�A����O[�S�6v��ܣP�o"�?���_,v���=�_X���i�l�%�1�p��B2^�|�qo^��xPZ�]�h�*$��S�`�(b�"\G7��n;���C-����I��G���Ɉ#6��x#���0��b|��jgfE���\p���oi�k����vT7O��4?��{� ]F�J_?�@FQm���af0^��`L:xV��G���y��< 	a�+����q��V�>H�T}i�p(�Vc�6o+�VY07U���/�{ه��ð� ��E�����o��u��,���z"���XTަ��ivM*�R#�F�o=��5��2���R�L 㤷�� U�x�<s.��ЅVcm4�4Σ�sQs��m�H_���e�Lka�d���Zj����P$����&[��`]8��JeAi̮��h���F�wU�tz�<[.m�xU?4}}�I�G��6��8��b�uaM���5$�\Fޜ���䴸[���+��v�\+�̯��F>w�yS�y�e�Q~D��?
��a
��5�(ޖA��6��)'NQ��+3�:�� e� �I<	C��q^��A�p���_v�1���h�!qz@�3�C�,���guP��i��E�cy`y ���}�"k0)�%�Bӯ����m(?b��?������O�L�J�����d�7�I�=n�4g�C�7V� |���QA�����IZ'�R��p�hG���;����o����̛�J�u�4K:�G��*yg�ZH��p��PB1��g�)B�� ��rzlRm��+_��/D겟�ϗ����!d�K�"�@�1Y��ן짇z�KG
��iH�eg���Q�����m�'͎ᑏ���J�ȡ�^ay�.�R�^��?��c�g�B �e31 YA���0�����&[��o����bk[38�IKb.�y���E��J<D���&8 ��5dѤM���G�)�vN�#�i�H.i���$���i�Ck�q���_��gss֚��߳�Fa��b���E3R��F0e�M.��;UFJ5�!�;X>�z�2%�$G��x�g��*�Xf�(�=�ӫS��~K�|x�D��Db�"lu�"���xBي��լ��pKe�q��J�eb�z9�V�	��z��w�pM@�d�_����������'<K�FW��s��w*�`F��8��(���m�M�v���9UG����rR7C3�3�F80[�R�=�J�0�`���X!�|$Nw66��~K
B�0�I�σs2�<wJ�Ʒ��R��c�ܟx\Fb?�T���������DlL�w�`���_]e���*/�#*�c�>A�!)�j��*�b���2c%}��3 ��)Bc���n� -�Uss�P���u#�� �u�(ͳZ8K+_PQ��F80��Zۦp�;3G���d{E��p�!�Ab�E��2"X�b��О�s�{���0��AK>������F���賍v�H�{p��r�Ij.�Mǩ7r2ʥ:f�.�aig���@IgMM	@���y����Z��D��
/*�s�oA�7�1f���`j�Qe�H���FC�o�K�����}?�-v��7�"FX�-��e�UEZ�%�N~�Z�+��V��PA�z?��i��N��px�����Q��6��w��3��"��B?��i��e5Z뼏�ApW�sH{�?j�e��q�@�n{}���l��1٭�^����=I��K0��:���,��`,-�2P�Q��L�i��+��{�I�7W��T�y�2����RR�X(-Q ��Hkxx�_ Omv\rV64�����0��t��
�����I	�Y( sy�)F�-��aG���1�S�9`��+U#0�->��	����~{/T�|�G��:��R�_���M�ZMJ����gj��pP�c���5�������9Bn�\C/�s�0z}�q�L�T�9̳�GY������΄\���a�p?�����g�1�\䏔!q�_K����\�/4&���Q�����2�J�Rb��8�n���	|#K)�I7=��S0����h�b�34�ؘ�T��~�m��3�+|��<������S���ɼ���n��9~�Gg���.����甲	b��[-���f���G���˵���+����n�ɂ"����F�c{�(�+��Yv��n��|Tp���G�[&,}���*��ܭ���M?�JR�r�w����8>�/�v(����Q���J��k�`$|�м�H
ks1�B�� 3gr��10K�o֭$@�㜠OP%���}�iɳ�lY�/�Wm�3WtޭEfVY��]���W��M�YX+a1��l�?X㡚8�>S#>omDL+,���P+? b�(v*]y�E��O�q�(�#)�s0��)�A��~��H�<�QJ|z�,�C:O���(Jx~ٮ��:�Ork:!J!h��Р`}g,V8����O�����.T����f�3c\���V���&�}�o�����d
ԭ4˟�,�e}޻)oty�S���(�7�^�6kA�>'�YD��c�t't`���k� �P	�J��Z�r�v!'�H����;kV��:lO��.��* 8�:��T�HG��1����
���Z�/�q�FS
i:H��^�p	a�f�ݛ�Eq��w�E�a��߉�O)W,�C:��6G)N񷂬8���A~E]��k~��vT�GI�M[/=-���� c�ϊ��$����oК�O���)��A-\qL9^�͛��!�ⵠ%m%�Ok~�-�a�����i�x����`�qzN�5ՌV�E�	�0��='q-�ï[V���)�����V&Q�A/��Aц�'z����, ���'9 �FL�&B�o�{�O��^���:�#�����*�1�2H�%C�a=�Rķ{s.�ғ��{]�Ĥ'~Eh�I��{���o��=)�Y� �S�����7������H��>]��H�N��Er�t��|Y+t�^^5K�Ŕ�WG<p�
�w�/�q.��J�����/G��ٛݳ��n�QE�]��DR��HW~Ff�iylBɐ2 ��V��%�E_� �nm�O��~y`x��yk�HJ�u�ѝV<���/֔S�m�s����J�KG��c����^��X�ȯEnB+�[g�������K��n5âvA8�"��ԕ�� �&�Ȉ��t����������V���2��g���3$Y��q6���"�`|̶QŮ2�~���R:�ɴ/^�zٟ���B�6�C�:��ح�QB4���P4m�I�i�m���0�	ųۭ��n`6E3�:��$`g)?U��:�q{'N>f{���*��1�0����_(*�S)$z�jd�B(4�k�v��` �<2��.*������hP�];�����R0�:��y4\_�94o�{̷����Q����}Q�6sW���M��d��i ���}" #9�'�`�P~:�|g1ųK���C��D��}����]�u$<E��`��&V�!�nt���J\���&�o�F�<�E�J�aG(��K7�� �⴯}c7`��D��hWu�S�(- DA��g�h9׿O-�Ij;��09�\\�S�u�lY���G���Oʈ����EТυT�'m0�����o�&�cГ��������F?��$��Ѩ�P�CDH8����|"}���w����B�����Ѹ\g�k!�.l�u����؃O�	��
N�X!�`���qz�_�7B7��w΅������ē��D%�wd;Ѵ�9�\�ꞈr1�/���q3z�P�1s������2�[:ط�x��L������:E�V�=�O�o�5��Ă�%��ÝQ��#Q�C8B>��
ʭ�p���c��Օ�R�.�=�8��y�ԑ��Z��]�S%��+Z�c����`�U������������f�9��/����ˁ�Ms�Η�Z�
~!+`���^'�j@�N�p�si"�y��k(Ub�>=1���`��1�A^[���L3iV]?m�>�ÛRq���7U�5y�R_��|6��d�3~V����u�y�-���~���\�T�yĆ�����\VB�(��Zqo�U�]I�.[1�S�t�e-�kQP�Z�ZgM�s�?�Z*"Ô�<��Ut��PYIe�?�C�u#��8c��ۅ��vsR�C��������}��E_�� �Y	c�hV/��'�8kY�m��4���h�l�'��]��ւ���E�i��:o�8i��9��N��%`u%�rc`A��S1�0:6�)7 U;n�v�^[ �9Z�FNq��B���VXf�4��Ī�f/w��V[��Yx�{@��x��_od����p�be��=��9.�>^P��U��[X�?C���, Jar�}��p�w�?j���Y�U�j���q�3W�܎������d�-e��;��v�2����F���6L�]���x�'�W�3&k��I�a�u�7M�Y�k����}M��KEbM'�hq���P䪵ju��^t��N��nz��}�a�`�b�[�O�������E�ծ:���UQ��Ђ��~�G����r�:�R5M�x�j�*WP1�7; �4�E1�@�W=���&�-BI֋T���R��F���s��e8��L{D9#�Pm�61t�2�(>_p%�ܑ�շp���sg	ԑ�H�"����'$G����|$��s��s��=��C���a�c>��YN��hY�8q`S�;�i��հ��9eo���+��P� �Ʃ�������(lpg�8XMb����@RrYy��Q��M��k �7�u�8!��f�����$͢�6_U-k�� ��\UR�E�i���m�zơ� Ma1��\}f�ab�4�ST�{����~����C��:��B+���x����-����W��bj�B����ڿg6��{��-���$R�imaj�{}�D�A_6������`f����%�]DE7zO�P#FsF1l>��ka�AC�C��T	'��A��uZ�|}T��D
0����kS[麂��[������>��N��c�o{Ġ���ޚY��/l�$�Al��1}�R �eOfXA2��� fy�X���v��I�\n�#�D�5x�bg=�B!S�n��C|�'#HO�: �2;��9�W2,
���"mB����oH��>:�r(hP�D���2�c��U�� Q��, ���S}Ou��c$:�[z�V���\���r�9�Q2;�|�*��d�sY	r$�����e��W�L��T!bkl+-�=O�j�$B����؈l㆖��U�:�Y��U��θ�4'��R6A	���>	b��A�H�Q�Fl+6�#H�*�|7~�-Y�^��'��]����;( �{y��RJ�?w�4\���&@0���K��M�Β���ɀP�J�*E׶=H�$E����&��8n���Ǣx�i����φ���N�4���Y�A(�gp:Y3| s_ɫ���/ȥ7��k1�K�2_�n��],�'�FbXH2@_u��:<��9qQ:��s���X=��o^�������\���SR*�j}��j�o�'S��6��,�	õ=q�"��"����%���&BѤ��P�3�  8n��LQ�0�e|���%�s��9 ���s�Ŷ�<7`1/sǭe�.� S��& �Hc-��c���^�$�G��w�S��� 9�h�?0�N���q���T�����7]4�a-/�T2��8������
������3�E5;,]`hY�hvbMZ+���F8�
rY�F��%8���y
����^=��&��c;�7������� x�>�Mt��	3�]'*�\F�����z��r�ʰ^��;�nE���A5�b�����@����k�s=��Ӫ����ݱ��2]�u�@2��hy '�n�C���骃Z������b���x����|Ƕ�_��F��j��L��U�R$X����o�"�/�q%+�����R�B
���,/$�#C�"j/�R'P]�����G�&���tЯ��t����˿�s�nD����7����:oS��rA�<�g�=����,�f���8�Ж��1�s����2�>oE&��q��`�fU������k^�]PyuٕV�Cl�B��
B�^�k�Ғ���PQ$�zr��u� ��=�a�����8�t����f��=��v�Tg(��@�7RP�~��������R�v��֝>�Z���R��$'C��m�g�#e�ӡ�4B�u�ʹ��-Z�T��V������i��~t���� Q|�0Ƴ�l�Y!��"�4\���^>1y����1�#tޞ��W��Q���� ʈoV��b�>�[Q�tT�U�!���掐�öe/ �W�o\��:yV���pZ���1.+�K7���V]*��e}$�ͺ�e`;!��]��	K��h�=�c��_�{��U*�6��x��c���|��K�����/�Ǘ(�&��$�5�Nw����� ���ep:G�5+�6"J�Ђ�NT���Đ��M�](%�������OwV=h����?ߊ�[C���N�C6�grX��8h8q�u/a���1L�gp�1��z�����Q��M9��p�:�Pmt�Re�����\�k�Jr���RlS��<)h��>���]%�ˢ�kb཈(���ko]՘�Qx
8 ItP�#L��~��Oz4�F�r��AbO��[Z���+~�=m��le��tU#~q�)��j6�����������rܵ��s����!<��������̲�&����
>�;c��`���*�M[�!Q�H^���/ۑ͵��T³{��l���Ni�4�ۿZ�]߁X�e� ʑ���&�:����4�?t�)�I*A�U�%L��Z露3O��:�������-�"f]YY��z����X6�^�V��`��s�Xx���h�TF���H,V�������91����M\1ne�6�#犽�
�&c���l�!�n֯l^}&��8�Y1�y��V�����J� ��2�=���'_�VNQŐ��B}=鋎�Hŏ� d'R#�y�иVJ N}��UhD���{/�^~���0-�F�ONM��/Tj���	��]��?�d��e�D]����7�4ۊfs�>Ʉ#�I)����Tt�9�ȉ*�����k"�p�Ί�HN�شēߑu0��<��n�坢��)�D�N���i%�W� ^�2�lc������Jb�cGX�A�s��Ʌ8)��0�V�Z��w�>�O���	fe'�$����[�X̬S���"��>����F�����c��o��v&OJ/��7#JnGZ���w���v;D�!D��$������y��UZ���A+�nT�1;�|��ӑ��Ț��0U�;/�M����r|�� ��c�g�̀u0θ������d����i����6��֥C"F���
�y�Ȓ�Yϭzp�B���Ų��\p���d3��Q��6����.W���dq̳��� *<�pzLf:����tX5���r��?�n[a�U�&�:���d�}/.5�l�ѐ��#uթ{��~_�m��ku��8|Er��$<9�c6�whZ����9�[g$Nɒ��k�����/�Ƌg���q[���P�3V`�7��H�Iܟ	e��� x�T��@�B�,9b��)*��.	� g0�*"ۂdljQI���7��!�4��JCaP�&��˥ʄ��z��*���A��\y�܊����')	��v�$;=�:��Dn������ �7�?j��=aX��4��9k������>��~=Y9��؉C!$ٗ:��kL&]f����C�ҋ���@ߌ���z�XB� �Ug�5O<Gd���E�K��s!�̈���?ֽ�AõA���_�⪡|�3��R{xዡ����6q������>ޔ-��&iF}"��a-iJ?v忘�c8���[)�!;fl��㞦*�c� pG���+bE~3]�p�kÏ��Q�!Z%a��t9(�r�,-o�uk'�{�?
�����O)�*a]º��dӣz2��k���r�J`�bf7\�Rb!k��a�A�G�j`Q�Փ!��qk�$A`O��!��.ӂhdwKB����E!FQ��R�Ԗ�%�sɦI��0�
���pz>l�j)OV�hJgH��bu��eBW����~Y��֨ה�f�S�(o�Jd얳ۚ���G/�/k������$]߿i�/�΀�ӿJY�|��Gr*��ƴ�u��
�ц�a�>]o��-��I�vbXO���GUA7�q��d��`��:�x��*�L��AX������3��ʈݙ� ���hA�Ҙ���W/��Ec�]�5V��!�
��_����E��v�'#��[~��p�Ω}��vQ2T%�dk�uq8/��w���Ke���-{�[ϠDS���> �.'q8��_�X��RL^<��u��_���]�۹%�v�������<�_N� �Jjr�K!Ռc+)�!�����#-6�,b>���^Q���Qb�TB�#XI"�-�'>n���j����t_$�?�6+�Db�5=j�`fQ�▙i,����yXT��G�XF(5Z�{�o�J��?��T���b��y�j�L_��8w�5h{��$=���\��<��/1z:�@����5NR�a�ī^Rw�GZñ)?$�aJF�j:M����#O��˲ʡ��ў���<���]�vGE�l�p���v�1j�Qg&�R*X�E:��E�D��0�Ye�/�>��'�:���Ʌ�ϯ��oGT��`� f������K�`{B��bl=%P��X���_ܶ���C��|FYE���d��A^	i���邸
q<j�t.��A6��[W��G2΂k�tA��`�&ںi^���FRڌRa{[�}x]Ѻ�kjK��*�u"ېU<�]���A���=絠�-�9X����P���h�<�H�g�j9@�<�?���X���l��/^�w�fh�~I����3ӹ���{�Dۓ-�N�:@Z;�}��'�t�A��<I2j5D�F��n�6��EU�1V��fn�)��H����\���W��ꀹ��T/9r�U=go?��|[�+]+��b��*��W<�n�M�-M���te"Cy�cl���kٳ��
�܅&�8�)G]x�.&��h�˽Ę�e�Sĝ	�h`Y���ٌ���.�����ƲT�&��&���*��c��qu0�ǉR�sC0��D��Z�yY�~�r���hVJ�',�[`x��aj�ݿ
��H��g|�(����.uZ~_Bo�*�sB��p�Nti�Τ<ڃ��qw?c�+��詫�����X
tj@>�]�͹2w;"�Uo#3 a��8��:�h�k'L��3��ݿ&����,��c�׽�Mh����\ϳ���[���% �5�A�`edt�% K������gֶ�6�j�s�1x6�f̳�����v��u��@E��r
�5`�a�ȧ�=�K�>�͸��";#����*x3����	h��� D2��ֱ5��BJm�'9�6�~�bcŁe,o��:_�%S(��{6�>K	�Pf&!;�Ҩ�iX�A#yJ�x���.>��)�����Zx11�o��c�R���ta��YHϵ�л3%ea'�UZT��Em ��E�*��:�s��>֧��|��DYO�6���s�}�s>��}Dj��qk�?������#�O��V@~I���q�QClj�����׍�8��*t֝&�O���.B�A��v�̳��u� ۆ*��/B�bz��A�� 
a#z��;�����?2���w"@˽��n�u��]\n� 8=k`����QH�V^�@^���P�o�����`]�e�ʦ�H[Q���ϰ�~n����¯0�w��»��_!�+V�'=K.wH7&�="��
ʇ�2hE���F�j�����m�֗?H� ��ufo���V��
MT�fL	[�X��R�1��&}%�LJ�x�Va������sףXx�88�O)��p��䋎���'�:ZVNU%�M�rN��ֱ^�c�埭}�Lz��vb@�z�^���k�������Y���A����fs����E���%�x��0�R��Nʠ�T����7Q78����u/�a��
u�4�$�΀uX�	�o&j"��L���T
�ԬL�⋍���,S�Z6�@.py%蝅���P�H���^���K��5��=�ۖb�B��!�R*�c���$��>�B:.۵ٵڪQ[k'�iAP�rs6�@:�u3cr&7�n���_WQ�~�J�$!�U����g
��f5�h��g2Zpi*�l�}#�㬻�j�����A��� a�ۤ�g$r��,d,��JwA"RټP/p�m���N�xH�o�o��.��|Yq,��^ ]��kG�ߥ[S��{+����&V�:�Hx�����|@kƐ9|� R��ʟJZ�%����6� C������d�����Nm�_�E�69�To��?Q#�
Q]�!�p����	�{��R։�8V�c�-J|��R�CL}W����۾���7p��,C)  S2�12�E�� ��	��w�ds�4~��4$�nb��#�7_D�M����ٛt}!���(/N9ez�lID���*g�?pTWϲ���6Ѹ��e����#��;"���p`h�V|� ����+�1�Ǝd�`��t{��#&��é̊rђN�7��͋'�G�@>ұ���e4����x��`�C��s�j�t~pV`9'�z3�@�ӎ>K|����������<�y�U����О�kX����l��q�hD;.�΄z�U�%ޒ��(�h0�o뛐�C������cIrF)Q(w�:�(�Y=1�}�$���Bqy�ܽ�0�f�_.בj�;Ç�eY?���k�~)��29_qFK�<�����T�����qp����o�6k���?i�F�v�����)?6b��3��{�����-/�i֚�V�@7�F�g�fl6����P/�~���}S����O�d[ӧ:Go�����7�W�H�p]���4�Bf�i7����ԍ7�bܭ��Ӗ;�Ux.����#%q;S�R�Y/���귫H'�=���m��B/�B��|[���>�L��Qf��h�ؓ��'�X@�o~�g�إ�dЮ1������^]���d�f���8_�+����c��"p¿~��Qf�Q�T�h�/tgť����pA pf�ݮ���Ve�ׯ�i��F�X�pPi;�=2�$��k�vb֫yR\��]��noگ�ecI�C�Rz!�ej\�y�xO8r?�@��ЊU ��c���N��@�3�4���%�+�%��ܖ��P����k ��5`�k�/��S�7{�5��Wy_
��t� ��[��>U~��Mz����G�5���� wx�o�D+�)d��ɓ�w@�1��"Ƒ�s�j�����>N`������1�/3�ړWc¥�7���_����D^T�<���H�:����q���2j�L�

�;���Oᘩ�Y�)g�0j)�9+�\�`&c}�k�	I��ס1�����H��]ݐ��E^�)!�P-�6���#��Y��?WKc��!L���WJ\�屽?Y�j��7�F�O#̓���y`R�|5�|[��/�"�es��� �g�'.���Dغ%B�����Z8q�5� %��!���2�^9]v)=T8'�FC��N�:�hU=5���-���h�eh�=��ófe����N}o�!��j*�����M�6v37�%�a	8N��~��7�:9	g���0<d�N�q�(ue(l�8�4�3�G�[3�ZBLl&�>�q��an����r���Kj��!�{��s�sf�n�L!���q���n�Zޑ^�֣w>q �i�RD: �c��Ԣ�a*T/��d)*�\d�N/�zD)�5�t�����j�[.�*۟�$+e)ء+݆ ���_�W�Z��l�G��dH,lX=�*T%���'hYl��륦n*s>摮��FZhus���{#0� ����~9��1P��>��x��@ �,��m���O�"u��3�Q֎F>��k��(���
w�K��� Q,���U��U��	�g���y5U��d��5x�0d��sBf��|S�*2
�j?)��������.w���T�7�W�����8��Ո����H�#x>_��0���I@G�*Ӹ�h�`����U�W�2�e&뻥/F�-e���� ���,��]��4*+�=4��j����xD/ܽg��Xr�L]��T8R
�=��5?��DyH��h��@����u1V��u^Y���=DQ�!�������
T�"R����Ӏ�d��s�(��J[-�qވI�;+�*U�C.�/گ�t-_��X(����1WN�'h����G�D^�BW��])ޭW�#-�I�<w�r#��<f����2�s��N�v`�~'{���|���w��]�k-|�&c��J�������Қ ���'��n���䞠)���U�n����$�|�g{�ؕ���t��9E�'k6��uv)9�U�v�P�޾�����Fݟ�v�B���Q>�=Ԥ8S�����7r�,�>�y��)U��U?����<e��B���K���ܧz��p;Ч�Q�������� J.�Nok��Ƈ�F׋�d��KwS�̺ZF�ƿq�,..O�=L��zUGV�T}x�0oy:�	�u��\/��v`�'��,?��s<O�u%]ÒAZ�o���e�2��5M��+�Ot��"IT\�7.&�� Lm+U`>zkT�$�}�e�K�]
3�5�0��8��l���!�,AW}jӘP��2$`{y�K��.��!<�q�����&��\��Ơ\����� eN�7��
������<N��Zd����/f,jq/^�m�%��xplB�
�bu�2[;@���4�_M9ј��lF�c�ii���c���������;������^�D�D��oi���)�������o}������7�2�=uea¤X�t����D�1�B�	�Ag�s���4@w����+���E�Q����f�����.?j%f�t:4r�Y���|o�s��'�1FD@$C���<�����U2u=\�ä��ø@��n!g4�[ �u�:����PF�N/����5������_����.K˯��W����YY�3�UlŮ���qw�aF��m�ۤ|�98�p��f0��st{�/��˻fB$�N8g���q�n��q{I��(���,SN�f'у�m�G^g	+�s�h�����.X�����Z��Z�b���y���uB�H�^Mw��XI�7ˆ 
�` V���kjq�C?e���܍^�IX��,�A&o����B��\5G�ζV��E#�Q�Շ���W�o(cV3����D���x��Iu��a�7ip�zH68�Gq�E��Z�q}"θ"�� ��$i0�sG;Em�X��V�*}��7C�	B�&cbt���Ry����v��w��z�mB�K��x��I��_��g��B8�m3LǏ��ߧD'DߍNX���V�Ee�V�oݪ����Ҷ]m������6�"E����SP��1�k&��y"���s h5S��������WB�v���3����'T������ʻR�`\�L~�U�a�f;�w?�cRo�����W�I2���c�����6�XC(��V2���i�C��c׃�p�2|ڙZ�2PL!89�t���J��	Lb���ު�k��8��2.y�4��K����
��jl�f���dK�EaƦ 7u`��t���h�}�f��_��mm���L^/Z-�0���'�a�N�yZN$n�;����b÷��v��ӀӤ��H='�nѭ���ϓH��/�Q�QB��WbR����_���$�0YV#��j���8��Mװ����3T� ϣ������l��n��N�p���r���Wp++�Öȏ���3i�B	�<�n���De�H�z�&\gS�L_ݻISY�ۘMW�Ė� ?$��bɿ���fd��A��� ���f�\�g��P�*`��%+^6P8�o���3^���z��g�{@͝�42��h�{���a�A)��Z ��e�]�-�}BҼ��u�)���>
�#.�\�lsXY�2_٢�v���?J4������?Ǵ�`G>km7�{De\�*њ5�ٍ���$�6@���ۖ Y����Ru���V��GE<��d���.L�"��*�+X��+����*R��T{��T��.U�|�Q*�3$>6t��ԄT�nC��C��l^��|5���yA��ݝ3%��ٻ
ۿӕN��R�ũ*L�ƭF�S-�{{'��)Ff#[^�L�G%����u�x�B�n��|q����m��� �t�@烋�8�����̻n9���?N8����Vʐ8��
v0�6anY��HC�w��:U�?�]�h%�$k�*V�tMF��4����E���Q?����/�mv�<%�_-�H����o�i}�Fm!�����f&%�z`�1��ck]�*�@Rܦ�`��g�f<D�}���&�dc��e�y �<ZzN�Y����U�gm�-��nn��o�2��Ғ�I��Q�hdL�<�/=,�$rUc��G���X^
��|��,��i��f����a��(�{P�k|�T	f��(�!O⢚�8�C~��2��`fʥ���~����F�z���T��+Y9=�]�AwJ��%�Aݧ�Ћcƒ�ޞ�=*��R:H��!�ZtW�5�R���Є�s���^�����MJ[�t���S9�������7���E`C�� �6R���*|FU�əu�:�������U��&鵤A��� ��!p�s��l�8�J�V��@�5Uj��fB��$���GËq����4��P�'��-���d��0�9ޢ�.0Xt��}���_�t���`rG�W�T��1%~B�-zq��@��<3d��8mNO�Q.K��]�,�tc��̑��Z�[����Z��U����w&ܵ�-�-0�F5��(���L�9�XML!����ɄY+���B����h&oބ������*(���m������kP�nZ_��K9��A�}�+������@�f��ҽ}�|7��Gi�ՠ���눘|D����1���o��}���8O��SC������A��5�����/�qJ$o�"�+&�nD2-1��J�	z.�*�}�~Yu|��0a�ũ��9��oe�͈��v��/�|�h(��7ǻr��S�r���ga�2�)���?'n���Ak�	��d/'+�o��k�r�sY��6*�e��3g�" т.�=��J�� Ā���"/>ѓD����S��tg{��[��>b�aF��^��U�7ժO���aB"���: ��ٹ��Y�/���mμ�	��"��'a[�ݖQ���~9�-��'4�6&�xř�wLL�U���#��we/���a��T��O������ ��>n���]�0��5�O�T�*`XnY7)c�tik�%{I�4�u�Y�s8A�s��V"^L�ԙ�XOL�_�sݵ �]�Ĵ�W���aM�@�Q:�a��EW��Y6>�<� �)�Ta*��п#m�ȏ�6�G;�X\6?�h��&0N�Hs�M�ɻ��Hi��Mګ��a���	k�����sm.2-\Jx�=[v�=��nc&�/��~�U�@XP��˼��/�h�����	��^���6�[���uD0���NDn��=Õ�Ĕ��kT%9�X�m�ɥ<��b_{,|�WO)l���b�X�Q��?޵�6,n��b����*痪H�8�\� ��h!k�փA~3	�@+���km=���PC��U��jQN��(�Q�3�Y�Ӭs�ыt\&w�&;���댿�6-�.%ɚ�ѓ����Z�v-�������x�r���+����v���o*��T�;w��J�K�*�6���u���( d���� ~5����o�C�gz& Yzw��?�U��oY��8��_�rBZxOoFt�u��6*���."��]������%M�;�*琰�BR"A�kT�;�T�4E�j ����"��-ׄ��H��B-M
ۏ�.5?�yг�{8��w��r��Y�^qBB�my��ԡ��R"���胤�Z��)��q����&S.�����~XՏ[c�ҮF}��yWo��mԺ�L��=x S��#���V����h�w�U��SFA$GQ'X �U���}0g�BUΦ���O\�)����x�`���I�t������;|G�a�.�p��w����MI�T�+�1��4�	5��yq'v��'>v�^:��LcuGAz`!�\i�y�|4Jئ(��}k��hʉ�J����H*ɫ�p�zE�6e/�^�{SK�FC?����MN�z���u U��z��G7��F������A^���q��c�K������{N�?��2���G=����!]A>S���� �ʏ�8O�\M|`[�.�&�ٸZ�/�P�l��7��E����S�;��8[@��	z�xg��p���;Z�K�W�v����F�MF��4:�aF*p<�a���wG#��;�߯(\�i�<����fTЄ�+�SO$��S�I��0Z�F-|_�4W�lP��3�\v^ܘi�#��>j����Ui}��h���tV�Eh�Q[J�?lp�K����Tw M��3�f$�OK�*{��^	ĺ��`���Y��1 �.��v<�V^g����bE��'k��M*��8��Aڮ��)?3���2K����%��`����8�/E�g�2����6��[3υ+[Q?[�.�~+��M����S��H?� I��w|A0`� U)�����7D��8��7�4"�䌤jd�C���]1��K*W���lK���32���~8N?RHf��d�K[we��_�Z|�`��N���i�P�3�Ⱥ�c)�2~˳"a�-�U�����M�$��������xĮf�Ywxx 7?ռ܈%;n�(}E*]U��OA �A�\�A
1v
�:=o�m�L�
�6�| �M9��0JV��Ggê�~�&������7���2�ă��;q�Y%�ݘ��T�xy����ƔXϱ�{����l��M�U��;�,R{O��D���|�K|H�Zs��H��*�$q��,)yj��	,@Ɂ�p����~��My&$m=��L�n��y	��:��� ����[����D_��nbQes�S7$�e4^�~��~� ��W�7J�?����]���M�7Y�[Q�|��j�;+W -��� ;�������#"0��J�Cj�������-Z��\ӿ	������bf9K"��}��>UkAZ����!�hu_�rT��%�+��Cay�{��n����\N�Y��ߎ�P�E
��og`��Bǆ��k��M�r�2�������v-HI��x�scT�S���]'����P�-��t����ky�Nk&���j��t�fW�u��}C�R�DL㣸* ����L����~�L���V�#���������@��z��
g�K�Q���-6�9oo���,ل���\w��C���\�1��{�� ��A4e��2���w<d.�Y�����a���b���˼u��%�$�m�KO�ė\�SLڬ9���O�j��9�?���2��vQj�Ӌ#ˬ'}�)�Ǐ7�q�#�6xq�/2l��mj�χ��n�	dYpA�ݧ�&O���B[�uû�ډ��hx)l����&ޗ$���R}�?�bx�ozp�ڨ�H�}�k�Qt�u�N�c�^5���4&
��Y�����������x��f�J\ �xH��B�fFl�7� V�1;�]K�E?�&�=dW� ���q�EX �&2X����Į�y�����=qn+=�+f��1��е�"po�Wᜮ���w�:�G$|���g����@|���*0t���o�1�e�������E�s�`,
�[������a�Rcv���<�E7	��sM/���5
 V��3`���@����Q?�tjG2Q��o��������~n�R��ś��*� s5����n��v.�% ��+���Ś������,,���r*�a.��\w�5�d_]G䜳�`���o���8YU��E��^�1t7lx�HN����>�S��R���ƾ��z��xh��th��pi�e%]��oNf�
x�� �{��_w��v���)��ň˗�,�	��tn���b����%��2�O81Z��`z���w��?jU�����Q'[�0я���N���b�5li���Z6r�G�V�I׭���#��T�
�wf����5�TE��C���� ]�8q���v+��3G��r,%}lh�~��2�]�NIɪ�bۻqAoA�t�9�L��02�^�wC�݌��80��'��8�Z�wtT��L7)[D��{��|��L�A'�/+�q�8�:ģ�#Чve���y�G�cכp�����΀t��B�of2�N���Y�9�>�ʸ���H��V��uX%3/��<4�����HVJ�[G�F(x��NC7�Cܸ<E.k�;�0���(e|�%-��Lm7����	]��"�W�fB���:�H��}E7�������"��i�o�%ֱ6_��j��i�)��,�8�׆"~�r�K����ݶ!�%�v5A%�$˴�4�{���Jo��v;�r�9�z��fY@���6Tƹ#uE�#{e$��:!��^��J��&@���{{9�D�����N(��zV.�x:d��^G��N��1�EXD��.�r�h�ȇ|c�G�u�6^A�S� Ϥl�%�ˬb�,$��߅5�_�"���cdqS�����@a�S��e�W�\�6dU�Hs�.� 2�wM�Q�Ҧ�D���7��BC�ͽ3ԴJ!_= ���ԗ���t��]B��������V�cً�F���ʴVgg�L�"�ϳ밾4����q�?ډ�8��*"P�vg���9����R�TI¼��k��+���T:��Е��i��	��HR���y��%���_�N��"z�G#qH���������^����[D��׉ �M��	�КPM�A� ���22�pի�_W�^E�T�[��l��eY=�"4D�g��
��iÄ�I�el��_�C+i(�������Y/��*#�ए���x�=x����#�Ⱥ �����zz~Q��B��1�&��rN"�c���3Cf�8Ϟm�a@���|.!u�v9?ﴫ��\����捾��M��$:e��^>(0�?�I����ܓ1=7B�S���R$�O �y�evG����i>���`�' ��7�:�Z^ǯ�# �Jv��'Q�"�fb�`��˫7Pt*�nq����w�0�!�,�S��;�����c��&m1FD�D)���7��)���z�-q6�����{���@j��VWa�L�ڝ�Z��1���R�5�_H`�R�P�_4y����,v)Z�Û�I^��/0�pI$_h�ȸԧe��)W�+���]0/���AЪ���R� B�
�	3j����KB�M>R���Ẋ��R�i���MH�%���(0
i��R�Qwjg��"c����.��ؽ0�s�2����q��Q�a�8X�y*��Ѷ_`�@6���G�hh^	����G��z��b���fnXN��_�C���/s�D[����(Gs i?�'h�̦}�`c݈�#��im�w<������'�B�e5�xA�(}��M	
V����~V�f�]�*8�i~����u=F��N"-���³������[ߪm.�? � )�L%�1L�=���م���r�^��g��|r�f��SvY���[�.TW�s����FpY\�3w��%%L�3o�}-<���(����M"R/�'�]"��J�o��\��Ja�T�S�)pb���ϰ&(���mӱj������I�~���2o,�k.Y�}_>BT��E���&U�e�A0�%���:酓��N�h��[���\H8F��&�9���b��ݟ	z]��NE}����đ=����#�Y��-�
/!�������F�f@��x�麶�҆�x���Ƀ	��)Q��m0�0e xZ�P^eI��ل^g/dZ���%�3a�m\��-��;D��[-J��'�B��;� �A�Nc��o�'�	qS�]�?�hZ�w�)���5`!Xz���k���R�}��p<�Y���H����JT�	��!7Η_Ix˝�|�[����ZXBSQ��Tm�sᾫhȪ
�Z�~
n�-�����a'.���� J�*���@��b�,�,������t؏9���V�?��/�~5�6������[T����x{I���h�?.��Bvpƻ�
���	6��$��6���0��x��j$D�G� �|!z�A�Z7}�?�L�vU��}�V$�u�B6�V��j����}�_(j�X��*%��I�ѰZ�<��:�N~�;ӵ�0�4����`�Q'��3��Y�Oo��5���P��cj�c������6��p���p�t;Q��X���u�U�Rw��\#�j��u���)͚�!fA7�<D���L�a��k��5'}{�9M����l�b��z��M��/Qu��`�~m<0VO�Uk�&���.��r4�iY?�JV�]+����� �p`�դ*�`�����|]u`fVnr[QqX�F�K�ӿ\��W�C~����BN��ح}�X/�"eU�����E�I1A�Eo�=��nB�9nk���&��z{g�	���!�&�!-X���=�t8���9�aY�AO��r�`8u-�KI��t����//�S!�cY(��+߶���*�E��7��U�>�z���Z�f�̘�q��ȗD×o��Jt}�V[�#���T$2o���0�t%�����tgg�!��o��P�U�N�Һ�g
�;�Zw�5��"��}��}Ѐ�.��ky��I�.����?��)��6�+�d$�E$�˥�0B?��{8ètW!(#�Ntvmy��sd��q�j�+�C� "��I` .9^|Q����@A\��O�v���4��zJ�]#�Vm` χ�UV��U�<���*@6E�8���}ܪ�gaҟj� ���^\��QQ����:�=�py�GN~4j��m�'���Q�づ�}��ɪ[���6����6d 6�J�gֽ����C-#��߸z�T�(Yô��5oAa-ly)D&��4��g�M��7K�E��w�@;���b8�]���o+K&�U�J*�m^���;��	���KU�~V���00I�">�57֜xH��Ն>��K� �w�(JNM��$�|T��ù�TE���$�~T��S��N�B��WC�_���$g�:����(�]�0<�D���B�e���%��{w2�1�y�'�T�ԍR��&��H<�����(��(���k��S�fB��e�R��p;}-fSҀ�ArG�] �d������h�C�Mm��ҫ9�:�8��e6g���;$P<���g|��|��%q-{Խ��lgn���hN�P��Q��=Q1S
�.*zb��C'Wc4��f���p� б=��i�����B 5o��u�l��	E�d&�ʃI�)���'���7��h5���W`��%\�t�g�� ��<x�s�)��9GB9���a�6�b���Nga) Ee�0"�\�p��h�N2�2��yclY�Ԉ���Fϱ�}5�A�*91�;a�0M��2�僉,(p�
p��^��t����dە�=����:��nD���[������킋�7T��v�m[��@�e��0�
���n�'�>�~��_\T� ��7����pɤ܇��.Nq'\���F�,��*~3w�*�����\�kꂙ�Dy��k$fM�L���,���1�A�cYsJ������jM�4��T���%����*��C'��hz�<�Z[�p����'�����JR�����	r�:�Sb��mx)���YM�)�F���8F�ľJ��+��(��7�'�Q�MeB�����g0�QC���>wy�9���?�H���ܾ[vru4
y�+�� c��~�O&�zfF|�Άg�b�a�]<7�o�J|(�_Zo�)k�U���U~��4=��0�#�2�+~E�@��|�y,�a�n�T z��-��B��Ũ9���D��SƜ�W+���y�`7��Q~��R�$�l5M ��l�s[�Dޜ��9����tE���1J�oX�HN�G«=�ˢ��u�)l�zL�� �o�J[�c�~~�E����갿���Z��N��H��~��-]��1�{�Ԅ��f��I�©��$��ct��Yr�o�u<�����V+�)l��!Z�w'f1������>Q����B1.#�ItzF����x�Ӯ?	<���c3x����{yH��kt���a�tX�<`�?�c�@g$�pH�y��,�<��
�#�q�אWGY���X~�s�	����QG����({�w�[�;��/i�J�8�l�9)�e
����t�z����� �'0�I8��β��W���@�y��Okդ�������p�N��w���Wߘ ؉�6=���	��Y��t�xJu'r��[U��e5��!�Lk�i��9@�U�L�U'��{��\�)ԅU���=[�P�L$'��߀}��Mi/>��>�і�9��=�X�����e�{���ϒM��y�;���+���
w?�W�+��}�J<Ѷ�n|�`�A��K���p�E�c�v�n3�Q�bƇ>���`G��|Z�{�y�W��w�4�(����?"�7����_��*?�5P�[��y&��gr�m:u&&+pb���'t���,�9����$��ͥ�T�e&u[娰����!��(!�\UL=�'�jË�FU�D&��.����:%r��.���=eA�BȞ�5$\�C�MKŕ6O4���驡�އ���,3��e_�>�[pI9�O�n�n��Q㩕i���@��@s	�a&�ޢ�k�f̻�==�Q�;�ͦ�-����z�%�{�{�2d*��4��f���#�����2"ag�����*K�c��Ќ�JÝ��H���B1q?�(�L����,>�c:�/�߄l�0XW-����F<Ã�Co����v7��2�U3�G�/4�5�z�t��g78��CmAˡ��4�.�+���0u�G�����#&�`;�1jK��I�"yٻլ�ܐ�<�.�<�`�zٗx�g��;bW����E�����i�� �͚ݎix���SҒ�~p��P�16�s�Z����Z�&���l�~����F�H$�H�#]�f�4����=�w����Q.e�}��q�	g�`�T�c�}�I��bY�ϊD_�B�,�J&1!Z����۬֥/˲�yQ��YKe�M=��L�~291�������ZJ"�{�,�C�2���Z ����0#`���Ɠ-�)F��B�n�\�~����sp�j�19LBZy{K��D5:�%4��i�$_���L\�H���`�>��6��GZ�l��b�,��'�ک�E���$������bI7��b�h�'�-4�lF���))묁����Ӏ�����
�{�!����ӯ�yU�����.�H��y�p�*�.�*�����E}���ﰀUT���	B~�v2(�:pZ�����Sl�9�/�V��J��Gȭ��*唍�:����'�[��*rIy�=�tO�S��n�M�L�9���H��uPG&l��@d89�H_�EM� UDD�Sf= }H�˚�U�%c���2(wo(�\�mU[B͇W<W�'25�T�+��0���P�0~���,���ǅ���;��ӌ)�^ܠ;�����bs�Y-T����""�5�,�3"S�߶�P����>�B���5�f�����)+%:�J��7R���36�m�:t�h+S��d�hD�
�.d���g�Ԋ �\^}��5��B@փB}���c�Ün*� �Y+�q�����Fx�0�J�$	w�-LZ�{��ˍ7Z Y˻��/u���g �f6A�AP `�����o��´)���kv��U�O����#*���e�;�?�	�� ���?h�h�N�̎���_A���9O�{������8�2~�w���	�'�%ld�CF�:��/��ϔ��l܁��}�|G#�gO����y�$\Gi��f٦� ���)i']g�d�<\�I�P^�m;�/���u��q?�ȗd]��F"(!��V�⹯hT}���Ze�'\",��bN �H��F��Fb�4��:7�m/���J��o#e��g��#T�"���T�@X�K=�$K̈́]�f��l�L�r5&^(���?�[��)q���j}�z���i�VO�G�}.����R�sL��� �+_��s�vV�o��b�.����D����\�����ך+�s"�5c�1=O�56u~�
R]�9:|��Z"RC�8�Ģ���am;�h���4��Ɨ�|�$~��h��	�{MX's~#��S(��W����u��M7^n�f�[�����X�bɋĬ�i�(��=������D�I�h�+�>��!�b�8l>me��bgY�����Έ.W�_f��-�=q0 n:u|?��Dz?��YvO���[�q�#�nG�M\���վ���qe&�w|�ƾ0�H�bVe:G��xϫ�*�cM��?����޾�~��,��%n�*���g�U�]��;�b�Rض��<��wl��`F�\�V�ڮ0ԋyj�ǻ�6/J���_�t޹���s�j�)�;�pӹ���v�d�o	b�������X��%@���S��.�� t�19�heI�`�q���9�+�.�e��T��ʁ���z8k�G[̧U���KD��v�`��Yꎠ�����2�`!� YD�=�=T�it�3Y2! eI�%S�QKb�:9��T�k��	KO�/�4Pr��@*�G���J��+KT�v��"Oү#�p>�>.k3U�b�{6a�A��\�Yw�t��ƝgR��P�Id�$���S5S���5�X�9l�� ��
XH'c�|��j(т�d/g�m�����B2]�x���_F-����v���-&��J�O�ߘ� ��7��ݰ��9d���!��^E������J�d���틈˧�����;!�xP�0� ��3���ќlL�0vrq���$��,���
����h=���w<�:����Y0�t�$)���{AV��I�"�%��m�!#O�T�����!��~�l	i"N����E�X]�٥ܦ0�R�����P�\�Q}��&3�A񳩃n�8��Wb���\<�q��5mA�T���xDڽ�[މ�/+oX��{������0&�<�@���J�BI�����a�Z��ӛ`2���ԓ-5��j(G���n�I��Z�
>H�/	VI�?�3�F!��6���Ոqÿk]ܬ���.��W�ZJXx<1lL��O�@�ucL��_��P�Orq��n������B�p|�%�c8��-F�!��������Js�����ԣ�p�pw���� vl�m�N���VZ��ȉ��~n[6C��X��E�����;���B����W6�Z�9c�oܱ�@ƌ�6�ܵ�n�9eA��eQ���cr������]�V�ص��ءJĹs������=�(Э��k��wG]t�h}ӵ�`H���ET.gw�Qk8l��2 xl�l�0B�*5k)E4��f}� [k=�R�emV�	�mT��<`D�:��j��sbVZw9&m�A:��4c��t�%�G�R%Y/�h�\�=1�jQ7D�w`�eש%�|�1�>񼛱=�zgѣ���4T�ѳ�����޾�m�;KM�g�wi�d
�đA�2�|�-�R#�j^ڬ��){�L���m��Z����P��z�U��xE�R���(e�'�+]ӿ"����
��q<����&[����:��tOG�l�����
��-����v��؆Z�kB�	��K8��UD!��3>!S)ʛa���k��C{��@��j(����'�eúv�5�}�o�VF0
i��� E4�(�r����*�J���/�m�i_s�� c�D�SQ�8Aw�!7Y��C!�J(����I����趮�;&���Z��0�K�=�l��O=�ӾRH:sGڌ��^�W��Ӆ�"kA�%@|��<�V���vo7�D��i���e��U����3e#�塢���
Pv?� h_���]�u��7=wzE�"d�tg-�?j�9���������0�kQ��-丹:�U���C�W<@b[e��uX�u�c#�q�. �������I��a��	�%�I�ؾ6z���Y��Ǉ�a��BL�BE��R�5�MAP�ո0�3��b��ފ10�l/L���{ثBZQ�k����t�.r�uJ��i��-F/à�z���*M�����C����m�s�x���?4�Ł�M��#�ժ�0m�Do�`����(��6�Kdo��Wb�{�Cm�@��S����G S� �s�2��}���VZ�lf� (�/�o��5x�o��C=�W�͛is,�^��Խ=�h�$���b������|n��΋0Z!�=����=ӳ[̺�rk^cN�z}$j����r��$�Ɔ0�1e a��l��◴EJ�������#go3ԯ�C(wPF\�:�dJ�3~��KR�Ϳ�{�O��OX�p�gG!ҍYm�̾$��OAYG��������}="�}�A��u`��t���t�N�0��i�b�s�ݩ[�m��Ɠ�,,O|�W;ʪ��ݫ�Go�_"��H�hӅ��QB*&`#ӛ\�{���]n[��* �y׹�'����F���ŷ�v��p���|�
f좕&B��PD^K�P���*0��p Ym�2K�f��,냨�Yp��Amn1��C΅��g� ��:w����`�'M��As��"��±�C�3�/��wk�±�>�,�e�/�2,=>��E'=��m)��':FΎda��03�Te�g�M�8�O�=��p��Iٺg���t��[π+l�nF��{��^�Dm�멍����je��)/i�Z���}�k���a��}�)@
dv����x)t�s�����Jw�8��4����6�&�s���uO� �����@�4k-�M���W�f<9��~��f��h?n�;�^H��sCR/��)Y�K�I�~j������$�I�QB3bqJ�wk��Ib��0�������Q=-)ʗ�U+dq��"���D�z6Q�b�:q	l�����l ��3ג�L)�q{~����("%{M:�B2�r׹�J~��|���M���y��|j��Y4��H���M���.��/��zgM�6v��<����$V��X��M&���[�֭D;��GhHo��q�~�NK��޻����6W<�إ7E�s<�\��%lU��� ��b;/���ʎ/v-d(#6�����\�DPeU納�
��nD�\aA'�~��y�u��jϼ��[�	8eeG���r�F�s�Pޘ�i��`9l���N���5]�k��>�7���҆���:ғ�u�NyoT��:�s[.�+��&	�R" ��L]G�'b\�<�4RG���p�Iqe�w�\���G/�EB���>Gte�%m���^�:�L������,o[�XH�S���39'+~��9[��Y��G�-+8{�2X�f&$��E!�~�vM����%m�=����T��%�����a,?4�ȁ�����.g��-��vogcr�J�o�/�Z����Ol��w���C��˞��M�Q������|6�˅xSAT�'��
&�3��r��x��SV����<�����6�`�e:u@���P1��]+t�Д�5���0O���o��>-�s�aC:/��s��?�N�?�y�-� ��� �#���.��"�j��X��g��^���b���3v1�H:0��q%L���D�닖w���=�H}�3غ�e��Ҧ�AF�4��rޗ�aR����UI��PV>Ǜ�1�x�%��ϋsVĪ,�\UOd�*U��v?_�ṵB0�-L,�l���Zєt�_�����B��� kB$�`�рf����6:�:���G��%,��UO�:���Tq]^��&jh)'�Y+��c��F��-�;`����,�e��A�����H7T�u��.QCq��T�I;,p�U��j���s �b���S"`�!�����!`x͉d!~�u����-��|K"p9χ����x�GLF�EJu�Yk$��z��a�2+9Fb%BT<ƨz�>Xsܑ��ih6R�Na�)������p'i�+"x�G������>P�Bj�!"�����t���4��\(L�^���j�N�-u�V��W�9�<��)��=X���!k&Kb+�nF��o�>���Q��I�!uK��P1�q�68
$�-�*��pE���n���Qh�%*j��q��@,��?�^=H�R����Obw"f.{
�4�4=_V!c�	v"l��$��=����4Zګw cۡW,�dg����`�R�|q7�;9UzT���E�Új�V�nԌOe��ϷY�~�7q��+;TF�Gn&��db*�" ���s)����P�Y�m�3�"}�3"W�a�.4��^�Q��[��t��@�S����ؾ��B�FF���:�>4�o�(?��}N߹�z��<�M�6ȼu�_wFؚ�b�����D����8�K}I�+�+F�{�:H.�/��i6ҙ�}���[�0m�z���#�5{m4N��n&�FR��gD��>��Յ���Evv��C�ᖟ�?��'ꊩCz��-#.���A6��&N��(�27m��c��+J@�7��B#ڰ~p��=ц \�K��0v���(Z�^�a�d�U![���%M�oj�%�/� ��Z�0��N�ͨND V �.���}���rt�
���T�
K��ɝ7���(�B�DQ�y��U�%}
б�PI�8d��OU/E��~��m4cդ���n�)=ުp�9Ӝg�Ik�+b
�=�??6���_o�$n{?�����'"I�rt���{����A���j�@���G��	�Bl�z�H�T;C���w����*��jO�c1�8���"�UX�G��%��zevx�T�_g��}2[O�L�1�9Jt]ݽ��R�*̐�ʬF&��t���E�i��1�A�i��"���� k85�q&���#�dH)���;f����-��{�]]���a<sS'��l��*4W!ϕ?��]���3n<����&gukvqK�|��lђ3���O�SA�f�&Q�w������1��4�5]�J9y��8@.Jg��{?�t<�uJ���5�G���"�[�\RR���%���Sh�b�%�Yh��.�Ǟ�z�T����\&t�QD��ԥ�L�͡*���@��{��6\�ź���Z� �96��^�l��1F�U,Pp@���˙��=o�C�q��Ů��.���ձwT!��F�����ٛ�_WW��-��L��$�>j	)��V?���B�R3:Ze�?���@F���$�:�[�ߛJǓ[wِ\4z�o�}`�I*Xr��1�a�"�;�?w��g�#(�o%8��c����
rf���y�Ϙ��-�*�# ����6PxEoR�pX��ơ�=ĂUIRР�4�W��6�g�D� I�,d�.-�tEE�HL�8Q�'l��C}��$> y]ļ����lix���j<V_���k4�nwG�m����g���z�h��7SQ�C����g��#�P쯢|c���nq�x����r�碥+B�$c'�l1��(���4�����;���U�
��< GE��<����ήN�1��UxKj���1��j����J�xa��!�w�湳'-j#�������f��t:��lkz��X����Ѯ�����%�xé�i㰎��ϖ�\'#�kJH� s�r��E\�Il�-D�C>$8� hfrG���%z5��r��98�;)B�ׯ@�ھF�_��\��U:L��0���ؔ����	�9}Әh1��bw�����tE��}ɣ����RYH>�L-(Q��q��j���.4wwL��<�D�ϧ���
���� ��d_ic��!I'�OHg�j��rR����^y�nb��y�R��^ه���2�[���7�_�Ur%y�;2o�:Pt�a2tH�Ԡ���F�H���/�/��$ǈ�gGB�,TN]�\�]�?�pJbc�+�N�J�I̪�����8*����(:F��� ���R��|��Ժ!`�)Bt�&W%�t�9�?�^<�:YA�	�َ�׈�p���"�u���>/�*!Q��,��`�|�	�#+']��vՂ�giX�:n;�D�C���g��9�>Ʋ[c����a&�t��I.TĆ���r�X�y@�Je�^�5�ɬ=��1���kUP��RE�h��Hu�A���j�L��gN�W����6w�0@*���i����j�|=�sSɟ2�_ChD����_��҇ y��m����sC��"C�!c�R�u0&�����;���G˭��)*Ie�=O�'�t�9P\首��ד�ȭ���t�;@��,�#�Z�e}52�ZH'Ab�����F;�y��,�ڄ�(C��ۼUF=#op$>��\R���f]P���}�G��X����8MJ
�օ$���0��d/��Nw����$��HC�:T��$^�Gg,��
^��$��@E����*�ө�K�9���.�W���Lʹ���S���:��iϔ=|�&o֯m��5KNL�d������ܢ��RcupN��K�A�<�j]1���ʘ ��(,F飬�NԦ�Ur��3��hG��qDZ3"��:3�Zg_�������*��.�T�4WK�z�l�O�(˜���!�C ��2��(��)v�%�be�F��(EM���.?GǺF�m�qp�]�|�f������A����W�D
2+)��"h|�֡Q�^�$d	��V���=��G���=d9��í+��{����QP��#m�h⍒�ViH ݳA=ft�c�>{�M�[���l+؛��l�Z�"��9Kʢ/t�`O	nN��%�goRT�.��ɦc��#/�,�]ͧ�G!)I'A�z��-^���c�f'�8������N��9 �a��b���-�E�J����ɐ�w+�:eD�)A�h�oš��5��f���io|�*L��G�W9���az�s bN���1�L5�n�?�Z�+�����N�����I��,���V�5L��_~׉/���k��W�V:�k���hP���hX�n���=��c�������T�?v%ӱ�+�������;j�����8��ضwR{vQ!�d�b#�Fd�V�~��b���|��.v�T> bn�0..�fr:�%[0���"|0�s���y*�"L?E
��B��t7�ɥ�I{��������/�;,pkE��]�s��Q��k�B[��XE��4��I������B����|�3�hn�(>5/��t�|�����84�# ��,�������8C���9RL�������;���AGh�7�0H�#����<)G��Y;��X��m�)쒨7�Jv�=�b��d������ҧ=�}���H��Z�����[�b~�+Ӄ���/�
3"�/�$��F2���iU=��E�*` �@��1�95�S�=��9�oCy���B�a�L��q��tv��/��f��LF%`�q�t�\vc�k��ʜE����B0�����kG°q�%��)�Y��Fh�i�û�`�iN����U4�h��������[���<4��#�a�$�8kAR~�H���M�Cޔ�YNZ~s�X��S��)�2x�#�@_t\��T�6,���p��%5
أ�e��*����qn���M�,������`h���Z���X�B�!�����oLεT�ו����+L	I���?C�x|����:����Y�z:�Tԃ�_���=%O��ˏ�D�*�JO�2^Q�C�����	������f�_��O��&c���;T��Jt�ae�Ι�s�e��b�J��X͑Y[��Qք"i��IJF��y<���SKu�j\JN:�_w�BbFolO��j�:���:�05��RM�e4�%Lm��MI��f�)O�.w	��'ʸ�jh՗��:L��[�n�*��ˢf�ve	���2�R��9�"��#���F��"�/H��ASIg���$h�/�J�~|����v�:`����!A�l���AT�9�D�{�9��z���)��]{���b]�QS�q�-�5���m��/�O64��}�W���O����ے�H�u��RX�7�z�	�fu�ܳÉI�Hty�nش����ӫ/���5Z�I�z����5�w��kd,������K2���K��B��ELZ%8�1v��/� �p)��-���`M�@�sIJ!�󋤶9p"�UX�0N��ReX���ATJ��t����]G�:2c���,��4in��/�,Oٵǁ��ϣd�o��������:�
'Lט���Vހp�o�Hd�\9O��!j�fn��Mm����s��@�kM���%��� 0?�P�ù������*TU�$����qG����L���c�/���J����r������*�=�\���ꦫ�1�_s�ύ�3���Mg�w�2��������L'@��j��6N]j�T�!�\�H���5YKR��'�`��p�M ;��7.V��BҾ.?i(D効_���Hs��C����2ma�vE�!T�m����!Ah�%}�/%̠�����=	�(U5]�Q��V���fz���)M��JH`�qֶѢ!�݆].8�%^��ޘ��Qe����CC����+�2��)G��gT����M7=PdѺ[���I@�Ya��e��t/(��������9�gN.q�� ?�}�f�5/;���jKjQ�g�ظ'������,RwA���$��w�J��q�[Xex�N.K�3����.�����Z]/m�Lr�	�ġCǋ����vd̒=���Ut)�������X��`��392�N=j�ᆏ�իd]-���;!aT��x������~k>�Ó1쒶�[�֦�3�t����jQ��	���N���k�8�d�-ɢ��ݴG�
`n��@f\�}�*�vX�x�k]T3����v�#��D0�M�o2<���&Y:�!����U-��U� �J#�u��"J7��� ��z4��Ʈ�t��<��J5�ؘi��������2=�$_`4�� ��d]��(��S�;<b�Q����0��b���e�R�V�b�˪ka��]_�d����z:��Jv3�7J����A���L.�&�)�S���Y�=��!������0V�΍�n�q4��\@�F%�O������<-qr��͊jG�n�Ǫe� �Sp�}�ש()>;2��o~F�������3�}��E��+�I.��:����VۼL�T-cc���^�3#����R��q��Nш+�.���ɓY��9�㒋a�����?�H>�O��6h-!-!��=~�k������.R\4f^Vk&�F�8����-�
a���9�p�7T_L�K~5Z�q�B�51��B��0��h�>�s���=�%�Q�{ÛЪ>@�ˢl�V��.(�Xyu�=�Q�rܮ�}ʘS��[4�Cӏ{�V�����ɲ�3��\]v�'�r��Ep�L]q��kͿ��|X�#���ig:��+�~�㍑Jrx�.��&)�QǏo�olto���m{��ƴ�Q�Hs@I`7Ck�Sa)G�TF򭅻Z:��� n VTyi�q��2�������ӱ
�X6D�~ZUR~��b>�k��O|�I��qǒ�)���ڥ�8'�Lܛ.��UbF*��zq
�C��|��a�ن|���>��رq��{~#�E��!��ʝ]���,�����6���C�����=�e�Kr�������xYA�&{��r����w���Jި|���YJv'h����\Z�c���Ϝ.�����DL��*�Va�U����ᵓ7�#,�XL�oG18��2�tҟ]٧����U˚U����p���t1�ms��ȇ�V;��:A8A@H��I�gM�K��z#�d�H��������Z�e��k��X$��[&��b�Z�i��]�ܸ��-���MdgeU���XΫYXq:�~zO����zM���+�|3���c�� �j}6��^�v��Q�nJҴX&J��XN�(�yxhΡ(>�~t��F2si!:F�ы�����?��/3�^ht��EZ��!]�j����?;��(�>���9��9a�pH���9h�Cy`OD��6>��c�i�=�(�StY;�� xڳ��(�������Ig��������<��y�=D����h�Z��S ��E�9��ST���������j��d�gn�֘�N���e�9�>'N   �����#	f9.��7��Ҿ|�u(�����/����T��뛟Dg�����;¾�Q��^��u��Q��h"�~`�4/�|bk�#`�B|+��`�?*8e�ɦQg�R�	A��}��oy(Z��aH���i�A��fP'�b+���>s���xa�J`ZF�뀆�ki�G>@����r�
���zχ7u�Cٸ ~z��!�|�T�t���_�0�05�	�+n�ܕ
�H�$�R]�׹�t���Iζf9���ƂN����Us���n�#Ю�{�j�a
�C�l w�tv	�i�*�-���'zm�[�f8<g%�;�?��Ͱ�3�(s+Ք��ܣ�G��aԺ-������2�lJo8�=;�zG�@Ű�4!�	�0�C<�����ߡ_�gGbF����|��Kܘ���-tS�'/�m���pn����0�	誮*:Y�lv��i��]�ʢ\�?�X.�%���M&��8�dF����P�e�)#f���K&�gR�(ݽ��*º�c��Ε��/o_7�GHW�we�ߖ<���M�ҝ�]{W��݆JK=���Q����&/KAC�_k�}�x�<�W�n�Iד����M��{���k�C)>�aY{���g6�%i�Â�L&�FG�P��5���)ד�]��h	_q���+H�{�7�!&y��4����T�l	��Q��$�X	�/EL�;0�}�n��~�'DS����=�b𛪘c1�� 1r̔ϱ�_ 6(���i�<Ϊ�4]��Ez�oy��ӁN�q�
�Ԉ����:f���,sZ&��6�rh���?d���xٻ�@n}��	l�:��@@C�)�ht��QQ�&��d��UxO��l���ǤxSf	���s6��4��`<-LP�_���Vi��/��С���q�,]G��#�I�Kc:�:�� ��\ضn����H+^��oYnF�m�?DU�6Oe����:ϋ����Q/��;����!Hp��73;�9O�Vc��5���Nv��h���c�F�)}�K'J�ua v�6�nv\��)d�#%�f����_���o�c"�.|��
q@�ބ�_P>�F�����̪#�d�5+r3��M�O�� >��I������41��^C1�!�7�e�x��/�{���X�qM*ܠ)�P����^uAY�w����c��dܺ�F�����Ԫ��=w��GUA�d��]�،%�$k/�3=Z�:��s��Lyuj3���X�DqCd$�I���������ټ�x��7��t�����f���qW�GL+�-��X�vh6��b9�f]���/ϒ�M�%�K2��P*�c��}r��Z�|��~�b����YyE:��J�A�_����������1>�o?��}VRj[B�0*�p�s�@��Ԥ���&���s�j^�5���ｷ�R��sJ@��Vjt��H{�ϕ�
�i|��,�[a�D�%�N
�x}D�����tT�,!���:��<���"Y�]� ׌���t�`Y�;ġKmF���{(SLǣw�d8�PL��X����&��[���Q�����{�è�*�f������'M���?6�_~��ʫ�f�[�q��o�H�䥽 ����'9�Z�A��B��)�gO34��~L��ش�� m���k#���ը;^���p�����7�c۹`�_ÃF'�I��$�ڟ�~�VA���W����x:Ca��C�_���(7#���g\x�PGbu?2:����9!�[4��+M�R7���Qy�v�4d��cɿ�Ğ��Y�{&���$X���ō�5��� g��@��:8���9x�'�vؕ�P^L�DX�3��IKHh�5����RDy�^q�E/#���X��������P��N�}�y �KZq�O/B��������	8�0hdɤ:�)b��zp��H�y�����4ΚJ�ը���W�C�-S��p8d��NYӍ*�ѐg:%T�z ���4b<�� �R���a}��%/B��)�Qr�{��ֈ��DݓH�ۺ����h�����仄�Al2R[�U�#�w;��)^QQ�HzZ
�g�/)-򂋚�5�nsc�vnG�m�J�.?E��!O����|��m<ķ$=b��m�LF���[ WT軹�w���+ <�`�?O�b��7�?I��
j>��e�O���F�%�Է����*�>�}6P���][�t��}���VXm ��m�O�8�W���D���
j2v*�tB���3��l��%n��3�7 ���
�r����+-*�j�U�a�duX1n�S�.��r�Y��x.�U�t�nada��Wd���~��H��ᑪzvK��D�v�圆�/�����7d��͵��+�l���I��/w����%0��r�)�O*�xyɛ%�]5FƏ��� f]�pܺ�ݲzcASB�C�ċ0*��0��h� ��%�QD�Ŵ�����!��-�J��5Wm}ZoG��'�]J�Y#<������������Bb�̮��b ���R��׶��o�ɿ�yE#MM��=@>�3�`z&���U�0������x�][[�	 R�8ۑ|���9Poɿ� UW��m;'Rg��A㪎�_�VG�� I�4���Sֺ6 I�����*{�+�y���6�L|��Xd]�;o�ӂ|8��A���"�)�4�Tɧ���ZC?��U�q/E��25)��!	�b	-@%��2R��c(�S�f!��\'���'��P�s>��OY�O�*������U�ݶ�����|8.�=���\B�=1�=�ND �}j��Y��8>���t�����Q�'Kt�5�*b���r��q��H������,9K�[�b��Nk�Q�q!+d�$�?����i�J3~��8�V�2���ov=p��.�7��1خQ_~(�bˁ�q3���I��兦�%�>jYE;�s�b��I�i���ۑE�ؔ��h�p`�hB�}�
K��ݏ�o*��dasb��B�^N@wMb���(��:��zЬ�uc��3:b�p����3�TPh��\
��5�D��`��&��~���9�xYW�?����U�կ`���bB�����OB4=�K�K3������ғ�|~����5=bm
喝<BF�)Ay����zL�X����~���veRV+�j�"�$�V?����9�u�F﬷�;6r��h�Ѕ:9��[3 ���c⚅:x��"�-�$�^xn��)�:���	�����_exc��=�U�>�$4~�l��2ik|�x������2��C�*����gL�ղ
��KD�ɎE�\��im?Py����i�R^d uS�{�����|�5֌�0��E��Z�#3��0�i�}ڇS���@�=4�ڀC?	�D#��-_���n��`0q�3�\�'.5��:f�|e+H�f��l<c}��]/�4��"����$er@����y��Hɒ�ì��Ѕ�G��i��Ӽ��5;���KU
`��맱sN��6k�S�վc���*$O	���Cv{/��x6�L?z71���S#;
�����(�x���$ݴ�i5���0����;�����)��H��u:L$;�ҽ!�����Y=�=w ���I�O�{��=|���s�l�r����{kz����
	ew:r���܂��\�h���)*���K:+�J���-�a/� R=w]����b�%�̝�R`R<O��:���>�������*��*.e�L2����7��>��n��������m��5d�*0�yZLXTl]���SLR��e�J����;�&4Mw��q��chh���ԓҲ��6ȗ���vA��f���fq���l����]@u�dT\>	X{t���e���E�:���N�?�ZJ3gv��7��5F�G쐹��tG�=(�K�yR	���a�����+_ƽ�(q�W֞�'N�"���*�G�M���q��>$�W��g�V]�Y �p�W2t��~e�hC�VUGy�+Y��8�k��<�7����]Bg��ԋ���lPry(T�����p��t'��]�^��gp��{0Xe�x�v���9ɾWA؉2G�D���� 1:��,��N��a�zὲ���>��)l���u+�[��8Vky�F�&Wfe�Vq��ٯ��7��e�r.+��@B{����`����t+�mӯ�]���&�TJ�ۙ�=}`"`���(�-�Y�A����`2`�a&��b8M��]$5,�S�����Y�Puu�¦w����#���q����]���jͨB�)Yo�E�����n'���F99���,l>"��-V�5v��E������L���.R��ޫe���?�}n`�t�orP�F` ��N	}����yXݬ|ʀ�*�A}�j��ِ�Pt��l+w�´��w���O��	I�
�վ��0��H\�קbw�ІE̱ĭc�a��[,���up�������؅�^��Ȗ�K̤�|X
�	P��\�YM����R���4���M���q�4+ �~�����9-k
l�(%��K����;i�6�0��v�7�e�ox�~L���u~��,�a�M�܉�́m6��d(ICRn�w��>SR�m�FY�d��5�I�Z�����st%ҁ"��2G3WO-�*�"�j�5q�s�ے!E/�\�_�S�i#�Ŝ���9
�㛙���U�����̬_n�wG�U���x\�*�܁�0���-V�!w,-�6��^L����%�xt j\��r�I�ٙMd�J)�W�Ng������dlץ�oEɑ�kbIHT�Z�E-�T��	�<P�E�,g��1;�5���5��t<��uP(D�ew0_�l�����k�k�C{�њ��P)$�D�{�2�jd֕�
з<6����N4�F/�D*р�
CIW�Už�ږ��FbaU�G#��>�Y�WVD'�����JQo�!>i�=X�9�+��Qt9�Z������gzD�
`R�o����[>w*d"&h�� ��3r�L�Á�5�~����jX�%�����n��7�~Xv9�a�֙�~��˪��n�Π�����^`?�K�ǎua�JW�LnOJ5�E��I%~2n+uN�c�':�ȜU�����2mcF.զ'�5J�fّT}�j��[X|�Z�|g���Ŭ�)u��9����!�-%)w@��A7�V���f�/���6�SdWBfQ�|a��I�@����ZF�XU�r�u�)\Ѵce1\ￓ���Fo|T�>���r��Q�a̸OeW�`�<����$�<�9����÷rE���n��3�ù��N�j���j�C�Dk4��4�A$S�]cYbi"y0�{��${�f^B=��)#�T	��o��[kS��#�B9KZֺ-��.��ɪ.� ��\m*�c]��ڝ��)���&�\Љ�=�UF���V^Hwi�?W�*U�P>ʀ��S�C!�O���c�O�4�B��V(�uyw)f�@^@����iz�hM����QÐ|D���z��j67n8;�]љA_�,�x�˩��t�D��:�NR��adyU���[��
�������}�� ��K�7�����?�E>(M�=��0ȍ]�E��!+E�"�1φ�U]�x��a�bd�5����Oʓ�D.v�o���%ӛ5�<�^H�}ʱ��fXvּ�����ڧ��+y�H=i��Pt�]�Pɜ�6��������n��c�v��Xh��*��g�(��a��VE`z�����Y�}{O$?�l�u����EB�̾)��Nqo�(,��Jw�(9�0φ�̔��pH��.�m��:ǎ�X�h����Щք'֘x������Nq5�4�MT>/BsK)X�G���$���O�tyixK��!.�1|���-�Z��E�T����`8���
~���yY�)hn�o��©�V$`5.,i�����_��.��d�Bɻ5���E��D.��|�0˒�v0��y|B��a��O�����+��Ð	W81����m�uh�U��9$E�TD���CM
(�4�(�U��A5�C�
���K)1Ō|}�y��4]�r�e��'[�@�k���+����~��|k�i�y@��BX͡<-x��7a]))��מ�n���l]��HjOZ�^��g)���I�_�E�+��H߻�2`�yt������S\��O�r�rb���ƭ�;�(/��;b��<�N��\����8�x��˜e��qoz�/N�����S+�S���D� M�E�M�:�Mz�'�lȘ%n	�R��q���^&IY$ES �5�$��<S�a�#V���Yv~r�zpq�쬔T=Q[� õ-�4�&����;����<O�MFO�-Y��Ԑ'�8�2���c���/�wnWLɣy�.��5��ٝ����L��f�[��_F�ΐ��3/���y�M��{�)�Œv�����g�1�M�_Nux�F���[�BS|Ƈ���ռ�����s��}�80�Pz����X9.|Q�J���M��hgiPPޢ$8��2�����B��mo�A�wY�?o��0�rR��P�ڵ��$��@v�����H@�7�Q��%1:%e�|�I<-�Z1e�i��3ALDߟ�,�ᛣ���y�ZM#���?��(~]�����wOU����� �>�,��,�D����e����c�:�y1���1���H��4߮�d�讽1�η�n0Dw)����C-�^�i�1j��Y���������C��� y����^�X�8�{�X�i������݆�7��W�Ԩp)g4��d'b@5b�4w80b���4�+V����c�{j[j��L�í\!kaO#�f�"#����.����[�ow�ћ��[�`C������G*��S54��D�b�����Yٵ� )Ѡ��w�MZ�qW�������;-�өV�Rc��,�l����W�����.iΪ�������H���;�Z�r+;[99u��-yj���esa��oI�/15�B��q�k�
0��p'����������VI_�ɯ�󕶿�0~����(���� �~P��ŀ���oڢU��e�ȰƜ!\�9�J��7i��A��A�h�8n�CIt��l����T޿h�m�H|�������w��?�یR�D�;PCB�}< f�!�Anpf����̨��V�]�ݴE;������kf��p��V�I�lR�G�����1�%������
�J��5���_���M������*_��B��/F2X*��SA�jJ��ۿ� ���w�\�x\��Q6z����ս�� 5 �0k;1CU��J4H��~|�`5}���E�Vp�;�T�X"ӝ��U
\��%B��Kۑ+�|��]Џ/�k�bD�=�#O�D�~͏����G���aq��-L�F�ׁoG���k0Vٵ�^~�z���`�8���۰vU!�B��`���n	!O^4m���q �{Z��G ����}�&.�s��3)]�榸�LA3$1�+�J1j�L���)���x<���R�-�7e�~�6�u��j��I�8�����Y�|l���Q	���^M�~���~I��S��?��,���5_`�[V��_l��\cz�8�T���`S��#
����GQ�B����O������*�-V�����ic��)�Z�op_6fP��%e�r��g�|@�	eX�jbAq�/-S����;E�{���LY��o�ѫ�������q�hcE[���ߣ�=�v~E!��
A@�_�j��r���0O��#_=��
Zf�������X����T������t���YZv�M,����ob�J]�4�G��*�Ŝ�C"β�o\�2��W���>~�w6���~��EN�{�E��e���i��3�|�s��օ,~;�#�k�,z�7�E5i�!����l�����KЋ��q�{�"�p��i�r��-����� �_�g�Wz�JG���p-���l�Z�����<_����'�&�	� �߾K]����Lw�K,Q�����y�W,�!�(6d��sa��1�M촻�ւ���*)���5<B�}���-F��Q�	DH�+;�Ȟ��u��*��/�4i��!hL߶�FԿs���-T��m��6��N��!-l�%�|���� =I�Jx2/���t`��*�)A�*��r���P����d��a�Q
�vn��Q�M��ϴ*��!eg��$��M^CRX_9�CA��pzh�m��S�'&��憛�?�Ր�k/3���9��p�"B5!��w�W�e�ë�ۋ��{H%��r!x
���s�Wі.��"T�j�������]ˌ?O+S��oG�n�7�y�������	j��@SZË��� ^q�+n�CFJ�L:x=�f���V��G7�p:3ƕ�S�(��;o���(*F��Ij�5穚�J��iq�� ""L�����
��4Re�9��]��[9�9�0�U�S+�%�ແ"]���t�nJym0ͮ�B���e��F���I��Xl<+�v����ą��M�wU$1�P��Y҆�ˑ�@�A����m��]`�tT�ǡ%j�.�{��P�	�S-Y�j\�e�C�c0(�쑺E �.p�s�I���#0 `�M��B�ZU)VF��3���a��,l#�w�V��b����fٸ*^���c�s.��G��;t!^�,T�}X$[Y�>An���/R��)��"N'ښB�됋mY4���*����n�;ᓭYs�`�f���6������U��v+)�^5��M�s���~`!�	��%;l1�ѢI��vݏh}�h�@�d�ᳯ����m�P�Kfi!�wϻ��Q!2}Տ�񩕬Q:��c��P�Ɖ�pi�g,K�B6Tae�@����j<��(G�G���^��(;���ـ[���.�O��*����f`U�gU��9Ϣ��>k��OD�J;�����}V)l�i]J��1�uI�'�pv��W��C�g��|��d��Z�M�[�,���h� ����>D~��1�_�{�,���yF]>��l�|z�FuD;X���(��u$��d�)�u�]�4�u��RS*`�54/Q� K�FCdu�h�
M�}/ZZ8OKՙ�2[(��=�YU�	�'�*���ϸ�ސ����2W��lܐ��}5V�L�g�m���ￋY�9���7(�~���W:k�P����A�ӹ�����D�H2�il��OP�u�|`ާR�
HĹ��T<�󯚧/U�<2sNf�dw{�b�;��&a۝ �~��z���� ���Om���f��fe����f`y!,�w��]R�lo�v?_"F�����ꁶh�/!vBK���d�P�j6�����=����+�,��� �;�P����MP�LF ٟ��
���S���;�<�	��a�r
�=����R�vr ��"��6��آ7�m�WWr���\S-�w߮U�$={�7��!g1w��̳��j������ˢW���
�-pJ���������U?�!?!�dS��W�qrU�WK)E�v\(�e/�g�7����	�JφtY�exŔ��*�|�g�m�����[���e=?6U�-���R�,�T�f�B�Åj�ݳ�.F��4/�]����������ِ��z��L�c�l�2���|��J*�=R���<���8"�yҟ����%��Af��H�:���evY���<Ksg�O�û'9P#Cم3?1��+����ŝ��Kz	��/��?����|�_Y`�Q��J�K@�$����zA(�[el�����u�嗔_%���j�:�š�A�!��,*�m�'���
�<��8��]�v���Vq�
�&E�<���6����$]"�����N>��8��Z�\=Rb:l����!�@o7y�fK�}�E��s��S7CuC��*B %/�K.�W�&z�B����z �#�
.S/�H�������w��l�6+6[�"����|����@A��6	�%��)}�p�2�*,���{4���q�X�hR�!cȷ9�ֹb��FO�]�NS�
n�
*�qmg,����ճeS�,|H��+g���9A����4��L�����e?��������;C�`�H&��X*���1o��$�ɛ���������G��	�x�%�x���OF��Z{>99q��PK��Ħ�"N��hcA����e�_��������M@�0 �|U֜TrG�i��Ru�fٸ#��SU+�e�:d)C�s���Sm���vPf�0�����)��N"�L�\�l��e�ׇm��H����m �w�=��od�@��W�U�a�ڟv̖A��fX�hb���$:��?j�lR-eb�	��S���_D��c��S7�Ђ_�9o;}��:���Y8��,b�W��ǉ�����h䗀�y="/W?"|���P��60pʃ�]�%���w�[Z�)�Eq絗�IrU���8��ި���QV[e�h��ѧ��ph����)5ѣW0Ou$;�M���aV��-t� �@hܛ ����-N) �w�����i��I*���H�L�0�f3E�is8�\Z����ًj� AG��@	�ˤTj�,8mP�俓���y�Pi�T<�`p�z�1���$w=|�����!��h�qHш���������l���ʢ�^I؍���L�,}� ��k��5�=����9�;N�����64[�}\C�:ʙ�M9���J30��#��[u�"x�~9�Cy5H�o����X�Ou��xV��F?*c��\p%��t��}&k��tC#=��`�e�]��H��`�/(N��]t�Hj������~�T����O��S�ϫE,oz�v�9�$[$Lů(18���D'��i�6W5CN��[�n>�=�z��HIl'Ԭ{r$��ޅ{%�G@ڔ�'hT[�lD ?`�`�{�k�=��#����vB#��Q�EƏ;�3>3���y7�k��̃m�_��_7tA1SQav�r�O	�M}�4��ʷ㤔��C�c�IQS�����4��2��3�d0P\%_�!�]��0�T�F��ߡ
Ҡ�x�����z�t�.�;�O��% sNK�(�����	5d�2V�+�V���j����jJ�.��|�|�FI+e i*�6S���a8��U�w0g��4��L�,��nCT_�ϧ̛>� m5C��K_yN����,5��5n�³V�f��#���>tfD���m���W�y� x��UE�'�=�.p6�w�&F��,WS,%��d[cc�%Qy�f��D��5)Jb.���c���`���D�c���a[Qڰ����M�g>�f��M�E�//��wm�����Ɵyo�T�-9�)�%CV�#*�ښy5�=~�� ��c5��1�3��v��4� �Dz�� ��VM�-3����}��/n��i?Ｘ����%m���b����3;�z�^S�����&��;[%��M�8�A��=��v\W)�
�����^S'�5�=,��dG�H�#ż��{�gFI��PvY�A�՘�����N~�pT Ғ��ګ}��j�x�AM:A�j�+��n��AMg�\�UXnI��as!㍦��drrv�׭�;����#NH���&�u��6�*-����C>	�T���e�g��-��tb�G�x TgA����u.b~ÕM�.>d��v[]*4!��
�&E�bK��ٗ.�x���D]p�ؗd��<���o�\��ݦ�|>�i�ދ��d[��	]�l����'��9�6�BKt�'�Ĵb��ȧ�N��$�n�1����z�-��Cp�Us���9���f���w:99޳�וA rҕ�:)l��!�͕sn�g�u�%�8�dv�߀%1cZ�s��s>xSiK�9�~zT^G2��sAvP �p�Y�H���+9!Yd�Ð+P4p@��'>$�䎕=ǾO�rJFĦ���)�]6~�te�s�Z��c���ȡI��Vf�CZ��R}=�ޗW�\������ξ�*D.[��P����(��<���5�2w�{������1��zH=�%�|�;d��瑜�O�����&���(�V����� |�x�ϊt��9�!����ޠ֣��GS��ܬx�9Y����5�l-��s���K!P��������M>���^��8�e�!�̞@������T��<"�����=���CR ���QkmP�R<�: �u�dTP�Mv0bX1��f��[p���G��w�j]�T;�F���iO��g���_D��Ѡ��&Gv��3��<��%�x�v�^��:β�U��7l��Ra�0{�d���]��sTDh�ߨ�f�f�'
�Pղ>�籖|ܝ�1�M�AĜ�b�*�{pM�@�	Z1��N�9K�#%y8j5�
lX(5���Twߗ��)��yn%(r�U��F���'�>=�O}�RT�KX`a5���vz�z��zR�V k���V�DW��<�|�G�K�, (Q���h�~V��K���el��bT�u6�a���e��o�?�V��	�}<R���� �H@��7��Ow�^5�0L�,xթ;Ut�D[�t��Ҁ�Yt����,ߖ�4�G�i��W��O�9�� +o�������i���p�4�8)�'T(�iFE,/5p>�
r���+� ��N��3Qg����K/3�ֻނ�}�2K��}�Fe�+s�����{΄A���6ջ�hi(��M�(�O��ʹD�T$bUM��2GƉ�9��̘?~�3ƶ\�v+	E�Uw,�$R.��J�Z�R<Ϛ��Öщ�=��?ᘐ�	v����c�I���%AU���3�	־��Fu����q�Ε���t�`p�A�c������:s��_����0��r)���r���R̘y}��Twȇݸ���st��x���23����&��U�G������_g���U g���1�UiEC�ᭋ��|�M���ݠ�hr�����}-,����f.Aia1-�{�/#��Ѿ�m߲����p�Kl��j7���Lu���<�T�(G���>�񃚃�E3����Gp{:�գ�D�e8���:� s�Z�Y6��C�ųҷH�#x*����*�|x�rR�m2o	:zLb��+G��U�O?Ű��;F$7���d��U�Jœ#Hڹn"�P��?�#T���)�0�]i!q[���c�r�	0�����]^�g�KӠ�ש���|�M�g���t19��c2#'j<��8���k��~��=𗘎K\���ˬ�� ��r9��.5(�%R�p	,�"��Ju�/���o�ds�1�� c@����!��t|���(��}7���\�-'`���&�m��rYXn{�q�T���H�$�T[��ީc�@�O�/ѝ��_����K�y�̠ajl�)n{ �mXr���Ȭ�]���݀�
���1�2���u����Dy��j�X�$�-��j����%�(I	�p����|bL��YG�IwW%�~��Oh������θf",p:>}�������[�z �`,��m����1�E��L�by����*��NK�<r�/P�kF�$I��KduX�ÕɆ_�h:��#q����l-j���L�5�RaZ�r[w��@8����|I
�{�]�g����>\L�L~}����Ś��Q#Q��F�N�ϭ���'�"@o7)�����}�6,I���u��<?%�q�1"oy�x�����G�+d%��H�'~���I¯\Z�2,n��E���L�Y�	�%dC|b*?�K��T�JDnW�4��&0����кn��*�&i�!�t��{*��g�}����t��ʞ^f�E�u1p�h�r����N����)��k�U�g���Qnʢz�d6lվ����^
����+�u�_RR��ʣ�\�ܣ��^���Ć-؄��KK�IQJ�'2`%�#�;���0Q�{-�u׎G��?4!���v.̚P��O@~/�k�����kك�$6h��a/��+����V��@4��r�Q��DMR1��Z5.gu��^Q/�,ە��>�;�HTQ�-�1n����	�L��H��*~鉦����f}���gC�u��:H�>��Q}�N;ʩ&3qo �P	E]�`�G+�y�ш�'t�Ɉޅ��N�+����ڞ�lmD8��C��g�k5USqN���j;̈�T������u�g�6�'�����0�C�o[ճ8-��?��1�G��,�G�a����Y�ߴ"SmD)t��s�K�1�̵Xv���C��/��K�_A��H8�s�}Ų�?����Lc��ڧر*�t{���x0=�v ��V��٬�^@.	��y�~�k�� �mt�g+-��ZA�z	{�����c
F.��k���Iec�sq��mD#p������5
�@���y&i�~E�tl��0y��Mz"~Z$hɷo��
�v�m�]�<12M����<�vԔĞCꤱ,�Dl&�N�&.��T�N?�?M�Q�Z��q�Yi���e�>�Gֳ����w�՟���F�ޅ�Ī�"��]�m�-5 K7}v���"�l��S��nj�à ��^�q��k$$����G)��,/�DJ���qKq���^��̛����z��6�PL^֨�2��-�(JO܄�ؘ�/ѽTԹ�m�4#l�#S��Q�h~�Ž��T�b�Z+q�5�j�n�?�.�H���;�V����P�i�'%�űiΉi��o��ۖHw�S�����wL�uI#�a[M�ȍ8�2K�q�'5����'-?4��nG�'��݀�QM0��7�n��W�,`	��d���,q�AW)!��N5������u��:I2��qϰ�[����#
�Z�Eh�](}��B��)��g8��v�	�����2z�r�$���Y��W��*D��O	Q�U�_����@�xH�H
��-��7��b�K�F�V�s����mT�2�#S��� =zIV�Cьê��6ѽ[,��R���౵�;$���|��Űjg!�sbAx\I��A<�k���a�r�9\/�0�Iَ!��P|c�#g���J�-,��}C��"D�����M��	�J@F|�FJu/��$���ݞ�[���?�s���Y��G�G-��N6޾i}C�7�Y�qR%y� ¿)1�4J�x.S�uօ�2`)%k�����oU斥�����z����X��6�Ȯl�x�O:����v��BZ�Ԯա=�4c�)�T:{t�!��Jc1q���[}��t�3Wh�,��}{�c}kŗgg@Ws�ʬV?	�ٗ�y�${�U	�Z{qA{���o%�����q>��6 ��Ê�o����^z��N��d�{����&.}��k��yU�-$�tV�jD��-��)��� ��Gu�7L!d�r+s�pJšG����Ս�u�'U�r�_��N�MRvq�7���m�P8�p�bb~��/+t�1��X�%x�ڜ&�)xM���r�/0Lx�Xi�V����M�P}^_צ�^�%��}��D�Iz(��X��rS���ȕ|a�Y�>�%�Nf��c&|@��"�H;@$FwZ��+`�T渌'rz.�gm�@�ޡy��mOG����BL"��hU�.ڻ0�z��_Lv98�f�$��3�t�R�ݍ����
Ո ��ųI�{��HL�T�mmì��Z<P$\����t��vFj�Q �D����1�Zng��k0����4�͜�y2r��%����r���q
\!5�f��b;�?��}�%�P��K&_�5�2���V�TF�gN���Vݍ��9$�������3�l�`���H䳫���qrx�q0N�!�bHD�������E�[�>c�lo��r2Ĭ����.���{L<��s���4^�_#����$W0{i�N�_=�A8����x��L�7�o"$�/�:k�^i���G��J�2��z���T�L�����sI��sp�̕�Ž�m�t�6�h�sSH7f�'@��L�B��3��ߓG�H�_;kyv�?���޲�3����=d��*��hE�����H+킨�4%w��J+c���)�-d�������-�X��r�?i��"~�����qK� ��0��{����p֭�"3+C��֩���*����u�B��b��κ̦�	�o�Ҵ\s�Gm�BƉ�&�!E�$ʭsV����!���Ѡ+r8E��<1%�0�^�J֊�L��ܢx/�Y?a�4��c e0�~�,PEJ���2�6�aL�W�����R�������ϨTrk��a��(pδ�<jQ<�Z��ǈ�!�k�30�:/QI,c56�i���W填R��w��iB����q8)V�6}sp'k228��z�����Rz��ў����D��oPJY���_0_[c��\>���/�Nj��!���*0����LMU��Fr8.`�˹����F�N\�^��d uzg	�G���K��ݍn.����)���������CF~B����%�g�(pj�,�-`�d"u�D���J�ˆi�v%{a�l�nq�f��f&;��ؾF�\-i�{�C�1E�͂�s1�t2�����};����U��㪼�:�*@�=��<�F����N�[�w^��dʾ�$�1��	{"���j; ,]�1�b4Ϻ�F���2ܨ�;�F�ӐJ4��B�~:o�6P��1m���&���KqTE����g$>ߑ�����w�6� >��^N��+PcS��ӡTQ��'��x���>���J�W{I"��=ܐ��jϾw�^�-�u�L��)���I�8��D��߀�jg	(��J��̬7`o�gBk�Ꮊ��~ �s�h�R_��<G�޼���I4&�D��ԫr��7�r2�ӭ,�:��	�\���#��ɧ�Cє���Bw��"�]��mF��w!���X� ��Q�n�AG���sc����Jh��� ��[�`��݋_ٙ�Q)�k\(�*�T�>L7��%�������?KS�N���_r����1�B����GL1�������-����1�o{O����&
������������g�>�U]|um��^&?����M�0�N�'���SF,mbϘ��:ym�45o��Ѩ��͆�,A����7����ꨠ��Ү`u4����(��Y� ���[1X�Rj���.���4��t�1�����&��1ZtP�=�9;P
�׽�a�%���������a��M��yB,8��6ض8wb�Ȃ ���4�n�xc@vco�՗x�N�(B� 0L�B��yH(�+��]W�4�(�*��/�X�J7���gS�%y�c����]�(�j����2�N��!�~��N�qW��%�cv[ϜFE�D�?��w.
�xþ QTbE͠T�V�ql���D/�G�q�%����i�H�$�·Ġ��Isʦ5�1-��Y��Q�zf_IQG���� \�gv�n5���yKGQ���s*xI`d�� ����,�r�C��GC��X���~|�9H.�+a}0��m>+r�j|�y
�q:�n��d��#�8�Q�e)��`�P��v:>����PEVэ�cH_���I��)��Q�7]xOe�����y�F��x�J�9q����Z��c��e�w��#��kr�sL�佱�}�{���_07�%��ϻm�qUiJ�E�S]u�CB�8�+*����γmt �p��H��d�$۶������G���O��)���L^m��@c2E�1��pr���*�(�:o��Z$(�x��R}y?�a��g�m ���
uJ���,��ݐ	���
�d������Z~�5c�B_|�����y��5&����j'\A!���A�Ny��S4���,�,1䂭}Ѐ�WN���F<�b���$�t���O����� 
�.��E�R��]��f������L��*j��c��r�e���^�-%o�۔�Ǡ�+������j���2�σ�x�t2ʙ��$�@�|����[*��'��9�:���=0
�}92y	ǵf��^��O&��$��f�h j>ɴ�*��XNe�:�������'>�CΝ�͏%:���4�< I~�~%�i�~ I5�o��O9+&.��s�(�n�4�*�����pl�ΒɅ$ҫ`�ڒ�q:�J�'6t��70�n��9��E�M�+#7妗u��Ȳ�u�ݚ�74;�l6� #^�k�1�?Q�Mc�o����Or@��a�=��
Ǣ��$�jKx��*��z�>Z]*�%����I!{��Sp%��g�9�����M�Lƫ1a:
z�J"��~\�}�U���"� 5*xΊ<�[JK�1U�����V)�LY��w�2� S��oR>��ʨ�������I�1�vCf?��w��L�QrdM��n���6�ħj���NA�WFj�};k~��j�{��.�м���Q�+4[4co������ �Y�Ձx���T���0z%���2�S��q����K,�P���nD�ހL����p�K�|s�޹���MXh>d�T��]��Nf�%���Ȃ�7f2�	�&���T����� �$�� ��j������tG�F��:f��};��%�f$�� U蘭�ג�}p��G��7|���nv��n�[�!�mD:�:�g��ކ�i�o"ĤXq_kU��m�A10�[��l]�}���9�'�o���m/���Z�2G���!�C�ʍ&�,����՗�e��C��f�B��@G�k�i�l�A���5��k��w��n���h���c�׻��/�;�1k�`�5���	I��}5J����s1U��umV�Yu_�Wot[E�rD������~�Lo��u�o����_�MC���YE�MȄ�{��3�AqU���U����M�E�-��3��ﮇr�I9չ�u����"3>
g�,#�zX�X&yK�N$a�8tG���S�C^�0�t&������Q�﹁#KrOE���]F�;_�l�����x]s�#4��$�d�,�ni,ߚ�K:�M�#g��_� ��v+�^����f��ף#G�/Tf�g���CM����"���u���7�
 l����w� R��U��r�p���U�f�5<�������L��F�s�]���b�G+�����&�{x���B⇪��G�U���*����A���OY�k��kg��x�#�}�=�g7���ұ��gxƚVMU���R�(|�f�b�R�X�_\ �'�����w2�/�����uw�F��#�=�]�rA;<F�}�AP�[��k���b��YFg�ڷwv���s/��<C�^�Y	�Fr��,]/�O?|X�a��a�gC$�pi�m��)1V�63����7i��_��yj��~��#�6"H]DR�	��R>����]�t���H5�jV�%�ŮcE�2wZ�{�����3�톰��-��G� ��!TUE���\=�y�$8���� |3�׵��G�2@�E���>X�?�-��xH��8��]�tf�M�+,,|��?���z2�O|���MU1��cQ֛̾á�1p��P��<�^f��˵a�k�dL�%���bnS\̪V�eB&� �W�RX�U�߻&J���M	$Ӓ&����ZꢲaH$R�~r�4
�Kŧ)f������DUi���+�q���4�����N� ��l+"'�3ۆ�evh�<7 �n�i��t	v3#�KwzU��^2ܖ#�%��H`[��2HE�P�=qޝ�p�v�ȈiLrQ����\%��Q�O��Npwf}=�x��#_:�67"36�a�Y����+���E��$#?���-�+�6�F�~�W��V�� �ֳK����جQay��a��˅��#B�+,���ݴ�ґV��1��9A�L����;Q��Zl���[q\9Q%����=j�?+n�i����޸����9H4���&�ւ�
A��S���}���[����Lb�w�x�G��y�ܢ���\�����v��%��k*��0��A�m��t��-�.�0�$-7� Y	�q�����g�K#*�2}�މ�ҥ�;�]��	��XE�%�� ]�kOԥ^xTt��'�S��-� q%�g���UJ���tFw�m\���6w��8��+�t��2wG����4p:�J�i��������xt�fh�2�6�ǋ�5������sq!�)N�m\yt��hf�/�6t�Y������o���>ޟ>�z�y�C�9"�E�Xs-xL�O��H���po^M!X�f-J�8�W��ڨ��}^���׭\��Rkg_P��Ov/Qも��V�^Z��D���h�����*����sLI�D�T��@��	q� V����A��{��Y񾐻�Y�fVc����U� l6?��u+���~��.?3�	L�Y*I���QN�k|Q�Jra���?���q��^�Y6���,X�2���X�:HU� b�L"WӀ��$���H�p�p SYs�F9��m@���_~:g�N�߁#�Xp�U�hJ��i�E���[}��$�� �aZ��`qw�p'7�=j��Q�\N~sWď�]���x�3���S|�����_�6r�xA�c�� �@o�-�sr�7U*G'��{�<�ĜPN�-ύY��cM	�£�t	t�K���"�<�~������IIl��p_o�,�^.,
>q�k���-N�6&���{����k�m�C5����L��P�i�����`���=� �%�U�5ǩ<NEت�QS]�B�YW#��iH�Q��щ
��wޝ��2�@3w�Vqм��ÿ���(��t��#�1�M#k*jJ�l�8s���"��í��m^�g�$
��G�#�{.�)bK=�3��X[��ǔn��������8�	��
��&�����VN�Z,H�K��Q�2;=���⤜�)��ٴ	k���=�6���F��u�
�'v'����U��F/ʄ�&t�aՙ���k����\�����9��Ƚ~^�F7PQ�|m���Y˛[���C���?(��m"�˩	��~�
����6a�|EZ�@:�c+�ݜ��38�9Hi����`�t���{Z�5m�����8��%9R�^X�ϩ�w�9�6��Up~�ޢگ�k>�����P��x�!]<84`��ou���Th�!oF�~v�G"�to�r��NjV�J�C���}	�ڥ�Ѓ�振��]��wM����/��q�]4�ɉi+�qƷɕu.�\��k>=�~w����������1�ݮU>e4Ժ%��Tǌ���ґ��+[E3�a9�S�S�(,�t��rJK;����S@�.vfDM-W��mb)�	[D�����sm��p�4z�R��O�^��P���:?��hHGJeuZ���G��	&��7g�}Vl U9�s�g�`Ǝ����G		��ي�T�G�M�?@����-
��_�A�Ɇ!y�H��-x��R�nL=�e���#�|;v�p�z�-�/�o��R|��
AC����.���oYC�d�KzbX�G�:����l)�/�W��rVd� [F<������'��g)T	�$s�=�S�m�P���\:q:kgO�&qD'6���g��������{�r��W\Tѡ���8�ëm�6�L+H�^C/�O^l�	�-���S�^�`0����"֐�t�~� Iz����	,��ri�@��w��ڹw���|�Y� 1�_�uP�P�G�!Z$�L�} �¬�������|�_]Hy0�7'd$�� ���8(��/ɉQ\���������X��I�D|�Q C��3
����9_F &�%�:��O�ٚmK�\(�77��SZr�I+��d��J�o�����yoQ5��}9�� �;+ƤZɹS����_��1%��@����]�t�U(�j��*��=���Lv���|<��5��:<�'\'�����A��f���Й�,��Ƕ�R�b�$��B|��"��)�庪'�gS��V۳H4�4+��H4��uCǴl��PP��pa� �J�|Gꀦ����,Ҽ��)`[�_�;X�5��nX{)�Vf�g�!bР7����,���4R���`���W7����QA���\��� �ZA@=�^������P3����j�<Q��YYY����z˜�r9&s9�����@�-�꛲e���ޛ��sZD� ��O�'��Kq��W�^�r�-X�.��.Nq�?ձ�L#��M{��=�'4KL�O�����>	Q�=��Q
S�R��֚LZ�K��z�0["�&� i}�3r���JprMt]����м��C5n�|QA�ơ��q�����0��O�.9��:�OT���~@�-�,(3����aY�ï�In���A�0�T��P�:�S��QG����zY����y	L==���F�v3�3�iwM,�a�m]�Yn.���r0�1A�
��,��ؽS����߽M������\Ph`r���ο�v�{a��< `�5�r3 ��Uՠ.ι@E0�m
w
AQb��C�b�nԃ��Ԩ�Ǡdc�m-5\+z�j	�费X�y�o�n�S�l핀�P�����J2�_ͧ�&8�я����y���KYM}��������j�(�q4m]����Q����V�~ڀRK9����5���	���5Ch?%a�� eO��~��+))� !��:��;�����fz4h�VQ�q���nP���!��*�>�����.��j�ݺ,�V�XHT0�8��GugL�L̙b_�~���xH(��>3tK���e�bɀ�C���c��x>E��<��A��\���Ur�,�� '�*L�!o�p�)*j���{��S���A�r1Z6�YHKG�pK��Z��E0�d���x�X�Vli���~ߩ���vm�#;��H(&�)�O�ɟ>�z��|����Z�0�,ݹ{zՠ��
{���v����w���C�@���*U��<�Q�=S�ߋ���K���9>mJ�h�p:�`�JYK�7Q@�c'R�rxz��eH����j	;�LP�v�]���/��<.Ni"+��:� )h��ZA���Q�>��(+A�_&���I�D��Wy�5��ȭ㧈��-�����#�ANA����Τ�t��f�{pC�1��7� �8U�F����}r-���/�clio�/����特��葭��ˮ?��[f)�a�|�[��Zvo)!��+Ç"b)���=�PF�u5��W��]K+"f=M�9��߭~J�B�dL�A ��X�V
b[���	h�z���V��B����ֆ<My����ȇ���Ǥ��xɅ�qIF+
� !(?��'�5��ak��:F��3�qi����5nF���`5>�/3���<�qY詞W�{>���2#�U��۬��F����c|� � ���,���X�&�ס��Cj�M�]�`���F���hX$=���wL�C4y�������{��u%=��`���ap�H=i��'[ԠK0�CS!�4��l6�\�����ǘ��O_Cmb����1(���|����<��6X���n�����u���\��D.�1%�D��	Gc�]@L\�N��9��uV̋'�\���?����*6�c(kl�> ��,�B���	���V�5�����'+\R{�j��.
�J���y�r��-����b�LmF��q{�.6����w�2NX)}0ø�����Y�z���T%c4���N<�ΩF3Cn�D?��Ԕ�P��i>�	)�7ե��( L{�Da=^vv���A��p��諧��a���֛�[�~Fh��z���û��qKvU��[vB������̓���Z��8^;)��1�c��99� �ȐV-�ɍ��5y��C�^|0�C�󊽺S�y��w�ZɒJޛ�{�XwV=�� �m�>z�Xs�<�v��|+��>�Oƙ�������1t�QT���pu�:�|�)��"v�=Ey1;ZʜQ���t�ُ�T�������(�v�Q�����9�3����B��h�C��n�uPAz ��ggv�+B�D��?z�`Й���!�E�FB?�F�����Y:�����"^"������rĤ]��bI��N�t	�I�<�U4}E)H�_����a�#������)��Q�41��V�J���D
d�R5���נT�kE~?�:*=%[�) XSed�'_e@��C�J�^K�@���,���&t���1li�se0�9��ٞ�Kl�,�Z9�U�r*�[7��a�R$�-WV�őG{��U�� ���6ԣ+��;a�;�?/ͅ��j/�;E .�vE�ȹQ��Ŀ��*k� �3o�F��g�a���hեc.C.��"m�����-�2�����3��g��+������0RJ�d��f��#5{�q/A��!l���x��˃i���\p#�n�� ��ͩs�?
��HPB5��B}j8�AT*��)��1y��82�;yV7J;�?'j��vv�����-�-�2����G�)6���:wsC�,Q�+��@�J���9�NK%P���ۤ��4�?m��t��RS�^%�)~����.�0��Y��E���?H{^���S��_<k+�ܾ0�.�<A��_s0L���!����c�lhdKa�/�tR�aK���%�ԟv^���6�U��U^5�ey�h�� �rzٟ�#���-ʞ�Ĺ+�������T�B(�h����G��eZ\�%3M��ZY�'&tX$��`z�%,��1��;��h��&�F[1���|2@P����Os��$�@ŝ#3�����V�cA_$HW�VpO^�D�Ǟ�R�1��N�h�5Y�<aa'�P�	�m�4�~��:X����`��Y��]����kj��%����:���ȷ�'M��&����jt�ٱ�z�O�D�c�$�\��+��m�;�ɭ�^f�F,e�1��Sg߄K�*�
�]��N�XuF@=�HfP¶�#�6�������D�
�k���E�������;kt�p{t��7�f>�Q��7)3�l%���c�Ⅸ>��V['�W	���TM�ŧt�̢���1J%�xә�Q'u�ʠб2��E&&�t�kM��uT�Ѥe͢��Y"?�BM�GŒC�@� �2A�
T�+,"󚖦	�c8d��� S+H����?9S��@jݲu��s����_�Q���"i#���(2 ��ص'��&~\*����s~H�����r'o�`B'�B �X�+��m`�5_���<����R}oǤ+�iC�j����}LZ15H��ԭ��"���Fw.���v���L ���&�.�A8]��YDW���C��ч���߃f"�PZ��D5J�n[��F����d7�읕g�b��*��Ʒ���eʗ�ہ-��Ŵo0��1\�qZNl<�)h�}Ju
�&��N6Vꢝq1���ۈ�O�i��z��6T|�vOe�-��Xf|���ժ�"�u$�?�?S͐󤕝"&���r?�u��[P�z��Zop;�� �M�������3�_�{k5Q��57�5NYpA8 �<�[<V�0��p[o��͝(�o��=D
8�!&-X�.I8�+Ʋ��d��܎�fRZ �����z3�~Yavxg��a�⫩����,X�H��NVǂ5Ê\�xN%~�ڲ$S�FI�q�]7A�!^��+qF١�R_�9����Sۃ��Sрhð���jc[�����ͱ�b�A�m�b溂��4y��P�vV�X��L�8�-�f��w쌼}t�F31��|iPͷ����]�$I�8�����W����?[eY��sA~_�ڷ��$nJ8'�h�ͳ�����FL} Ag����5�-v{i�1�9���g�*s�)�l�� P�I����7�v�]g��}��y�����;+\rZ 7e�̮'L*J-�}���p��T���YV2�ht�� pw�(�j�;�Oy���t׉�e�֪����A�U���xّ֚�oc��>��ȹv��
72��Ux!�����lޜsHA/�4�BR1YP�䦼1��w�ކ���>�p�RH1D��n��^>\8�L��e�Ȥ��j?��`�ݠY��N���Jh��1����%��&��+����5Uw��a�s^��L��M;��_c����_�Bʯ�Ҷ"��_\���R!�;�*R����AVVn!��`�����h��v\s��ۧX��u5�nQ�oH�*�Cj����8�I!��8�j���f���pR���������� w�V9&ߘ���nH&PEd�9��������\2~�+I�1��ӎ4�^+�Y�/Z��H�|r�!�ժ�ϺMl~��ݍ�A�x5���"��0H�!t�cO��K����{�k/v.��9��h��N竅�*�����O|(�@�.2F�Ʀ<#sE�%�H�K�>v���'�{Yc��ǔ���ӑ� �U��o�vhAmx	[|�%�t���^SЈ�ޙ/MZ���S��	�x�,/�\��TVi�>>bp�������u���|�V�fV�Tb�<������e���#G�m'��Dw��*�1�аG9iN'Ԧ��[���v���a�G�Uξ-���1˩�7�J�/���1+�3��TD�!������(�7���s-7�|&Ґ�]�IO2�,�f�aaMx�2���خA��i��:=>Ŗ��x'��U�EYJ��F<������qS�;���g�a;��2��n�~,c:�![kF캼�Z{S���U��B�����.)��t>��F���E���R�)�9�p��_��2� `W6lHN⎪)#$*����b��`{hY	Z���<���uGr	n�M��0�;����:����2̺��� ѓn�#A%X����+w���IË����b�����X;�^i8*��,�<�y��bk��Њ%�\��~�{7�S]�/\|��L;i���РA���h�ŷ�u�_�̲�X������c��l�7f�S�'���75Ul)��"�r׆����K�'H5f�>����I���u�e�I�c�����)(�5�*B��Y�\X앎F[�w!�K~(���oڮ�RF9�Su`��M7���>�
R��t)`J���`��mT����j���5A�OyyO�Aь@[O*A��;�t9�/�xe%�`@s�:�0j�h�@k�mG�RM��*�`䂮���T�����+���%��}�SS7ҠX(�����;�F	��ۭ���r9��;d��M�v;^��>GqI��y�A���i6��Lj�2�MD��7l��l�6C�y��IP��=<-�#,/D�|�*IԶ����>S7g�x�@���	�e7�$� ��t-��h�`8��Tr[�BTDcMthx��*k\omo�}����f�)�Q�i��H=ɗ>ag璅%v?������h�x���5����EXb�?�*�Kv LR#M��vF�afMW|�
�f���V�	X]���ԕ���w��D��]�����6��[u��4́c�7w{D����ڷK黩�-�$���^�PJѢIщ2BmĻ���7.&;���&0D�d���e�C�?�b�՚�]�ٴ����>�m*o��P�Z��h���lRY?�6��<�2��yNu~b�5�%������ �(�� һ���c�����'B׃e�s���P�y=SE>')&^��8i�?�1+�`� q���6"
�+*5M�vi�I���D�͵��dǇ�^�>���M4���JtS'�ape[���@��Hi3�
�_�.��9`9�yc��Tb)�h�ş�~�����='P����T�J�(��~�/���Ԧ��F+OVl�f��lS%��c�	�t�s�q4�>%���W��݋,�x�؇;EuA��Jؘ���N��U�`,<��8����]�7�|'���rSz�c�g��~�Z���l�yh��9�WA���]T#�$ZwC'�� �3�r��ab�ٔ�g���A�x-eؔ�T��[�~�EN3���'0�|��)�C�Wr?:N��@���ERp�)��/���Ǚ����=W~����0"�7O��n�@>(M����0�@�Y�h2���lyY�)��2��pD���L�2Q*���cp����OݦP:�b��8"!y�홷�>���f1�$��q����/�C�8���q�)?^�_�BYq�~��}���G�!����+��5�z�Ф2�n<h�n{�3�VԴ���� l�"���j���|)�a�6bgV�ԡ!N��YD#I�-ï����d����H�j���h�>��vB-���GM|S��h�	g�8V�2����������V͔.�	��R�ׇ	4�����Y�,�-U+o�K�������f�Č��b��8��]�~���V���pG�U�~��M��+��#��c�'��t��׏�JN�<�gwn�����q�mB�9,4��CHU0��b��溝#���pX#6�}�����j��k��~;=��`D2�Qŕ�����OΪ�I�?="NP��s]%���ɎO5������cã7O�UC6ɴum`(�e��	!�+ �u��f>%�� 8Pp�#Vx����:u#�9w[���8��@��C�HhD��G2�E�wU$-p��D7���Вܛp�jb�������9��"
5��g�}��c �[b�k��P�*���������Q�f����T����H�QH΍$X��TT_A/ꈤe
�F���f�������ݢ`�����I�o����|�����ۨ�CHQ�ϸ$?�}�MO���7�m�� ���OU��z�l�.c�~Xl�]'��sE2y�;�"�z0��\b{�E�Z�X*+6�w\q
��b�͐�߈!��,;B�6G\�'(�]�lV�l��qBЉ@>�>���\~ʦ�K,F<�w��_�2���Y�X��Zj{g��{O��2���=�mY�[�X���g�(�z��F6��غ���A���$�"�$��Yu��~�x�Y7k�-�(��b�z�������L�{]��(L�n!�����M.}�H�;�*1{�� ��H�c2�ʁN~$M�XT��׷�IHtGD�ѡG��m,нAo�7����*��゠���(��#�Iδ�j߹Q��$	}&r�i3�ٶ'�f�:����+�6V�!��8� J�{va��ܞ�9b�s��	*��Z�W�9t¹��_Y�N�Q-H��_w,K��C�!(,B���/���n�5b�w�A^`��A��"�ՠ�?�gq	�6#�v�JD�sk͓&�������c�z��1о_�?40k�D�y�([�v\�D2QN���� }�	�'��D�W89/�OJѻ�y%e�89b��?P���~z��6c�a��>�ʍ�#J� �(�.���u)�|_��om��Y��b����p#���g��s���yM�BiH���o�bPʧ���rh�{� !�F�'�%�@�}xw�>_�������rd!B�1Zӑ�����Y�؜}�%Z�6ʩ�r�uL.]q��{j���ևT}e*��6�����0���2�P���^����w�DPh����� ��G�S��/l��#��H
6;NYz.P�?Lc����BZ�\��f�U	��%�6R*�s�4��$uM�b5޳��\�qȬ;8��k������'�ixn�cZdG,B���9V(�$�4ԫ$<�h��W@wu"��܂Y@B�X9������t���;Si?��1[~�`[�,hY�A��M �O<5o9 jrE�	�Q��|> ��Y#���$Ѣ���$��>42(ղ[������|�����<���@&,Mh���f3Pf5�����l4R��:���Sr�My*�B�ŷ�]�������HYs+�_�(�{��w���m�"c�x�4�!A���)�� ���M��0���pf����D���+tX�$�3�J���q�� R�*YW�� "�{��/�(�=�ҩN�E*D�B3ÊL^u����qU��2
����������+/�����D�S����1@P����	�`#��'�RtDbĵ�k>��0)�:����ZX3�]��L�J^v��!Ɲ�F!�Eo1#�zr����N1ָ�k��BS�ib��9�����Ђ�	�<�X���n������4p: >;,:�M��}3'_w��B[���ݺ��̈́�"�q�Ć.�e��Q|����Q'f����>�C�BFyU���2�X%e8hҭ���]Z<���Ռ
�}%Ӗ��䩇��
!3ۛW}&_}���}RҔ����z��J��}t��ǵ���FÛ�%����	×\[(�Q����%_���.N�)���c�!�gc��[J#F�5*��<�����\[��ΔIU�ٕP��*2Z�<e�<lf.�ɼ��_L����VqW1U�ق�<�\Ou�Ї�Vp%���X�[q'�8��E�@S��r�"� lۊ	�E�[���o���<$А�"�~1�zRP�d��O�^`��]����q|DH�C�E�q-��{�y!LЕQ&G�3I�r�O�
"���q8�����i�+��(]��$~ɣ��Z�(vm���"��T���*�`�3G)���p�X3�+��$�Π~r��|��VVDj&�W�ynC������m��\�T�U�>c_-�z�H�.( ��I�$~��n��*�1@���V�z�ئ?�#��z�Lg�� |��|��z��ËHC8����;+J���m W�K�Mk��aۛa��4�A���IS(��Z�� E��W��nB�2jY?¡�v���H��zS��t���_W��iqnQ��N_<=����� `�v|p ����V~�i�_BᏐ��W�0���C��u���)��FH}�Dk��H'�H1N0I��;LhZ|	��������~���:^��q�7�	�JwP�KV����f�:lt�>芺axz|���OG��+r+�+B��P̪f�j��'��ro�w1:J���I6������ 4���d�Ś{���Fԩ�������'���O��u|�7�u�dk�y晒ib�f����Ki�d�����#�i�2dr��
4Z��j�S@ԯqGw#�[y�]ԈA�D�j�.{�c�b��@`@�k|G���P�FQi���ˈ��M�Q%h��{�r���2��X��W����4�^�
�ġ���\m.���sؘr��K��c�أ1zv`�.��C�i'}'���TO�c�>��pk$�蒮�Y���%8%��~�z�K�κ���ȈW��T�#
}.����;��
G}���6L͕�8��<�=���c�ex������!A@mD �%m��et�N�~����蔋�ZM F��ٵ0ɽ��pu�����!a�ʳ�;mt}م9ؾᶇ�����e����+�
�T��@)��.!���y���n	���ZW(Yכg8_o�Ik��0Z��+��G�URL������{->O���ꀭ:����iy�Z�r�n���^ �l��
�1���"��<�f�h/��sa��p�#9.
}�$ � �gg��n���-��R��<��Z$@�{f�{5A��:��q���@�����:��5�
��< i����/w�͛B��,8$B��t��p�z�۷�;�"��~�.L�-U"fB�|1u���TX��A���C�콰��^���k~&�Q���)�笶,�<#�0��RWú���!i}G����iC��&B=�	%�� )�ִ��~:d�]0�$�ڻ-���X�BF��D6cD	�l1A+6r�s�G��<�[�*��Z
!dm��(+҆�P�NCN^��IDY������P��e y�^�G�X5�nם�j�L7�.UGf�;B��prK-~�ao�S��W�<#7a>1��d�:��ⶏ��#}H�J'��T��:��Ce\��)�%��
���$!v�R�R�s^���v6����j1����M��vD9���r�_����z3A�_b�K�U���K��N��^���`�U��Y���42�g `�#�5�Tt�V��(G'5�4 )�	�)%6`�~M���X0��q�Ğz�#�0�u;�$��'�a�(B�S�|�Vu^���'2u;5SX!_�>����;�8�q��+(`}��[M�#�e��W�e_Wo��h���v/ Nk{rC2ֽE�at����!�4#�j�O��drB��4��8��� 2:�b}��v4���J~y�]���}��b�y���Qfc�r�.�%�g����n�ܐ�� ��ֵ`�Gg�q��ع���xΖsxz���ҫ����ŕ��LͿ�>s�T_�	}�r�{���2����;HQ���׊~V1��LLx�X����F���L���q��+�XPsbjv$�r�7���ޢ��gĤy?�7�#�o[V,v&��xճ�t���G	�T��,3Ǻ��5�(Q�����}[+[�P��J�J�Q�G�vb��#�n>6��O���
~q��Uof����!N932�6S!}��2]���Ӑ��h��0� �r��X *PͲ'� ?�ϔ^e5Izs�e��k�,;��o��p,�0�I�r��8|��)r��]��p�#6�� �W�����T�!~����vھ�Y>w~��ר��Q�I����E�D}M�"n9f��  �5�\���.�rZ�[iDP_�y0�z{
����[VNR�}�۰�O��~�)K�/�P��,1�ו�H~1�'C9�������� [L��Ƨ��'�ۄe=��O;����Ȃ�p.yE���ԏ���HM#⸋������Y}D_-�iq���?iA��;�{B��"��z�H/cj S͊(�;�uU٬�a`_����|�D��"cݜ�r_�6ڶ�1Х�-]r��>C*�9V�ѣ�$��� ��n J	l��k���{-�3{�����$紞�w. �D �ö\��~ ���Wʾs���Aq����xd+\�,�۪k�&DҁQH($`�x�q�����������n�bV0��$�}c��Mi������}m=�MV�:<�;���4�:�Xl����Xx��Er�V�,�|��z���m����fY���g���A���w�z�ʘ>NG��+�
�ak�:������e.3�'��B�5EhZ�T,�5���Qen���c��Ċ/B�E�g���?�&����#�}�+�X��t3=�վK$��j}6N�]�f^�pH�,��
����F=�u����K�ס�6�&�u�G�ܠ��䜫~���p;[H�1���&���^�.n�p�hۤ�'��7<����,wZY��̚�/��v#Ө9 8q���3����V�w-Kze�2_���k�5�N��j@���o�[	�o@�D���zsE��6��I��B�n%Z�?B���� ��sG�e"sRA�[O$ׂN�s�F�D�d�V��!��x��y�s�W�%"�+)�XQ�r�j����7�k>x"��WIe>a��=B��7������8���4��|���Q9xz�g2�wȼ,�zڱZ]�4�7_�����O��|�J����k�oX	P���~V�m6�����7�v����6�~O�L�i��7P}�ٹ��]yj�����DE�a�ֹaP4��.��=[o�#Jz�{!��T�ظE� �����y'Qa����*��u����u�
H���z���zܟ�uJT��W^��a���߲����Π���UG����5�_/�e���j�̚-N]���Zmy�tM�&U����7�e������c�Z=!��PM\�Fn��.}'8�x�<]x� �y2KF�Z���Ti%!�un�>b"(c`N:h�L�����s��%CH�&HLv�[%�A����C׎=�y��_�ah�tjdLw���7���"g'^��B����a�RE�̿�?�**т}r��X��Y��)M7��/�-2v&n���D*Aغ[�Ż�4�	�c�0�`ޥ�������e�Ou t�j������s�J�	}z``������/ң���Z���݂ı�@��Bcw��~�UlV�� �7�Ꮪ}��wmtSAU��)�|,=�"t�~P���wB�D�v��U�iKH�P_��M�[��\J�0:�W���=�̗������6O(�����;��e)K��>���^�&a��ىe�^Jy]&\A�c<(?k4��Q��6^
ǨW�z	4ݘO�
B��D�	�Ȫi_��� ����8#�H�3���������<>;�:��J����\�5娀�MS�m����'�
M��;�$��\�\���2��-�(lz���0E��;�i�M�j ����b����&,�Z�C��׺_���$���X�d}�[[3ͧ�$��xN�Xؔ�dU�*Fx<t ~���P�' x@?v������h���1Ul�}=/���3�'��y�<mZ2'P�Wԧ�+d��Z朩X�%f:�y�D��کd��^�Iݟ������K��y,Z���[V�Y��g��M��.?0����XHq�[�KSw��#ݥA�e }�B��)�#��:�ڴ�ԧ4s}���T�I����R�Ò�̄���ևZ^Dj]M��w��0j�����3�?H89��͑ƵCD��np'z�X6��P�1��=����נ����8H� c��[��V�� �M߿k�$�|����XO��J�<� Zr�ֱ��
6ʏq<�ۦ+��1Q��b��1�w���f� ��4'���e�h�m����z��(����8�Z�&@���vU�߉3�T�8��7�;Z��8�o��g�֦9p�������K�^�2�,�W{�z����]�g�=m��~�-��f_�P���X�2!���9�NI�d[$:h����^-��M�Oj��aJ�4W����F�������������Ã<g葜exCM�d������۽0E����:qP�VE�"�oɓ��0���|��պ�!��X��H�h:M�����]��y��]���rg�-G$hY��k�c�䛆���zw���o��"�S21Gi^��}�]��K���
wPEH|�-���F���Y��,��a��\>����.�/eX�i#U�^�\�T�W;2p�\�W���Q����%��cZ�����<�s�˦g��A���ǯ|���l�zK�S���{o|�Ֆ��,��Qo@E�m��ޙ��@@��b$\B�0h��5��&�!�tj3�E�u�m"(Ą2��u�X!�����z��V�u��XQ��k��} ~����i�'#�,)�|ϋ��aH��
��5��a�����%���0�%(\{,n6@W�~A/I"�l *�(Ad~%�;���	��1�x���UE�{��.�p�wT���g�� �k���Ei#_���r�V�~��v'7��$xL{,[���X�f�>)�͛�R���{�ق+��{�6GA,,A&�� &8�em�;���^^���~��2�8/�B��ْ�J����v�k9�s���S�%�����Rǳ��ƍ����I�x$sAH���(�s��l����F�da<�uH�i3�	M�y��K���y���=�0��5�����N&�N�Ed(���	w�Ďf2���̾9�F=���d�z��Z��Ԉ���1%3��{7���&��������_k(�e�8��??m��d����͇3b!Qe:+����>Ή��t@��5�8��Q2�����~��(Ҙ�{ �%�Ȧ�5!5ؘ�9Rw?f�7�\��p*�֫���/��D����Z4v$[#��(�UGV�o�bա�[���d�w�j,�����v���<j���Ֆ�����Jq���Hm���ŧ���q3�w��~�>��YB-�L��ï��V]�pdIl�$�����{�X�=8�X��x HȎ��{�eN*�
���f���P%4ez<��Ll�ݪ�d�r9T/�r<��2� ��2f� ;�Ƹ���:?l�u|�&�Ċ�*��\H]�@P��	�F��φ�ڒJ^��d3�沭���E�Gp���fI>blM���䵱䦖Z>��d��"�F0a�]#dR���������
v���i?>����*�.��	�yX���IR.:�gN�v=�v�qQ�D�>�܋��?L�gJ@�ݝV���Z3,�������H�0���k.p��{u��0t-�p��p���&��>�Z����۬7����4rbn��Dy���R�iPZQ�&�R���7) �{�W�[^��;����P%P0��R�=ULP��s�}��l��<w�.1�k��lo*sefD6�r��� p������\N�:���85�3�Җ�x��B��>d<�P�bVۘ6?��u)xqv ��{���ׁs�," �,���GG#2ȧd�{R���Xi�Mt)��A�Hc�~�=�J�Eb���p�����m8$�;7�4�x_1�"�j�l�4��x=��͏VO��#�5�M��p���+���A��v?����b��7���y'�4d�X�%����,EM��w< ��	)ǗilToL���L�L3����ϕ�h�Z@o��zm��������tk]`�	9c���KZ9~q��,���������ԛ�1�B��>릣2���!9��G�yd��L�d��8TC@T ��$A�[|:]�~�૵�9�C�P����"
@�g��K�����^N6��_V�
��^��6?!cL����2+~�2����٨}馭l�P�>C8�V��ҙ@�l�*��Mn�u��v��<qc{�6�j_n=��Aњ����EJ�W�=����;bO��n���0�99�-��S��f���N�̅�O�˲�y�"���)�����_���ߌ��$�a�u���~�;��|�`�7x���a��irlXڞ[���8cx�M�V�j��rs���N-���x�;��~J�L�Ō"�|�b{q��,{b􁌀ͬ�dC�k6@r�,�7�9���1��fx��'����� ����V����C�K02X)p�h��gQO��ꑊ�yqǁ	4;H�tCk)[��,Y�0��}?^���
'�yz�|R�6#z"U%8��ɇ�������)8�QnUt�����8E�zU�$�U��a��D�o����u/biL�{�<F_8��}�-u����۠�,��\͛�2A�����-��Gj�)��"<%x3Ï>0K�kbl����=AH�
-��r����o�HPiF]�>�3���#O����Q�)�g��I�z�|c�kZ�Y�ޜ�,y0�i�
&�g1$`��i�VL�o�`z�0�B�P�`䕳u���H�T��X%��8���h5�G���H���|x�G�h��VD]�5�����6��VmJ,\����������_O|4��ș�{�u��"ʖ�f����LcEy-�Ӧ>�>/e|��
c��ބ���u���Q��A�J
�٪�j���������,+R��x��u�ȥ-��|J���t@��Hԗ��pY�a�kk|�X�(d� �3Ȼ~�x�� ��Zh�	�(tN��� ��=ǋ���MȂ�: 'xs�ٽ����+���+��7E�1
!�@��x�Q���q ����hx�.D�L�����S>�t0��+�!��Wm����ڗ4�}n�)��읈�[N�m���eà�ıK�;��� ӯ�x��]hơ2`඼k�'�� 6�uOx�a���r=�ei���{f�u��Xzzɦ~��eF9�"MV4(�����Q@�n�K0E=���qF�7e�N`�;��U�������bk؀ ���9�΂ԣ�L��3��8�g�hZ���؈� �%H��F���@�aV
��H#�J9���:����Kᴾ^ܭ�8���b��!�%�w����@�3��G�$��ITr����'� x�K�ٰT�0lVeuꭚ�
3�>����c��,�z�BuAr0;��z���r���d�t�2�
�_�Nyz���`f��<�g��W����i��@���P~��Z�_�[�6�j���'�4\����C��q�S�9��3yS�OB(�)��$��	�X�с�JV׮�Y�f."c��D<إ��(��E_#��{\a(��m���$��a+��xɰ(��4�rc���i��������<������+� �'����I/'��]Ncb$R3���z���9G��֦/h�����5D�PE�%�av�Lc��c��5��������a����c��T�z�ݍS�e�����){X6�у���8Xٳ�v_��F�t�ZSö�*��$�G�^��b���XI/�5T��o\�B&�_��z�qF1,ۭ�Y��~2\c���q��>:�cB�=�r+�(����(����!�L?0�S1tH��m�\[/
}����,N��Hۉ�)�%<r���D�G�9�B.����3#Ŕ�1C�L��l ���h}�F�P�>�W믝�9V�l#<"#�2��(�[5���vd��d�T�qNӬ��*'��m$u���$�+0���)���ٛ	݃����1"E��4ǦeA��'?�ʙ�|�SK]���gp���Eg4����K	r�Mt���w�R}��LzX0�����	�\&9��x�"WS=O��k��6�<�����Z�cl��m>�Q_�G���䊩vU�
���vZ�R�`��SR�J�tݰ1�;[z �w��BȌ���M��g���F�S_9�@*��͝�sZ�����2���v��FLЛ�qUe�o*ip�<1�~������d���E�t�؁��r�!�����UW�w;pQ�0YPV�wF�Dg)�7.y۲��?%d���FT�u��l��@ �f�dx=p��ts!�4G����*r{8i�W:<r�Cryctb�[U��@�~���x��c��H�8|�!_���-8���o������C�'�e㺫=SE�k�f����mL
�x�4N���ݛ����t���|�g���]����	�,���ݛMe-(���dd��U�Q���n��5Ѿ��M${�B��Tz����_�f�6����h�w��3ʺn)"���� �Yq�y��ڨ?�	��,(ػH��$�"YPWb��1 B�"�[
�2|��'u[�P���YYf��o��{�H��9 PZ�Hl�n��1�/m)��Q��)��X�Aq��)~�$ص,��n��I�(������+餄̏IF�z��븉�gI���@�������4h��N}�~��87�亙<���zl��DI��U{���wW��wD�(���L�@!c+�UX�	b�,=�5�+1iG����]/݌Nn�2�.U�! �ԃa���}�����쉩�#��L#l��j �l�Ebwb&����9/�J3�|�x�n,��ɢ
�K��d&����`0z@R���h��o9r�U�P��$�H=����D�>���ن�X�ݸU��\�����r���Fn5T58z�p<##��P] څ�@(r#�v���� Ji��G2�vB�Zz>#�9�č-�g�3*����X��$/��s�S�I��G�A�9�T��� ��Kx=�%xuT� p�,@��Q��mx��ڤκ�Zws���x�SA�;i<�X�d�qA�ˈW�_���WA�HD�|(�/�Z�V4����[��&.P��a2�oo�E�%�>�s������t��ͤl����|��
�Ѥ���ک�T�"P9���l@���e�7�eS�4��̩�SD���2sK!���x��_�Wb�%�֏�s��p�a���k�b5�Nш{�A�C(�y�j3W;��r�)}��9^�e1�
h�鈣�����]��<�G]�3��_R�p��ֺ�ů�~��!�u1{[�ͱ��nm �_��f9T%�}�g�2��8�a�9���9hd	�.ەZO����[��C8��C�s	�\�7ڱ,ya"$j,�h�s*K�/�19� �]�l��'h-{���g�ڴP�ɹ=��sVAᕷ���kȯ@��
gڐ�Ӱ�t�PD+�?�]c���a�Cuz������夵���ҋe�4��?���8'� ���]��D���3`Zt���M E~�d�,���`��Ee�m	��P�h�r�|����T�^ W�@f�&}*={ϼ�����J-eH#W#�PGuU�o'T��;���u� ��-4�H�O�ms$��N�Gȑ�v[+PZ{P7��Ѻ�S9���AZy��moU �YY��|���#�j8�y6ڑ����=2���2��@ˠǸ��Z��Jq��±~�����8V'L���y�e�r�JO���70�Hr4j�:�K_�(�4]Ҳ��?��,�Pd����Α��&u��ƨ�d*�k=�t��D��	m�En�*��n��U|�4.\ZP`� \�¯���h�"�c�p��p������@*���8�W��"��r�0�J�"VkL��������C��FMO��J	��ʞv�	�Vҳ1�nLrn^V��R���=��گ�~Uڐ5�:��v�p�Ӿյ��Bʡ�۱#��	 L ��&S��r䷒$6�=��%�E�6Q����'�C@�B_��픏�v�Y��'$���Z�ȓc��N���D`�O������ q�in1EI�WQ.5eU4�b�*��{��=��I��ǫI�GB8��a<�?�|$�w��!.u{�6/3>C�S߫�7o@�1��f:6��5Y1�/+�)�>��� �H��حl��d+��~�T�F�Ǻ�R���oe�_ʨ1��z�^��W)"�qa�*�6���IGX���6��]��c����}4+���j���ġ.���8 ��P��jh�����U\ҡ��@b��o�1�$���0�8|� o%�6er�=K�l��Տ���F��})$sƃY�ܓV��>�o[o�|�72yt���w��B�ع�}������t�C	�aW��tF.��k�yoW���v��9$ (GÆ�.��"G�D�Z�RRD:��?]�H���l_P.L7�x$��[�� �`�B2[��~�z�S+9'��r����1�� �O������M���`�Ӟ�|�c�wl�>�C��Ӂqج1zj�2��5iҾ{l���x	b���bA����K��=A��pƃ��w�І�����Ȁd�����۔�ּT�t��#ϰ-���䃯���7�������w���d����0��5۸J�ý����*\�ԫh����&vro�J#K�cA�|I�Nm�׀e &c�R�����Ό���6:S�&﷢������P���ȁ�[`����ڴ���۶/:�Em�2B��w;�o޴Z�"Y$���#G� �=��>4]�d2�I/З*�
��UJ���<���T`n�zu϶P����I��'�����Qn���-���[At*$5,����?w��U�1]|5�횑�k����!Ť�} 
vjP �>�-îƼ���39�5
�R/��]�'�Tc���:�K�?����;['nҰ&lJ���a��=���. �}]`��-!�
�Ѻ��A-r_��A�C�Hr����9+;��;�[���}$P)����F��2v2V�B���8��fJ��
�O\bd7?�����o"�?
�1�k��J<ޙ㒩���hsG�YK� ��o��	���p˘mn5�*��2��@Mw�<S4Z:X$�ňW�e�������z��{��������h�zƦ˟�\�m��� ��M�[�Z�ﭲ+�箂�7a��w� �_$`���f�rH�$��wtIK�� �j\!�v��έ�������ruKO�_���b��=/"�Mf�����)��K��c��H���H�=��\�5�>_�Kؔ[�qu��jg+O�G�����7�IG!��r�&(��k��������y2��i�:�t�j���)�_���Ȓ�%��E}j��=�h�r{�y�AԈGu.g܊Ȳ���6�]��߭\ů�e������_��SO���ں,bR66�&�`:��m�+��H0���V�0���jA�Ҽ�^�"��/��=��t�ӯ K/*^v�g	=E_�f�)t�����B����)?���3~�
?|������GU�^m�Lc^A:�5:xػ'7��?�Z'�-��s�M"L�n]���\�R�)//�Z��H�wG�#(��1�U�y��0�ӡ
�!�� ��3�<q�b,�7&z.�9��Ef5J4��b`E��,cIW�����Nz�MdMlC]
�r�78��~:���$;�����z����N����k���%���E+���ǖ�E�u�Q�\�`#�/Cf��S���tN3&_�Wm����f���aO�L�#��|�d=%������~D�o�%�E.ף�%����q�]P�������<H!H _7���уWa|������n/u��Р�Wr���Z{�
��Mv�0���l5��O�E
�j���i�K]n�{Bv/�8���+���Y�
�7��D>tr�����M��Lg����¶m��<J��B���!�����v\��lh��G�G%��lT\��f��5� �\���z�
��Ȥ(�E<k���Zt���7�m��8���9q�YWB3Y�;2��ɘH��V�7	�o��]#��'�����X./�x���74�%f�ԃqt��������0k ���|��D�ʧ���$P�{��x��5�V�|�{A�oa%�4n�P��r��X������:�ڸR��	Qh�����Fc����ܒ���'Rπ�9M����ڶ���,�KVS�)]�&5��})��8�[6t���� O�L'�P�X-ZӔ�Q�庲{O��6m]��*}�<=��5������߉�#�6�,��o���յ�k���h@e.��1ޠ�Cܣ��ŋ�0�ت5�s�C/6�>[l��T����jg"v���;
>�GM*���rs�v��������\���$��M���NhY�W�����?��Y��r�����^�'�d�1{܎mj�#R\�Iy0����]�s�����H������)����d��4y��	m��~�n]��7��B��V�2�~nW<)��ق_��h�߿�s����]��2a*���!�:{J蹉��,~��bv���2K����%�L�d���on�r���OE���+�伪p�aQ�z+�	O~�C�������"�CC��WT(�;�D�+J�L�~���4���D���qjNY�����#�k64�a|����i0H ςBB�z��*�G/Hd�Ur4/a��Ncai��S�,��.�������0�l�j�q����Vr/����w@3�tˣ�@��n<BYת����
�Fvߩ�ؤ���	%Ǝ�5y��̰���I��f-�:C�{J�ء�i=qU���1�#,��,��$��4!�� �(�XV�N�[;�#�iN6��:�ݫN�|v���$H7�t�*b�3�M,�\S�uQ%&� ������T2.������ɒ��'&���M�@*9�s^⹫�hU�fB��Ku��5X���g��d!t�s��,>=��
�읳ʩ��8`��N˝y��>hsz�=t3Nl�_?t��a���$9%�_���|Mx�l�~��-�W_�1��T����}F4g&q7�B^~�5��ऐ��K\����]�,[��M���O��	3P���o�ַ��%Vl�����W���u7�����)QF;̆ZQ�C:"�@�7����ꜛz��FI�����SSVo`�KбpA�z��~b2G+�F��S���,~�����q^����IFy�A%�Lp��3lꗍ����}�;�	�L�W+
UeV��|�6����(��ߗ���{���],��������7.Z��Ј4u�������<0���Y�����D�M�`D���9�젇Y!����j|�U�6���Y�`d����^ڬ�I����s_;\tW��^�J.�N�uH�/wd":c
��f����-�·C
�B��	8��l�e5����[KWm�8�^�$�;��O�b�T���}&��-�P��Ӥ���� �����~�b@�b�CkZH�$������(�X�cX{O��,Y�r��GaL ���J£(Bz}������B�6N##�1%�9�,��Ǿ�~e���h�D�u�D��]:�`U�hƂh�B���S�~�h꣗�N6����<���ڬ������Hⓑ)?���Gd��VBN��%=y_.5J�a=�R�Q�7q���Y�9irB7%�,b�RGВ	��֙���Y\s���#ϥ��G6�`JNzg/Y�������T���f��z_H\���u�����7+9�{;w&sY�e��b�l%ə�BH|�F�S��,h�a1�=�D����f!l�W����v�h�[u�7g���2�D,�/��@= �(2��ʂ�ΗL�������h��W�$SM�í�?%�X�%1�%�lh��V�GLOr̡�]������b��db�}4�����_)8�j��na�I�ߗ�y�*��%aN���ު�tPZ�ͫ��(_���a5�4:"sE�P�۠�U��Z	UX6���m����>�$E�$U
�4��'
�(��G�ht����NZ�����LTԖ@�,1� s��p��w�Gw��)��W;���5�]p�Mkq��k�z9�)�֠�v%���r?� ��e�r��S����d<�7ȗ�l7뎥���j"i�Q�X����8=���F~=�ft=v���:�΁��]��Px� d*v ;�l���6�����y��� ���D�-�����-1_!lì�`��b��UZ����[5ORK٘�Tf�CE����-�	���C}���ɞ�!j���)��84��w��v/���h�/�O?�� �u�'�<�	K�����~nJ/Jm�� ���?|�����q6�7p7d�ȯhT�5���r<ً�9�iZa�j�o:�p�/���S�΄˖y�3���
�e��2)GT�/�,�T��V�ま�|LtY�/A�{�ޖA���|�N4?/��2
��2�u�@,#`��(�� �����崺7���13{ʝ�p� ������q�c�mʖ�W��1���U���\��<��t�3�B�9Z7�O��ёӯ$Su�W����`ܮ�uL)�1W��4���J������/Qg����=�C�Vߥ1��z+��޽�+O��ec���������������L��Qj �MɹM4�7�:��5�8.��[�?sĻ�X�y�iZ�j�$� 4o�Q~�L#i�0�r����Ԡ4C�t��'���Nn���󟃷�.(�i��	X��<�9FP���q���!�SWqpa�����f����_tߌ����K��a�
�
g�
GY,a8�T,𳐖)��a��i�ml�>����Czw��6��ٜJ>�g������~������3�����d^;���&���N7��j��׍\�Ʃ(��Q�*�ɼbF7H�ii���t�6��z�j�6v��ΉJǠ��D����'��*G`�|����8(��:�|䰺�����AB[h�#�k���U}��1a�r�b��N�&^@��X��ry�Q#�=I6~�cۯ�c��}P��p�g'��?�-{�x�Ѩ�^���р�Fc�J��j3ѝ���}
�`��oG���qNZ��a.����ۭ}f�8H����xR�1{x	��`���Ls���DnU��9"��QQ�$-�jG81��N�	�)ilƸ��&�h7�Ø}Jl'�bN��3ޢ+U����ɩ�I��_�x��{�մm�Bw�_���v��s��a�M� �W���}��qr2�#4����w�oSWq��Q�͠��NyBE���".�x�aw�D�
r�%Bi�p=b�>q}h�i���$H�v��ŭ<fo�����Ό]�ri�,B��Z���������C{�����F^ ����������~"�]ڊ��9�x.�-ԼE�x�ٵ�~~��>�Ȕ��m%�O�z�&Q��3�qL�Vhs����k���,;�G�����H�i�O��I��-��N��W?iȳ����:龪ڎmQ�e�����@��*-��Fi���}vt���h�,鑧6ny�$���Κ�]���y�-�/���[��\�BC�Ju ��y��uͫS���g\�y/��1�aH�@���@�ڎ�ߊ�	��SؗV*��V�S���6	���t&�Vóu)
I�r�K�᭺$�!?�n8b�9ێ�
�2fQ���2��(�n��g�
�|h|������]������"=����B��f�W	-�(ȁɦ�R���#_�3NH���U.=��&P�4ڟ/0Pf0���A�EM8� mP!��� �L.��S�v��K��g�B����Ba��>-�\�.?2B��
����wizM:B@h|����nb �=Cخ0�����u]~E��JT�W�z-ؖ�j�71��*5�֐3l�Ƀ�z5�PB|<������� ��4%ƚٖ'�{J50�l	�~��B�8i����3��NF��8�#���^���T�S�u�]��>�� =���
���}�#қ���%��LG	�b�f��oN��\�	�RƜH�E�%�cf�<Y�9�zГ�"���ήg�E��ơ�������u[w��mB}��䈺UU/E�^��{��I���2a�
����������b8�b��D~�<o��8劽(���V�"%�5o�-��G�*�X�9��W�j�Y�a{f�zw�t�z}� ��	g�e�p��cd���i��6T%{be��/����o�b�˄�<~�K�I���f�L�D�y�	),�ّ��x��2D.U�%���8��y����g���6�ݚb�j�m?>��7SU: ���ڄ�{a�7�[�'�IRR�S�kϔ������x�躒���V8a��?��~���E$ڟ$y0�⻈9/��vhǛ��Ə<A�K	���W�d[��X#�qC��F+�`E}��x��5�r�e~��s» i�׳$�D�D��m�~�}�P�S�m��Q��[���Eŕ>[��	c*���$!�8��X�����2>��A@<a'�2V�U�m�Ar�����H�Z3�?��79�TM_���3�����
�����Ĺ*��&IR�s�#����9-��/��$U��f�!(da��&Ϙ��7_�	��2��]d�5O�����9�@Y�_.�(�Q�O��[��·11t��$<C��A�d��+qv��Eǜ����Na�qD����2�v�{y`:�O�^���y���%��Q����*@G"�b�$D������ 9�*�[0���ry�L���!*+���yi�Vz<�A��H�1�m�J�d�:�~_�U)��}x��q���/r],�a��X}R��淏�;�GƷ$���M~���q[��|���xY�M�~y�z���U��+�����1�+���WM� D��C�灤B[:���#3u&/o��K�`GW�R>̆+I3� ��C����l&��CW�ۗ;�*中�����&H�����z�ҳ�Q%���X}s`5i������W�ɿ� �i{6֓���>��"���r쀺�ћ��2�ݷ,�[��ð��[�� ���F����F����iY�����>�=DX�JHz�ؓ�pm�;��������:g�N�&A���_M�-԰>?�v-p8d�����p��@�I� z���"O��W�� 5N҈[��e� g����b@��PccW�������fGb���=nX<_�@�I��yfv�2CD"���[�՞3D tv\{��� ^*�V�q��:0�f��ʃ�E-T�l��D�p�@�tUI9)M������tu���eX�n�DA" �+�z��z`ӨI���'�5���>,\����@�$?�%�����1`l���y�W�?��sR���L�Xq�)�쮓缾(5�pع�LOs7�\_>���}����sS��t��{�k�d 
���e9"Z�������N�ѧu���w�;�+=����8��
�h~��e�R�Ɔ��$Ў<���]�i��'#��1wC�^���d���;hy����i_8�yt�e����E���C����X�Y�����P܃1�wә9��_���R���"��#N�,ɚ���َ
A<5ކi�L\](�u�$� �:�!���y#@�,��$!�f��;���F���:[�����3�d�G�F�ܵ�/�FA��%�.���D=�{As̡V�W_c��18/b��f?*xu�����B���Y��ݐ����o,��~�{+����p�l�zWZ¾&�}��{S� �I�|N�����-�b��)\��W祝�q�9�F3f���'//�A�|�8�� ��%:��{R����_�|H�pN�fG��
��,��B�nH��Z+W�g�d4I^�?)�u4���A��UA�Z|��N(���xr�ZP�<	u�J�V�<K\�;qa�JFI�u_U���ρ2��<�ϼ?Q48+3$To���^T?�	L�4z�m˩�]��=8�|�U�Z`�3���.ό
�I�����z>��|��O�)����X~��RδĴm-��i+�"�K��Ձ�<M"�d�b��Ar�/!�n4H҃3��#7n�·���Ѕk�0�UG\r���Z���3X/�fr�ދ:fY�BK#����뾶�GV=��n�cm�*x�H�� �*�2�2e=���v���얒Hl�ħ� �AhS�ʬ��9�}��>�Jv~�^��=H�����L򭟵H�dO��?Z���P"Ģ��b�l��A">1�16��ԍ9C��p�0�GƘە��w������J���`�X����R/3C?q���:�ƌNfEI���(5n�hf@��x�Z��v��j^�������H��	Q������x�]����$J���DPr&#4)�^F�n�4��%pn�{^#i�4����	F��)�&�w�]$wR�8wv\(F�F��.i�0BW
0�h��0�he�!�u�6o�����4Ad��cNH����r}@��a���+P@�l.��=,� ���Gv�;��c�֣�mA��C�|n���*�o�X]��-����KI�3�-�<��������	?Z.�C~�r�����E>_J���#��Ҡ��B�+�U6���U\�v2l�o9�g��,���D����<�+�Ϡ��܃sH��Y1)�٧qĜJ��|�`���׷\@V�����!|��I�Q���E�t�*����Ǧ�kd�s�=��B>�[� �A4��=c�$�M����<�	6y�/8�$7I��S�'��#<C�h�sD� eޒ��F@!��̵�W�-o�_���.T�SG��}%B?�L/+OB��#q��ava�Y�OI�c����)�)�pƐ����au㕻����k�{3C=� 6���1]~c�V_-9Ƌ �6M�*�B���vz>�'*nY���`���80;�=��琮I�"�o�휧Ww��A��]521��WƎwt�MQ/=���ݞCrB��H�=���8[���T�X+���UH��d�,?�؜̣^3���8s�
|p���!J�����BM$�;&N �ܷ�A�Py$~^0_�����cm���Jv`���C�:\\<pf���Z;g�����'�f_�B+�L)&�Bs!��O� l	*�7f�<ǃ�,�"����+
��r�J��[����n��.��@\�n��|+��]T��$�����[�/N\z���EC1����A��M�#`�h�ў[�8i����Ǖ��V��Θ�'�!hBc���=(��q��N����!v�M˴L�����^.5aF��u����C�_+�����݀UH��>��-H�H}��葛�*M}��s��㜼o�`x��b~�:����W�c�2\��|�d)�2�㜶�xS�$-nمxm�Ql���J��=���N���}@�#?��_�:��'���CLf�W}y�[�<��*A]�� a��Pߍ��\�U���������.f�ƫ�E��>{�N,q��⹱V����h׫�X�֭ ���g7T��QZ��N��̈J��y���zo�E�IZ�mn�z��^t�ٴ#�ȥp�eU��{� �ľP2ڗߌ����d#��q��j>lw�Orڨ>Ō�*�d����at>�ͥ�~C���v����*�>��Z��ː�j�6	u�L�āޙτ���"�P��"�'Q��jl�0����r\����Ma��~�rKj�$�$k0��މI$����T��׻3 ??�c�d>��MWkQ`\�k���0��l)B�-�j�7�{k������r @����b�WD2�r��{^'!yS�.����{�H��{#�K�<�}��9��Ph� ��[�2Ԃ\�����Ѧ��/�U�Ν��&���гCQw	�B[�x#쑡�q�$z���L�p�a�A"�61���#d�8>�H�%�8rYpn��u�I*�įX�J:�Ӌc`�~���qbã9���>�ފ���֓��ٶ�� �Sj&,�@���� $ �Һ�Sg�|�U�xt�d	6�^U�w,ʸ�u��l�	扈�،�o���~�C�F�'�4[>k��Pg{�:$�'G�#�����뷊���ǡ���M�����9ǥ�?2v�����x	gX�o����CGWl�#������$CU6�tp��K�� ���հ�f�EU�%��!�0�c��LU��#����!R�QK�/�C7�>Q�sn>���R
��#ҳ<��������T�ϿhL��|q�b�%��BT��m��N?��j�L��C�����.�t)��bq�/�}���A���6!޵�޴��c���BR:ڻ�:6{.M�ϸ�5o�=ؑ�o�iO��p��Z�vV�&<݃r��d!��ǫ�\�؇�)rn�D��К޼��x��3��7῍�S\���-as�Ĭ�!�[������=��K��;�����2�e����HF�ϼn�-xCko���y� ��|>�| tp�T;.|�^�&�^��4�[G��J�����Elm_>57��uCV����u!���)��+r$�,4ی-��9����֎�rh�Y�6\=��0F޾^Q�m�1D� s[A�
�]�� �_k��]{�����9D]l�Z���.���A9�%��)���#���A����ђW~(�莾�1��,��%���#�H�qQ�{oq��tʘ �aLW
.}3����0��"p0	J�d�%����E�ԑ��,E�U��
k��A�GX5\�����8��U������%�҉��*t�sWv�-�l]�u�W�$�x��m� �o9�2E	G#��xf)����$�j@f�Hb������7���ƒo����y�����)Sw�5Wv�+��p<����叁�s<�7|����� ��i>�#O���rly ��0#<p�,vE$}�~��Z�����ˉ6�X���xP�U:�&S:*ժ���v7��^A�y�or.&H	E����)H	�$' �⮁=0����46�E�eT�f#�g|#Я��*r�ĮOaf�b]HI�r��k������c�=���,𚱼F�A8~�cTq��թ�݀8����"�U�˘Wor�@�LPĕG��Ǡ�R���PG�r�a�;nJ�X��Z�0���{���!�s��e"Qw��ʬD�
��e�!��-�W��lT���61��sW�Z��y ����?`Њ�Q v` t̺��]<��&ڀ �B���c��°F�t��[@��D�I�-S!���U`}ˊE�G� �h������E_.�`���)79�B}R�8r>=��撶�<���Ύ��WR�t��+awcõ�c.e(��qz���rZ_�5Y�&��p.�[7!m�����e�ꍙ���pY΋�+�`ZI��C�%�_�bG6��&�d`J�8bi��>
8\�fz떡e��EI}p��KH�BTElq0'����_0ʛ�ʉ�
j�-,I,�Z�\�s扦=d9��[߬?+����%,�#O&iI!����]���bj�.��~IY�{��HM2=��xtN�j�h���,�ӟW�;�]\�z�vq7��z���L">���C����'��uK�3�&�Z����4?��g��ox��W�<�d# r��'�<74=r}($= a9���ozb|G1��O���kץ˴bG����GSZ�ju��6������9�a��a�+�Jx����@�1���ZX+7�^L�SC����+Ƌ�˵%i��z�������.��ʡH⺘�iO��A0��lv�����n��@]��s��[�#��L&��0��h*�t�	f�� �Y0Z��!�� �&� �$�0��h���Ke��Z�i���gU��0����ق\F�T�p6I7�/���u�dDT����{}��I�T[�*������O$�#:Cn�?����;����N�I���V��0�t�ԙ�7�i�t�++c� ��rL;�&\�����? �WeԲ�� @���*�l!�|�h�M��4�L��m��i�9�ߓO^m����� ��w��T�^����%���L����E�T,���-1��$K@���VXJ���QW��;/55(wI`�ys�'����5���]K�
���y-��*cX
2xx,kM��b�ڦ���sA��S@%M@�!z4�.���1�b�ᲣU^{	�/l��!46�]�]���7��B�U���-:7�l��I/lyRe�l��o�^M0�s�V�<� Rě�.�v�b�M�!�&/���x�n?���o=�(�o�VSO!Ku�ފ�c���þ�/����*#j�'j�:c#nZ���>|�æ:L����j��B�>�����;�͝'��QH�R�|g+�gB��ґ'0����=w�*y6�g���_�����PĮ`d��UT� �3������ݞL�������p�ԭ��Z�����*�y��3�eT�_��(����X0ݘ�jM�lo�'�.a��8��v�)�B��̈�°��a���ܺ�{����f� �j��v���)�zi l��@�lvO6���T[D�-��$���O�ׄ�e��	?�S؇�6ٷw)0� |���#΋�u���y�D�'�Z�Ն������f�NgC�� �Ym=�58͎��Wĭ��h~�!�s(�4w�[�tJ������3C�$N�_��)��2Z` ��O�cG�Q�Q{!Ӓ�)�����4��ٽޚ����O��x�Ofd�+��@�}��X77��%���b\#E��3���c�0 �?z������K>7���t�-؀�]9*<�&XlQ)�5	�΋V]�����%�(�X�֮�=��Y�V�P{�ʋ1�Z�����B��]mW���'���:�>��J>HAB>�R�
��t]��Ў4g���h�� 7n���8�H0�p��?��\Y����!��0~�!�Y�m�I���Y�G��H�Fd�Yr��@
����]��-��ƪ�ݑ��bCj�6R��(���vs���	�ZuA��#�D^�J�Ⱥ4 �b���ā*�Q3P���$Պɳc`/�A���b3X5n�)�x�腉f�6�ě]�t����R���L=Kڄ�!%`U"'�n��X�3����?�N�h�u�#�4���ė7����MDNLKL]�9��+H�pUj�Y��>i�C����!A �>�K�<�༏�h�Hx6 呌�ω5�4������M\��Č&�A����,!Jwu�f�%˅�`Jn��g�~N��q8��pwL5�J�U�5UF�q����O1�ZC1�=hp����Q�1[�D7��H��S�Q���?�
�Y������u�|�PH>M�pzy^��aC���:�d�r*S���a��L47
�k��8�I���x�D�x4$��2Ba�MK���E�!M��3�4�߸瘣%�~�/�,�77� 0>F�D�ҫwm#���V�!�
MܪbS�;��;�Jۍ�\��x�4�7hD� �Z�p�T�\��Pʿ���R���^�=�.��B�PG��C19�\'��SVp
��=�7�%�2%"݊��3*�,���RӠd�k��D<r�RU�=���'j�h�!W�YD��1_�v�������U�^�aU	'�R�J�Mt�Kf\����ç�<�z&'%7G7���U�:`��97X��&T+b{V��2���*��Y��i��a4�N���5��������h�
���&$<�sϭ����5��f�����HO��|���[��$fu������랺�-5��5������R$�0�����E���e��[�ѭ�z�R���h$�\���ٱ�L�(��֍u��&�v���GP����vH3*����ee���0Hgڡ�� Q�tKԢY$D{��sk�o@_���V��7(�Ha��+��;�D�>�H�^�,�[�Q�IZ�֬��ʡ�B�XXh�%2�WM]�f�s1S=�S��@��{����1��F��j	� �aO��f	)�?o5f�'h�D�Z�ŉ͈<iJF ��xc��SrB>�!���.�%?�ť�":�j�����d����sSp'�G��9���*�	_}����j��W�\�m<a��;^�C2��؞�l����
�x��~�R4��خ�$ o4���.9��'���O�˾�#26X3�50�q�� ���AZ������t�)�-�\Suʿ���� �'QP�0Ʒ��"�x�ͼ�Gi�&�Oȯ�^aދ��is�n�&X�M�.���ڌDrY%���X�FiB������]Mv5K[�v^����1���x4�-�o Q$�~��Q;x��3ʧ�S�S�=����~�ˋݶ(���{���&}�l�K��Y��)<�%���T�b��#�.Y�����̻�F���y�3�,��:��cUN�@aBL�i×U&Q?he��	����(�Q��M�bY����o�Lt���Wb9���Wi��i��BHy��k!�n5Z���a�,)��������X*�7��k`�|���#�
da2Plτ�j �O��.��\2�8fe}��t�D�'�*�� 3��q#���#Ԃ�w�'_d�!�t�8��U���s|��2�d_�v��j�nO�X�t�����l{������lԈ)Z�B�Y�7��1Jq�.�á����5<�2�������o9��I�u(�k�*�+���M�P���m>������
Q�1��O�p>O��]�˚�3}#třv\\ބ\�e�ߕ,C���9�4rR��	�7���3���$�������G-?��;y�k�|��o�[3��؛�f�l&��`ΰm�yf6ۄ�y�*����k�Ғ&gH���s'tɁne����[�@��U��Tud�nX�݁�n��! LyG��b�S�Dr��騫f�?�7�i��{�k�F�=(��E�ks�Y��n�>�Rs��L	��`�J�`C�'��T8��t���9!c=��m� �����+/�:�aHi����6�1���o�8{_Ydg�x �g�?B����6.�6'��IGb3N�%Q0gā�? 1��k��aO.�e�2�:n�g���4��ƂZ�ψÞ��0cv�� r.���U�4� !�.Af+}I�-���Y�=�GM��f�&i�N4@ܞ�M$��$�����j־9�LiǱ����Y[��Ͷ�$�)������^oM��[��uϟ.�?�5���BZv�u|���T:�:c�g�;�R��K��2������Q��1��1����m�kY�Ѻm��^�����%�Z����:-d�u���?�  iY�k�n.Z��^bavkۮ���iw���m�S���Jf�Ũ|B��j4�2��+_�#]��1�]�dIk+��=��|��=)u�"�i������F�ȭ��c"�B�ųʅ����qr%H�V�t�S�g�"mД:w��0c�sz8��#$�C�i׌d\i�R�Ir�3���3�L�n7�q巿�/>g����;<�o��aQ3\�,����Վ�
��YKû�g0��!��*�����	g��\Q�����!Ƅ��j�'+Wb�c^�"�����)	���Zͦa�m�(3 `���#j�Ɯ0`�:��.x
8��oiQ��u�T�!<�9�H���ن>�#$��F�3��'��+��X����߫tم�k.�i9��h�^�8G����>�����q�m�r1�?^�92��TWy�jDF��~�Ezh���%{�z8�,��qŒ �_�Q�u(؟�NS��]�ZXzG'���Ԯ��W=���t��Z��?�8� �:Q����J5p�9k@��v�Y/v#�����Y��0 �`A��U�(���T����M��.��Y��ŋ��#�p���ӂs2�դ�����?�nE��%��
�u�	+_{�ɴ�����P�8v�lЖ�fB��������e�:�4�~�ؘ�����8�d�"�&FwIs��*�`��E��s�q\y��w�fx+�㘱��P�L�Ws������1����_���}�(��q����e��;�`��i|�����p�Aw�ɿ�ԙ_m���Y��KS`3�4�����9�Z�֐��+X�(x�^g1-pg�(.y%�8Zb�#���qg�uRQ��%��7MO���;_����|�;�$�B�
�pOYT�,]�^��S�8�`lp�{�����d"��D���QB,m4��u^y�Y"��Pc�=	nL6�T+�/��V�y:�Ƿ�v��o���1:oI���1w�廒���8>;XT�#�Xu0����$�	���}j-���0�u���bV�ݸ����VOl�s�a����ex����J�S#!+�fS�rIt���� ��*�i�����5���z���磜�� ��IP8�4����<?X�=C�^���i��#V򺍢Z�V��l�b(�9YH"�1�㡜'���I���A���SM򿐇4�Q=�<(�q�Ѻᐚ%�^v ��O�k�|��t엿�$k�2�,��x;X�UK�b#����8�Z'K��u%.�����*c}�Cu����,��GX��M֋��-�}V(3'sh�_��b��AH�� p@��1eќ�,	\��a�0w��"d���	����?�.��K�O9_��+`2Z���aT�u����b���}g��Sp�N�N�~"���qq�m] �ˏtGP+��Ã��"u��_&j�.��,����<yԶ��U���6��-[<���C��R��8Y~3͖g�ri�X�O��cd�s,*ịBW���aĉ�˞���ǒҳ�ʯ'����|k‱�g�4���X���a��'<N�͢�>�Qa�8�x�����C$:�c5ZןŃ���~2Q��d�TG�Q���������t��a�Mڢ������ZB��ǚ3� %�>=���km�-
3��q�ļ�#�LF�D�c�&r���Q��LB�����x�u�L%ߋq9G���4�p�2�%��UfW�Uy���aWS����QQ��k:�[Q4[\| {�oBa��G�d�5�v�y�A����tA0�m>~�2
�BUR�a��aO�(�w_�
��q��q�th���|�KD
����L�����3��������lB~�L��^BS9��_E6��5r�u|�o�������}�ٰ�;:��W� �a�iL�ڝ�L�q�i�p����D��<���}�(��L��o8��@O�2��I�k|��n�w��f(@N(�g���E%�L9&�a��.���QƢL���Џ�7���g�{�DI���җ��Dmq?T���k�G��MTąh�L����K2?P9�@��>�V�k�0�6F��k���*q'_�E$P�����u �S[�k[�����ج�_[�� 8 gV�;�A��>�_�@4nd�(+s(D��4�?m��t���<Pg@���������*^�y�uz�&Rj�#v��$�̄<���E���(E꙼�A> wŨׄ�P�]��<gY��*�؉>]pͭ��_�%0S��I6e���]`Z�G�o��O_��9�XG�Ē�7|哋�9}��C_��[��\���m��|D����Ab��6�L'&�G�����ſDN|��Q+��ɫ����LtqT�R�������!ިMu�dH���2��^'�I�24Y)����t��7B�����*azHƄ��^��!S�� \��LF΋Ԃ��_K���9��wpƤƺѸ����sڱ�c�0���`�U*>p�Uw�c�OڗF�Y�����h4��}�^�V�����/���*�E�A,4��|LC�Jjon����J̘�_%b�u!�X���~�^P3��#2�.�����@�y�o�����h�1�ni*���k�/�?���ɑ&D��j�YK &\[�u|n��1���ʸ��be��J%�f��,%.�O��:8)h�&ͽ��:z�ٝ��j�c�rv�2���z�`��gE�n���/�!���0H�ۚʥQ�9*�˲�`Q�[p0��8��#�9@H4"����.�j}��5��,і?W�����Z*u&z�&�9S��sjW�R�)gmI�S'�v��sn��}��~-�~� :����K?ʋ��Pܜ�:���x�o[{#�H=2��莧�$�Q˵S��N�@���\eh���J�<A�#4B1�ntH/���&�4��"���Em�Y(5d�S`"|_G�������F�d[3�{ji�� �Y�0'������:I(�B�A�"	�	��\<�t��#����^�	ؖ[��{q�3q��چ2�z��(�̽�gG��@Y)�v���L�h��厹_�ts#�71�Y����kYg��h!K�+�Ao��
�6���HV8�& z�Jˌ��y�d�!�0 �K$���t^iQ@K���6�)�.��%ES������}��#S�R*�s�ѧjn[p��Q.Ն�j���YgZ�x�7�h��n�{�J�ߎ�?� ����9�ׇ�
���2�~�)��=�䭨���D�8��3��CG��]{��#���lqc֟��S��ԍ��Ye)���R�i"����qQ�ׄ^A,{�[6�șfUh������<��[�CBy�,=���=#�FbKc4�/�*�� ��5������K��e�FL�G���T/�g@��?��WYE��v��V����H��t����^ڰ�
ct���#��GŅ�NC�F�<kF!�s����'����&�`��2�t�q�	HZ�}R�j��}��V����N���m���8#jP��Si�i;�s���K�_�b6$��PGW@��ӎ��Zh�}́c�1d�^�n�	j<���f�W҇�T#F��E����M�\�����r�s��p9�5��E_���,M]1(�V�:����45��.�x�F�$=/�o��jZۜZ+��!F[<GE���>�EۑsO�j��c����aS&F@�����u��w��s]�4���:�q�� Ss��N�oB��{�g��F�g���Hｧ�x�<�j���c�A��pA�н�Y�n��U�H�5�XZ��^Fe0Vo���N_�G���C�ڋ#�	�Wf�C�c�Ɇ1�q[I�]��HW+ g�+i�������j���Z`��4�����H�fC�>���$'����,8��J� vb��e2a�-b�>Y����4x�Á3 7C�se����{�@�**Do?�Fߞ�1�c�P?���{N�y�ş�h+'���5�5S��`���]�%1}\�z�����uT�zz�)�)n ����Ǥ
���3�P!�~�Fm��E:����� �0i�&��߬1�s�����K�?���"@�lK��3G��da�8����;a��a7�;���o�R2����/J�ٞý"I����֮�'a5}� ��p^�?���=�V��#��g��vȓ���&'zୄ�6!=A]+P�Rt�)�Ys��½3��čx��ٿ}�K��R�A�o
|o��.�d����R񷼂3*�z��}���(���E�:������- �m��4x7�@(����)���)�\���X*���}�*yCE�|M������~�y�r~*;�͠�������'��Q�|	TK���'����H`�39�9���I^IW�����7��r�藧��F$1��6j�y���1���^����6�f��<��<.݊��CV���\js�u��ő��(rD������ܷW�_��h��F1�&�a)�=�Iʣ�<H��'�L��g��4�E,*t��h��H�x�����Vc;�
 sg/��,��m�ثL�sV��	Z�0����ܞ[FP����Y�V��×Jl�+b����eسӭ���U�@�t�7]�#�ĵ�Mj��ªEZ�����-޶E��I3�����F_̟�_d�w4A��)V󔹛�=u�b��h&I+*��g;�Tw\H'�W�5�5�m�+�Z<�>M0�gm�@6,�nZ����/a�As���x��t��[f�jH��R���5̊h�9jp�j=u�s����'���9����9sȻ��lZ��vWư�}|X������A٠rƈ;w�)#��qd�ˇ���2sѮ!r���Uvw�P#c���!>��8�\"��nrJ�ƅK�+5�q�
�Ж�>�d.2嘅�i��/�-�d�B��C"#�X9��*��ʄ���+v&!�K�݂��(��+��q�d"��{���b#��+�:��װjN*�ᬃR'����!�V�n�E���]��.Ӽ�`F�<�NSFd4�uA9���{�Ņ%K���;�j(tgWFō��z��� }���f�K���A!X�DoR�'��*}+n:��:"I�:,{�9N�����('4Ӵ�����.2��+
���Th�=�| ���u��/I�4Sc+G-,��P�.�S�	�`}��1�M!�:��&����<�@|A̡���䯭BM�f-B`�y>G$�*�� ��!q���Z#�FКC���U��y�+.G�|B��{D�c�A�}�[�/�G�3�Au,��m"i|Q.��,Y|&��K��\�N��B>�$�T�����4�ahN��jbX�S�f��@�JNO_J���sR��2w;��ji�wR���J�.�̇����b
�˓+��_����ϗ�ұ���	N�a�	V2$�$��6��I���,�ٗX�{5D�Co�-�k{l��G�P��n�:���p�8��$DF�5-Xoua��{�$!POnQWCF���`��I&-��G+�O{ED�3m��ƽ_~k���X��Dtv��ƛҮ�vdR_n�9��);��W t������s#^��%���l&���"w�\(���ܞ��i>�5ƫ���Bϊiq�S>���'��PI��IG'@ߡ���⪱����cc&����2�1�hI�t��ʦ�M5'P��.�}=�2��|��'��M%�׽7�P�ψ�<��C-L��K��i�(E��xbL���?�č\#���Js�(l�1��Ϲ��3��G4ưCt}HH�>��s%�������!O|�_�2-}�!"�2�)�	X�ؒ�:��n��}�����e,�.b��D��0'nq�!muW[����R *w�7�h�ݝ�zZ@7 (j�Āړ���!T���(c�[f�7k�[�7�90��F�	7����@��$�6�;��W��ҵCI��G>��5KS0>��0Epw�����|Z�̋N91��O:�T�8��N�>�h�w�&��ͦr�"�j�~�yj��������(����m�LGo
Ha���)�ˬ[��*nw<��Bļ�S�n������!�3܍[����j���Za�B7��8F�E�e��1��v�S��}��6dM�a�v��m�B̖���d�1�{T��þ�%���"�U;@��'���).Sh�����3x �����9��}bQ��S�d�u�C���y����-�i����MڋWR�nV��W?è��@�o�:�z$Ж��/!�!y�^ ��BV�Y�4M�Y��*��;5�D�������3�����A*RV��3��(0��xql&�:�������/.[Z��4�+��#�|��5fזp$�]��/�n�Pa�\�ek�{hk=��� ��Z��_(�4�}���U�����.*�yA�4�ɺ�iJ'�:��o9�|�+�[��ի��1(�\�䷌=5�|92�K�h��z^���X�B��J􃄽��g�{i4�5��;a����M��9T�ӘgM0�,����]�����/ޠ�z�UX��q������{�t�^�3�`4U%E�U)F_���W�?� ����'��*=���T���7�x<��6I��xe�?�x��+��;�ʤr�{1�s^�ڝ!|���,In�N^���B 8��4�V�RE`�p{��C��v���k$I�ԧR~=��fYȻJ�y��0�~Ycؿ�����]Q̓b��B,Zh3r�b�ϙ<��0�a��fJ0hE� 6��mh:�^��_0}�Qe�f$����-��|������W��!O�ߡU��jJ��{�iz?����"�؁ ����{ڝ�3vFn�\�j)����0��;� �< Y��u��Ӊ1��%�M;E[�˙jH�\9��[�R'v�g�d���	�R���1�?��ud�����Bt�]Ӣ/C����$&�LD]�@/G� Z0c�vXuec����\�h�"ښ�-���V~ܟ�򪞲7[�I��_^wV��GJ{�o�RNn��e`Ϩ"��P���+�E��7��?մfo��fk�RW�p>�3��׾�臹,�_�)�U�(F)b�b����x`�16��b͹�W�g4�*�8��=&wk�����x�A��w�����[oK���K	���L�fV���W�z��#��n�pD� �M
̟mm��^ 9-�l� ���޴ĞܓG�����B��Y������"I��T�q�gE��N�R����H+�*岔��K�� �ly��o��P�Oo��������O��.�{w��~=��ǚ�#Y�6����7���E�c%̂�Lu���� ��4�R�R��	zI�q�,ْ���j�^�Q<���Q:Q�V�Sma��6�գW����	(Zؕ�\�oN.��;�*��?�ͣ��j�
�� O8��o�4K����đ� ͩ�Pz��AK!�a��'�������g�,�W�@�bﾳB8OH�>�C*-�wX��1�r��U*�S����8�ǖ:�<�?oko�Y��K��C����ո �%�ʀ��J��k���]3��HY`�"����e����/�R�ha����[ڄ���-��[�5�^s�b��a���zJh�|�{B�Z�Iε_'��U�HRs�0�#���@6Kׯ����'�aE2o���=X��X�eY�o�Kd%=}F�N�h��߷<a���)�S��	�Q2=�{�?�*!䕡���!�bѰ9\q/mP<U3'7�0�@�E\[�a����˔�c�6 ����"�%A�,�p��r�c)�����-3�;,G�[�P�63�Φ�0�ف7�?�e- h�����\~�q�{p��-�c~��*1�rh�,������ �rG�;��!���8��W�<a�i��}�=�P����'tÃ�8�`�g��2.͘&��/���qG�o1-C��N��s�(�6Ti��?�=�s�0�n����I5��]��X�����Հu��!d�(尅vø$O�;B�x��,q�C5�`��o�2��8"��k#�7&��59}��M�a��S��l�:H���˦F�ʔ�j>�1�'�eYPs5_t<��n�/�:	9ͱ���$;��m-����K\�9=�1Oq�p3��ջ�3�؊c�G*��*@���;'>�~����w��q�$١��X9��-���'�wC�RS��)^2�_�9�jt+����Iw8�dyN���
/]�9F�����j�Ï�#gUoxdNd�m�=2�׋��#�DQuW�9��@�%�YIӡq%w8iң�m-3�v z��_�Xrd��E��1�������,N��.͕�n���\`u�J�\+���hN9��,�S,��2Ns~�uE�'0M���k�f	����'�j����?T�x��N�k��Xz���U��YM״ů�#�:6��s�YG��6t"�������з9�(&�R#��`K�.^Ɗ�������=-՟�Z�Ȫ`�m�1Nk/]�7^���g#� O,d�f����w�B9?��}�f_�T�Cx��[�q$9+��T����j\�,L��˞�S��A8��.���!��s��F	�����mE���N` ����4Xp�$0_���Gba݁;�ոQ3�m��E|A���7����˅B���țm�u����wa�cl6�q���Ҩ۞9�z|�ѽ��1��
_�n�r�9��ik7�r����hڑO�C?֭��^��6��<��� A�i�����W���G_JW3�[թ�LdxS'���
Ε��$��3*�U�t:I�s%�ۇƫ�5�X�7^��HN.	������ONA��қ��Ƶ�9E��ơ��y�8#���l�}����V���\�R�a�+hq�GgO9p��ozH	��� GT�|�W���'��$�ny��藱2��3�,EC��\g�!z���qc�����8�������L$�'�+���z�
kt���9���w����k֐���փ��2�tg�A�-�r28�>���)M
����H?B[��Q��Kv���� �B�#�C�Lh�bA4�;hJz�L����S"����]�yd��D�y�Rx���~��U���M{��6ܘ��n���;�΍�����WI�5�����r�i=�tt)����ށ��u9O�5�Y�ʝ�Ef�:�s�Mo8DZe�������b��ב2R����,�A�Hw��Z�"��7�:2��j�6�G�!�[����_� ����[?�^Ɍ5�ԥ�Ts&?�����`�	�$�IL�S[�����2+
敖T���֭-(�����JB���8@n*9�蓾�����s�2����=h���ؠ��m�I����a���i�+�x�@}	W���&6*u�:K��H��;�1�,@X��\-� ��uF�+&�b���hq}�讔�!U�%#��'*z�-�c�6�7
qr[
��Ƈj���y�/��D`�O�d2�?B]�EF����xyh�kc�p�z9�-I+����wᦂ��\b|EƸ`s��3��l�,���"��>	l4���1��^G��l���������ae0�ʥ]ܡ�����+@��I�oI�HB�`�ї�%{�F�ж=I�y����b �K;E��c@A�U
��B�Hr^��G�9Ǳ|�2w�)��U��*O�dn��ҟ�H9~*D~�9ij8D�����	�]e�yy[o����+ړD��Ժn4J5J��
��A���� �1U����I���s�R`a���4��5��
ӌ�K;���G��;+=~{��{`XYA�UKY�1������xc�#�-Y4�G�R�H�����a�$����y�$X(s@��Coy�P�M1~��9�m���4�`�j�+�.$O�)$Z�p>�w$��9�?k���"YC�%�7��d�QJSt��INr
t�����T�@���4�����D���Tdi��걠%��cC�{b��p�l"��b�|:O6��ż��-�:�#��f.�/�$N�Z
�"��m���&�t�=L{�}����u��1ud��5� EݭUH�e�kv�aF"IT��B���D��2J��PﻧS�y{XyM����!���p\~	M�"��c�?���7<����_!���jr<�[i��Q��hO�(�*Uq��2k���m��:н�ߗ�Rp.�#D�<�����H��4VX��w���wr�j��c�~2���y��j��5�)�l(
jo��E��v@m�fD�D#�Yu�lZ�՛�3� �1}}s?��	8.�r`��tzB`�3�+���*l����j�->б�)z��t�S�zǏ��@�ٓ�����K(��Aͥ�fΏ��I3��&��"T�\���%����౹=I<��Lw�]�T�zv]�X�HWڈ�V{�&���#ܳ����y�i0��MTfhb����P�.뭝��߇d�^�v����~`.oEA�o@�Ā���2�Yz�G6z�Sp��Z�P�X���x!.���3��wF+�	%۵��\P� 3Op�
������"N��%�?�e�л�V(�q�[TCA�%�p��j�-n!���T1�+�̣6
�MzP�|{�1}Y����"llK�}&���R�(�&�N{R%���S8�$��X�*�VZ~� B�����-�e����hr�~���}>�8�M�x%/@П���/����&�"M�>Dl��@�o��[!�C����v�'�7��fC����=g�4�w2A�6Z����#����^cj椞��hh��~������N�ŝ�s��׉�fH�8<P�L6@
���D�`��@��;s!�z�b��#$�&�2_�t+�\���/��/:8H����m����,�S%X��J �Ύ�Y�Jd$�Q9�QH0����\a�>쟒1�}J��m�0��B��k$��S�����`�̖/J� �1.ƅC��j5��.����w�:� <���@��B�Kpr�B-Q�6HŎ�!����w/K��닗�0f�U��y�|��&	�H�c�_~@����$մ��w2��2AȄ���Yq�/`�O��f�{�?(��-�u�*@����N5]��R���!�<0�d���W������0�&v�J&=�ú��@�,=^����no�B�X�ʲ�M~����d��q�@��lrh\�l~�I�W�N�=��E��R��2.�X!���0��&�c��[����߫Ek���6�HmP�J~>N�N�B<�����Ȕ�Jv���{����[БM�)���v�`�����7{ㅒ�;h		�B�l���6NX�l�Cf��%�v_ކ��f�Ȍ�h�����$t�'�z��.'�^�Z�)��?� \Q�}1B�J *ow[�60�P��%=��^�8OG٥g�vA�����ы/���P`��p�{y��,AXW}c(Ӑ*�����,
�4m�՗�҄nJ�BƝ`�d�q��h��3�xq�Bi����8;�-�X��V�/����~�a��JA��Ѫt���0h��/B�6��Kؒ f̸��Gq��X_К�$}��;�n?2/��|D��M7OF����uZzTw�#�����b��6(�	��4O�(������I�A�UEKt������=k{Z!�9���*~�����A�rS����?Bj�֟V��;ݶD�5W@E�A�4łj�m�.؄�|��G��d�{m}M d����?~(Qd�%	9[��yv��E�R�
z{������r��*x3�	�� gT�����yq=�P(��@�j�,�Q��r#�S��������.8k��Ʊ=���g��SGZ��p�����ٙ:S��M6R-�*@zs����̗����4�Vi�V���`��ݻ{#c��|d�\���O�F�X�ϬN�������d��lܾ���d���L2s58)H�ð�K�	�@�C�xh7K���;7�)�d��m�qcn�D+��қi����S���}?V�k��䢋=��"�jEVI��|
���w��O��a�x�nU��17�zq�F$��S=�:n�2���ѡF��(g#Pv_�!�Vz���EV�y2��w���Ӥyљ[Y����FL��s�lHI֊�)z�'J�J\6(�n�ԋa-�"�d��hϾ�7��A��f�OH�.�^� Wz���������"\Xu�Ŭ�i�$��T��F��<Ƒ=㕢�|*+NQt�0CS,px,q�եp9�N:�`�G&�V;	@�b�?�����n}���� t\��#��|�����[t���#�qU������ʠW���. `��MB��X������0ߴ�1��=W�m)����BZ=� A��=��8�+���Q<o���&I@1��{:f�H�AY�8�+�.,�
/H�ԿC�r�?{:]E{�Vq*�-�Ќ�.�d��2�VĞ�}P��PE���B��G��F���᧩Iη��!1CP�j�ٞ�k�V�_-���PqS��{���8	O�PN׏�� `m��CvMZ�t#�x��U��GKc�,������n�l�ů�6Q7����J���4��8���I2�H��)L0M!�IJ��>R�/��>����B?nk`����C��*m3��_�
��W�;j%N۾��b<X��Ȫ�
�����B��� i�d�'Hz���N���=�1O�gQ�j�˚;���1o�����fb�Έ�[J授��Y��l?���n�c9��{����M�����g�*���ރ�o��{NnXD�f��b��
�zd]�ԗpϤ�;�q* ��1�NP�ȯp�ȧ�����\K�%�W���<�� ������Gܬ�H�0���:�ļ�þ��� $1K�l����z=��;k�[���M:�?ݱP<u��ٹA�'��5FQ�JJ���]/�ћ�C-+WXEݪ��G�܄���Н4� Fz���_�`�� ǆ������ h��������5�$�e{�ere�o���ؑ餛�@�M����u�e�dY��X#o��H�,q�	���*A\�E� LDl�B �i�V�Ӥj�v�s�f�}�֙:�c��V.�c�Ć�	�f�$�,խ�����ش�6�.�Wb n ���;x �����u��f��yox[g�Պ�*Mq�I`�O�f�l��� �:�_R����}̪'��ވ�Kk���������:��!ieH��Y���� Ս�"l�{��Í� ���H��w����-�6L��Ċr|�?���a��;������C�GGe���# �*��0���^�C�'��'<�e�خ��Bd��.hy�i�5�q�VHug[����x`g�k\x�!���Uy���DbL��N �l�{������,݉��l���EI�ǁGksd�[��LWd{�е,Ch���n�h��~��.:Aܘbۻ�Uh๋P4���*-�Z�f�19���G5
2��߱�Ą�uf�D�?��b�3�����*�����o;w�_g�Ӯ���e������щ��D[�6�IK�	+u��d��:h�&z���o�DW+�CO�b)�Z ),�[����h>s1���a�d%��TD���K�����$�ѵ��n+5Y��T,:7�����a��ب<#��}#m�y�Dͼ���{Ò��!$�-���j_FLp��RY`���
7�KK�T�WB�cy�qbf���������4��d��Ү�?$QrJ��C����׳��b��}����5N�ey�^�~��=)o��v��7�Gq�uǬgY��
�^���C�M�����1`�/C�n�ܘ((��)�V�c~��9�#X?���0B���t�������%�ǈ@(x��.R0f�1�'�	O��O�k��)��J>�*��k��Ff�='l��!��	�?�������J��(�[�Hٕ���Ѹ:�(9����-\������7�.�O��x������eZo�o�?�'l�������4�2���aw2snC~\2��lb����[�4S�*y]煺A��_�F��Bu�)�۩ۧ�X�x�-ͥqn�'�1j\��I������r��|�H뿥����u8�e�^𡿰q��t��;Z�0���˔ͨ�%,�7��Z��������9�A���~�33x���$w��=ռ�ɣU��^xuC�XO6��7x��D�,��2��_zot]'��5��)���{Z�T�A۪O��g��> �ټY�28t��X�4$�$�ctr>K]��hv�߀ ��l�K�	���G�D�A3����p�� �c��� %�n���`�l[���(T%��"po�M)�e5��^�p��-^T���k!1V^i���#�Y�V0�F���W�*�m.&���P�XM������ZN3)[�G�vعJ�
���O�PPE��;��Kp��	`C4���6r��8��*Ae���A~�x�J�k���j�l>/�s��Փ
��c��a�Ᏼk�xK>T@OEE��}�&L�*�Bt��W��0E�G/�����N���c<&��̣P|��[>w���5&�Ρ]�L����p���вe×�n<��ۗ3\;�%�6�?AE{Pm��~Vû0H��}�!Z7ڒ�`�DB"a�l��r�����ؒ͟yV�A�f?��	��&���|������/ �*)D��o��3(�yr�/�?�SpZ��=$�3�]�,���Dg�D��(C��?e�G.�&��^��(;e`Bb� ���n��u�0J*\ &"![��A��m�F��9p���It��-LW�7�9"����og��L	$�O�G�ݱ��5���������h�h�'�N>����W���Ad� i��w� �\���� ��C~o��+��-��F�.+�/	qж��Kd���Q7��B~�b�� �������p�/���%�W��,?uXT�L寈���Z��$C�*��[e�i�>��ۻk��@�{��"9�SU��%=�J�������-Bh��4$��R:!�E`�U����Rs����b�a梻wɄi��H K�����)<�=�������
6͢z�h�k��m��5$_2��X8,�!�S��],28F��n3��[Cݙ,)��� �%�������Bx���t��	����+�+����� �_������"R���M�0h��w�UAxK���X���+��XPՑA�h�86�%�!��zJ��?I����O
��6H�)�Y9����/Q/�9���i��{s'+��|6$,1lʚ�
z	D��GB��GrWs��� B$,(���{���5Q�',��I�I�3��-�[T�A_�{. �J�r�]
�A^�G�G�,�pg}eY����#��۫At��c�h��w�]�/F��-%m�o<�m��E�Z�u�S���c*8���$�h�QA�Cv;�$��yc3_��Xt��,Q� �{Pz�+�-�'�&tL��=�i�xzq�o�aBFzY�11�����-����$�Pw�a�Nb�%ڻ��o$��Q��7>��no�4�>���{����vF;t���5M���B����hMl\.����@�G�c�C>��ע��9H���k��p/?y	@�i�
V\�]�M��o���C7�/����k���b��`�G��j�L_e�ZC�F�z�-�	�ҽ��@#�\7���U"�i��:'�A��-1�ELPn	-���͉��02z�w��+=�/�9�O?$z����JO���h�u����*��d�R��5�XZ�c�շ���s��.e&���ں����0 �:����=��*��g=��D��=m����l��LQ3 ?E����0��H����X�	�u��+��Y��tC:j]�c(�:��U��'d�-\�+�d�eK���X s�lW�VJ
c��CXV���#7�[�x�W�r(R&kB̕�ڏ����dH@��L7�g��NR��oU�GgegD�����pE(��Ǽ	�Ǥ�]Nb0Q�r�%bsᢗ�	�l� �V���\J��\1�H~�F�~��%_X�%�O�@,̒q����C�.���� 3\�	8��B|��,�D6g���+�j�%J�`�f���>�`��� ��9u��#�:h�؀��)�K�Q�R�^�߰M�$���5�j3�Zm��д����U���&��Xp���R/M���5i�NYP��O;1Y�Qj�m�+����֓Z/������ba�<ϳd��DL��Q�F���.��[�,�˻ 	���G���+���+"��Fz1[> ���K}vc���Q����_���ܽ׭���,l�lk3�o�eM�R��.rFֵz� 4�	�}�x5C�x�G��sV�]Ƕ��\�m��o�|\�:�d'F��:�P�u~�07[*Z��ҽ��(���hv-rǨ4����n.��Q��H �rd�,*��r����e��B±�.��\���g>��R�D'���v���I�4ɲ��Td�1�f��2�rOV>�(�J5����$�4�p_<�������h�C�p�:���-H�X�s�ߌ�@���o<U޼!�a�u��'DU�k�x��q�^�E��Eb���vV���,-9����Wę�8�#g�$&�N�y�;H::�(��:�ܲ��d�V�dvA�� i��������BK�dnJC\��ш/��M\iPJQX>�@���f� �f������<n>֋���ٟ�`����=�%�����	��P�df��ߚ�K��n+��Z���,^��"X����Ǣ�9����Y�� ��+��uL���.d�'�;����Z��I���m�5߁'�e���9�87��������{�ӧ�w������,�{l�y��{��޺u�A|�1�ٽq�7Ss7�u�g7bGqE�,Ұ�ҹzfU�D3|�8�s�!lr�A��y�d3�'�{�I��`e!��~Ѫjv>��-Ċ�SI��_��;���y��agl���O�@�_��c'cxt�l�V���ɡn M{����e�K����~Z|����u�韅/ײ�!����ײ�8�[pv1N	��L�=�C�L2�Q�HW��@��as����W�Ƒ�~u�W�ly���j߆R)��ц /f���C� ��vfNl��A�ɽ�'�Y�(��u`�}	��۳��00��μ.+�vGLDm��8��/�'�_n��A1�=5�_�B�ل����ܩ�>U��^����lXAT�u����ؼ��B)�zV���KU�u0�	��l�'2 �"�3����uϦOӊ�:�2����G(3X�I���bk4�sn׉��³�Ls%,5u����)�[it�#�%�␙*����� �M��O�%x�?���׾�o������= �f~V��&�������B�E �K+��۝w��?�qW�9W�"�'���"����0u`5t�#�����2�	U�@W���L�-�HC=�=�Uy7�i�x_��3���d��{B��� ��K��=%�Z6?�:i.W:K���r��&rP}��ps���.�}�T{��,��C���*����Q+rR�8�R�&j���c2���W6#-��S�k�;�!�0�� _N��#`��4�/�@�hU��ڭf�;Bg�6����y�[��I-�?�*���C�Ʉ�p%�)��i��)N�.)A6�����g˝�ۨξ�	Y����c޻��D�p�ޏB����{o}�c���]_,-"��q7JœF�Ć������A�u#�P��\�,s�!�au����<�-}S��c֪��;��<`�=g�@�m���*r�����l��AӔ�4�2����@i�%ۂ�0�l��а��j����"�/��np�9B��ϓ~p�z8GR����2BĒW6��H v����})8�,���8�$��Y�Am���V$�9h�{cl_�ڄ-��3���z��0�� C<��(�38�<^.4�)>We�+�0��}[�Չ�*�.�uY�q�iju���#)��[�y�\��/#]�Om�k�,������&��k���C�S�P*�2���@���TraE����Ⱥu�{߾	/b{)��[���&^A,�Ӕ�H�Ƀ�,Ᵹs�n�_4��>y�4�6���}��6b��a
PR���� W��}�#�]0��r��t�귤2R����nVz��W���o��wK��[K��\�*T����P7�-��L=�YcD�Fٚ,���Z9���4Tn��o7����L�s�>�|����Fs���$V���H$�������=v�W#�Y���4�t��)]T>��X��L��w8�X�1|�J�ӿ���)�N�{!��~�N�:7�B �~p֨��U�`@�v�m�4*�����]5�t� ���E�?O�4��Y!/�j���k�}����A��hȆ��gU�C�A�X�}:��+ؤ�~�����"}�A�k�^����>>�x��uUKd����m���1h�B�GvfS��Пq�_T�-J�)�cJ��~O:(�Y>�o�ᕖ)��
�E�.�ɦ�n�!�sE�J����=x..&"O)��/<�vp���z�����kdh�q�à>�q1m��3vQuEW��/�r�֝����̊�e���6�#�򵽘�����R�|b�E)��ʭ}�����O��%x<�N"a�Q��}����7�ۨ���f?��<��Ӥ�Uɰ�l��D	>��A4�n��58�G���8���6�r{�� Y�6�;��kD5_X�%�R����y� &o{�nROC��.r���ӽy֌�r�5�gt}�!G�_)���$���b5�H��=�/q>&IMc\,4}���Kj���s�So�˙bC���q�?���hjnA���
_�v����ik��y%��A�p��i�2�B" ���d�G��A6{*	�<D{�.�&�F_��4t?��3��G�
�|WP���^n�9����" ����@e�/�%��3������ېu���V�0����W��{���L�3��� ��z��B�)��~�)�c��}�Y2>W�}�nG�wb�I�	�s����_��hb��01���Y�w�#�μ�����D��nT[�I�#�+�ʲ]����5H&����W6��
�ҷ(�6���.����7�4}m��`�ŷV���ṊH��o?sH���&ݷ�I+"��I����Ҧ�uDύ#�r��fXSV���zb��y	�ӹ��ZWq�� ���U�H�5�'�`堕�&ļ�e���h�=sh��RH�ƢQcwQU/��Y�����F���N��>kBf.ɞ7ⷌ�ȘȪ�����$U�Cv�W�;��V�v�q9*�:_F�Q���0�|v��|�I�$Ĳ�deΙp6�F�-h��5dl5�r�W&���q�:#�7bxt��]l�a�8�u���%߽U͆�$��6���/Z�+���9��N��;��F���\���k��tnV���a�4��*>�ؖ�Y'�~���[#T�:���B����(0�T��<}>��VXbL�?Y"(9��t�)�gS>Oq�)���f��(};������,�:�3%�[� �R�`)�@�Ag�����zlh�A�pvoU!|�����.��m.�NHe�E�p!`�^���Qn>G�v��R�WI?	��2_��`?},��kF�G�LY�`��lM�p�5�'��go����.�l��W"�R܋O
~��!��9�&(s�D��t`T޺�}��%`t�aY��]�h���� O��l&Є�0dڧ�T���j���BU�뇜�5�PR}ח���}y�nhjQx.o������Z�\*���pZߕ��6��x���؄�O�:r�C��NI�b�ۧi؍�s���ko�G��p��߷ND6�Grٯ��{���h�Y��z�ꋥ�xz
�kξ�u�~k�#�D��m�ڇ����=�Qr~�1P��sP������0w^��,oIL��{��?Ӝ8��W��A߇.�1>W ���N�݅�T6W����y؆`Z�kO��Њ�X�H�(b�+2��Tzb1��w'Uo1_Ḷ��`�ص��6 }{=��C���e����k�e�2pE�4������+x�ߓ�WXd���;g���iT�jF�J  ���o�K���/e�~��⤮�����j+��CX��ZT���-�yĢ��v���;~=:^!�v@��������-ӻ����A��`������6�b�.�t�Fl�|>�1z��|�N��3�pk����y��-��Ф����^��V֦�>?�mI��.�MA���U�}��d�5Я�2��z�T��!�A��
��W$�^l���4dɈ��~�į�G��e����>:p����K�@ �V���5�jO0�8R�ˁ�A9s
�b�ˆ����"���B��P�E����"�?�����6�7~d0_D���}
�X�O:��EZ�t㪯%���2.���׵���{]�b���������a5�6��P��p�6�Iv����F������C�����l�h�7��|��٘��h�N��f�ys�2R��*-zA�֞p��H߉�d2�B�|{;[&Z+�9{I�@۸6�I�M��JU@��wj�c�g9�W�Y0��_�)3h2?0;@���������g]S �4���q�&H�(;��sbn�ǳ�
j�N�`i��Y�D�-�K���Ƿ��3X����FB~PzC�������Ȯ`YԤ	�3 �&a���Lz�+����v,J����X��Sk�����;�)*�Q��E�.2 ���ܽ��c�qw�anT��r��E|�7�]�}������Ƌ}�����r΀ƩNȚ�=����"?3j�� 7�1^X���-~w��-v�~�t4����v� o�)ln�{�X���5��a���vn!d�F�y�ݩ��آ�t(1x�~B����&�簗���2<���(�§E"�u�?6�[���XteɄ1��1���s�AF��KF!*~(TK�,.K7F��:?��:J�v�{�-iJ`$UDrv��qg��ŀ*(�y��BM��V9�Úo�ך�5�Fɇ+]��gKɾ�hMeǪ��s
�N0��ǒ���GE�\g ޥ�ЅdF�5T2�����Sc '��}��%FYN�t�H��a�b���u���Zi ��𺒻A���� ~�$̍o� ���FN}&�n.!c�Z>����z-<:�p����Ia���6u���
R�k�bĴ���ݹr�5'��orq�eKe2�U8b���1d�U�j
ι�K��W/(?�)���3-�h������
���$(��&h���f��|�,��b�zN�C�����ds�W��?]�n�#*���p2QXpg?DWi��`v8���#2l�hƐ�T�+C��F�&��*���&�WvϪ{P��*����o��}Q�Ա�Y��һ��M:��ΐO�&7���������E.�@V4�'�����;�S	�U�����{L|�����
��TW+���D��)�#oэ��#V_��;B�D��P5#��C���5y�����<�Ppkv�G -H��SɅ�$�Jb:�n��)ax��4��Z׊�c��u�K�)R�.�����Y���0W��[���0(G_��=�� ��(_�?��Wd����?9:Q�a\Ϳ'�)7��C���x���ܣ
��X�>��ǃ_�5�t'l���`��`�������s���D��w� 
J�C���"����LRgT���>���t����~��\�3Q�o[B�C���A�aH4I"�,H�?�m�C]�@+ha�}ԩ'W��vqAmC[9�͆��i1T��L�9~��KW�б���[ؘ�!_���
�v!�<���%��dU�?�Q�c��8a�� D%���Ͽ=_�qpFh�-�:����Y��I�bRw���]Oɘ��w_���rC�
�Z�I�&8�=]�>�o4˱y�����<��MG����hE.�-�9�Q滤G�R���N������?��U�1	𰣁V8��v��UFԹ�� �7�Շ���V�D�q;q`�_P���8D6���'�$:��ޛϪA����)e�ǅ+u(�M����v�'"ш��pq�����;�і�/F��D`B-G|2�!i6�B+o�궁х�ⱏ��0mB˱Z���w�^m���	�)��1�75Am��E%���Dy�\h-[z@�����e����N��՜4Hz�`��M�S��! ϰ"�TpK�vv�c�apýyz��X%�+`X�ԊР0z�)M/��8�c�SL�Q5��~��R�ݻ%#�ߧ���㘚:�7�Ƥ��o�t <@n�qdj;dF�դ@F 5�c7� �\ba�GA�௃]��뉝ʁ3@�0���?E�`]-���������j�KE!:���x6�6�9�������~�M�lY��_k�Q>|\±��"*N"�D��r�N�߶4��̚�`�ߛ+��Z�d��c{����M�e�G�۾V�Q��	 ��C���v2���U�,���Wt�vq?F�JKs���X����Ԕ��*��"�����&GN��XUH�N�.����K��N�U�գ��an��:�dVr"2G��Wp� P���j�ї�'d��Ѩ_-Dg�j�فww�������H�K]�#�̳I�~$���x�FtE��j�.���r@� {�έ�%����f̆�����03��ؘ cP*��`��S��?qM�k�\I���<��Ք|F��E�*b+K���49Zŭt3:�f������Xӧ���}���gv��J]�|y裪��^G%A��Is���	)������>�a{_��ü<�ٷ���Y�&�ʧ�&r�������ܤ�`�����.��}ڸ[���1Z�r�(ܼ�ֲ?��5xl�,8�/�3G5���<W	�x뻩?��`�ڎ�VVѽ
�=W\�UBf�Q�3���AZ<1�F�����8Nb�\.E1R5�P�v����<N�j-�p.�}�Ǳ�\Њ�����Q�	��d=p�PV� י���pΤHq�t@���&ո��#h5oQr�)���ׄ^��<z�R����fۣ��\����G�[�o��*�n�̌`�Z���X�Sء�̑zq�D"p�f�r�ͣOi�\�/�"���D�G���ԙ�<��P�ҞR0��:}U�"��a�`�vN���K'rvߔ��"��z���Ũ�('��>1�[���zw����-���s�.��'�q� �Y<�ŋѱ��(,��x=52ト�+bݏ��Ț�J��3-;X�L>@s�L_x YA�؆�#t�X�ǒo ��0�7'��0K�`�T}f ğ,y՜�,�<5�u}�j���e ��Ţ�ʐV�߅P�
8+vo�r5�BM;np��6&�LxstԚ=P�S,E���Wl�hi��4L�>H��TF�@��?�Ͻm\7�Ӭ�	��})�T=�[�C�{%ڛ�j�� A�o�̽S��@f6r�Ị�^���о�4��"�6Z�oDѫM~֪�]����JYɀ��c7GZ����5����ħ0���_��):��n��-���u�^���`��fK$g*�U{��;WLdd������FkC�������K3�u�}<�J�2��W���W_�a6� �!����%2V�ӗ�Y~�t�̭��D3��|߁�s��jnO�N�v�ڻ7�W�9�U6�0��?���.[R@�m���3a�z���PgU�G���,d,�o&6�n��ي���4�&P6���  %�@�ǝ�*o;���A���R=�p���H=�|٬	�U*�=𼜩��R�@5�R�����*���v)�8������ֿ���ґ۹8�{��KjP��ŎS�?�y�a-p�� F�k}*hW`%�\uPd���Q�(nal��r$�z����pe�4N�Ջ���l�������[�B>c���[�]�&�Rn���:/Z��7=*�"�s�o��wZ���x�C+��p�εR㱖J���j�*�4���R�[3���d��J���г��`�dpwJ���(�5��'���0�܁���[�U�p�!�)?z0qpu��MO�A�ۮ��xm&�:J�f #6�)���n3���L�@Ֆ�X��&f�_r��ܹ����л����I�23���	���I��/Mh��*���cF˞&/ȝ# M)?1E�H�]ei˲�?��G����/�*$l����v�Y}�+�w�F��n�ۤ��R�y�J�[A V�A2	bozk��-��%~�Jb�\�Fs��@��4� �3���f8K��r�OZ��i/�%"g�v@J*�3�`fQ2J��a���-��[1`Ǔݳ��6-��(�>��;�z��������$˔y�	�d!x,��W���X_��41�h�6���$-I��3Xp��k�w�2��ȶ7<!_�vj]��|��IG&�K(���<󾦷f�����k�_�ο�5�6��ѫ����H/!:��+L#<1��H�D�q%D2�4����g!��	����`�+�Bj�;�J��8��؁�ؙ�$��`>]��]�P��(e�/�xس�Epމ{�nr�<�;	y���dU1?��')_L��19Fu#�A��Ci�?�'!��EXBA�M��|�Eܽ��b���� #�1�v�$~��k�;u��m !�>e�Ⱥ�@�ѫGx������)��k���;����i~�=g�\a�Т/&�Ոg�S�6O�h��'a L?�Id�62���L�+�������I|r�<\8��sBZ�Xb�TIĪ�N������Y�F�7Y�O+��m0�s������3�!^O΍���!B-t��uUh�5mJ�9~a���Y2�'���;\"���-�Ʀ�Mů�(�;���gC5��P�����������G��p�CMVsq!#�Y�P|�t���C�n�S��{`{�z
��=���h�$A�Tq��\1Z��M*v��bzF�� W��yҐ�'VvN��Z���\��C��t��	���'���/�I���:�|�;`ŔP�	l�79z�T��_�4Y��PXL��ڐT��֛��>�'0dcՖ�(�+~6;�9���O{^��*�Sq9��z��+�~�1����,��`}��=zPT\�j�7�(c�FݒTO���[�E�U	�l�*6:D��0��<<�����J,%�
�[\�"bDξ.�v)�G�	�h�kڋ"v{�U_�B�&�)G׫���*�?(í�V�mf����_/0_�R�w|Y�Rʘ�4��*��� ���æ`�����M|�b�#I�*#���ݹ�O�u�4��vH\��-̮˽<���G���W�)`h�����%w�j��Z5#c���S~���x�<�.�K�SM� Dj<a˔*Q?�-�T���:Dxs����9Q@!?�%�7,�� �(����h���P�[�����ٟ)ɯ�֍����:d�8�j	~�����߸��X��x46��������A�؎��~+/�^�M���uQ-��3�k�F�P_>�]`b<���N_e�Y��??MN�eP"g�W���	�H�~��L8�68B͔/�H��#3�&��Č�	`�L-�ʳ'�VQmx���-�(P%G��j�����ڸ�H��
w�1X��S^������'��fQ:mL8ʨ���fu4�\�0������&��w��GP���ސ��}�k�U����j8/5��	RϜ6so�E�¬^����j�e�V9c럟N��F�*�Ct�G���{A�t4��ͼ�u&p�v��X�����#����YX>�Lk|U�Lsf/[��c�_qq������cv$K��>�򭸠x�:h��ۑZ&� ��eoW����#m;��%+?K�B�S���G��*�_�W������vFv�7��h����V��p0o��d��R��(��4��_�a�T��$Zn,y��S%�?�	�ܠ�vd��[NB��o�����sb�S0�ل�Á��$��R�#�y�i#Ip��H�2��h$��{�>U
���T�����ޤ����8F	�^D�ab��z�����̔��^�����$�Y�d�)�۲���Xc�7�:RQ���O������ Ҿ@=�`̝���w�D<�I2=�|r��C�s&���u�=�׉	���{��/�%��Z�]i��.���yةR�����A0��!d���3�K�c�!� �[a���B���V= ����J���ǘ�8C�f.zt	�c���_�1x��u(��^�������g?�^���ԅ�1������El�EI�9h33nuyq^��[7V�R�@A���8t
��լ�ֵS[U�)|�`�Hn�`K��j5���+V������7���,�ג�F�j?b~�
�'�N3*pF3h�ph�1MI��P}L��ɜ� ����{��"Z'p�q|�����W$I3vr��6�2�G)�y��hI}ߪ�FB���@��_������2�l	����A ���(�rߘo�U���l��R�e{���1򰍄&��.˷A�.*��7�� 1W�h�I�';+\�t�5��7����d�A\2�H1>�j���l�25]����v����ֿ��#��* w�=ၯ4z?��j��ݳ��`e����D{]��܀ߧ8�����4*��aa��s�������o�-�ч�	6�R++� 4d�0y�mj��]�?�Rz}R%nj�+�Ũj9��(�E2�|;P<m1X۲chR^�$�K�[�p�A5�pR{b*2p]��?=ԭL�}{ql[��PĨ��̃
�٘�S�5���n����/k�>��4�� "��2�N)�jK�{��=�Pj��N��:Z`��n��<@�w���)��1n{�	4�z(ރ��"��÷�
Ѯ�Q9��7ߐx��d�'�'\[��^��u�{�Ze�_���0�ճ�{���rNf]b��p��o�Az�l�Q]����2�o�`n=��=#i�]@�Y�61>j0d���v��U�\��� �7�D��y�a�K�`NC�0G��5�/}wHN1�u��A|G�����^���ɨ��fG��7�>��]�&Vc3}�@w�0��QLp�?��hۂ��~]fpb�ٵĂyT⚋fK}�K�ĆU	���:��FA�A5�͇����ޘ��~>�l_���oo��$��Cد����\|'5P���8��V��X��� �X��Da����_(�3��5�_�'�o�rt1/R�9z����w>�jL>�Oaϡ;f�R��k ���,�*����Lϖ�h�ᥤ]@J�J(M^z]�H�U9E3ܡ���w�83i�ʱ��3�Ro�����c��%��P�b'�HX� ��	-9cCG�4":�)�x��tqJ�ޖ�Q������}=��Q�N�~���c{�Fӡl���U�����������5��x�%��>����?�Ͻhq(C�t� �������4���/��E�������>����[_��U��Q�8Q�.��MӜ��3�4��5�,���bx}�3���'��y�k ���,�?^�V� ��l����?�W�,Zu�5M(�J+�>�����Iʲ�i��4�+�<�0L���x�O�`�>��R�L��_������t�g$p��G6�s$��������y�F�n�K���};?;�ߗ6%|��r��/�D����VfDA�+�#��NU?������"�j	8�.�x�{>�I���$GM���%�DEB~���	s��(m�������� �Vp�����6��ڀ	/���*�`U�6a����=��N��� {\1���v����zֱ��:g��і�"�pH���Lr�E^S=nvX(����S��`G9��my�:��
6~X	��{��O]tU $k������zmHk�{��h���-���^�JH'T��1W�̒�y� G�>��:��jP�F��ωȕtb^ҵ�o��aʟ�W^ [�^�d�+�������ޏN�^�������ntH�j������1#�`���y��h�&�ٶb܄���bYW�l|�G�{��(���3X��f�$r_$����n��9�����s�!����c���@���פ���8��$��<�x�7	�P}Jﭸ&.���+�}喈VQ�C��T��*��p׫�1/wq!��|k�'m��kU�CbP���'S2DH������\wۗ,��o8#�ٶ5��{ݯY���9q�/��^ +�Sȇ���־E�$qy߯N%���e�߮�"�Y�)�*.�&.�v��%`��<�Zsg#l�:>J���j�D���X�?�j�pa�)���9!Az)q���_����]�f�>���Fh��[2�W��to�oY(OP��t�X�z�`����.�����Y�f�~���ѽ�4�tUx�Ð����tD#G��a�HP&��2c��V$U��f�XgY��:�y�I['�N��^ٙS��\��I�k����& tJ�9_І�-Z	��Q-u��+[�)����ǀE���=̼��g=�=�������� �bWv�0u��
��Ty�8,�Oֻ��Ҧ��gX&��`-y�m�R�:ay1Ȭ�XU�zt�'�a��8��D,ۘ�� Ԏ?O��.�4�Ƞd�7�	us�UJ3׈���{��'R�?�!�d6
�	b���Na�c2���k,8�R����8���4��d�xNds�|U�b����0��e�'kU��u�X���(�-WaT6S-��:����m�hC@{�*��@[h�X��x3��7ʏ����Sʊ��6s�	�!��aq���b��Z,���X0�) �L,p��C�ג�X�-�.����Qb��k���0�e0b��-Q*��RTA������@�gV�P�/q̱�V�p�������=�NfT��XqN&���6N��o�Y ��W�V��]f٢&
s�����VЈ��@0��r@�Õ��ϔ������w����;_U�\y��DT��p�]#����Faє4�W46�S�����/�>"�ma�5�MuK� �0r�C+�����5YE|�}!V��S�TJ�l{����Mp��~�<��sG�0��oF����;��	pǬ���Sx�{�yd`�@�[��yj�,Z�[V0���mJ�
%H��� B�&��x��������C��<�;wF�L�.�ŕ��/T)����)���������泜_�X����6�)S�3IдA����S���-��uo`�6$��;�Q%'Ev����ҕ�[�4�k�:f1��0,z.w�Q�9�
�ج�vsi�O���K�!�/tф�����V:c}!�\o8�t�_��i魟h�t�x%���-���o0l�sooH\��D9���m�N�I`�m���5_�Wĥ�vr�7d^�X�s:9:�eAy��e��6L6�^e,h�y��Vְ\���eF89��\��3��&Z�c4<����j��
�Oi���/�^��7�	G9)��� A��h��f�5���ĺj���1$l5"�����Ƿ��F���";�+K�٧e�C2�Mo��#�r~��uŉN��b�9u�f{2��.�Y������ҕ!i�7C�	��Z��l��_��.�q��צ%�T�e�6��I�<����A��sOL�Hy�K�#Ս��))���!-�'���Zɲ���S:9?>�T��chL�����pBp�jWVdN�	��� ��sR������@�_�.XQe���	lt�0��۳;2�v�%������Aw�#���4%5؉�}�4��QT/M":�)�촓4�Q��w�r�X_��5��� �*��."����G�l��.=]Zf�6��Db���l�����a>��-	|`�r������(%��^2���~3�H�,�f��sđ�(�_�S+l`�#J��g����^�@��/�	On$K%���g�@�zC�<I!�S�W�^�L%8O+Hh|�n�'rb F�[i��b��#��c��XA�㭇�g�ӍgXqpMԊ��g����UeF���
�ؙ,S�+F���]��6]���v��N���E�K�=�sf�v�Q��{�a���n��xڔ��^n'�����Y�)R��-z�dY���*�I�_��I��<wێ�c���f�������[(\�?쫢]�U�ھ�C����b��g�f�G�	f� .���:�Bx��׳�%	���T��*I��@�0���-N9qBv1`s�e��N�ɰ�Ӹ���#<R�I�%_��'⣩k%��C��ļD�|�1�V@o_�ՅKFc���j���}��m[>�g�v
��A���ASd���j�5PC�;������oO;�	8�H���,8Y��ط8E,��Fq�O�.�5�x	fs�3�����V�DS

^��3���&��\�y�ۤ5Ë&��Y�ъ4�s�j����RW}?���A��!�$>(�S�;�hy5�[���v���?�T�5��-[w��UC;�r�
�?��ʺ45��=�H�)���X�k�%��V��)-Rw�z2m��[����G�hCo����f15��w��¸��.��'9�p��)CNm4���A�"�x��)��|2�1��^Z5i�Ԫ����m�o��.��q(ލ��%��4L8R-�pI�Ga.1�Kv3Zv+r���۟(qT	��7Z�ZIc_����������D�\��Vf6C)�eܩ�;��X{���XL)O[?�q�������xX����a-��D�Nٛ��+aW��*�_��Y��sw�T@S�f��WA�����U���aM�0�k:t=�ե�:��$N�`�1��;g���J;Q;����楘���j{%\n�8z���|��z�^s���I��CZ7�t�1S���e��S���.ɳ�l}�z<`���B�z��i����!��mP��%�p�Ct4h�kGt`�J���Qߛ�������/�9y���qp�5	r�!/(!��U����P-Q��q��MA��ҴU-�B=w`�X/x�3�$�����ſ#au�X�#u��(�����$�< @�@�;S?��.E�$�RjJb�hP=F���?��3npj��|�ƙ��T�����QV��y<Sy�p�e�N�<�*���8���X��^#�\
䛹�N�l@a��rӵ`<���WN/���(f�-e[��[�fN�:�$�J!�#HW�=��eGB��H�e0A�p�,L#�5��u	���"؃�\l�%�q@�ly5�6X���G2�0�o��[Η��t�' 'Nz��g�VB=L9�X�>0���
�ΌL�Ğ�����S$+%kMЫ��}�y�x�)��{��T�p<B�X�^��Ň��%lpY��F,�`���11�@�;���������~U�����z�%�=a<��KcXg��(/Y=*��v:��k'�#���3 �K��<�����#�I��!�[�+3$��R���FgH��3�RƱ��꬚�sϠ�U��>H��5-��ǁ��c���_cNt���Țz����aD:-)o�*��h�Pi�U�,M�~Z���#~�	ӑ�v��+	'� �����G�w��X�%r8^*��
��wfZ����o�w��M���`����g㴁�4.z��Z�f0� ��J2w�4�.VƖ����
��]W�.$Ę�|%��q,���� 0��[����P���ᐹ�]h	G�ݎ�s#�hznV�oCu�ڥ�Ɗ cU?��"��:��QmEՆ|KS��^ه�z�]Nj����$@1��D�����k,.ޔ�������X�"<�?����Ϯ�N����������5�1*����ig���nC?J�;ؗ�Y&52�/��>Gڥ�z�J���Ѱ��큉x��x�+�/���SV9`
��62�go�1x�z1�'͒X��uVM��2�'���$�E�xo�H, O��v�3P}W����\�� &��
�s���jI�C+�7���78�P��������4'}.��&��������:�R� ��~r�y�3��f�~��xo�'X�h�2���#����׺�n{:�_/խ��M�PMyz�F1�xDt7�t%�:UK�>�e'��& �9G�6�F+��p��]�w�yC�ʝ>�^��B[���t_	�#����ڼ'L^�xu"��k���pgj�#k�uY4�͎H"��A.������.��J�(ل��V�O�G���ls~�_$=0�^d�(+S��+܏�a��( S+�B����{���}8�TB�颾?�M@���̈́�ۋ˶y��`5�IUw�kI����Ǔ��B�t(y���F�'�q
�rٔ��x���+F��s�I\���V�y�w��dI.t�T�0pLf2�]������|��7�� Cp�����q�d�l�ݏ{*� {n��U�F�S���{&5��3z����\vx@��6��x�9�5s9�C��1W����h��U�I�9��N�Y��%R��t���i�c��}O�d<��<����k���dM�	����Cv�m��ѬX`���0OD~����a��u�rS)�z5��읫��ރƿxv"�:?���:����c6HJ?�,�QP7t��W���W�ޣ�����&�N��&�5&{ϨC�cAbN�W��\.�2�4�� �����=a�#����rH��ۦR�ίBh��N|�0;�s���x"���{��{��%/K�\D�R�|�?k� �p��v�%�8j��Sі����%)�Yro�;�kǂ [�[A�yS�#a[^R*��o��@wx���T��n�y;��/�l�w㼮 [����m$�?�21�M&m�~�>�/<Q]��ɚ���:J[�N���U@�L�.��!���v��C��g�����v�|p@�3l�G�x��i����Q��VXPg*:x0`'&�&0�� �R����M~G��C�W��q��_�^9�B��/�ʍy��׮��D?�L����ꡘv�M���6��S0-c�q���� �������/(Ü~��/T.�-��d�	z$���)���fH�n�� Չ��g�>c��p�^[#I�b%�W�m�<Jx���U^��F� G�͑��W�߶+-3���a@"	~
C�)Yȑ
�L_���l$co<������@��67���{�1��ڸ���E{������wu��� ��C�vIߎ>��i*n��I�W)%g�n�b&��1��Y�O�� ֶ�n�C7H��a.�B}��7�D<��\՟q����ŵ�x
+}8���,]ODuy�!@FLh�2n%�	z�c���c���$ \Ji[�)�;5K�v������̵z�_�y���끊k�\����	ג����Ot�t�s�.&��R���V
�FLN#X��;���2�\!mߏB�ʎ�8�;��K���k�nƻ���ό�����X��-����f7��S8ɕʋ=��"��'1���z��o���T3��#E��x�>b�"#�B�E��w�n^�-��-��*��zu ��j*� -%�[Ӧ��˱��q�R����mޣ��Xުi5'��J�o��I��~Z|�T]�pN���h�3ʻ�T� iq����ߕ��EWV�A��dN�&O�ހ�:�A�v�dL?��D5E_�p����i9�X�p��4h`�����;�-M��=D������2A�P|\����x{�ٗ�dQC�3��,�>�1�~��Tj˔��%�o�RMd��b?Ṉ�2��2�,�/�U���s���K��`+����)�}o�[1B�q�员�
E0�m���Dx��K�?�t����h�=�G��*:gF.���T2���Q|,�
�A���@c[�3�/dJ
��.�[���̓wÓ���8�!4P�4R�̬�"A��W+�tdq\�*X1dA"sPis�3�B�c����ױ���I����bTX��-s@��n��x���Y�H�X�s��9/����]����>Cr���5B�P��f�W9p�gbS��qo}�V��v�G�c�@Q��K�P"�B{Q�eQ�������,���:�a%Bw>�;�@�b�ư��C��~�����Y1$G�>��
��i?Tǻ��J�g�����p�m��a����M|�����qk�C�h���a�R�7�/(����#b}�2}�+~�ʗcC�1b�����c@�eb4,�H�����mb��6/�o\]���Bk���.?���[���W����u�M�P�y�@H|�Gb��9�-Q-����~	�kj��f,c����4�r�U4��$ꋳԤ���po�J�FPdy�9S�7�$����w?���Ĥb�d�����8��;�0�����4cJА���A�66P��"v_��t�k��m�p(�$��^ќ�5�A��F��e�U=�;��9�Š[��m��`�eMD�0����՞�ۑ�q+'��!M���(I!RBR؂Y�8m{d�Jy;b�j)����Φ$~ůUT�$��7�ޚf�+���_�%r( ����ܾ��z��]�_ߞ缻��[���	{`��=[�c�������<F�S_2��y`�6�DK�1H��L'q�	�@���JC�ln^���r��S9,[f���M�Qw# )Lm�$�����?�@����p|�_p8��ydv/�x�����18V��L��|��m�(�r�VWb��ӷ}t�O������m��c�So����7�/�a��')�U;�:~jq���V�I���;����0HK}~fE�]�TqX�[��O�G��4�B�ĦO�(��t���@�<A��ʽ`<E	1q�nS-�������JG ��i�A[�T��H�u,��M�}d���B�ͨ�+^��{V!��o^Rf�Ѽ�������h͘�έ�'��l��6����`����|�$�G��;R�p������o��e��Q_�����;��J2&G�� ¢�d5ꜞ{9��
��	PY#M<�j�v%��%l�'�b	Nb���&r?�<W8C�K1-VCh�q�$j4k��+�D[wX�Ʉ���JRR���>*�5K~"LI�߅�#WJ��L�YZ/�;�!#`9�Q��t&5�R��\��˽&��Y����׽�2�`�h�F��P#����H;HE��o�t�%]YQ{Ŏh��f���dm�/���6E238�R� 1S�<5����&�@��������$)�����L�%�g[��aw^��v�?ǒ#�M��Ʉ�st�I��sB���}puSw\�M�Y�|��.��-����ȣ�F� ޳�ܷ�G�@RGhC���ǼP�]T�Q ?�cS����ZϾ��3��N�`��F6njB{�(��T��G�ô\_�wpuL��Lć���,��͵N	�+w���^�� �l�YB`(5���F�
�֩��ZDU����t��	�4����;�|#�a�Q'Z��Acz!��d����0\��#��)�Dm+����y���|�����;��7VQ:�k�3҃�/��-�*�`�JV���?���.��Ҵ��{��*G��9|�Bޭ��C������b>Ugc�	=���U,�ݒ���z��վ����Y�U4��ޗg�kQ��gdxB�}�8
6���{���.崵��Z�(�U�}�>v���+�"D�	\q�^=p��Y5�LP�v����z�����w_��^�gϕ=A@x����(y�7P]�Q�&��{�=�ǖ�7l�G6`����9��uN
���K]N�u;�p~�khx������lyYt�y��X;�=c���z�%�aB3�%�/.��_'�~�)���p0}�#�b�gY=�@�1����0���7���������*�}�B��C_�Y������-��h�m���t�h�=���[�@$F��@��>�"�K�u��h���	Uݦ���F���vB����lTz��vJ�\~��6�kR�߯}X�q���6_��X��BU����N�~X�С\�L)ls���b��2���7G̿�<0�!:���B]}�?	2�������H�i�}�W��wUg��3���'��b��@�����������U9�n-⁶,j"(���Y�(	8o�ؖ
��	�n�l�x���{���I���ezk`���&��F.��Y}\�OeV-���K(�`����g5�!��}]F+�x�tZ~�:��A+$�-� ��E�2�t?��=c��^CߢMé]��B���B~ti�b�p�2��Nu\���f�'�~4*-�\O8��q��8�p/�ҡcz��wP6j�%X��WSe�Ae�ک�z�G��k|�	�$�@�?�p�?3py륓d:	�!8���Pa@+�$M�{9�O�ĹѡQk�_�Ψ @~�<i(�c�G7B����,V�̛�"������*&�j��/��$O��0j4��������)�s���q����7���4�0B:�����8Y��l-��W��9�ϔ��O@_2`K��F:Vtv��ôÒ�~ |�{\h�(r�Q�-��L\��VjJ�Uǫ�}k���T�FR��2�,o���m�hnet���s[e��6`@93r�`c�&�>��D�#l��kv���=0� V5��g�b|{�`��ؽ=w�Y'����M���5(?.�+�3[h����n�C�Q�Ia�>���8d.y����;�>>�$��э��V�.%��u[�8*�ǻN�p�i%�ѳ�p9�I�bۃ�d�d��Q��{O�<^R���)9≫р��
��?&ӳ>�\���#Ʀ͝VEe<h�G�NP�&,7"�+�2��,y���2Q);�y����{�%� i+��,���&w��� �_�����u0$�ydD�N ^�Y7�����!�::i ���Df�)�w,�Xi3o�B�w�Z��Yy������>Z�[�4��!��3&h2Jh6[!�V�%�@#�Ɏ�lmO�7���fN��d��]z�yR�Sc϶�[�m����yEDxy}�m�H�>S����§\���$z�=���n-<����85I]�L��������E��$���8�Ɔl>�H_`3$�ŵ!�}~=�`T��׻��Gr��7�PfY��w��5s�7��c���u
��c�� �C"sf�Y�*�M_}��^V���E]���S��D3p��X[�`sٴ�����q�FX-f�Y���5ͤ�m�0�3L<I�'_J�n�^�[Si� �~��@AU�I���R�80�F�J��^�K��i(e~iמd4F4t���^fj�}������ZB��ShYB䢆M��BaP� w"i�K�;�1X��[�"�&s�7�	}'��іg跋I�`���-9mo>�gm2- MsU���pk]u�����GC� ��x���9��XV;R[3�
����a�EI��*G{�N�z���r7���Pi�i�y�󺟺���1�?����%X��D4�׀�4`�7��"J��(�-w�Z��H󬍋�@��0G�ZY%K�#I&j�r*��Q�Ӄ'��RE��C:ᩰ64�KJ�����U�/�&K���H�i��'�0�[h���Wʳs����Ӯ׽�B ՆZw|�׋�H"��ˆ8ŋ���n�M�5�Xad�r�uAO@�p{;s�>FQ�oE؂�1�-y�r\3z��%�'!4a�'됝�?S�ۀT����2�?9�g��$�0r@��#N<������qT���m]�T@�L�O&?�����'5��@�Q���5���|��v���A�G��x[�vNp�/��x����2�v��k�y{"@6�����k����"	"�0 tǽ�%_���zTs�4�}ʜ�����3{8~Az+�-�.4e2�V����C���3����ˤ���)3*�;
�Q������b��x��3Ų���8������p�d 'j�\c�J����Z�*>�j'2�G�R�^m�M���f�
2�g��hr֑������օ�dPD4JI3��OJ�Y��q�ӁS�$���'	eu���r���uO�1!]P^4���ɷ<,�2�.����ct��ӑ>�D�"j9
�sY��y���:3�0��ހv���7�xH���i3�#6i�8���zc�a�,���U��d迼���I"�6���t���P:�& �h $��3�nI�y�N`���U+u{˴��k,����	��$���$��"���;q�聋Q>S�3�ٹ\2�\H��Bb�)�3��uls�p�PJ�A��|�I�c��UbN�h�\9� ��nc𙵨�s���w߯�a~�+W�Ut2�Mn�V}�w*ǡC�����z�:(QH/��yZ�OM�-�y�Oc��<^��1i����~K	��eP�2u�7k��m]��vN�� ���
'��i,�9��Y���_��2���&i=�z�u��3t�t���Q�,F����q^�:8��6�� Ϋ�����{j S��g�����璡|��ѿ�{טh�� �`0��uhL��u�
����h�N_۞?v�m�)¥/\J���3&.�y����;�5�-�tX�Њ�S�M���� �|;	�T�ڏ���i]/���x�\a���ǚ������g��{��r�i�,�,=+?�_�)�ߠ�~���1@�9I@$������ova���n����{�c����*\�F�,���P;��Ճan�lt�^>#I|c:ݿ�u�/�zI�����v�F0�!�]&f�B�t;�P��c�4-'�| 0jY�`=7��Q��7��?�
��-��˜P;�$�s應K�6�QP)K�W�v�f�R�$ؒsh׺c<x5���D��T���*���RZ��1�k;�0�	����!ܐ��ڷĴ�Ӓ���3alJ��׶^��9�ʪ���E�9�n�0���r���l�����B7�H6�^�tm�Ҁ1�	�ص:�W�ft� tw�}�5JiN���L�6�Q}H}�#;ؕw�/�VG��7�p���eu����G�^Cw�Z����k�7���	I�ࣂ$ta�/'�`Gvk~0��'�7)�J�tެd��_{i93����)Ge'		vL��vo�xq*��Q
�W6LE���@l�{Գ��Ъ�}@
���tt��S(͝4���]�!�xcO�ƚ,�*I��s���4-6�Ơ�}�.�M*�Q�
����f-}�L�[`�bm|V���-vQ|�D�����>�����;@�SJiTO(ʋ�N!�_�f{-��t�Q�1��.l�f0��ڤx,n���'<��v���e_�c����}�����p  �!�J�7nNV��VH'�Q�����d�:����df����*������̩�9�S�<iI@ G6t�h�\��n� ����'��_�Q�lW���E� B�p��[Ȍy6p8{��x0oO�����=�R���q~�'�	?8C]2��>`�	�dڭ/�?���� �˯Λ�v���d����r�P�C�ÓEt����y'h��Ĺ"�H���7c������g����3~�(ǲ[�z�%7P�ř?�c�D���q�[�V-_��}��S9����۔D҉�LB�]��e��(g�5��8���+y>��U.%��z�@��ab�{�=D��)_Ш�2Sn\�@�`��9O�������I���bz1�^�c�z������!Q��)��)묗��n.]�ړE�����MH�8�s�7��ZD~�h%z�� �����a�l^�dE���I��FX��ҚH=i�!Nү1ߜ6�]��>O7+��jA�p��Sv�t�DKЈ�}��\����H�e���R+�n4�cp}��&�_��D�B��W��6��L���Jf�M�	B����(�j0�t_8�N�u���a�i�,�f~X�������U�R��n����t��r����;R�2W%WW��(��{pĕ:Ϲ�%���8@,}ø�\��S�c�p��R�t����a��˄0��M�IY�]�o߮�yÐ��1�T�ӗfܟ1Ԇ�N�;��:��k��v��� ~���.�]��e G�����G��l3����+��5�l8x������1�=e��/���S�[q��O��V�CM�`�hA2��U���F�:��^��wY8���2Y����ቇ���tE?��UT��Ʒf@���q�M
H�A����UK�b(��΅�����j�I�b1 p -W�\�C�N�2��*���HH�>y���%2<��	Xl�.�h��$I?�r����{O�� ~�w�7.%:ա�l�Ae�x�Y@���f��É��kU��H*b7��4Hmf��䈵S&�j���g��oܞH��Ep�Yg[��EJ
���͢�x�e�QQ����	L%jY�Ӎ9~� ����2~��Pz-7���Cq�<�������{���\zD�L�C�5�(E��-���/��'I*�&ĺ��/Ew���zN�qe��b�2��'6�A����Q)X��u�"<F�e���K_ߒab�_|]����d�E��m�2Z����-��P=�}���U5�j���K)}'��z]6|OЂWj��RN�A1�H�6f�%�z���D�\s@��*;_l&s)o2 �ٟy�ł�&���4@/��,�s�^�;<��O _i��~w�-
�բ�C(:�]?�Ѥ�����h���uJ�>���p�._BS:(�^���24}��9�=fq�1�H85yz3آB��(I$|�<*�i�'�JU2��(,�}��<-:=�}vߢ1��G2r����%�p5�H�K�My�ގ��Ud��"�hO��3��rh!��dǡ4�����b:
��6j5�N��&�����ٽ��f���Nu���yv�ӷ�W,y ��D���v_��I�>��־�����X��,Va>4�H�+)����r�Xsoq�MD���r�)��$���[�
$��"�I���v*8$姲]���Q~��t�I"@FS6�k����Vx%��gG��� ����GG$Lg@dΜn���6�����kA-Y��U�Z����0�y>�(e�:F�U4���+��?��-�kdF�A4���8�uH�B��J������X�b�uA��I}ja/P\&tN�1��tIx�.o�_��T�Y�M�ǃ���W����~;��n/#���/k\�U�.+������p8\X���C3c�œ�ξ���>��p�l�,��D�-7`I��twsw��R����q'.*�=��J�v���y��`������
�L{�����'Q��Ԇ���p��u��JN�Lb��C��(>	��$У=� �e/�Di� �� uW��Yc� "y��@ð�����!�L5��(���p�������}s�JmCj��W�Y�����&�pFy�s?�q�L��<��B-�.�wz��GW,���	�`Ǉ�n��l�wT�o�~*�z'l���*6���Z�m�nS���P�J)zH *��)X�	���p�Q�1`�9KI׉nlٮ#�НF�
Mn�aFS�����*t�����������I�Cb�:a�2�bs`����<�j���*�ڜ��Љ����uq�S�~Ը�R��9���H�W'���G�߱�e�"rű+��/W��I�~"T��Y`��e�.�+7!p��͘uZN�z�y�/��~�s��*��o�����������m��q<̾G��T�.�c|2(����?ףЗ7H1�0F5Ǵ����iB�Я���
�#��1K���Ҝ��ޱ$�X/OX��m2�7��Gj���P�!2���'o�"�r}�/1�f�ؓ+�f�������N�'7��dLYv}��#:�6��8�~�MLΈ+8�\�q<P���̞����_LS-G�Ю���#?bE�q~B���X@��L�0�C��C�>W��csXWI��UŽ,+"�$��v-V�E��!���Qה+�pF����F�>5�&�@3!�{R?��}L�5�K������m��js�N ����ȉ_O�YB)͂b��x��f/I����
ݎ ����^W���Ry����
���!es���7ŦywG���?F�KCdQ�����(�ΦY] (��eI �㵮�!x��Ƶ�=�0�v7�,�v��C?�u[� N&�C7Od��a�(���Q����K�zeD�8�DOPElaNF��[&O���j���<�^�XP2�u�	�S��18��l�GC�\O�G�k2���^p���Dz�k7}���m��{i�o�) �Q<7��`�Vf�
;��"a�&�|!�Ֆ�`/1����g{��_e��9CLR�Qq�(_��cu��m�2/����%��|.�Lo��Sq�E�Oܡh�r�ϼ-u�ݔo���g�ba�����N���UU����N�D�?�/�K��s�w�׀)�f���y�z
��-�&��>�����r�R#gn��I�����!��o��tp���n���c'���`Mqp�&-	���s|q�{
��tR<2	%R�b�UȖ��빺��Qx4��:��Qz$���7q?�
�j�&����*�E�jD}�j�0c�����ܫW3-�����2��jH�J��5a�
4e�R&��=�I2����,��c��9��(�M;MͲѕ�	/"��"%]�	D�=)*���)��N"c��r�����Ko��H(�b��my��e�s���%eA��3m�9)�j	�tLAa9��2�pւ�aK��K��K��籏�1�IM�^�,Nj'>>����'���Zk{���~��T��)3���X���-�Ϥ�k�����f�XBL���G<�Qkሢ0Xkr��$�,qzۤM����0]���(��`���w�|,��W%��I;w�%N��X�ℇ��,�����80*�K�59����`��� �Av�6�̧K	L�+ɪ�׎ڟ.�*�x�(�9?��e(7ǃ'�7����_VO�0����V�^�)H�܍V#yy��!SPyg�J��,毬��m1�-qQ`(��|�;k3ĉ�����M3�c1<o�t�'��L��u��'ҶB5_�AY�=9�>��?$7cv��Q��*�7G���$�9���-�3S��ᙻ;��ݍ����_$�����o�pE��7Kg7$X�X�~%��BR=���Et1N��P�A���!��E7J�ݭpi!�+ݿ����[���tk�m:�
_��t�;R�s>���0�d��ZE��Dv�����;�����d�o5}8S_�*�6���Y�&T\G�E��g��"=Ŏ�}d5$;Ʈ�DH����<s'��,Dz�Φ�N�w�!���<@�yFە��{�'Fq��Z�)�%B5rj��7�Me�)ͧ����)q�����n�����L��IEҺW)D�ц����4N��c��&������28�M(:���`�HP��+R�v�ѷRe �i�!s4�v~!u I�9h`���Z8\ot&���`�nk�}�D1sk�Chi/(ʍP]�L��o� fE�T�E��'���ZkT�)HW���^������p(�j�b����C����Q�9 �	.���dO���3��u�z��)����{��:\��V�����v�+*�3����;eaM�Af�$D���4)��ju5����u�9��L@�Y�6��^��WTg'N�=I��_r����/K�!�{�65���)�T�N�/J-,��R�U]^�[�QŜSAA��9�k��P�Ǐ��n/%��zw�iz���|z}����]-	t�*R���l41 �I�tWj?s�A� ?C�ލr�C�{X��?�C�������R)�gΤ�����M}-�>�b(c���w�9~� �≡��v��U�[l��4;���sY���&̓�?�|� N�=k��a䫹XpM�����.� :i��=Kri�����C�Ƣ|�?n�5_�F����M?M�>Ї�#���$�>/��<
��H�?�N] � �(dƣ�yu�-���:}Q���\�������V�$\#u�vD�HH	�<�!�xi�.Ŧ$�E.�Lt�
'��]�-p����H66���Ǜ_��0�@�i<��uTZ��;,]�m:mv�h�s��1���`1��J�ͱ )G��b��I�nc���Ze�kb����w[�;گ/�8hT*ߺ?�A}6m�����5o���]��2O؊�Q�˖�@�J�Sy}>b.4=,��^�}*)֯�T>�T�d������1��u��5�T�X��X$}^Ⱦ<�s�T�Al�vu��w�n5�D��g�Bq>Vܬ�����^4�ie�,�f��]�� BsRZ/=Դ\J��a�vz���5(��S�F�xa��{�m%�a�wW}Q�������!`J���m��o��60�R:����.d�PC�&;��o,^'^�Ѥ��I!ܚPtD���)�Z�+���Ϋ��T?�u#����g�K2��0V�w3�r�l*xc3�_�Jp�	쁕Պ
����tF����:C���VK}�F�����>�<����$�Q�6�.�"J�dH|�O���@��� FêH���$|]Ym[���$�ȣ��W:�s�{ܽO�����m�a{@{=k�;%�{<��x���Kw�|�&x�E'�����hQH�����p`�V�mp�O7��-u蠾k�F���-��]�Ơ<�� ���S�E�&����܂f]�����9��!���:��� �F���0ŃB͈��Jĩ�L3[��:m�$��/z�ә/�9�i+O�;�����������5��`4������ ><޻,)�k�Y`!�����`�g2���P;��.�\?F��k��R�19�z��9���-�sQ	�	�|\�UQ�1�l/ � ϟ�}�s8|�3�F�6��z��$���;��WdA�6�7�<]o��dj/ݍ���Â�R��bB��%��2�TIo�;��{^>׬j����^	��C�S������&������M߯�v�s!덨��
-_/p �������mt�-+E�� p6���(-���W0�n.ǜ�P�c��2�<����ܣ�ꈪXBq��鞵7;��Ms�v�fK�zi�Ϥвg�>�cF�6�8�)H���8��ǉ�h0���B�:C�*ABe�Cώ�烜A����>����Vl��F�iQ$�~=z@�lb�����jU���K�Ht.��n�oK�ޒm�~7y�1;�
�����s��y���΍�\�ee��i<V��H1��E/	��ׇ�z	}���Qʝ2:�y������ǳB#ea�J���תB��+����fT*�k��o�о'x��<c�(g�Kx�ېX�O�ݝYt˼�tX��T�27�-��9�g2d���������%�)�o����q�?5ݫ�+,<�+l I�No�T�<�pz��S"�]�>]��N_z��}$ tz�H��d���mU���}Y����o��y�ƽ/b?�&|$�!Z�}=�}"��,���N.�0Da/���tL+��"i�g"Ȋb�L���x-@Z�O����#P�n	T����\3~D��-��	�?S�����U3-�K�Շ��T�S�U�]Fʶ���0�<w-Sn?��������Y��7�M�!M�%�,�5FVc�U(�jVh�?�=�/C5��޶)w�ɺݿQ��\c�O�6͜��6k��E}�� ��%Qݺ#R��Id ��܁C�H,=�ڻSC���sn&L��JpLh�Vz&�̕TL\�.����D@��C��!���H�m��R���ϸ�#��3z���D�,O1�eɡ�Q�~�^b����c!B�P�=>��JV�bdpń+[�f���BNK! ����"L�}8�S�X�L�$����4-@R޻w�ﶖC���h�ԃ����1{o�B&;WZ���+�:Lb���4���a������(28�L����%����.N�El�1�<�#(t+�hTW���XF��1�Y���L�=GF5eE�$b�=�"�1UBYQ��X�r�i��+uO��]��2�.P�'}
���KaQ�	��k	[p�~G�'S^�(\�Za?~ǚ�j5�,�w��sD!E��E�U��j�
O���M] "��-8*i����ChY����!�u�
��V͠�g�Ѕ�O�����h��l\��QWk��Q6D���+�RÊ����lJ��en�Ȕ��a��HJ6�൫��3��W�%Yf�Z�Ф�4���u���<��x��_��d��Rzg�Y5S0�%6��~� �b�Q�J�4��2L�5h��j�1�B���:|v��T��~�+M��%�s�_G> Q���Zl��7���η1[G�s}�� !�����P�f;��#��Go��˻ޅ!�NKU��ОO\� G}b!�9�MgVs��Ի��	���3u���^~V���L��f��Vw0~[����������!�S����@*�g�)3]��*�Y�M/ף��R��B�i��@!�P�I�/{f�'O�0����EQQJ��Ui�i��s��v%ks3���䤐��MĢ4x8ķ��
*��"��RB�}���(舂?	Z�����(�����,�_җ ���)g��	�d�y"W?�TM��>.YC�d���cV ���R��1��G4ׇa	�w'̩9oE�f�Y�)�qF�����an�8���Q廪�S��kb��c�l��M�]He�J+m�#nb|ڡ�H�7�t�Z���h""9�Sc�#84m	���q��0Y�tM`y~��̴ϧdʞ�\U�����K����%��S~x�� b��M��k���v�Z�<��KHg.����L�Q����Ճ�*�8�P;�®�����Z#�S��˴дp|u�P��<Wy�Tlُ�c�s $�7wLaw�9�ѧ�MR���'���[~��<c[`�����2�jO��WH�cdz2��o� �G�����ټe��r)�O�_��v�0|S3r�4ئ����Nb�ǂ���X����	e�ƻ���36��z^`�~%�m��}e�i���s9�_9�������z��2�������r�H�W|{Q�$�x�cȨ��m�H-����@C��ܭ��~.��k����]� ��B���-:1:H�1SF:/y����%9����`��0a9V�&�� M�������zv�Z�2��Rw�@mL��m�aLu�� �W��@\
��ڮ��%��bm��AU2��.��2n��Z'��IGO�:IG���H�jY�3�zp�t��y���Rk������}ܗM-�;^|3����`�p`��j�3z��i�������2b�^T��O��L8	��q؊��8߶��}[v��F!�HrK�c�mf��F�y ��N s� �u�$��gN����v��a�d�)Q���0Ǔ�#�m>�Ҝ����k���ibq���a ���̫ml%��u&���|WЇ{%ԓC\��X1
��W�~���w�p'�uP�<�jT�j�EP�R�MNh6m&L �Ar��g� �4�L���ݺ�����nK^`aȧ55�ؤ`"���[ U��_P���pe6^O��kЋr|%��o���n�\��o�+M���~e���2TW�
2`xz�^ ��ּI�\���)7'=�׭0���K�:g�o���n�`�vb�Q��g��p*�c�fӜki���gQ�bi2�i/�lI�Jhr�4��rSWx��h#5��2?�����+T;�F������q�P6B%�(�������ȹ{��]1��p��<�蛳$�f�k���I���Y�vE6�2��%R�K�!'������Y�ef�a�@v9��k�[��7�K�d��SY���y��)8�N��#>㇯���𫼶"G�n�Lp��c/��Rή����K8n�=ꁯ�jp$�-s�^���ĩ��ؚs���$?gT�b���m.��#LE�9F;	33�ˢ�P��+��z�*�ը�p�efǄ3��-RQ���&�ni����a�<^�5����U,
I������W�ZꤿJ���
�h]{�����_���U}�W��_>��!����A�u%��S!W��������Ͽ������7P1 �kQ�+���Ȯ��$��Q�˫ҭR>�foF���n�a6��^x��4m~�jߓXvĢ�5����-�#V���̍	Z(��<A��95�8\��G�����P낕���-N��|WA�y0IE1��."u?=�ZO�y��e�r�ݖ�k��uG�����ͦ�ojȐ���S�z�ޭ���&��![�z�c�0�-���e��ς[0��}�`�׋3�O�dϾX�`�V���A������ut�9��l����Qus�TWq�-U���[�0�&̹�t*5�G�u��x__u Ur
�<eZR��b/����u�'Fb�my�Y�?�b� �昚��eP!��`P�z��n�U}��fi&�w�ԡ�~�xnK}�4?&�mP��@R1��kB5����t��K�m�w��,"&+(��w�� �@�J��:q��,�D�4K5��tU{V �h*��֔H1 �m#��� �;����D�Ьg8<�J�&.$�:&�-��7�y��bVמ9��e�cc.<��\\�!
m֑���р�^OY��>��z���m�ǡn��R,����$��
��4�j#����BB���K �H;���x��N��&���Hy'\ųD�EKV�	��[A�q�е��d�
�ӑ�`+�Nr���%��c����g���x7q�8����M�	7À����Uȵ��1�U��}��8V��$N�}��6L�5k��w��lv���=(R<T����
�V%�;^¯n#FK��׽@���R� �ܘ�ȟ��Z�/�ܡ�R�v��
���vp��E�H�*��ۑiS�r^���V7(��}�i��h���Qk6H��MsͲ������]�^�����27�,j���i��T{=]���Kj���.%�v�Ɖ��5�i�$��f�!rI)�<W��2�E9KG�&�+�>}��S������-vGvG�Y�x��a�u�OְQ�_�"��G����Ĝ���f0�9A���YN��ׁ ѤؐkMS���&0eyQǱao}/�ϸ�5~ܗ3��FL �Ƥ���ywM]<��!q=���gqNB�]�1�|qJE)zç�i���C�}�f�R{ydZ~��b*��q�[A|)���#2�u��̸�jj�F�ED��z��0��+:6�Hӕ;���d����Ha���C�Fgs���]HLsd�G���TT(D��"$)fӻ�|�%"C�:U�s��5}	.�>�R1�ؓq
�cz��^ҟsѱ��%h�"1�sw�<�8
Nݨ)��0Ym��ϥ���5�N%��z_6����[;����۪��e���r	�"z�.{5�ҭBR��*���v�f��݄vG}��p����a�3&����.oQ�Y#�E������Q��/ab]�����h~;��R���\��Y5�z���	,��s�{�f�G�J��w�_�b��~�~�����[j��)x��+�H��Y�g���O㊂�ڙ�F��UŴ���9b�����MsH7{�8��/}ʼ�_���i�"п�q�7--���o��8Q�A��i��� �|�f�����#̱����LB='F�z��Քx���Pgj����A�]��R��@5����%��q�K@1�2A>��ՓLh�63ԁ���ϊ�)2�^������h���yɸʗ��T]����_ނ}Ǧ3U����7�W?F��xY^�S�Y���K `���cr�'X�N�Jx�*Cy�(�tz�,2@	�i�ٹaǜ<'�z3?l�;�w�����'.Ez�����^��'Ƴ��H�k_���P^*�/}�Rsc�� 1鑥 oi�E�9Jb
�_�/X6��ttT�"�%`�<��l	줃Ѽ=B=�|$��y��懐��P0g*���Ϸu_	����u1
"���;�����a��w{���/����"ˮM�axZ.����P�Olb[@�VL��^ù=�:9P��"Tq�;έ�� <��p�l+@��z"�� NH���5飱APX{�*�Ӝ4��n��m]AӜF:K<�/?O���Q&���������JD�`XW5ד}�v��.�o��Cxtȿί;�\��-�c;i�lY�?.�X������#���hU-�߉җY᷆&:2�JgQ��j���s�_��e3E�=�!��96���������J>��~�3��?�d�f����Q�S���j n��~�Ǡ�i� �0��Y!��<* �[�	��]Qf�潩.%�O����sQ�	�M�H~�hK�>t��ý�fhajmv����C6�֓� ����"���-��a���/[�FB:#K�%��ˣ�t���E���
ȸ���L�]>��o��6��F��.����`�Y�ֆ�)��{��0��Mn�`{�x���3�o�,�[@Uc��4��goVT��$��h���� �EzƔ�g��#d���"��`S�1L;�5��T���3�T*2��G	R�p��[j�};����n��$�2Q��+�1ژ��	�Rz��<�Oh�k<p��k����3/���l���/m[��%��ɲ��Xo�AM�����~�!MO���3B�[
M��f����β�r���Q��Z(z3��o�h����y��Z-�Qt�X-I�r��we�_�O�1�����f8aa�CW�{�tZ`I!�ւ39����=��O?99�ƫ��P���kBjG	� m�mk�8��#1�1�:A�yh��ږ�o^���&�z?�(D}[r��WV��J��^�m���GK����u �����&���oS��+�z�9PSj1�-�|p�4�6b���<nN�q%�zQ��C���I�O����U�,U�"������.���Јl��'�m�q!��~��׏'�Ŏ��fC�	�P�7����)� -�X����\���;w��x:rѪlB�	6(Y�:&��������b�Y��+�ڒ�;g�YQ��]��>G^�����n�W�e��wA,	ßg%���,}�|@�(*���5K��%	i3�vg.�I�dY�fd�#X)���� y��kџ݉+blti�XD�>�Vj���;Ԑ}������X�K<`�W$»��ִ�{5�K��W5MR��%��j��Et6ɲ��:a�����_�G�vBZNnxRy�èXK�X�4�1���թȧP�������������)�.����T�h�,c���̈�j�l���K�N:њx���h.T�����EڕC��,MBO��,�p�k!�-�斞�::ҿ@M�p��Ơ5�ó6�]�2���-��#�V�U�쑍�ҵ��&M�ܸjt�E��A�����BB׿~�b^m��,_tƀ����WA�7z��Ԑ�CRJ��l<I!�P�}�W����!S���ڇ��oI�]tʊ:��"�&���)~�y�ح�8�-;����H��0l���	��۵Ӱ�&��i���r�$�ȴ%١S���p�C^��n<�9��Ϻ4rE�/�bC>%J�:
1��H�(]1F�R(7xT.��6��emj���lR�U���2rP�xK�*��a|.036�S��
��=f�Pܢ��i��>��4���`s�8k��5(b�`�w;�!�$#�z����'�[,��}��c����^��y���<n[����aA~b�l����O}Kl��M�<1	�Þ��2���
+�\�Ɲ�u�v\$|{�4Ԅ�w�����AiƳ�ތ$Ë3!T�զ�y����U^H��KZ$ۈ�y���<Hz���k�P݀Js_��Y�ԶbZO0aa*i@���_�<��$��*�0V���yM�z����A�^���؎�]P�?ߣ)�X�	7ϑ��,��E��۟H��iݕK3����K��?s��(���ue�� ���;�Y���/>��K=	�'��C�?��#t;ԒW��bLз�W6*�1\�C!P��P�4n�y�nO��j�)��.ְ`�&�ּ!Va{V��:@0�?����\s6?m���Aʇ=����Hc�c��k���hܡu��v�v�	�# 8��˖�����0a'æ1���1�I1-rRm3��s���1>�@��7;�m����K�&~},��	$�l���F|�����l�I*~����X�l��.��i���=-rE�&Ks�ұ�P+���ȯjZ��	'po���,&YjJ��wqa*���wk��Չ~7���+p�[��:^�I���I�b�x�?�Rn���~��z�[Zυ륫f$dwC�t�&
���X���6sV�:l�na�W��<2R$�P�����8����&�����;?s��2ho@S��*CȮ���U���G��l��9�	��=����$pw����z)0�_��)4�D����(��6�#H���d ��Ҕ��Tk��Ų>��?fF5u�i,���RuMa���m�����L*��H�$y$f���x&��'��6����5����х��$�mk�@���pµ��BN���ǩ��\�~�*p�o�y�����>u"5B�C^�'��ϻ��$����)iT̬+���3�e�H�o
����|����a��L�F-���������WY������OM*�h�RC^y�}S\���ڂm�6S�W=�5҇*M��{�cFYɣ\����.�H���0�ց���c��ʁأ�Ƽ'���<+J�e�C[c�-qO�"��lk�;�׊�7������Ž��D��=�x�4��a-c����p�h4vՐ���О��=��T+#�� ��I:=y,s����u����g�݄��~�L�Abp�w4?Bi�����*p\��<��N�󟄔WP��k��ֽH٥���3�ӡ1�)ykrA�����{g���^�z"tC�8U�7i�t�!e��%?E��ǩx����.G�P3�+X`��i���	#�K� ��P]��wܢ�"B����M*$bRM&/�r�T���V�����f�B�����6�11c/y7yĠ�2�
ap�]�k��E���a.�g���la�	I�$�Ft�b;�s��ؑ,�)�Kf��)����ᯛl�.�Cp�_s�������fj@�\7*��R�3�S�Js��0��Vi��2�:�t%uX�����d��������}~HYo$u�SP�`=�ji�v(�?�U�,o�]2�b�;�:uEO���s ����Fz���KO�<��G�暟.�J����nў��+�Խff�mb׹�=jK��2���G���j���އ\��Ƕ_�A3��$Ǘr�-`��=���ѧ`5i�>%5��6C�MM��T�6�ij�Ř�_�2~vz,�E�I\�J�o��϶�{�R<�E;��`�R"�ڞ�pI3��e^�%7Z79��RD���eT6�I���TVg£���cz'��g�B���A�OҘh��Vd1��1��{W�^*�]�2+E�S�	I^�>c�Ҵ�W(�~����+�d�g�i����<��9bjH�j��H�˾;������.}J�;����5����b��������b�=�,-Lvx�3izd@�����ԧ.[1B��^�W�[�mC)C��߾u�;@�L�N,��K��3�٧%Q�_·��pW�z�6��D���8�I&�1h|��&kA;�#K���!q��������Yw�eY�D&�X��#�||CT��ѴI��m�F
c���q���`��:|�2�ѼGK�O��x.���� �n��BQ�m�3�� ����'�'��g�JM�e�LjO�qY��A+=Q4��&�R~���kg��<֤;����,2��#�\_�T'!ХDpץDU[3�;�_bX��>fH 1$n�]~� �z�������8�x�DIp��Ϭ*�*�Fw�|���Hg�zr~��R��w����R�`<�.�'FU|�F<���aq��h׋�G�3��4�)�&0�:0��y�v�ŏ��0gk�b	����`9�(�A+n�qw��6���8�>T�o*�"W������[.+ir�veB�ʓ�c�/�Zº3Q����������#$<�l���2]����J,����1��r�O�0�dU�"ӄ��I�nή��+��4K*�!�Y%�+=ä�0ѝ��������Յ�o-�2R���;��q	����H� [=���"�=t��e><�~�wM�B�C��#.���)4�!��4��^���n�#&�d���؅A�7��_��Y�B� tHg.�H�2k�<���ք�fB���EG�B2;.�镭���'3{(�[�N�����H�p�����$�a篜|FvpZ��>G�E�l{`�$ �xII4:��|�_��E<@�5k�\!2Ԧ4V���=LNX���r�g�W�'�v���g{���W9�����J@N�ܰ��vJ��|{��8���n0j*n)��J��	\M�����K�hZ�_ܷ�!۪	J|j6�&|P�ڳ�_о���7sp�����cɀ=Z'T��$7�n/��YK6��qFdBZ���L����n@��bRq��u��Y�y�0?�I"�`C�ȁ�)WN�w$�vJ�b�Tc;KU� ����B�S���4����5N}>���K�&���p�L�Q?�V�.O��o��"h@V3n{��d9�KG��8XQ`+��=y0֞w	�noG�o��_{-�Ͼ����H
�Zg��pZh�[HU�.F\ɣ{���&!+��0�pKkt���j�j��BF��C��w(�h�ܣneM�SO��>闥ْ�S�Ź?XV��9'�bF�1��[�76)$�*5�-�8�B4�`��"+\Ҡݔ�O"��u ��PU�I]�YJ�n�k6�̆dc���̔�~�Q�>Ԩ�%#��' ��'z�)��R���m�\�j��,��3dH�MnH1����	����f�K�1�@�s�O��P ����Wղ2�j��|�K��EH����SP{h~���H� ����VW<�g\5�'^�֪�Dcܛ]
|���u�I^���h�48�֖V�l�1��S�<�Ȅ j�֊�͙Ϟ���S3׮���VsyٯFg)��q�%�'\�tj謴M�oيZ&:���KB���vSN��v��|���cú?��%�p|�4�Z��/¸�4OC��
��/�b뜈��@�	�el�*J�=��iNue�.P9in8\�#du�%O�����$�y��ǁ3в� ������sv�o	am�w���O���9$57�跭��1$��o

z�Z_�&��i� ��$�'2k�����'�`쵈�=�����OO;.3�����TZ���r������V�I��(�M��f��BR/K;'	�f/>kD��R�w�18� �Li��x��2�E��j����)�/Z��{��Æ>`Se?W��ET5vYH�e�5�G:�K;BYU�.������c�/ؓ(�&�P��ͭ�蜤��֓��(6?���i�̖����b0��*��y��,8����b!� f�x]������l>t �o�,и�P^��uߒ�nXr�`pq�8j��B�����r+����Q��@����� ' ��>!B�mtcU2�?��h��<��2��>�C�7?yLw>@"r�hs�J��E�1dh#�$]��B)��D�%׫�Qpj|q���0����x?^�����n���K:��C��8Ae�m�;���e�"�x>����G�Lg*�:X��rX<
T���p���\�Ɏ�|#bj>�zc>Ir�u�g�
z�B|�D@��d�u�c�����cGW�;w����ch�t2Y�sG:l:Z@U .��5���H�?�#���|���C�z�x�\f��OmV��a�d��So00�5����Ny�-�8��]+��:���Ҕ �z�wH%C��2x\p���#��j`�q��8ŪHlgo��ҎU�@�U�:$U�O�B8a�Y$G��X���]�-p�Wz�GQ=)�6�Nȕ�7#�T]n%��'?V�:1Km�-m|{���-�9Cb6�����5��ԋ�Lŏc˕�o��!�9:�8��X8mM*_��������i�g8g4��t�3���~�w��d�5ėG`�}�"����`�s�c� ���D�j�{U���7����Ls����E�������	*�&_�C]M_���eLB�)��X��J'b'/��[0����6;�()≃��U��]��Mp��6׏�t����N��!��æ�� 0>�%�'�n����K�yP_i��NQ:l�z�V֦1�:�_�d;����'�ȭ=��d�k|��k��������	��l����̷��S��^�0z����^����&K�|'�G�)�Y /CL5��t��Ox�'��4@�)�w�\%�6��{.C�����Ш����rɬ(j��_�d���F�nKfID�D�~����8Cr�#QpI���:�´(��=O��A��޵qH�3���r+N�q���k'�Z�J"D�� ~�+͎�N|$��lt��֬2��1���]Í�-�W�6��L~�M��j�>2�G����1�����I�Ep69ڬ�2�Ot�%�v" sgy��.wܨt]�����>68�S�
K;�p�0Qy��Zzc���sT}c�%��/"���Bϲ2g0k�q�>�r�j5�H�0��t@��>XMA\����+�W-S�j�|�����m!W�kK���ș�����]��.�5�|����Vqn�P��A��Ҝ����7*�Ͼ���1�)�0�716�|��n�g{�" �5VT�z���lTp�����?�#h+�Xt\��U���d�)��=&.Lg	3-�<�)�3����o�1��pĠ1ɮ�yGS�&$m�-~ई�c�O%��K�~U��L3a"UK7�ͥJ0��.���K�{*%"�i�ZP3�ˮ�ûsHlפ~�y��3�3�T�N�|���o4/��j����F��ɪ�8j�=I�k�i��^���k�#��e���ld�{�p��0\Xю�` �u���V��G��\-�����Y7��J;j�kDBhc��ϙ/��=�J 5�F�^���=5���{Tmz��K6SN�\�n�?���ٺ�RhH�H�>�*�8`e��Yx��df� ���[�B7�Um'� *�!��g��E�Á+~��W[ܷY�$*�hȻ���E�^A���9��!�>��/8�C7��˰n��X��bs1�Kk�*;���-�J�Йf]T���l������Y�9a�JUK�/z����<����LP������<Y] ��Sa3[1a�Y�W~�u5�گ�6�36 F'��+=ܖ�E;�����\�?���UŹt&I|��v�_���[H��<�h_ X;SV+i>Q�I�{��`Y����/t��-P)�9}������j�p��*r8���u0�R�t$O~�̽� ��\�zg,�ۗ��ָ�5��"�oH�$=Xv�����E�'��w�u1]%~�����[/�>��V'e"V����Ĵ�a����ǉ\Jy���Ԓ$�h�A��~t�ǜ]��uC�ԕ�;P�'�b��n�X���\� ����_�#Y3�2����d�J�$�wxt�l�p��0�Q0V�Y��U!:���ƱV%����hr7*�I�=���\�G�J:V�?���;iS�#�_�jM��w�[������?��븤���`�6 �kor��s���3�U������+�L��@�����j�8W,���D���ҿ��̊RP��d�����[q�����}��(�X�ϛ�~Q�iv���!�E��c�fi)��sޑY MV�*l�/�p�[�aoi1X�-��G,Ze�6+y]-�-��Ʌ���Z�c�@5�(��J:��A
��V����U�Sr��.��o�Ϲ���c��l����>�XL�K��$�cCK�+my�d��_�Nձ�f����b�����R�ˏ�G����.�?,,��_��zNh7�p�o���nw���H�p-���P#D�/�I�����N�p�K�l;c�{'�8�LWlK@���/��	X��'�.��-Y޼iH!��2�ʺУ�.w~ۣ�n� ��$ٵ�D���s�=�b!ge� -��*�>q��/S��Z�������Y>�8�E4F�'#o���l��mb.����\L�h	ԚRV}����Wb�ɚ�:��m�a���^���>���i��n��h݊� �t�skj��E\�;��f�,������� ߠ0�řM`)$E��r��
E�E[�`�%��ˑ���}r���On���}�llo���Я���L^�G��bcUVͺ	:>A�I`��v���=\Ww����V�4�0�-�a��׸ު�;��E�S�>��NDsY{d����7���
Ȉ|Hllk��g H�����u��i�6">�K�D9�P����}_0;7�Z�|q����A�y��"�|�P�H��#�qqm������<������j"��!�٬�Dϑ~�+� ٚ\�2��A�#����Z�2=��N,x��u�9gYE�,�Y�K9��R����(P���)��eK�}.G�QCz��3���(jfj��d�|�W��<������i���s׬F�N�FK�%��Z�"�g<�Y�E{Ѕc�a���3a҈(��� wv��Q���zT+�5뿟9]X�]�o䧀��pS.���Q��#�
���G3e���e�"H
��L��� �c��K�Hv�?`�����D�����$���n ��F���\��B
`��kH�����rG��4���o_ih�Go[��h����Z��C\V�3h��1���ڛ����05�c �a�
H�]�O\��X`���f��چ�v��*��ӏ�j�r%��u¥��P,Ӣǥ��𢵾$�fG�"�'@c��ٝ��!P^�j�/*�D-e�H�������e1�V}!
�n�w|m���ogĢlC�w�G��"�H�t�3�4�q��v#3�����8͠������0����M�EO��C�[<��ƈ�i@K���0��٣d*4�=�9n��v��8����'���:k��Ǉ� ��4\�IyT��M��8������iE�Y�Q-7
�굮�OO�8򝋞u���dStG��!P�q�#��g�,�v��5R�ȣ��	Jt�t�)��쨢"�}�.�)ba�fI���li�2�(�;���	q]�i��A�TL�QD �5�נ#�_ػ��jne�p����>�� �9<֬1A(|�P�> ���-&q��<�u�ԩ�ȷ�j��4w}����[P0��M�ب��E��ϿP̛س�܈�����?�
t�h�=w[|urH_���]ةޔ��U��;����ㅠ	B.���t�Rͳg�r�3(�O:�����n��vQ�S��즏~�4ܩ�%'�Z�l�{�[��1%W��n��FÜ�yeY�f7Y��?5���Z��pb�}���,ɯI������X��ƉJŲ#B�>^���2%U+PqB�D8�%�R)���NĘv!����n/R�\bNl]{H(�ec�y��uG�,3�<���;�E'38£��%��c��;��)�Ӈ����u��#qS� 2��%�<�������FͼҌ�	5�p��F�'VDʱ {#ȡ F��l�lN��~�Z��>} ``=�A�H�����m@��IR��t�f��}�k)��V�Ŗ�6{�q���k%A?�Mۺ@
Κ��iY|�!�*�wUd:J��Q/.��:i�;����^C�2iASl��)���3�	3�-�b�Qh���1�����2`;���W�p�.�i������i�#(9$�N�t���i7R�S5Jn��ͪi'r>�6��;�в��Y�y��˥l��e�U�7oV.i�2������u�xG[3�O�1�1�ȅ�r5?oB���(��L�go.�v��3�H��ʎQF^U@��Dq	V��8U��m�k�S�]���\�|���u<V�P*�5���A���͡���iu8
����s���$�<d1�)Kƍ,�H2T�,�����I�k�1���"���32�6���f�����dp��J,^:ڙ�Aa�[ef |��y%'ĸQ���1ԯ�~afM�찘��%^Ba.�d��g�����oMW���B��G��Ǖ��رtg߼�x�}O���!]��zoWY�`e��H�by#7�R����J�C�)t�U�{AG��ˎc�C{U�OT�.Ã�L[�0-��g��Vxqo��Jɝ�o�U�N�n�q��ܓ������FxD�Gz���M��ey��;V6���C�_�L���[.��ެ��d��*H��Y��ÕJS�[|	��4ߗO�f�6��|���va��,Wb����)H<�?)	j��D��&q{~�Ƕ-QB�����T�Z]�$h�c��O3�v*Y�^��Ǯ%Ks���tk�Fh;�D�k�%O)�H��e��	����$$4�)7����与�)M��v����Č(wO}����4f������4���yl�9�D>v��	�/2��3.�r(�兵�ʗ���#�����,�_�����(���dz��$��-�'b?Dt����#��j;Zf|�|E���|Bkh<��ʥ�'����'�Pev��rs_ww���$ީ�_	���!�f���p��wN˙ZE�6���M�Zx|Rx� ��+:�7�K�c ��i����ԙ�����`�\��[_����Oy]�3�A!k�J��_��G�Ag�CYnϖ}�-��V�Ed�AO����\m�� n��(����CPyy�S.,>#LW/�&�`}���]�ʤ���� 3̭�"2����p:`h�,_ؔÀ��9�Q�(��:)�3�K�g�������
ֿ����A�;O�n�)/�f�JZ��Vz�m�u�@�mv� qРɳ�-n�sd�������Z2��E*i�M����H�y����鳗����AS��M�+%��vp�+@g�l՝e�]�۟^b�1�I���f����d�g$b�q'��Q��
�x*i�.����a�u���%^O=S��#H6e"1�ڄ~���=Z*���r�����dt6X!�_4�P�jDץH�(�2�G�q����a�'K�vl(���9�f�ɀ��aM)�9%�������j��,�7��m����Q�Kce��S�SC/Y�|�1|��N�z�og���L~�}�Ш[sp�r�11���
�3��6�����ao�A����x~#�-к9"�;�:�;����0�k�<U�*5�%�cd�����m�O�%^�<��y���4m�5t��]yRƔ�uC]��dM��	A��M�^$�Xx�:���tv^�l/;p�g�:9]į0E�@�6�~�n2�]�}�t�����ob�����?��Bf�Q�Αfä3^����k���rTl��
�D)= ���: ��5������mܿ_2p��IW駨܆���J���o�z�-�GQJ^/ʼPm�.J��d���Z�=�d�L���ֵ����C�dti\�� V�[�\_s[�2��T_$��t:�_P�HMG^=�][��(Y�9H���(�ށ�E��-�94����_XXX6�YS����G�O�sg_��J��P��B�n��bG�$dyy�
�X1���lE�ߠC��<r�d�G�����bAs3�M�Y���PU���<��z��5�~��3_�o�&�{��VL8移�陸E��^+ԏ7y䷙��|jjYr< <`݄ݮ[1��4�)�[_i�vY9X��0��[�<O�B�:�+e����P���9����UViG�����ӢQfd���J9`K'3S�2�τ�>���N�w�ay��8K#:�
��\$~����Ei&c������#t����U��8�	�Q�w0Ŀ����ܷC��.�TD�/:�F��dj0R;(�5�h�u����y����AO�#�Agg詭p#ڙ�Ά'ڴ�b�kU��5�2�pd��~�8�����Ae$!��z�EY��B���GG�S�����I1���@9{�	��G��lc�Ż��%`���Y;���EsK��5�RV+��Uwy˿�u(t>yW�pV6D�lX�O�>n:h�%�z�U��j�O��)h�֦�SRsUt��4���g������ڳ�� ���nsC'(NH�@VcU���W�x*#���Q���F�i���tH��ϲ#n(��	�-�1ʹP�
B�������J�xޏa�u�ۤ�=����g�4�����#�jX�b[p~�\l��P	3�GvA� �͉ �:�݉�+�:I(�)�jg��-��ƪ�e+�m��C�y4&��"�؅�%a���	���Q��Q���ȓ�OG�`�z��u�ۉ�޾�S�H~��&N�."�F���)��7Գ����2]p���%�G��UlD9��f��Э6�f C����Y=�(�+F]]
�^����SR��:ms*�X�^mӃD��'T�M�W4�vٱ����C,��f�;1���P�E2���IE h��z[���Dz��l�l�|^�?�W����sP"���І$�O��&�~�fs�\'�6��5�L���$��pE?��B���:�4�?��0��.�!���7JD�\���C��{��#��u��iw$�q�S.��6�䣛_w[.��X�W��ܽpе1����i�3�G�fJ�]��܇�;��C���05�*\�)���6�pU���ϋ�U��<ŬQ�~'E�K�:#0\��}�/�`�������.=`��Ų�ЬL�Y�+7�э-H
��k��xC�#��ly�&ܓ���(%�p�} vl��ty~����׽�8�!d�s��%$D��`A*뢧�c&��k+-5ǎ���b���/�ۧ��y͂��}� K��S �g�6�qń��6*���Mۏ���'p�!�};%�T���N*v�E�ا=$7\R@#熹���5pJ���iR�Z]6ٔh�����
d2��uTy�!�QZ���K�v��i�r��J���%�.�����[$ⰲo�V�d���he{�*�mH��F������s�7��+�d���J`��'�e���i%���#=Yi����3��q���O�Ŗ_N=���"�X	@$N�C~��\�_�;<Kl�B��w�4T_�m���s�̸���<���G4��&9DPP���ډ�8�&O���q����v����J�lxG7O�$x�_1�%x {���|UZ���	T2�������L��׋�j�&���]�f�����$��=<n�(����h��Q�}�̲ҿX�u�
f����	i��c���e����zBb���2KJ�R��iL�͠��lv Yj.�x`S�I�'��2c���E�k����wv�~�Y�ִ-���=fLN�`�<2N�?�T�{�%꟰
<k�J����Ý�/�a�M͕�2�O�ྴk��J�hU��a��2�J�~t������h�s˜.�6�	ՠT�y�w��ӈ�ZrY=���Բ{��싓FP���t˨�g�#6tN��s���'��`��; _��vJ�i�Й�UKM����_����z�$;�4�h��w����(|,X�p���>�������mt�V�>I򾼤�YO�s���0<[��ۉl�׻�ڴ:����z�}R���K��Ї-?!;}��DO1�!�X���N[��M/4V�n\6U�dC1M9�j�s���cqv[z��]������E|!�b����6�>���d)G)K�ԹEb.�ڑr�輇��<�nz^���\N�D�BA��Lģ�$o�!.<�QJ'
�-�-E�#�'Mi�]��{mD�g�$�&��G$��c;��L����n����)*[yoGV�$W�A��p��3o�(�fbEb$l�^��F̡	�)�J��3��gS7$�I���V5���UQ\�0�-�l��R�.|�K���@�U�d+~���Р���+Jjr`
����g��r��b�����x &cE��&�J��f�;���@q$Bi�R�,! ��݉q�aĺ5�a�K�(���_��5'~�Sn$��-���&P����N��̨�ٙ�d���#u�$�w���n70�|^�Je�p�ZPL� ���<&}�D��3�E���'�5"��>�jyJY�Z������a�Uw��Dۅ��Y3���n\�&�=dK7ϩO�,i6���_��a�7��}=�GԤEb�j��١�1�J�_�(��:\��(-���\.@*��.�N�P�J�j܀����vժ�.�ʣ=����!�!X�)�n�@�����7��A�R^�|�-�b,�CI�U3nƨ���	��3xm#��5��.�0n!/��l!BD�y�~C�
�U��Q����t/hI�R����6�sa�7,ar�xf̎���@���sE��Z#pp��E�*��u� xC��I�<�1�7��{Tӵy��͸æY�O�쪾1X��<#2�7'P\x��PZ��$$�@�Y��cGI�W��޼���d���'b����OC2a�;�!��q����B2SJr���p�M�[��&+c��`h)?�3��C����*vA���Km�����R=̨4f�ο������i��J��>8�{��=b�53sxbQf�\I�;�T�H{҂�ݎ<��K�����J�P^��	��X�k��·C?}{�{@���H�=8��t�k �u����K���i��T���x�N�ϊsU��5z6t w��fy�*��6�s�JA���B�W0�)��c܎k����6�ӂx��`�N�{+�eV�P�[��?�
�C�;���x�g�9�D'n�pN�D�����Eby�s:�O4��ľ��k��d}9�eM �q�%�!yL�hE2��'�� U��11�m��(��^��X�����t�M?��ߍ���\F�	m�̆:���a�*>3�%ׅO�!z��\gn���pF�-�=dԋ���g�f�����؂t���YmO�G��rM��tv��@d������{Y2T`*)Z�<�*tkPG�d?���f����u�4���-��hN���8&Y%��L`>��u7�+��"7��S��w�vokHHh�G��ds�u��|�@&�=� �0��])	M��� B?�d���єCB�:o�����hh��d7� 7���:�7���tasd�����������Bʦ�1�`�F;���5CY��W˴8��k�@�|���Ug�k��SP�A�
����اk��%D~e�ٰF�|��KHi5�U�='u'����j
�H
�[jQ㍬9�'����;�#�S/��,��5=��r�YA@l�0mp�܃�rOGُ�~H	:]C�,��R=��F(�$� ��]Z���dc]�.cʇ^�����!%ou<��2��ۡ��$4�XȟV��L����cS�l����@ϓ��t��'I��A�q�P�A�`����q>V������@�>-�W�`_A|��PK�,Im�$�s/���$m��t;.؛��RE��~��ކZ�����hR+K_K����ޢ Ȣ-�<O*���� �tU#~�� Pk/�3�U �h��O9:���D�Lg��o�f:.�~�ω:�����`,�M��1����O��?:6q6�6��_#��5,�F��S/^ݓ?ȵ�Ŋ�6{�
ū���""�2�5'b<Z{j�x�鋣%r�y}|���~�VX�����/�jѕ�����_����,m��|g��{6��� iv��ʔ�R{��6�~�݂��am��Vk�iK�hj	t -�2�>(��KT0L%olg��i/����pD�����&��v���s���F��9�t��T�l�d�����P�
�JJ�:�y�T�r6L�w�Q؇���K��yc~x-�=�y�"�����?ȫ�^gRˍܭ�?+�ַ�!8[ڏ�_���������'���8�����)Q�az�w_�JI��'�hI��m��z�h���b�t������@�T1~7�_���û��uemL��`7�OX�&�-�u�/��o���"3�ՋO9q�c��iD����[��欰La�4\ W����:�V!�`�ds�Si�Z�xKT���t�v��XVz�z�nP8d��F���Ʉl�j�i'��n�2$���8z��4�G/�ŤC�ʛx���v�꣛���GdY��ΉD�B�ƞ]��IA����,��o,dj�z$�@��׬3�ݷ��А��'�-�'z�a�� ���[[��'����|�呋��qW��l��H����ve�n��"�{�R��Ǌ��7kv9 ���D����d5;B�M$ˎ�u!�k.�(5���,�Pd���繜�P�|��O�kAMr ���$�&X����˼��0�{6�j[s�E[̩r�?�~4Eo�7�t �_KQ�!�]��P�����U�DH�cc�"lp�P��,���&�K1��)YSf���@s���|uw����C:HƼ�k�m�(�=���83s����O�̟��t2(28f!�ޣ�fH���8������%�3�)�6wJp�t��?��M*��@��\�T�'=$�/�xl^8��#b��,6{l�f�ðK�)��v�LP�C��+J�Z贼�#�ۆȟ�݉�h�C�ߏ<|A��v���B����<�w���jm��cg�r�^ńB!�0 ��s���	>�7���P���3��Z��R��H#��3��Q�[:%0y���Q5x���s9���]���y���� �1��i}֦R�CiĨ��L&�bJYL�D*M�{j�dmieS�($�z��c�d�*�m#�'8���5�����玴�x�;ĝ&�平����Zr�&����2u����T�D�)���ȑԫ�dFY��Cn�}uX|Ua�H0fV�b8����=2G�������#(9��mț�x&a�R��m`��(�/��B��q6+��	��(s�8�vY�7 :8��c��HRR�����@���B'=h�����L�(gNn'�8[�^�:4Ϩ/HT h�+�j)�'K��`E�<Ζ�g��.c���fא����m,=2�v^�,�^���T�ޕ� "h���H=X� �ib�L�*�a�
�f��������U�6��ɐ�5�"��>���J�,��sL���P�����0��'�]�k�D�X���,��_�]�-�I�8����N�v�<꽪�[I��o�O�DG������(�^X�]g�3{�;�&F]<�`�����B�	���fڝ	#w�W�ل ��	U�����|Z1�Jd��&��t�MڬQ�=	�)~�����~ ᐏ����BVS�#�#�5�g�U���x�<��4��zNA��R��w�"�q�3
@�D�����ݜ�bR��,��������<�x��+X�Gj�����oM]ȏ�\W����B(�A駭AQ'�U[�u�'?����X��7 �c��f2��[��un;X�k�� �Qϣꀕ���� ����D���ܮ&+p��Z+8���G3ˑ�ߠ�_<M�{���`�m[(�D�`���|�̈Ƴ�(z�X.d_b��w)�^�U'ܪ_��;2��d4Uw�D>��q7/m<���q�ag\�0��^�~ �3�[}pl]�$`s+�a���nJ,c����'߸��������# �(���7#{�*���!�%��q���|`2s��'�u�sh"Ԇ=�}�y�7P��4$��ܽr���o�(4�"0d��]R���l���Z+��7U�6u��	8�q�W�2�R�2������7������O�Pр�vh�W�Ow��\��������>_�lp;i����r��jp�PM���S�I<�gG��z�!sMƠ�l�������PQ�t>��bхn�Q����|���1l�՛�E����L�Z'�?/�k$?z�A��D�����4��[��#�eب��0���IH�l�h Yi5�2��=s7q��M^��а� �1�����2֡�.Y΍�r��5�����S�M٫�L`�Jf{t{�c�P�(��/M�	,�g �Ű�x�Y]t?hm�}WLs���ku�HEG���[]p�1�j~9���o��H��2B�+�e���M��#T�rA�8� 1	 .��d�{I���G�)���@���:{6A��1�	����4��7"h��_	��1|//#�z4ٞ�/T�H9Db,F��fhǑ� �� G��&C�ɦ��R`����Ek���Ab��=�sR����A<j�F�[�hDg�i��Tɭ�t�%���n�ʞ��%�b��H�F����F��E���ryR�t�U� P ���F����&��05��``����L��Ɂ��h�1ﶟ�2�&9f*�L�ҼT\�T�b��}�1,i֥f	ʾ����逶��O�eCu���|7�����5s�xß}��j�{}Lt�Dr�e�H8V�zx���GՃx��G:	�	�[t��V,X!�Y+nV�F�"e_��6�:LT����>�)���XO�2]��K��a�.9J!���3v[L�A����_}���6Y�ȹC6]Y,�f��'���1Ͱ������b>�7<k�Ϊ�ˏ '4�b��Yl#8���7�T]փt�K����9�+2�z�0*ڮ{���+-kc����a���P;�õ�Gao	��~3��&�kx��׀Ƀ)<��C��$����zB������[����h4\8ǘ2�?���O��}O��`xۚ�z�HVo D	��q������?��u��� �i�b��m�)qj���P\�w���^0�r� �s=���( F��/�q#��c����?�[�3@�9/�%k�F�t����GC�aXu֘�.B*�o����ǝ
��#uE�H��b���Vm���9��1MH\�XG�i�BCMS��c%���NՊ���L�f�Y�����>�r^*JT�>�C�W,0#]����"�j�T��4LݱKt~�i5 �Ta&�FJ�¬�p	�V�������n����]~l���o�4�����u�M��ld������r'�n���3��tF�H`e����& � �ROr�w���B>f�0�/X�낸�t��mY�xn쫊��IMl3z�T𝭨q�Ը�;sUm�]�	��m��d&>Zi�H1%y�c�7���!"zge����F���Y�.c'A$��+�9}N_���UDu�WzX�v}��O+�o�����CnE_rx�ʒ�E�8i�]s�b2sPJ�2ܪ� g̥^:M��.�VFC�$�F]��x�B�W�)�b�l�s�4�׾��k[��-�i��El�.ZE�|�2x������pjy����6����7��mU$��J���cw^ ���BrE=8ܞ?������B｝�5�!1�ްWs��օ��B�� 7J�(rS;�h<:�55�:��Jk�/M�Rn'$Ni���f��񡞽�����-v��iP�*ʟ�H2�?p-�ׄ3��g���Um��x�V���}�"J��d���#ơ�-k� ���d:~N0�o��s�ˈ� ���e�_�F���v�Ռ:�
�������%�!i�">+�����V��r?	�W(0gA�SN,.)��9�C��M�g�rF�tt%%S�!W��":}؅:j#�A����K���@���m��rE����S��i���n���E��
E�"�+Q�'/t�D���+��8y���N�e͐�{ˋ���q�0�g~Y,1�N�[�&��a���kkK䰆p��n	��{���\4< �u��/��u>_�>���@�`B|e�o_�냂�=<[��o,�C҆o��MUG�#��{�6��Q��`�1�&�`?�;5��O��"�9� ? �7RI�1�QM]�#��"�D��g|X5��Cx(35躙}L��f� ��N ���9�C��L|�&#��	�WK��w8̇D��)f"�|��v���yd��"9C5*�I-�GC~��_1-ͷ���A����v�;E�Tu=\�K9/t�e�j[ܨ���?z5%U�`��8��O[\QI���ݹ1�F ��銼��=�D�o"��9�ݲlJ���y\KgQ�,��q��"S]��`m���7&m܈"m�}��.w*�RGA���G��։��[9כ�ђ��
���	��I�r�E}���0����H˥Աv=��М���b��r�ry���}=s���E�B����V��}�7�-\���fR�@��9��?����@5F�U�͋������#x��7]qTM���|��-VI�����g����󨻞����&&�	0��n���i�KZCtl9��	T�|�&h���0SIM���R]��V�C�*�ny��WK�ȄE�����Lm�5��;S�ܮa�?6�=ֱ�)aG��՞���W����l5���q\`�.�gĺ�����CZ5Z�Px��+�b��ڮs��|�;��)&].*�K�]���עd�2���'e5��=ya�(�Ibq��'C�c@*dg���,����f�����F���^�SC�g�� ��E��X0�@��yDZ�,K�� /�> �;,Z��C
�ńU�P����^�����������`�"�&9��Y�Ϛ1#?^{N��j7�4��%�0D��	���H�!�Ȕ*)g�D�,f2���=8)10��?t�_��XdhW��Ê���\��Y�m8�*8
�O���A� "F3�@�0���<oO4s�[,a�9���[����B'�N=�]X$��V�܁���ˈ4����"�-���t�㜘�֣J�ĵl=�(wk��/N�J�|H��xQ�{����3�\������]M���E��l�h+�6�X��;7 i�c�����<L�������6��P
��p#���!�OM����z�	�<)��Z�d�S�a�{n^<U�^�u��Dn\�A6a���]��1����H���������#��Jg��X�@�����L�}�]�y�%,5�>�Q4F�4?���`)v�0�{(r�]e7��^�!8�1Ee�w��m��$1�$=��5�00&����r�������JX�q";��^�����ov�-�\�Ӝ9( H�D�;\k�d��P �����[��r�fV������.�\�a9��7�:Oy=̨Ed%'�,�DL~��-'�`�>x s���R�rDD+�hr�ա���F�@8���Q�p��b�r�*І%Gi� �oA�O�0?���mQ�L�L�8��u̻d:�7#��mm�j��'��~v뙛ȟ���I+=mT
87a/�Ɉ?��J�f�%�i��p�C�,��Z�k㱛5S��8�}�V0���k��&j�͏�n���rl|޹�_��@6M���LVj�/Z���C��ù�&�	a/{��r�0�l���e!�]��{|����(M���f��� ��0�� �"k��q8x�[c`"��,��WˏZ�Q�M#8���ܷ��u�� ���u_�a�����?"$�3�1��]���2�������������϶J������gb�C}8׆������>e�#y�i���Q��q��h��z:(.�d$?�K��=�HH��u��՜	��[/�^��A��TaN�E,�I����/f]�*ű������YN&3�0��cxq*+~�г}vQJI"X���d�QK X��M��Z͊F���� �DZ�i11:�X�x��co���2��$��8$�-��l<�Q�W�	yP�W� y�z
ן>��r�����ĒJ ���8ҍ�����u6���+R���n J"��3W�EgP+���V�#l娀c=$�/9��fw�`ł��hM.3�7�c�"X��Tu	"}�9�r�{��-����I
q�Ӫ&�9�:m�d�G� Sc���`-���2�R�j�� �
��hX�Xl�hK=���r;�q7�a�i�m��+&�5ib�Ǹ�c�����WBL�y|P붯lTl��I6�$N;U˞"�T�{(00�Jq���m��͛=@m�&�5����@�5�4�������0���N�։��pUaB'�q1��lr�{� ��;6�4�3X,]b��5�@@�8�b	adGms�'�<|eF\��:s.gL�L���0B�|�c+��]�V䜶���B|R���L�3��4@8��2������Uy_sN�0���i��V�oo�E���@��;���E��^.��[\ۢg ���X�)�͜Lѽ)7Y�sЛ�H����u9�Z�`M�y�pR��/WK��˚�i�P]��`w���q���Y8�2���\�)���z�*Z:�vy����	�� %R����e���K]l��L.9s�&@@�6l�b� �1��j�Y�����W��J�"������pEM	%e�VNL���lՅ��A�
�̮l�A��dH��C3���f �y?�29�f�F�_Ȯ�0�e�[��*��K���҆��"�{���9-�Z��IIQIH��df�����I�'��Wġ�SG?zruش���_�T�R��r����=��%�����y@b���WVݼq��Eߊ�����Cj���f]1�/�7ʨi^0��ZSB����<]g��=�z� E�سu��͂��¼}k�cgI>9�k���O�՜�_��Y�K��4�D�Z�=�Y5���)�X�W��굈�;e�
�Q�̈QZ���X*���^K� /�df_�' �w�I��s��=B�`j�|&�Y�軟Uΐ�~#��0^&���z�̳�^��G� ���7��A9eks��#"���3Ú��@.}�a�ȣfP? {6��K\�5���]�>n��!-64׵[j���80����(�p���Ȉ��;ň��worf�9N\����5��%78y��W8�|�(�OH����`�Y�`�Y��3��!�Z�Fع��Έ�?�����἟+t;��)3�L/rW��.��Y\}��\QEd�JL�@a��O=jp#o<���&�1��)�,�9���θE��=N�,�?�X��3A �|n��;���I���V�S����-���۟���g��ikl��� V}��5�`��'O���Q�:6 �#�N0���w�un,�=�ٟ��pX�to���:H��x��e}�/iƤ�Po��yG�Bw�ђ�0�\f �=���ႉo�ē�Q�/�E����]��
��� ~�yƹy�M@�sf�V{��qj���%�3�9:e7�iP���q
x���(�1�i�k�;��^�����֖# �$��8�Հ��L����^k�}���y`���m.WXTV �/�)��{�k��?�B�ר��ϐOzD[��E���ut�����̈�=�Ѽ����1��,��wdhD�w�62I�=�*��6�������Q������d[���E�	�h�	�ݭ�2�����sQv�r^�]��ǄIm�7�!N_W�OLݾe�:�!p���o���k�J��$���R�P��o39-��,���U�`�k��7a�m5�T�P--D�T:��G4]�oh<|7/I��E�H�M��Z8M��,��=�h���Ā�MY�xh������*Ό�	!(�O�Q���Tp���!���k7��̪| =��o��W_�q�=��{(�YEr�8�n}��
GTۘ:R�~�Q[�[9SO*s�ַd�}hd��������� j�LA����^%�,��Y���tT�j$�"_`'xB�){4��rD5��\�f���=�9GI����op��b����WQ��a��]�t����H�J*8���C��d��b���n�%�y��L�qP-XP�ށi���E}E��Q�>���O���&�A�v���ɍ�ݖ��;[]��v����W��n&Y٤���v�� 	>�XY�$ə�aIZ\��^	�\L���{[�|t�ά�����?���1���5��a*��p h<����⬘�T�������/��]{�� q�JN@���f�x�]4��X�?��V�$W
p�{T�;��;qivr�ՖSh��u�Brʹ�(5F�
���"�5�,/�1T��D�$H�m��1ƜEA��dhD���ܷ�\ hd�l�@�ʕ�v%Q�*�ή&#h?��j�k[�~_F	�.�S�	�'
sm������m������=�vv�wq�^h�gD��$r�ݎ��O�F�kr+m*��{SbJ�"6�W�,DX�Y6�@A��?S�2h��n�,�Q3ؚ�x�^xT2/~S�d����> Q��eb�h��� �~F�,�<vb����V�4��c{�Z��ӥ
��O�-f� 
��vT�,k�z�ik������7%���8	b$ K?���{ri�+
Au;`��6U����K�i��i:����-�?��G�#�Ǎ�$=aj �[MJ}�
'hr1�#�e	xpY����!��n8Dy��ꢶi:����<n�{�Z��F�
&?��h�[$��1S^��owz��s�� ,�]�>��I�T��<�L6y�R�9��8����k?�x�<�٣᷃&:��Z:���L�;ĥ:�q�%|*��F�@z'�����$�t���&�
�����d�I�ǳ����bo�D��1@��5��`����z2�fk�U͌12o7s5a3�NwQ�`*cv���DS�cBĜD%Eg���`�6�� �o⍊q�T�}#�v��igczC�8��s��o��(��h�τ(�����'���Т>���V�Y��C#�E mI^ޮ)Ƥ�נ_�M���_ y�����!�Z~?���q a`�߽W�| ��k�mO�Q(0��]t���1���Q��j�;�mN��?!+U$W�X���Hwv�'��/��Pe�Y�αh��Ԋ�:4���$@����#��?���JZ�A�E..Է+�F�f�ej��`B���H.5��%�oi'��&�#�	�ѽD�-8.���5yo���R����zx��v��FS��R1Ꜣ\����o�b��m�l�ڌ�A�f�KL�k�õ�;�A�9o|}���p
���V��`���80�ױ�&��o���?���X,λ-lb�kCz��*I聁`9���
��H�zE��y��fg��UjQh��;7�FǶ%��O���g Z'&	�����Ђ���XTj�r����k��� �w�|#���>�O:c�4[{٤�r�5�=݈�=_ث�O�8K��˹���+��
�.e�^$��.˯�3��]%��HS��@q��x�ճ|����F��h<'<NX �.����R��-�|��
#��&�?���� K�L��t]���i��8�B���i@�=���B`�b���.�����l��>3�oB�~�����k~���J]�Lہ]~�8�d-3�h��|Q�����2d�E��s"�oO����6�m��@��
�7�_��l3����5�x=��GծF�];fJ��0P7i+'-��!�i �(���P@z\�I��Xz��OxFZ�CÌ�;�J?}��nQ�`T�7��Z�?�t�q����	w�f��s�{!5,���|mov���uA���"v���`�Sڸ�#q��o�G��r~g��t�SE��4v	
?p���f'ܦ�Q�NF���W�K�9s�~2|s��m��h1�E2ٻB;㬗�W��t��}"#x��y �<N�f���z���5����de�~dT{�-�w��c�1�0��#z�OO�A�4E�H8��>�h���V�������|#��J;��DͶf�Ɛ�4lB�b0h�Җ���kX�X����*�si3W[�������q�L��g�}_Lo�
5zM%�<��|Z�K
�d�q�c(���]�F1�ϐ����Ei6Z���-��lV)��g��"R�����P��nJ^5Rn��O�L%l��ч��U��K�G~�@e�>��$�g�Oɒ*xC��g�m0�A�����.2���#B�qb��}�Ě��_����sf����x��i��w�xvYiED�4�X�Ey�՜�����;dc@���̛������5�TjP�gzX$�v��g�k��[^�/��>��,���7q4�!f���R:�W�q���|,p ͉��b�F��D۫lZ�u�
�LR��\Y�:��'u	UZ��&u�ܙ3A�/�bnUI)�;>Jl�c�� I�͎��W�$]k�PQ���7��P� {,�{\� ys�l�&�B"..�����V�$@�K�����	#>젭ΥՅ����1���O(��J.�(��EW#�.=Z�=E�-�����s����;#@�Eq�hr�� +��r.u�"i�d��g����M���Ed�
ˠ$�`�B�����M!���'��˚Ju�ũj�'��ɽ��o��IQ#3�9�c<HE��i�i$�2{%ë�Ε�[�NX2��w>i�GR��B���S����o,ns��!Ԉ�hUp[��$�!#.�S�qӊ�G�px�YDvc)�p��.m}uڻ���1?�����q)�t�8�W��}氜�'�(GP�#����@�d�q��qj��j"�,��T�%��E	�۶ʴ�#��qY�tē��퐙]�>��>�˼듗A9"�?%oY�KP�k}�vp�B殥��V�B�{O��s��=�ce/��{��ia�R�̲J��S�C�?���6�P�F��u�����:����2��)�Y{��^��j���RR3��[�g���:�u�0J��w�2m~��G�f���(�a�a�'�����i?��BB�U�20������֨�Մ�!��h���ɩ2�<^���[�D�<� ���t[�ISA�NV&�RF�ޏ�n� �H�#������>��V=��yZ|�Q�z'�B�IO7��v�g�oFl���Ƅ@d�SZ��p�_���HP?pPy����.�}�#���;��[�����1����w��$�Oe�Vg�9y m��n	w�8X|m�T�]�v�g���2Q��w��BM&�[��K�i)�#1P�&ޒ�vza�J� V	\�����L���/�ii��QR���~V��҅�M%�v,�b�C>�&��z���	�L�$O�v�!�$B�6<�7������#.�Ӳ��"~�|��f]���K��6�����Y�X��_�>[B�~�o.��*�_�����&��T�p�Z��A�'�ξ#C��.�H��J�,/�>��e?�O{�@?�(�zQ�d�K�p�e@�b�~�a�ڧ!N��˜�lZ��P�2d?	f�n�����N�=�����Ъ�wn��R���PQ�"B�LW��^/R� ��\���Q,^�_���aɹ��v��&�[^<�8!�5��'E
Ҁo���%��C�;�Ju�n�8 cR5P!��<�:�μ�)�����+ �rP��#~5�`�ӕ]�\�"���cLd�h��f�/-q˄O��ú�#rZ��-��Vg�:2 y�Iش����q�HK�QՑh؄�}�8'EM�b�#�݀�Y��W�R�����.��%��
�)�U6@"kc,�T�*���SV���x�5�И���)MO�Z�{�o;�`dїWbT�g-ԟ;�y�� L���i��w�jY�]�#(�c���Avj�+�%�RY&�B	��&lz��� 2̖���Qo���̫�d�(:�D�a�� Jr2]:��d��2턂�\�_�K�"���Ě,(g2���|c��`�\�����ݛl;/�&����ż[����-���*�yL��1(���t	��"U���sar=,�A`�8b2-A�b��߮�[wԤ+hA�B' ^��
�POB�h)�ml]}G�8�s�ٶUb]���#�|��H���ﷰ U�����Z��P���E�ϗ�aVɸ��i�)G��1vhs4�=r̾�v
���&��C�	���a�y��i
O"�C��k2�$�׫����;�u���������_7�C��V{i��7��[	��b���ѡ�O��v?����-�*�D��3$�-T-�m�ɔ��ᥕa0�E�o�!���I�r�\n	�K�V�Q�P���FuJG��B?3��z��B�3����{8Te��z�S��w�"�`A��l~ý�5{�t[~YR.���5�*����It�̾�4&����x�T��[�zb�2��b���f�$���7S+8bk����b>j?����;g�iH�_
�p{�����#�e�3R�e�3H��W;H�l��ӎ>�+7�8��dئ�?Lh��Ak|zJ�,fs�17#�\�������R?7H����3e+��*����c�x�0RI�8�ga�/��>�T�4�K�)������=���0���X��� [1� �K��<q:-����h�b愹�@i��F<�W���\�0x�s<�q�E���KU���1���v=�[3:����;:Stm�߈�2Q��S�$[bW6��tR�E��C��T�
�EwF�򻗎�6�c�y�֎�6�K���NR>" "U;�i><�"/->�J���S���N�m�/l��^yDau͊O8��S��[�f���hJ��d�i���Q��mu�!Ђ�� ޮ:�|\"��ʨ�k�"���n�`E��Qii��]2H3탅jC�w��=�����w�B@��c�Pau!J,[,�׏��J��!x�S�|ؚ��ז�F��6�'�-r0��5	���u���ճ�n[\Q(֗k�$�V�~�i�7@��)� ���~Op�YH\B�r�q�@��ե��86CR���n�9nc9�,�N��RL�`Yr\���p2��{�A[jk�+&;󵳙�#J�Ien�S��v�N�jT�	H/A��ګS���9����w�
0���V�y2O˷�9!���um��ӞCܕ�F�l�`(]�y����T�����i3"�t-��ʰ"T�ܕS����,ۍ+ ��3��*5���)�>��jd�[(��1�n&�N���2���?��r�8c-��s�a<iĲg�{����/����"��
﵄-ԩ[�ߝ[�#��"VY�����o��2, �QF�.1|�!�j�-��륰���](�v�4��� �a%&�?M��6CJ�e-�2�CP�Hy�G�����<T��N���:HϤ�=O���f�ߵͰ�蛼�Nw��aa�I�����z�7|��c(�[�����|R^�Z��H��!�l����Wĉз�`�G����La;IG��K��(9�MΎi�t�1XƜ[�K�A�+�5FS��7�?�Dq�!g��F~�.R-;-A�<���jN^y�#�-�yYfv�@ ��#_�>2�?����su�ǩS���7��YِY��'�γ�F:XT�^Lm��˵�F��p5��Ah�2 ���&�Al^��ᬰ?��9��0u��D����΂KÛ�x��O.�S5Ƹ��z�x��b�7\6$�5
E�-�)A�<t]5s�e�X��K�W������Z�k�<�e� ���޳��À��udL�I��}N�󮡨�s��� %�L}���yŅ��r+��7���%8��U�K��AhQn������-�eO�dn��ҝ�I�9V+��k���|͕�Dl�[&�J�#����t���ןT�ye��e�j(K>��=�+�&P��)���k�?x��p��T�(UQ���֥xN��T�Hj����j󫪃Mr_@�@������)t�Ѱ����|�,e)Omc���7��b�3���|���EC &'#S �a�7+t�rѩ]4#C��֐13`�m���P�q_z���ښ����y[�`݅yK�*>�a�U=�k�yvwQB�oD?Ƅ���>��GJ��$�ޚ׈քC+0�s}�@+|����5�Kf�7��\oN��ϭ�yd#CZ��^F���<��a����9ܘ��t�΢^�z#�s�^R3>DO/�K�m�UE���w��M�ܡ�`����-��||�E�U�Q�z;��}:?g�����Ѳ���R��R�5�$��;b���.wD[��](��ϡ+���@M}9'a���-Iݕ�6�r���f�� s�P�!4���#��C����`糘Y����h�>�4��0t3DMx�bZEn�{G����ag����Ǉ�G(Z��UBU��!��	T���J�;���Y�z������Q4�0�����ٿ�,lH[;ݟ��U��Y06��8q����pbn6�VEC����N�A�/q�uzDv�zmH��o�ժ)2�z�$��η8Q'*���x�3*4��@�0�46��vK����q|��C ��� ��v�4ȁ�w��N����#�C�X��nR�;gcy+N
�Q�ʛ.�v���x��������
��d�0�	;��B ��9�'����w���lBR��-����Ί��q
'��`|G`���w@��1ؽ��t����(F�o�r�cwu�-���4:f�-[���G�R�����z�^����I
Ϻ��ࢃ�ph�s�����^�$�(iZ�˖:���)"zD�
��e�W���
���
�h�QƁ�����o�7W/f�Mల�O���3���ɮ�>�f���;q낒4j��ɱ���
)��)rW!�U"�hN�����_@��6X�E����#�hQ�1o4���"��l�5�^���n/^���?{���ʷ�e����ni(p�Z�z�C	��͵���a	K�K����:��)��1��~"�B��\;]�5��t8���\����o`�4�9��z�
���6�~l�?�KT���eƿg<\�q��1剥H�<��"s��GYg�	sS���[ fLlW��z�ܬ�'x���0������E��6hu�5����C��8�U���G�����t~Y:H�7�IZ<�˫�r�x��^��RW����}����{�����������M�(���Z�:zl�;�m�Ю��d�R���a9΢H��oůs3�#�R'�:z�ɦ�L��ʑnCJ�-��nTĹ�G"7$7�n��>k�"4��.  �;�>��kujzp��C����4�8@{R@�ou��(yKVA ���&Ɏ�����xΠ&H�ʒ7%D)�M�Q�K�;�U�e�b�8|9��e��E�k1��r��D=�IR�d#�m�7V�%WZũ)�J �	$��@7(z�l@:�jKc������`@�n�
ǌq�4x~G��[>3k,L��ё\0�u@e�o� ��J�;�9ɻL��� ������
���|�R�wF�a���b��D�a!z��j�,���N��II��{����[��d�|'8�����^J1�������L,�s@�mP�%��?K��p��H3eWKNDr�������=<@�� �����x��1^�|5s=��V�+T})[.+�����U�Z�X���M�"��6��$Sv�җ�\�
�����ư���w5�1�e��!
�&�qWY��ޏ��M���M*�<R%��6��!
K�ٚ�{A�ֺ�ٙ�~o���faH�����[�S3<]���s�̛��@,>'������|��&�3��R�
�b$�gޖ!))��c�h��ج�=x��ו�������2���6k�!.�+�C��z��@�{g˂��L��+���P�oj�&,Qa~�0v�Dӻ+��s�_����lf?g�-���~ҸQ���>�&������{�	#�ox��j7t�X�� �F �b�����PǩC��Y#|S E�H�2���,�<�Ӿ�p�/TG?�*6�vP�g,�g�-��P"���M����b���"�i�e��j�_��b�I���S�f� e�C�d�D>���T>�o]k�ڋ��R~����k�W�͢4����B�{������DG� �MS�UF5C\�G�i�W���޺;�3&S��sP� SmN'�_��իB����Bl�*;/�޷� �[�ƙ�e+�o�����pS �f�c�/s��V�����	�V&o�R��D$,ƚՊ�}��k��p3.$p�ː_�+[s�[1�l���$3��
|�]�)�� GW�}z�=��}�h?
6[TX�	O6%��\v�1������H��w��P��&�#��J��֙k�s���<���F�M�X��+�D�[, ���;vE�K�K.�j�V{۫�ǣ ,��"qQ��.����S�(e�dj}+����N�)���8n�?���b��և�(f�s��7_��17�ڲ�
B�u,Y���W����`��r�c� a�62[p󫂶�e�ȡ�^�i�ܭ��"���-���}����!��}-�?RS����ƙ�S�2�0����[Ӝ�(?V&��$�h�<JJ�3�zp���IՊ��	o^h�d�rN�r�J2%$b[ᳩ��`i�U3`p�'�i7ýS=�mR	�ť+c
��
���k���Q���H%g������Cx �iMIl�{Ay���"����
|/:��K<�+�j�T�f3F��O�Pҷ���.�<�[���12*6���}P�u~��-�%���wY'�!8Q����S����+Ƽ�����u��R���؏e�Ǩ�#ĕl�'E��(+ԝ��}��Gs�\�DT�|\��#^�r��_"��/�5��/���
E�<DU|�{� a}Ƭ�C��i��ݛ0�z�l�]�|N���;�MV�.�6���E� vJ֔{a����}o�2t�x�g�OfL��9ݍ�&(��(�+�m�D@h��������G��:B�(��)�׼h��=F�nNя��	DO�7�Գz��K�����I?�dV�& z �l�lØ~��1�6h\�*�b^Nh-\�/��|`�s)v��F8tz��aVSosc={����P
�Ɓ�t2yH޹�o��7��[3ց�n�/A_c�KY�u��)��t%[_�W�q���~�C`p��$,���[��+60��"���'��d)��q����g�@�z�
��raw�v��9葕��	+E�*_�����,T�Q ?���}����sdQ�y���� H�E���۬x���(\��)����[�q��ɘ������{I����`V
��i�t��'[�@�]����'.,�S�ث[�I�bx�3fk0��b@���{�=�>���%!�T D�ܵ���@#$��B�C}v�L�D'���4�$��u��z@��:��쥥��-�s.�t�`�N(��k*��Ri͆�����L�gf�̄e��Q:k_l\�a��ϣٿhTs���6rogd��*OȖ��������h�*r�D�����1��m��T4��jvS�5A^mg�ϊ�2�� F�Ѽp�[�N���]��$�Ճ��T��6Q�[��=V�����wOD��'�4�b��N�_��M��f_]���J�*x%k�t�H�M�,ʇ��`-�I�ʳt���E��>� ����>HV�������%�����+Q�wK�Fp5��Q�$������=�&���Xޡq�B�I�����	d�vr#�\/���@��>�uMS�1�B�4P�l��ft5��������]�[����ӒN��*�F���l�:��ժc�u��X2�
nx����{_�/���'�=�6�.�
ц��;�iu� ��]�-X�8��`7$�����j��/�t�P���HK?��&�^��n���0�����r3�ɤ����b0���ԝEl��^}D��-	��@t����T�-��	��Z���p_�/�U��du���ə{3u,���}�A���׽�{���'N�(޷������=|��X�������A[��?��)Rl6��gQ9��P+Q~�i��1U)kJky��|����8��),rm~�E��B]n��R(��y�2��y�FY���!M�?f�;Y����O(�#��I�>�� �	�lId��l��~�`���P"��?&����5p�D��7����
���3�3�ŔpPA�ba�iRꦇ��Q3|��� x�類�;��@��nP킃>S*�I�O�௜VF"�V�&��
�CJZ�'Ѣ�l-�}D�������j��:���IT^CD���h��G�Ʊ,�q5%i��뀴�w�WP�ɀ>��8�h�i��zȶ��b@!OB�Ú�[D��	!3w�A�K�Tu\��c�@���U��(��Bo��m�4W��l6h�ոg�k�[��ƌ�-͖���DÐ E�2���c�so�,�JQ�v�d�~��]�*����u���Z ���(ҽ�9�#�WɟP�<K�M�p�[@ʏR�Fm���la�̏|,�A�b��H2�X�6�o��>��`��!�f���8S�sf��]��SY-���3��]=�+j`�`��������)��wQ9v�3��a��h'��� ���S�z,3�+pAg����!��=}������
p)YN�4�: �e%�Q�Ho�&�7N�,@9�c��EF�?�{�z�^�7$'��&��*pUɆ$�ePPǿWé�i�=-fI8_�������x����5���#��rN��Z�g�6���tR�N���@�
#Y�ӗ�� �U�B�lC*���6��r��}�pL��V�����}�P���,"�����hs+��g+7�3� �7�M�äʖ0n���}5�-=QnΈ�Ӳ���mN���q=�5��f� �@�.���pG�>1�.L��cHatt9eI"Y�����3�����.�7����[zI\�T?�����f���_7���
7���^U�|E�7q�L����.�wz��R$4O��vZ'f/�?
c=K���RE4�KK2	���z�]G7�Ιl���X �7y�iZ���c�����k����Cú�}���Mu�7=�jGdS��H�S�T&h��Y�c7�#�0@�)��"Q�|X� �@�d����j� ����Zĩ�[J6
�v��$��Ɯ�ff�ժ2�)�L��)��z:�.ӻ~2#���g�P�p؏�3�t}�v/yXt,��8z����q
]�P�ȻVy�$�o���e�j飌 ����WU�	2�� ��bD��bc	8|tgG<J� ���}�gdO�I�R��F_ehFQ�b�qL��&�,�����U����.�7b2~��A~	�GbA5x�G�S4so�����)�}X۝��B�N�p��6I󳸿
�2b��U�v6�.y�:�LX��<X�D�R�������2@|Xpz���Ef�������O���y��Q�b��i�cM�{*`��I�C����Vl�}�#i�E�t��~l�Sww��HV+`�H��!�9f?w��e=)Cz��O�	�{C�%=yW�}z��@V:�y��~�@Kv'>&�6��fm���c;F{>��+h%8�F�߆֎�#��,B��h?�S���q�ת=մ���\�C��6��RͨDݱ�!a���6�e��D	�%դ�ԝ��I�y�q���P�8Qg���������@�z�Ew�rCD")w�+�(�ۊ�O���^�6���V	G�������R�h�I���HhQH��_Ԫ�]�;b�B���'w�&w��f��[�"	7�Bf0ۙ�oa���6��(7	��V���m�
hυ"��% ���Fh��>�
��=���e�WO�6�W͍�_�Z����� <X51q�7�s��3��8�>�ڰnѭ�N*�7����G� �v������X���%��{�ɛ��A �5Jc� ��;�0`n���S�m��9����<j���.��A{��(_�P{�pg���E_�6��t��|��b��tA+�9��1;�:�fz�cQv~�aV���R���NB�oX���jzT���%I�I��p*|��'c-E>�{I�(r���|˭��7��
�,պc~�������<�GǄ�p�{:�sp�t�qPh��X��@|舛n2.��nE�&��ђ��w�օ8�&�{�κP�$���#�P�z-�w�"1gPb����N�<5���6�'K������3�K�oJX4����>�����s#�I>�eM˙r��\*k!���J�_�`#��K���D�x���e(٪�1�
�Z�����)b˃-�\!Mh����~/��G]�CBֺq&�������$��N�MN*�S��(���]�o��~X�s�X�6�ծ~�-��0�`+"!�b�P"$U"�>XO�� ��HQCD���3c��JG�uu�.pL�.zc��q�b��}�\���)@YJĆ���9�m�����6$P��1 D,�� �����~�wN�wߪ���~3�E������!��i �����@]����P��E�aQ�i���T�0�DV O����0]��W�s���C�Pm �,��I��.e8w��l"
�;���F
�H�H?��h[_*L� ���;ߴ�57��I�L�KH�V� 	wc�yf��8"a�V*��?�TW��2R!���"B/K|�{�[l��`ݩ��~�!�2Λ�b�/B
��Co����#k�Hwg\9p�i��p9� oQ.KԻ*[
��R�Tz!r��\�
�3I�ynu�N���0dʩ��;�VW�1��_�a����[��O��m�B4J���hшlM��,,��Aej�8�����#�{
��I�B1E���ap�7z���@�l:E���_)�	�ݿ��.�j����{�u^�d�:��1ًR�ElQ�,_��5���y0�������-��� tWe�[7�Sl��- ×���Қ��)�5y�e7{7?�4��fN�u>.����K���ɸ��vF��G|�Yt�_���=�H-��
P"t��<-����@\N������ڨQOO��t�c1B��f\Q���l�nO��"�g�
��@sF(Mai����$mt�n��A6/�rJ
�Vm�O�%<G6�0��M�������'�D�	���%��a ְ3濪]��&S5	r��@9]}�v;S�_��=�v�b�0
�V�v�B�C�.��,�遼��R�Q�p~=H"���J�n~�f�f*u��s>�P����1pE$<I�)��9J���'����ې�0��j�ϲWD�NkoǄG�v�B�T��frPƶa���wE�h����蒀R�H�?��5(G�s��,)�Ĵ;<�L�zi��@�L�S4��2�a�9�A��R	@?7��yED�:e��ٱ�)i/��������y$�^Ae������� ܟU��
?���Y�c�!;)g_3m9Ԁ�>=m� �~�qI|���n��I_�>��4���ĤeĦ��2i�u��" Z0��.C����M�l�|v�}���`p{����lo`�T�Դ O��7G��A�N1[�k�s�p�a���H�
���l/��LO�ƴɽOkV��;�(��{,�-��v�IEp*<��0�2�Ѥ1��K/��V���	R���^}�3�����?�� */],�oA�mG�T\03ւI��Ȯ
�$y��MՌ���kד��U�4��� l��"�n�/�P�WW��8)�i���j\j���̸�qԂ�;2y	�Oq�[�_̙�r�i"tj5w� �<NNh�u-���M�߅��.5e��A�s������0�'�&���;�G���e�Mm����Ĵ����S�S|j���0�O�4Zu�Z]�S�j��b�>`S����w=}��g����l�1Z��|��7�:.7qi�}�0�	������W8|����CيD�"t[\m�{gH����nJ�.�)B������.fεh.yW�vq-t��t�~�"
�mg	����b�CcR�%�6g��)/וm�	����l�5"Q1w$�:��{ᘞ9R���c��w��x��9t2 ��Y��r'9@���Ar&�Ǡ�Ip��܊GԢ��Uy�l���0GR`���4�-���K�s�6��\�%�h�NP
,{vY	X��K����O--��+�6�J�z�c��A"��A��kCDfn�(��*�u�c�B��r.7n�[�CJ�.e��Vq�˩�+��fpOhT�JV��j���7�_���Bvx�\�?�{�`���{�:�{��/=xϝ�`�g�p�m�M)֋3M��Q�%�S�,� ��r���h�m����!�b��Z
_�[�镤.�'����BҊ��z��3�&sep��ͦ�y#�_�.�O7}���i�-H�7�<�~#z��O�B�պ�=i~>��e_����J��s���Y�����t��0� ���KHw�+E�� ����Áa��}�	)~A?�QeOwk�Pd^�[�|B�v��^��4JBvV����s
�A/���M\+N��\N�n�����DF��J(���yW�0[)��D�VƋY$�xeI�lɁ�H���3�H�k$��%��,�T�:?��a�I�6hM<�� �b��ep>�2��8nNJ�L2��6W��/=#�5�q]�z��H\7.�H��Q?^�cA	��,N���`����>��.5W�+��x����3y;[��_s�Yi�m�m�|l�c��g�������K]�����W��9��_+KJ#D��߉���H�:�L�� � �l0����2���6�u��� >c_^����F��i��Q7(s� E:6��i��aѢ�: �t��)/"�,�X	]ͻ!����ib��{����A�幄��S�D����	�v�k�4�`;�=���\�̈́\}+�kգ�L�Ļ��?3���z8�@�PaKvAWy�wj�k�ns�mD]݊/z�C� 4W
���d|/
����Lƥ����s��D����g4��v*^�t6�ݛ�x�#���$"��A�k0y]�B��́�7��A���k�a�($�&������Q&mn�tJ����xv/��r���t��ua$����Oa�N��Ňr�V�2A:0��&0/��T�Ot�U��2F�
Y�a���Q�ϚW�ݡ�$;��fY�u���^&q���T���>�\��,�	�nY�I�9���񬌸T���!���ӏ*� vq:�*��~�8x%n�h!T�8�|0�S:rg�_���0���H����~aPBq#��&��[�U/t�[\���5-��J���d��^�u��d���,Ə����]�/��~}��qF}���`��?Xư�C��i��ko�ތs���wv�K�K���d� $/Ny��-Փt4.(x����S�g�����W�������lt�T�8�W��Y����ۉ�޲BG�A�6�v��<<�����W;�xBŊ��og�<���;���E��{��QGZ�h�'����[(r%5��rI�Ћ��e5&���h,M��(�S
�&zl��%�Y|�G3�c9����`_�����ä'��w�T��ye���N��A 4Dfo���t�������6�_z�ݓ&� ��:��(��i���Y{ߟ� ]��>wE.}P@�A�-��o�θY�q��'���L��Q�����n9���۸�5Fhl2����b�(�R�\���w��t�%����j鞢�!����vN�T52S$��}5�"$��ke�&?��@)�a���G��������ڶ���E��AQ0����4�6voAzX������t�!��������L>A(� �:�Tb׿9��^ۢ ��������5l��BS�]dק&���{b�P��'��~d��T�MpX�d�W��x0y$�e�y<��~}�yS�>��3��c��a��Kl��5���	l?�}��ez�p�9����b	Y��i$��C��C�RY"1�I�G�f�9�6��?L|p P� Ay]�Q_�`��_�r}�ʰO�HSDV��|0��"&�kUڧU3�=Z8�m�i�U�:{&��^�>�������J�񺣲�Ph$߄	�`�!��nn�"�~��a�i���+f��#��
k��<+W4X#T��tP���hsM��Mp%ob�
�#7��t����RK"�F�>
�n�םm{4#N�!���9X�1�g\8��h%F�����2�S��ey�Fс����*7Ƥ��2��HE�K�;\�H�Y�^	�uj�(b/�U��#~�z�0��,~�%�hh�(�U=�kVY1����x�~Η���!�|\�,w)b)hgv��f�u�8�b����WOP��`���\�2c�ɞ)���\���g�a��^�7nv����Z��K3f�oi�
��Z��$�asۛ��,����A�7��y�]	f�U�U�,�{Ņ�U%�F��V�
�Kw�`0o��N�K��J�+���C���,�5�NP����Y�#]���x5��&-�<����y���xM���_���%;Y�/d�-!�y>z�kx�����k��yr�����]H@����$�q��OK��i�=|�Q��=�FFg��0Ƀ:�fL���G�lL5�:NI.�{Kg�u�+}�;c�6���q'�Mz}bD��&J0i��������P���\����Ze���L��F[j��rф��gly���85F�L�'@�����q'�یg62������)O[��]��f�@�`a#
O���MF�nW��˼�ω����m�і�|o���e��7�m���,�:&�dv��'�G섰JP��H���xY��T�5�-E�k��:F����FNMآ&Kk�dM�8�X�o,��Ԃ�16��<z"#a�-�4�u������s���?EuϚOTT9�@X��&�*D�uS�*�%�.�v���(͔�J�49C+]�O��)Y�l��_�p;���)ٹ�՛��H4�d��WU%��4��q �T̵�W���(��n��)�
���5�����F�A�� �D�Ξ����k`0 �vT�=�-ӵ��c ��2e0I.̚Jτ	�̮��SS��隥޷n�ߊ�dr4E���*|7�Y�mK�*[�"j��4&�h��Cǆ!rV[.۸b�:([����ѡ(��aI3o��*o�E��?X}b�ZG��JL��o/	��]��i�y����|�x�h�Z�G�����|���"���:M�����N"�|3/�m;׆����V�ub�@�u ��ָ���є�D�h��	lg�`A����fN�x�j_��tLJ4�v�2K(�PC(�;�o齱���B���a����=+��ہ���L��\;��jq���V(4�HHع(=K�o/WO�/�݃Z0ՖFQUS۰(�D����1D�^�o��l����&[��M�lI�4�*��	��W����~�x�
7#W��QO`��2� 
��i���I,3��YZ�_5����0���W�b2��`-���ѥ%���Zd1n��2���I�*�q2n�_N.S*�п� _�3�=o���[� n�oS�9�Ȍ�sӓ��3%���T\�K}��j�`v��Rֻ����>N��5��pY�	/r�[*�22��q�i��Ms2�o}ZǪ!��� V��#2 	�ۢ[m
�~�|v��r��b�5�L�,�Q>�Ph�����X�<��8�4m���n�޵��|��%���4i�np�u�O�y��g��T�7��͢c ��:����뼞��a�>�F���^��y�mw�mȕ]���m6 7|OҀ���gW����0)C�`��_��u������捹�Q0@4Y^�/�I"���TEE�������ҍ��hj��	I^Q��_��_���m�צR�W���+�ﱑ�F�-"7=�I2�!���a͇�S�n��̬�hm��`�6`���[�U��]f�3jXk XqL����]s���6CJ�n�.u7���ŕA���hN�b��a�[�嶞?P{�X,[7��E�T�/X��%�5�L�e�����K���ɖ�Y��U���@��B@�6c,tT6<�"���WR�K+��ɶr ?��|�4}�"�2�ܙi{+"� ~fL�F�E�G��{+5�u�A4����Ȁ����{jnY�*��~7=�� ���ukl�_��s�y�»+;:c�g����B��^CA��[���[:�G����X�=���z�^"�r,Y�}��*�!���yj����Y�JF��V�0	C����{�LFG��-�mvOn$��Ǣ6�	�7�����6�CD����|!]��8�fo��1�򊵒Л_=���d&:���g��g��ךn�>ȍf����	ӷ4�Λ����^�ّQ� t���>���bͳ�	�p��zy�g2��=������ۮ��5Ӽi����c/�L����|�������2��)>,]L���RR)��5����~�`�1CH�g�i�o@����vM�hk�&�W��!\�ɯ���d�H����$ɼ9��Ԍ	��`�x���DӱlP��hT��]���h6t"��*s�BI;P��1��@x�fj�B�9��7\-%=�s5m���C��q��X���娾>��q��"x-���_Vf��2����jQ.X�[D��:'}��n3�(�C�v�0-:�}!���*������D<���:8xC��:h��!�`�Y�\�T:�oh}��e��H���j���R�!�
ߺ͌#~�)MF��t�
\CI�:1�MZ�)��+1R���h�px0��%�Oӊ�Qeg�eH��i(�V�x,����p���3�\�P�=��q���-SZ�����rrs��PK8�A��R����c�wY)�[K��S�6迧8���Ƒ�6��*+����R��āX!�w�P�F����uL�o��=j�[���h}GY��"j��c)	|�Kt��"J���'�o�@.�P���Б�S�kx-6swO'�u�~e�Jޮ��Y.A�6���!)M�^�"V�&����*��{������R����r�<���s�I�kW�a��`{�i��ULt�E��g�R��O�i�0S��yZ�i�$E��j�f��Z?������ZPhqֹ���C$ɥ�m�*��|��u�r�6AB�Hb+4���� :�l84��w<��	��\Þ����w5/S?�׹5(x�\���4ǘ��d9�'6�N��9q`v"(?{Jǿ��mP�MG���]���P�Ϭ�j�UV���f���@�z��;s��	G����ߡT&8�ѡ����Kh��X��`o�"����C�5�g�è���:�#��T1�����aP4Nf����	�{�G�oڼ��dq����]�B�Y��&:nfğia6|�*��A�#�ѐ������M�'��L�����at�t!���!@��&��	6�k���m����aH�[�!h�a�!���Ĉss�٨|��C��zہ���Ƀ�"d��J0uz��]-�˻ĭ��8h`v�k�#������4��Q��r�C*�pm�*x�^�X�n`m�A$�;L�[G���S���@���L7p@#U���,;C�}:�c�!�"F�8��j| ��騠U�,�id�t�wc��w}1R�ES�JV�6:I�^.�} �ۀSo]~,Ƞҽ&��#���[���v�̂9����/0FK���U�p[qěY���N�VS �"R��O� ����з�\e�/�8�ǈw3�4>n���c�FLz��ьq�".E�*߃9E�
��%l���D��$9v�HHD��m��t��"6j}�7����<�f%�ji"�����$b���;cY�b:2�t�M͉KZ�p����V�("G ��ch��ʕ�zD��7S)��	�T��͐pz�:� 8�ҿ�^?�I�vF�R4��H(�?>産;w,��$d��]��&����\�Sx�����Э��:of0qY6'=8���Wu*�ȓ�Zӟ����&*��p��ꞓ��ϰJ��@m�~��>w�ܺS+�\���vho��n�f�6%z�n��G5ϩ�n�v{��Vj56�'��z�`�GU���:�ޚoNc p�Lӫ�٬U)/�o'��U��bub��G���xg
;Z�#�]R��L��q��^�`�6���*���.Mh��<�K�/qP�*��Õ����l`�DQ̺�f��ueM(J"7��P�1��CEC�F������ ��ڟm����X�Ƀ�U|I����{6�e���=.�N����b�w�ߕ�@o� 7�!��nZǃy��|�[��5�go���X�S��5���� !�V�Rw�+��_�D�C]C���vU�w=�<_�
E7jQ�4��ك1)?��.lV7^,ߗҎw�X�hBȴ)$�u�.^|Y�'Z �_��;�00C	�8�ˡqlo�^Y����?��C`����|@�˥�B8�;�:�vP����i%I�"�K	��ؑh<�[�<q#�]"d��j�h`���<��6��� �(�q�eF��T�2̸y�,ڐ��}��M$tJM� XKfF*7.�x1�Q����O0��}��B�W�o�b׍�{7�a�^}K����r�ey%�
?@����seu���l�cv�}?�8tr0�h���}��[�fL�_w���$�CHO��o �7C�a0`x�J�|~a#7��F�|�^mZ�F%��o1�(~�pC���h)_M����C%2�"ͲE�^��x^I����f��!7�Lr ���Mu[���@��[�J!��U�/j.�X"N =�C9P��ȉ�]�dш��|[�/�@MLb{��w�&�Sr��.�.#p���rM�s�bV0n��/P�[M,5mE��,��� �!!s�M�����p7D�x������-� �X� ]���(R%����\�b� ��]>�}�����.�'�<��U�6^!-�����q�JLq�u�o���z�.����d�	]�R�'�D^9���YQ���K��76@�-����UHj�i柟|2G.���������J�\.Ŏ.��W�M��AF4V�#^�"�+�n�Vs��� ȁ�#�o���e��Q������v��?�皪�b K�3�����d�~����˧���`����7k�e����+"moj�FްwN�c&9�3oSK��7�u��6��_,��ᴆw�AR;�������*1ʊe�@ΆQ�t�^�#��qD�f���Q9���:�a ��^�E�OX�������,�Oߕ�[,؛E�[�9��8��NX�[1��kR��:����V�䪛;���VX ������@��I������nq+�Y���������l����5:F�U�81���l`���w�-��JF���L
�%z2�:����iև��)���~�$}D��Mt$w��X���u����>o� �>�B�ے�:yN�s1F�'vwtkw��\5v����%���<9�	_�/?&0�����&T����[o#��*V�|��c�or���6�{e���u�?����4D��SNY���@�6Ԭ�q�- �d7���Gߏ�ڨ�M�#[>N�f$�?~ꆂ�Lp��]XޥpP�p���t���F32�o� �J.o�D�	�����567���}���he�=�`��6i2*��N����e��������&�=}��\b�{0�e�8���0j�i�5���)�=��;�(.tYݑ����Sf	�@��'�iw��V&X+�Lp̅��*|�k�52]���GZ�g�A�`X��?��<��kKu�i1�T˭?HJy<�h<���1���������$��%��"���[�3���I���%gG��̜Qi�q��L~�݇�{/�����f�Ø$܄��h��!DZZ�
�d
��w��1�"�dH�9aT�s��|��qj��>���Jh�v;&➭�u�;��WX1�B}���0���Љ	�����"��-9�#VN��jȉ,H�)A}
PcW�[��5����Mlj�S��f�"\��Es�u�n���)��0)�h2�c���tdĶ�3��)����\DCdz��0�Ÿ�@7���BȌӁ�uL�[�_�?�/�����#����R��e�փ�i6򦿃����ij�x��
�������=ly��P~��u�q��fA�-^�f�pw%ܶLP�� �w��nU5Al�g�}�︧T�P�9Ed(�O6�KĚ�F�0��I��E�b%wg��ˏ�BpXᢦjog�@Zs�Y��KAH	< 2Ї0�|����R�-��N��<�EJ��3���S�T�/��Q��R���?_1�r�����:�E�@ɷ�"h�|�����%O���}��p�ۯY��e$ԃ��}P�xbg�o
��5��m�?��y �z�y!�`7��u �g����љ��4l�m����y�7����<{�!o{q��㮄f���~�T��i��AMYւ疫m��.w�Oy$����M�	��W�� Ӕ?i�OYPf��c����U�����ğQf��I/'��g	���MWր��N�7��Z��N\,zo��@���"X���G2���4��0�$Z��B���e�bU+͒���-p�^�g���NZ�;���n�D����fh�}Q��k�	^��0���&:�L�Yűٔ�.rC��d�|�Q�(����-�ڄ-��M�w�f����ȑ�Ӽ��LI��Յ�׋������sK�}�eJ�o�b��b�WPA�YQ����&e��؃����|�%"�`^��J����1=��A�-��0���s����Լ�@�������_�!F@Oϐ�ܭ7��vjD���Z�)����T/ �#]SrӴ@�U��W�bP��N3fX�l'�ÜT�3+3;���Uԅ.��o�f�0��3`A�<6%vH\м�4��}��]!�����;�?��� @�/n�g�_�<�cQ�@��ݩȗD��2y��!�,9Q,��0�Q�;i7��]�o�-?�}5b��k�5G ��4.[zv87������oq�_!Έ�x�)#I�e��x�&�0�V[ņ1�Hg�C%'&���8=��O�G����ck*�)V�q�*���1& 	膐��z�N����r���.+d�c����Z* ]�������e�
��k��ZB��W����C��ln3`c�Fz�W~�c̀7���pw������.4�JO���Hyv*�7E1�+�f��zӃ�m�
�m"�7<��(&�$cꘔ@�	���F|�"�z,������ ("8'���2���a����3�M��V����ttx�qO�?�Q����3t��ʒ<Pp�d�"���7|l��+�f���6����*妣� b�)���f��~J�O������n!�;�䛲B�k��vY�0������[�)
�[E/���5醒9'�M��Y]�\L2�P� �:὾�K����E��jw����\ Wdb��'/��@�Q�z��%� B��� �m�趙шĊ�����.U��x�1�_�2�q�jD��S�/	֦��/N\s�a�=���/Eү�M*Х;CQdy��+?��
!f�<>JLr� 9����.�f��uIS��N.��*�֚��?�8&�,�yso�	����gF�t�E�xZ'�ޮ�*<����fSg'�ޥͱ�r=�e��?*�A��l�f��[\�:�5 ,>P`��v�Y�8=�@BfNŀ����u����XMR\Lp�!���KМlZ��Dc�B0�3�>9%���A{��H�A�� �{c؟6"��k�t9f�lS��1my�@	x�����nA�JVm,��e�,�q��e�싽��R�bY-;����E�R��t�6��?�F�o�5��	J��(��$ǌ�S����-�T���t����fLm��<�)��U���:7�神-Hd�%@��G�����\?���	(p��T�����)�p�5b�/���^� ��x���|O�OCƳ��,Ji|��
���tɳw����J�&��k���(r�+H�>�?q�ϻ6%������3��_6_���"�u ��c'��~ӊM1�):hdkO��9�z�u��!���V�TV���Kr�����a>�V��"9g��l�aD�u�@��&<ɑ>'�E�]Dߏ, ���3G�݄آ���u8U�?�e�ܶ����:����N//�&�&�)� mBo�ZUL�r��
��� ��7�c(������T�~(.�qE5^�5!�h�Mθ|�_^�h��k�x�lX#Z��(PM��<����-�������#䃋HP_�|A��_L}!���?�4yS6u�E"4>liK_�t�<��X�n�/"ȏ���~yq}l.׏�wc����oy�WE֖�AY�d�c'(J��H�/Tf�u�	ቂ���yo��휌~�	��1���Q�$$�O��m>&-Q�� FCR��H�^�Ǭ=�圭&=��f��A-VL�?�P�j]��螢�rT�H�*�[�&	0��]������՟D�����*G���r�����}r>v�l�C~��k �DC@�8�x=�����{�'-X(�X�ݴs`�ٸ��"���Nc�6(��VB?������Ŵy&�����Q���%��-�����C�B�ޮ�H�$I���/�>��`kDSY��z
1���0�p�_��N|��-};���.��Ć�1�#�7�f��b<�,
�pt�X/���pRMn"��kP)����G��&5���I���F�^xpܵ�W�vh��LV��������Q�%��&���(���<3$Fi�&���g��yf��������=�$�ձM𗬵����奯n0��B;�j	i�F��AQ�%p�\�clE}s7�� ��ur�[�t[S#r�����b�
�F�ߦ|m��@HH�F�F�x�Q����ws}�c�Ԙ)A��M���aT%͸6�v�fv-�!�%:j�]�����뷀k}�2)+��W{��丗8SV�?��hc\"�'��N�!�@V�
?�&(⩢��:����lbV2��Y��L�,��
���iK��y��X�C�K�W�U��S�@��D�)�T��E�8TW/�������k?)N�u�pY�]~��-c��qX��vO�a��l��>��b]�U�[��5C�B��1��.��Dm��8d8����	�NM��zypf��/�����<Ǘ�v�)W��m�p�P�y"ϼw���1�8(~��&ak���D�2<��!�z3�\�fu�PZ
���	u`��\)zQ���b �zmJ%�N{���&����p�h�e���#ݺ���9�a���΃�^����+�{U�p��F\��j˂~^�A���B�z�����V�^}Z�N���X���rn�5B��~�3:Z��h�gp����-9�ğ�Aƣ!���V��M�+�D��Cr�?'���h@d;���.+k�6�'���H�5 �+�
D��xD�%��������}�፾��+��N�x/N��7v4�rG�x�=��Z# �AЋ��I��7�ۼ�ܖs�;x)� T�i��:/������Ō��{����l���]����F���G��z1�U�!��k����s�K��x���~33������l��[�Hkȷ������`��y�#�q�t�Z4��L-4���P%���oð9'F{!�itܶ�Dm����s�J�/��
u���s�'u�R�l�����p��(5��x�"��:��5��^1l��u����}�*``�"#%(|����x?���@��Ele��͏Fq��.�PIҰ`v�c�Hg�	k�MQԑt�El����x*ZU4����m�wu�'��<�QK9v�E!]�/����c���)C��u0�����Uk!�i�a��5��/���=���#ތ�H:M�j�KG[qI^�5 �P���Ńl4���<�I��V7[5�E������=�f�f�5>HCf�fki[n���Y�t�����Sa�m��e(: Z��
�����x|y��!�
%!LSH�1�:l�p���e7�6�s�4�c."�qކvIN�U4=3�i�<��B|>*���n���đ-�_/�aL�a�4��ԳJQS��dr�-�=<�逕\˴�UdKd�8�=|��x�ȷ�H���X�<�1)���!{����;n��}0h � �Oڠ��f�3W��u�' k��R����3�&�[��/b�<̊x�$���vo�\�`��`��_]�d)/ �I�[��}�EY�Q�p��_�=Q?��WR�E�f��v1�~,-��7��wCogAq��u[kk3e�J:�w��p`Do~�*8T��(�Eu�~��}�/��������vV{�Ȏ����c�QiZ�����c�� ���Пuh��'��=�J��G�b��M�}Z��S��7���Y2?P���ef�Ӛ���Y����K�-���Am���x� �A�C��w�
�N���z��]5w�[h�E�o���t�i���\@t
f��o��`E���;�\��X��}�V��q��'R�VZȊhD��I��*+�(>�30f�� A�Z�!����)#��E;u#b|Kj�$v�,2Z"��5���3x�}��(]hd9��7��'X�pRZ����7H����*�z7:�Ft+��+��C}�X��s5a>,��.N�5�bV|�g��:�JB�Cӯ���5���_�,�s7��G�Y�-F��YBñ�d�r{���ͣlĎ����<Ⲝ �;��c�B?�:w�'PcFl7 nþ�e'zI{}� m�e�ѝ���Tc��*���b���U��"�*!ؼ�\f�P`�o;2*�]E}=%�`���$�,�b�h��bܷ��Q��=��]���8v�f���m���5�]Ĺ���kaQ�C�gq� ��q��T�;��Sx�Ggz��*l�X"sm�ޓ�U}���J����[I�����"�,Z�ct�?]s�>���iu�8��0�>�]0����9d�$b�	R�s�X�ԑ邏q~/�}lz&���{�J�MzJ��G��Q[J�Q�"�w��I-y��f.��r^�՝�j�h��Z�=����t�}�̟>��j���.��2d@Ys��T�	��ώ�#&�YhISu�˷U�)Y9�H7�r����_��ß�
�]������ʱX������L��M��^�i�z8F.�*r{�Q\�;�J�����F����G'���n%t@�16dk����%	��r�+���BF��	�V���Ξd#�4��邅�G�o&b��r����%�_N����A�M�qq��Vꑍ�x\��Wڬ���� XY^_?E�J��+u4�'"s�iM<���� P�d��ꋕ��ml�>S�-j���;��Ç�?�Ô��,�w�ԁ��{����L���^�RljWQ�ep#��v�	��l�$�uCH�?#Ў���Z�3b�1�"U�:Hr�%�M��_�i�Fg*��3ڪA�/i�XZ�g���}Б�Ph��Y��W�nn�k��Wڄ@q�l��(�Ǵ��^�������z�	K.�Y�H8>�nZR�ȅm�@�@A�6�Ћ�Ë���P7�aZ��0�a��jn�ho}�cA�B	�V��҅��C�Sٓv����rF;i���X�o��b�&��6����l�kMԦh���+=���uo=���?2`4_��TS��ۧ��C��ae:��c��V�Cɇ�v�È��t3� �5<q�K�upb7������awSvx�u�c�EX͙�#�Zc��0Vwi5�8���;�G��&\�݂9]U��ɍso|\�TR,w�GCa+����gژ:�Cv[@Bf2,���No� ,5�k$��}�v �|�.��@?�A�IN��au�F,>`��d-�2��s���.��XHp��26c;�oIֿ�h����^� ��Yc	j��7,�A���µ0w��L��P�C�C�l�1ן^6���%���h����r�h�q
;G^=p}(�M/��CX� ���x`\0����@������,�~f�=���++����c�i`L01w�C3m�6��0�޺��mQ%�4�D��r�U8�����+_˴8B�F)�>N�#ּ�<�9i�=�NH��U��Ͳ�-qj��2��Y��4(  �2b(ͼ:��7�h�mn����R���4,)I�5j���`ϩ׮��_��qA���աn���k�6*��I'}�J����\8�*^�`+�0	���A�%1��8s�O�ߋ�n_U�-�7�$�/��<`ZTG'WX�&��]Yе�&�Q��v�9��fv���Z�,�%�A�fwX|�;��d��o�?����{O�O�����
����,*�B����|jȌ�މG����Q�;u'Ȥ}O�YK�/@ GU5v�J��?�[PυM���Zw�'y-*p�v��og�7d_����e�q��,yv����x6�i3��3[�3k\�_��P[%C�����4̬�0bw�fCu_SOi�ZXl�����,aK��4/��S/l��Y{@~[=8\��V������vMuy79���'�����f���4�	X�Cђ+8�����)��+"(���T�&�<�3�*��V��i8���#��k._�?��Yw7O�S2�V�%��]�Ę���!�!���h}�/g�670�]�,P���B慎�1���ҧ�9*�`:_>g��DN�8� 0T4<x�T�-�|d��qxr���䇸��-g%�C���G/7�S&��}�̚��o���x����uk���#����~�����0�)%]0ң�))�А%9�{�
��| .�INϛ��Q� Bvje:%�0��W�rd��I	gАZxy;T<|6�7E�a�@�UA��iRV8[��
�U����r�%D��v�U�I�ܭ{Vq`/�m�3ni鞞`݄Q�c�ܮk�<ӟ0�56���_��G�G�e�p��H�ؒmd��c�fe�t��BvT��;������f�ԃ�3 ^qn4n�R�r��Y"�TX]���҂�ZD�ʿc�ߜ5�D�¡��t����//3��G��IAh�d��W��:�9�A�T�
�/nrL���� ���Wk�A�8�*�Ρo �;�M6:[LaR�tD�5YG�i!>%�!�:L������}���6<�֝0�{>�Z�����U�ҿ�
�/� c�زu�w�m%i���6#Ub�b*h��L����/LqSf�Y���Jj�[��ֲ�y�EtK{�6I\����X�6ս ����ҫ"�����m��Ts�3dY�6���	9����������Q���3"}�9�ӝc��}�&��P��ũ�X�{g���t���k&P�mu���[��``�����?rΘ� X�r-�0o/��I��9v�$gK4�;l����zf���NY=�y�(�����I���R/�B�,�8�r�,h<6�=#��se��n����B<��Wo���N��X��ĩ���̐~��Q������^���L!��RI�+�q��	�L�Q2W�!
��-��n+�F������"�17�aAظƔ��j��B��&��녠�RJ.�o۬/Ъm0D���O��E��C=P8:o����u3dCs�����-7a���!3�O{p�B�p8��́�vǑ��4x� ��&_D�?Vie��=hıY��'J��ѼW�{ҤL�z�ώ�J�ЮM�#�P����N���O���F3x��z�{���B#q�D��+۫�}J�z�KS�!v����#�Dj�v<��::���1aG�韞,[iQ�+	}<���� 3��#���	�=x�}��<�&:/�y��}�M�J<�Wf."$)�=�%�	�~�OD�o�W���3m@����Y�p���O��u��~7(�(�t�N������%�\�'�7C��,I�<Y�8�o� �n�gy��4�MlQ#@��&�:�v6���DX�~غ��~\X:][�z^F�T�:TT0Z�+��`7��F�,�[���k�m�yh��w$B/xy~�Ș�<2-�L-H-�e.����S:����Q͔D�&�8���C�  K��/1��ԫ�Qä���]�?�bR�k��g���N>^���|�D��a����|c�`>��Z�3��]'�߅�r��C�X+�r�e�G��ԄT�ë�,1sU�@ϬG�f�E@f����	@�ZF#�8A����=HjyS�^���V-|3��7�f�u��C�4��*��K��ߤŔ��?��-huL��%��G�*X�(�"g��wV?�`���H����H���,����w�A`j���mE=Ӗv�QŢI��%��&x��I7 U�@��������.%Ddѧ�R�R%u�/2����i)-!E3k0Lx
��ɋM_��pUO���Gb�Bw+��Y��J�wϮ� ׍�v|"n�ٷ+L�� b/����>;Z�e�V ex��a�nE.۲R�^��}"6�Xvͬ�U�9��L���dXа�hX�Z`���mb
����dG*^-M���S�}�E3�gڷص�=$m&�o��/�z%�w_�p�)=K *<p�����۲J���<Q����YQq_+?K̆�%]�Q.\�M��"�C(�w��M���F%��A�����&���	QISuc�Eea�����|�����OUvI�7"=���������`VόV>%��YP���y�g�Zg�PvT�t�����b�0v<�&`He�>.<YP�Эt��w���z$(|y�8�W
�n��z�*�b����>�;pm�48{�3���JQ�v��hok�k�?��`��p1S3
q䷔�K���IsG�H��B|h9Sn*����ʕσc�|���D��w�|K�����r�7#�>H�g<�Ar \�Α��3ZX/9ˉ|l/��E�xmYe\R�S7��aRu��SM�L���A��G�'.�J|��+Ǉ-(�!���B��cVCt�(���9m���xUӀ�0(0�eU����'S&g���'$2M̷p�-h�Ǻ�9#�@ �X�^�W�,;�����B��1p\T_d�U�e�N�r_�������f�=]͕I���i��d��%g���	dG�sr��TU�SH��wt�Út�-�PT96[��=�Ȁ���<�te2�7={sT +��/8?�*�t0�����g���
�'54�/�I�I���pg��F��g1j@�4I����l��;�����5rs�w�h�߆��P7S�)�P��p���[E�à͔�.�"d��9�v���z�o�Ğ*� �V ��R燛{p�TK�+�6�����T���MW�f�l��G�9�g�,\���u�'��b�Za5���{�U��&t[�F N�Mm�Ml����_�#�>���ߍv�R/� b��Z�|�����νi�(�#P�c~}��`�ɗ�����jﴄ�ٞ?�v�w����.G%f3�.bx^��Hv0(�+�����+3k��� k���1!c��1
Vp>�@�K��;�R�e��ۑ�*c|�������%��jZ�2]�A������p�P��a>�i�ک.�d�%�s�v�� +�?��]
)���pFw�H��P�\��؉���[^Z<X,5��Q�&� b,C5��[�*��.�|V���_����>����0�Jk0v�8a?�F������<��)V[i�����v�z2��*H;�]��".IЯ��d���Q
����p�^���N�.,�	�fY�	���t����a�WU0%�p�`
SO�(�
e���	��kǀ��i��9�� ?d��	mvJ��K�,��˲�Ú���"��R��$�Mt=��R3\���}�1��)?�I�v`�גr�#Rv�@�;��Ս݄T,�(�>����۹��2U��c�pH����dC�T��aM�~���]~t�+�����lx=�����[X/I�f�>��%�L�.��:�|�b �bOX�4k�>���1;.L)$=���oB��"m�F��?ݔ���8ŀpPR��k5n�;C�CZ9������D�۪̿5}ՈK�+fC	j��/��v h'��ya��%�c�k���M>����C�0�����F���<3��E������t�@z�!�(n�Ł���ӊ�.�����N�-Y��^�XD�{��D4�~^��9F�M��u�nE�������ʐH��
~��G:>�H�2L�mj��Ε�w+D��&1��`.�on	�����3���d���$��-<�eH��!^�)`�)*N�[~��w� Al�/�����a���m�sQ��6�[/k�'�
IH�+�|zo�H8���tAS����х��PCȁ1�KJ�B3�d� �5�:t�Am���X�����-����r	 ���U̇�Մ��v�c�jH(�yu𣕊 �H���f�c̋��a
���N�F{4x+���U�'ܵB��?�f��i��Dz��}g������ZF���9	��1'#s�@�p�~Ӟ�@�5N���f/���m���vP�H�3k7�:_S�9�	�̧J		�h�{C~�K����t��c6��4���z�]��/AF�!Ҕ�p�o�T����zS�#.Hކ�tN�ә�ȅ�"�	�
�S>����+~-{�A�R%���ε��-;k�⠜�(Z'�p�扦jAuZ���Jw�D%{L��+�u��c�od2#����́FC�	�@!87���(Cw|�R�����~%~ 	vi��+��BUp��Ɔ�|�D����$O��`�ok +� ����5�%�l-�/ǆMdD�~����o�?UJ�����:�hU#��Ч壯��=|Ni -�!�vw�� \��*m���9?B�B�9��>,�Լ6E@��C,�b�\	0�/��6 D�s�A���L��;�`r�*��1�:�0igKx�d_x�!�~�*	�ޏ�O��}�KX��i�&z� /��T���,
H��H���������5�|Jk����)ۗ�١nR�p���7�R��Rt]��)�}��1ޗ�ەW���������c�OlZ��|� �9��w��|%����oY�n��.U���(�]�2����8%���� 
��R�5��^7s"������a �vk�}"��J�Y��r�ҙ�N�A����= /z��͵��ގm�kN(�sp���]`��@�Tķp��o����>�r��r�	��կ��M�z�G۬�(����S��F�2g90�ѫŌ�&+���Ͳ�M)*���=�>��(IM|��J��ynצ�A�t��4��5+�� .�an�yo�\*����������7(�u���r-�()э�>�ګ~���C<u��vI��^#@F[c�>+��BQ®3����Ĺ<�y� �iB	�-��B3)�]�3������{	>�l����^M(�u+��v`C�|cp�'���U_��\�|��p��c2��N^@U6����_N����Q�e&���T��h=�4�k��F`|%
"6��G$dJ��Y�3k�'g�r�ez��C�K;ל(~݉K��PI���ے^H�k�|L�f҃Ax3�W6�H�?g�]��������#���(O#��yU���U7!h�P�g��������cn{pw�Hjv�+��y��RS�-�W�h�J��^��jE�G�C�E��/�¶�T:=�p��<��t�l���yuCz��bd�R�~��K��I��M	�"�U1ܟԩHrvۙzJ������Z�p�(�:0�R�`/�Q.�k�K���>����q���f�ޕ
e5��i� �J)��9�/���x��M�܊�
�S�)A��Uf�)0젩r�?���)���+ �9�2�U��bt�cm�5 ��k{7��/�ۻ���
O�C�1�I06��|`�����+W���5��j��u��z��S-o��UBW+��-x����S{k� &G�K���^�aq%���d)dt *�e�p�ä�g�b2�Z�9&/7I��)9a�ʝ7��M��tZ��s�Bx�n���|�$��[�Ӆv�74?!y�F�zߏ�	��E�o��A8�%����ɤ���*w<�"n6n
�Z�-�^v8\�B�q�%�������U*�{����N-ߘؑ��-k�~�����0���$r]��ɗo�����e��q9ß�V�HZ	�ndԍ^�pmqi-w�9DrFi���S� ZП��2���0-�����;g��)߰����,��P<�t�l�g-�K�96�R��Gt�k�� �ma�m��5>�iF�:7���SmВ����$F�׃6.�s�����I`.E��Jt��Y�#��V���mJs�	����B�r_ U;���v�FO�F>�v7��l���3^5�6���+:��_���*����.'�+㑝��I1J� � �%��*�W�ľ.5�Iҿ�ވ��nL����p@'ːG9V��\̈́A1����f!u��
t)�җ���ɧy���<�T���"��l�~��G v����|���`S��~��u10�b�*V(rX���3z,Sw�>;wZ�zF�:pұ��E��;�cBOx���aG[ 3�Td���:M��B�>��5#�@�
���N�w�MB�Υ�u>d.7��Pږ���st*��b�������
.��7�X�h��w�׽�I�K��L����\����HD{E(wn�F!���n��n#�����ʇĩ F�Us���;� U��*W�\%%�ni/�o�J˥Q��S��~���,��c�y�ƺ%a�i�օq�L^�Y_9y�U�aoב^�ڣe�3m,�U����ajV�	�Dt�I��saH���s~���Q	��ZG�m@�y��F��r�@�]N����(�y
k~"���9���@����d�(�=HE�i?*�l.<�@��v���gm�ܹ�x���Y(su:����U��kza}��
�<����pû^e�B#����Z*��H�&>��5�|�ww�G�-�9{c*������Lxr�|KI�1���&I3Շ���3aJƔ�M�<�E!�ϳ�CZ˲_
�������$�B��31�ihSp�<�����^)"Q��b��(�Y���֐ߋ��h�:�.��C��$�oN�G�1���|I6n���@��b��cu�����(��x��n�>X�p��ku�S�b9u��^H��WM�<al���S�2�^�8�	�1І5���W1�����O?�j�C� �O&Do�K�����[J^�]���|lM=��I�)$p2plzs)@�:�T�d.Yվ�&3� �y��(]�h�����K �_�0��zk5��'<ۃ$��Ǖ'T���O�f"ꋢ��w�݄�W+�Y@T�.Z�$S&}>���g���69��t��%$�)���-iX)1���/"�n�z^�U����(�e;{�Ă/�E�-}¢���gфt�-��9+*�T��]C90ř�M�J9L��T�H�顄�?����F�{�\�-�l{����MapV �2�����9���}`�N�}�9�}�5]΍��~5�,G��a_pqڑ����YWMM9��6�9&�R3�.^�9PwY��:T�bX�f^�_��J ���X��^��X.��7}�7ꓤ[���i�K����� ��o�hPN_N�l���t�YO�ܨG������v?�n�͆c��6�&[��+H�vw�	�M'�iZ��(�ҩU����ƣ9�����E�\�_�s����2�(r��{}��ޙ@Cm�9�h��nB4՞��d�Z�C�m��J��|�g���]����K]Z��Qfܒ��G����0�>X[�h�!WbUnD��z��a@����Ó�>&elz�[;��% �K��
:���յ���*B*q/}ݝ�]���a �(�[0��rjSA*Ն?�w� v�!a��4�618�(���U�� ��	���ې�̑-�2p|�㓙�me�LmLp�W������C�*߆в��,x��=� "�G�}��M��~4�i�P|J�-�b�K�(����7�sBaZ	za� ���|���u�,�(�x�P��qF-Vm߅?��kК(�,������%/)�
�
j�H�a,Kb$K�;�?�i�Vu��2�fFSdC)o5L���X��v��BG}�9�������xp���!�f_�Z���_�Ut�����Å�E�ԗ6oj9��f�=]�/��9m���t*H2��T��9�Q�x���� �@nnYս �5�К$D���O��b���������4��u[^���I"�.!�-w�����ܧ5E�%�ɹ�Wj��`�?�c���d�Q]��r��d�z�z��v���_��X/%�+۸�< Y>@�>j�nebd�I;;�«,H4,q<�l>�-@Ѻn|s�l׃��M/5��>_'Z3KF�`T�h�����[�U���pc���5���!�đ�Y#tc������t�9�-Y2P��d�����:�b���56�w�v�: �9�8����PƃƏ�47���%��a�RqM�~���;@�+2�Z�.6U�&�I�2G ���d�v�9/�FX��4N�qlJ=��	)%�h��N=��u�0m�~#/K��$ۊ��F^�����)����1��:&[��:�t~'��� �j�
�ox��	K^��g.f�_3P,U�a6L��.rJ��S�S��� _��	J��uAT�L���{��l,!�s@'��}�F����������嫿�KLR>H]n�l!A %P��/��jAve�"$�����Ý�ݟ���c��V����G�����C��s�,�i�c�B��z��VzS�����A�2x!,ׂ$�z���1"�zǄ=k����2l��ȿͣ��l�E=WV�DW}z���F�v`�Yn��pa��wD���D��J*���8��^�=�6��|_0J8W���R�#����*D߷u�)8@�7W����y��^���.���=��yF�!����^o�H��Y
/�E%��(k���	�f��D�V�E�zMA����K2�C�pB��r`1�n�ڰ{��y���M{I���ꬱ��+/�ơ�V�ή�u��?7+q6q�LWx@K��Ǵ��K�m�ʆ��0�$0��`A~���s�F��}���N���ٽ�����w�V��>4;��C�>�Xo1d�Z6�t��� ���#��P
s)SQ�ڗh=������׹�w�.o[�>G�^�Ds�?��)���X<�q����>�~�� ˏ�����yT~>gq�a1���ʩѾ䭩�N�
ʹXNIǙh�ΧX��������K9� |���9�ŽO��*�7�H�!s( �i��f�J�"\+�AN�v�5�������$�,�ۖ\��I����5�P�`'��k=�<Bqk/�b��Sq����g��}s�'S��}���_T�P2���x��6P��;��\eK�J=O4��yR�/b���&@��F�[�i+��! ϝ��u|;ĸ�t�&��a>�t�i�$���/&����0������j�fQ�s;���s�����
�WO�����؆,c���[�������s�oȄ�Y�����4!Z��`'|�{��Uv݂����Kbp��2���U��к���0�Y7�n��T�1���ĭoD��>łj-�x&�C�iI�_q��s-Zjn,��y 3���O�`��q�:՚��ӯ�?�:��WI���y��M�W�a��jx�.As�����C�y]{'�+Ql���KWz~�h�D������MQԥx��g�^\'%Bn�ً�
���.,"�p�:2d��P���v%�sD��T��� ���yxx|�3�r�BA�im��4� kb_o� �um�4��N�T�=�1�@�L�����_, �$y�X�:b�~|�l����᳙y�
�˥�q�_�C=y&��t�-��n��)��rvl�0�y$K�������`�FӌmcN��Ѣ�@O�
[�YQ~t0�+ۅ�b��SUmv�c�xX�^{d���v���#)�.��9��� $�����3��g>EfY�JW�!F��������+)4̾�r�b7��a�}=So���̦�62�`��Yt�~��è&�:q�fq�k%�Z�&w�n��EŐ�������F�)��4\��"��}md*7Hއ�o�����>������W��)�\�~���B$[`9�|ӳ	#3T��R�}�D�X3Z��O?�p�t
3+���M��&��TxI @�_���5�9q!�þd[7Tb�p|�	!T��\X�[�r�ȁ�'�q�0�x�Ix�2�C�BC��	�*�6sE��ws�'��}�N��!�B�O�?��_���dl��
���d���-��߱�f�0�`��o���Ӂ��X�r�;l��o�V�)�ѪppA;i��� ,�?!_@5ab���A��J�k�r5?����.H޹8%Y���O��T�h��������~о�>�,�ua7Hvg�!�*f�-Äo	Ki�>�_ U�S-	c��#v����8�@o�W߯@sގm�D�_y���E �3c�9��).V~���ڡ9w]�!&�	V�: �`��U�*���U�aY ��d���0B&n�e�Xʿ$y����w�n�J4f��p������ڜ���Pe���8�iE�0��#��D��v&�C�%��A�k��&�@t|��k4��>��������^�<\�a�9̫�����>}I�u1����B�������[��G��;\�内Di�g�~ה�7Q!o��o�HתE=3���:�vp����zg�Y�k�.X����ú9
�RQu?�����oɅa�Uv̰;��y ���O=Y�x8����]����y'k<��U�,�|�ټ-��rI5������iS�:r�urԽ_�á`'�Y���S��qX�����!>�䮱��eEC)ĝ��k4�Ӳ����E�P��>ю�|YGlARI�m���9����ϱy,������k��S��a@��r�k����	S�O+j����A�d��@=����Q��9��j���O
@��9ĄݬfVރ��
6��k�Ep�*TO'����*W�1Yڽ���3�9f�R�/�����ygY�E���� K��vM������7e�m!�O�	 B�������<��"�I�i0�Dݕ����[��a��2�l�*9��T���C��6�ѿ�����'�����y�t�H[�鵊H�p�d01��G-�T���	��U�
�/W�!�����+�ͻ	R���d#��jjG 3"	���T@u+ӦoBx��%�S��\ 1�!z�A�ŻHnj�vg�  ����\C���a_�A���̊-����_���S:�Xf���ւ��4������I��;)t�#���/y���Ϥ	��Sy轑�R�sD�q�i+gɾ��I0d��{J�t��_>� GO��%�+\؂`v�m��Z2ۋY'����_�������sQ�ꄺ�*����� ���~~���{��GߨD�N3��/�*�U�#Bb���[��&v�:�X�"m�^��S՘�~+�a,"�2PZ�!Y�h`NZ���5�Q�K	� 3�謡[� ��	/f�	��{X��{�>K�"A9JU.�?�~L@"���3C��Rc���K:	,���?�Xm Pڤ<|�A���ݡb���;�5����K�\%�5��|�ܹAҚiL�8�r%&\����1w�?i�z��U|`j�Z����߯�`�� �1H�O	�*���ۀT��vK(k�'�q���Ή
�^�$H������0�*ɸ��N#f�:p�-���~6�|�ׯ#^� ��� ���s��;���%s��p�X��+��̀��٢�]����B'�����풖;��� �ű2�X2�pN������&��zs
��S��UTbA��7"!k�n�@8]4"զc��r_?��d3�*�W]����1�D�!����[�A�{C[{(9bx��\3��s3|���#�[��-��Eԩ��
k�:X�5��#2�_Z��z��)P���^�W=wr����?�=f���e�7��%.�]���;[����L�t�c�c|v���!�d�˻������a!���y�D�7cxE�_��v�HCFwu���������_�^�U�ѶԳ���2��%���G���[��}���>��J�l��xj#�a�P�N���{zʭ��ؒ|��26�"?r��yu�������5f�~�z̓1gS�"UR9�&�T4c#*h�Is⊷��nRN:zaf�g�@����c�1�tNt�v� m�ꖓu�2������p���Ɩ�Y����Aư[�M�&�.�V������zf�h#:�K��{Ixh��;�0M�l\�ܗ]A�����Č�[z��k��S���.)�XG��VV�H>M�0U)ET��� �?џ�Wϧ$"�ͼH�mC�2�g��O~t�`���l�6��8ؠ\�][��~PD[�!B�Bp���nW}3���I�>o��&��E��`�����V�C@�G������j�mQe@�th��{�L>��$`$��m�����Mk#?���-��K�ݷVْ�r��3~�i>��~�I�14�z��h�VA�&b�X� ˨N�.��+���M�'i���L���M��W�J�H+�Q�O.�T��켕Sw��^��4����tc_� �p�{�%@�jj�N�7�*��.1_������*�.�C{���N[��GjR��K�v��+�?Y�YF�@h�0��-��l��C\�"<��)�3�O�;'�~����&~#H����_X@	���+�|�n��������5��U�=d���������U7%K&D7hŭD�-z�A�Y�:�b0�V���f���3�hj{c�1�,�Ĝ:n{���ܱx�㽆Cwv��@W&�s��{ޘ��L�.Y�N�����l��k��7RR��e�΃y��S�~�����X 	ņJWuBU=�Ң|q6�aR���5()@��g��aB�����jҕ�Ӊ��v
� )����x�YRI�#9 ����Uz?�Å�`�+&.j��`����p�?�^S�7��M�-^8Ұ���.v�fj�:�¦R'��\�l�A���+�5H�����V({���d�,�]�q*����y�=RCe������y%��~X�ຣ��].��F�6�1���/�/�u9�j���M�B'��R�-E����p�:����J�������'��l4�Z?���Wb"��	�Rw�3N�\�ޏ�+",�>ف��d&fA��|~���
y^��	Сy�;�6��T�AS�Z:W�m�S�`a��j������z|���A�_yﵣ��N�=j-���h��ët�#�N*�y�8Ī�.Dn[���t���'-l��$n��-�%�=����n�s9Umb�A�#��[�ar�ݴb�fD�.����_�'㑉���B�F7X�F��X�/ǣԥ4�W߉�++nx M^�W���J�e��&޴,���N<��Ί䑥����5�q	ޞ���S������s%/��2�E�ư��K���4T�9���sBW1�,��.C�^O9�n8��li�"�����7 6�7���q���.e�1)<�KN~���������L��n]%#����'���nX��~dsp�f~tHK�����]
�Mg�Z�pBE�<��)�)yFh�)h�
�:&�߸ѫ��8�������F���a��* �Q�T�ʌ835�U�U������u\	ɋ�f(բ�Q_�!��]ZB
W��A��Y	��q�/��jzN/v)���}Z��)P�� �xM��a�G���ɸ\�GO��oQ�����"W"{e�ή����W�hB�?�\&�g!Z��}��'��;xBV�9�"�B�W��!':�������P�g��0���w�ܲƎ��ka�j\	�u�3m����3 �x^m�����=��]>���-�Y}�=_+�"��r�[�Ů֔�qc[�+d�[m�0 �������J^�4&7�u�ף`�N�C��0߼��"�EgE�����9۵�;!����
<�QR�G�/;=�>g�3�"[ �L'/i�D�3`�\Y��SXY5�C���ܑ� �¾�B�.I��kn��������4)�RDr�f�N"��nāA�  �e
�Y��
���l��G� �5t0�M�a��a�n�����+��0;`����;���v���KC[���s[$ˋ�}�{˭��fm�6���w�J���O��_zfb{��J2Q�U�s�O�i��b�M�;j#L�FV�bEZ��t �S ��Y}������S�x�u�7�W�֖@���؝��+�p|+<�q1���M}>�bK"r�R�^���Bc���x6E��D�C�ݚ|Ζ�~���΂��O`��{��$�r
�Vѩ��X:%6�c��4�3t��_���G�mڟ_�,�6�"^����5�K�Xʎ[%��İέYu"h	H�x�q��a.�F	�6�lx���/�ӷ̋nHuގFiZ;�9��Z�(�rԊ)d�2�>'�������\FKh+��Io�w"+1ĆS���n{�7�/t��py�3����?�V��/�#8�����8�m�&����}�U}�g� ����|�o"2��][��������ռ��^��z�M-1)�Ҳ��w�FL $ǆذ[�"+˂��j�0�A���0��a�:�*�۷��l�v�'_��K�!S)�D7R|���y�8�>���3�C�Z�8�k1y�p#8g:��\C��MR�o�Q���*6;q4�Ԛ�~���V����@���� ��KN����N5��O+�e�ϙ�*0G�37ޟ:�#�i��׮�F,�6�^�����TxE��7�EzPT����Vc�C&��9��F��NhN�^X���$DK6Ę�� ��c"�F	4(�����sg��Ix�4ʦ���\&�;UƓX�"��:�22*��e6\�g�y;�<�Æ�^���I��+�'��񷰀��� ��ӛ��L�OJ2S�_z�b&�UK�+��0$��k�ȵ_L�*2�IP��x��/�7�(+�WֲZdN3�p�j��5�`�6~jN��8.��M�Z
��d�IK�lO�j��qQ=� C��e���b0o�M2#K]�5�nLY�1$%}@'��qS�HP�j�V~�z<v)�SP���?�Z�|�˯\û��@EDοo� ����V����+���G!��:�,~��\��/����FF����J���i-���g�S܇#��3q�`o16[����>�g�'�v��͹风:C��~�0��FF�29z��)3�?5x��J�0��\�Ȱ������^2Q���SM�C��
Ҟ6�/_�P$�� b³��Y�#���)�o�?<=&�,���s�iUP4yF���o�ݯz$U�j��M�kl+&Ph�]Y���Nԩ�N��P3�Z�6�Qh<'Ʊש��s}ܫNr���O��H�fI��FX�0Ew�8�ZKOOƈї���O�u^aF,Y4U���5��3m&I���B,g\��.)-V(��·ly��(�)�W~��o݌�¯&!$�cʱ`H8p�SDgcؤ�����lː��G�q+l���t���F�#�s�ĠI%��O�jrg�
��G� #*$I�<�����@l�9�g��s�I�Q���ԟ��[g��<���P7����$����(��й�� J��=�ȏݒMJ �稨�sJ�w�*�н3���kL���֏���	R���U�	�� �0���(xs/��,EŘ��,`�o� h��V#}y>�>5����Ӭ{�Ƃ3��*^[T�r�>o^$#6d�Ϲ58�L��p�s|i���1��Ǆ`�d�x�E�GY<���r_�� ���f}��W�ñ�ˑI.�1¬��;�۽4�6z��,�}5Q~f
��{z8<��vd�����_\ f,@����~uU��!W�->�}�7ja)�3��l�z0%3��i�O�]{_�)#y�!�1���\��@�]Ύ���D�����H=������
`P�O9���?�]�G��K� U�**S0Ny���ek��� �ՐCf�)Ï�Ic�KO����#��Ji�m��G����@v��BH�L��mP�p�MpW����74m0|=�vQsaq}�م���sf���Q0"+�`K��̒/׸9������f 
�`�t��q�I-�$8z�B{q栴�A�
�k��أܛ��f�mP:��l�-���݋9]�!�=���Oo��x���h]*K�G �fv��;���Y&�s|+���-:���.��,qM� �<�K|�#/��i��oGk�{�Զ�@����!ۮ�H�5��n
 ��+����ז�V�+�3L. ª���(�6��Ϝ�S��,�vN�O�51���_x�����P={lg�)&�j,nsg�Z�S��}H�(N�����N@4��S�9z0���+Q|�o="�I�d )xY��'�z7'���� �w������x��W�l�,�Į�T����ke��V����9U�k�/r.���p��FD����6�=}�Z �P���:&{�>�	��:h�	ʼ� o��/�G�mɵ�̈́��E�뿚�x�/j��D����TAS!��.�i,����j��Ղ?�c�	���3���{U��_=<+kT���it5��N2�e�$�1���2E��qRI���������D�C��.zg����~Fr$��;���>bU�e��\�����C0C���/F}|�PNhG�fP*�ɞ��FJ��L	X��F"CayG���=j'M����ۺ��_�>w�HDl�2����{���gs�D���X�@�	�3��p����46^{�Ơ�*	���e��9��sY�T�O�=�d�O(Β�aqܿ�6�0��Y�cA�h�?�(��j+�C[v��%rP��V(�u�����,s���F������;��d�lJƲ@� �\����-�P�'��}`�_�抧XL��0��fE0��w�)si�W��� V,c��9��6N�Z_������NHo���FJ����:3�k�(�`N�N���������%`fo���[+@���i�$�������fR-�6.�I��tk�n��I&ŕ�D�:Ε��������J=t�q,�(��MI�)��mF���畠/�D/�j�,jn������_ϡ� �-͋Օ[�4�w��������HG�~����Y�M�2�L��yR����1�5[_�;ܠ3%(e܈��SE_�6>���m�p��_-�$|[w��E����	�u	�]�]q��v��ou֘�9m6�4�H\�7��+��{��I�]<����"��p@�7���@����^e��4��r�z�X#~��<<�;�͔jVtK�d��P����3������#[��	v1Џ<b$ ���:�*w��Ӄ	�%��+��c� ��=.�jy�/���/q���3�Ij��1��	y�cٌIH���ٓ+`5%S�|	��tBx��s5J��wHM��3������ՠ�!�J�;��M#�eȜ��,4ed���C��^�<�ڽ��t��F��!Z�h��~[�]н��ȼmM~�uq��t96����i��;��y�0U4�$F��
[��煘�$�*"�P������$1\{`1^�]k���#�d.��1��9YF�KŞW�]c+v�y��!p�t�$�_p5D�������ggj&(�M�b]īB�@�VR�`J0 �[�E�E� f�6��� �{�hr�^_���Dbkݰ�t�?��{��f?�a�ʿ(�d��U��z�|�$�ŏ�ܯ�]7۔��Dr��Q"�S\�0�1.�T�Y�~6cߊ_���
 �($f<V��9���H�T��b���c�r�����P�0_��m��c�g#����ˮ��!F�sV�h0�l�${�|�,t���n|�4,�\\/���?�u�絡[��a
�@"��a"��2��Č�d*�c�5b��Jn�1�O�ya:9�"�۳G�J�:)������/,�\������f%i$�M��XG���(�Tś��m�9�+��=��pi�|S�:Թq8)�[	��VP�U�����Q�R��{�<��O\����l]_��n;z�50��=^j7~[�� ����XcN�V�#L/�U��ѿH���@�ʖ��s~�>�
�a+��u�����Uػ��]�L��D�"��sN�;<SA�T?S�P ��4��w��뫦M���
���P�5�4��+Oc�i?4�o-=�9�|�#����:BF<�Iݧ��d�}pl�'��:v�ts0�1y9z�C?�����dL\�'l�}�E�uR�B�n{=i��J��%�6g9LW�\�i"x,f���l�S|!���2;��ߧ�c�(A7hN�c�k��'m��蛋S��h*���b!0��
��R��̾r2�	��=>�RyT�t4�^�Q�̣�8�C}�/���&�y��w����A��z�j:���]�0[b�9���h¬s{Էu��L��6r���+�������?��P�|�����U6X9f�@����lD�Y6ܓ�7�8��-N4�TN�Vմx���vp�,���X���z��o<�@:W���IJ�^	�G�a���X�T6fnK�H��� >jO4&���߈�������` ���4w6>vc�ݏm�$EB)�7�JЛ�S�-q��T���a��^���ɱ�����YKĈ:�Z�f>qh�JP8�)���R�ͬL�R܀�� �@.�BE�s��焳�c��s������E�h�i����:�b�/oMR�yS��� O�|�1 ���A�l��V���jɩ\0���Џ������h,�d�[�R���26����t֫��ÚAE�S��O���[�`p�z��kmH;@��D���8������3Z�Gs2��8s�N.,4�p�"�+����MH)�� zf+�#��P,F�D��=���������jX�6�6�C��_��B���Ns�=ar)��Y%�֓f�i�@�2ϧƂ�2�Ce �"�2��$z���X2�*���f���%�����i5rZ��yػ�ׂI��/Q��鹾Å����L�Zb]X���ؒ��U�V�~�{7,^�+��Y\ѓ�4��ޱB�W�A�,h2�����E!7�nZ_ŉ������f[_�\�%ڣ��9��0֘�}M�l#�^<�jE��~�r7r�:o�4��%�P|��'#�nG��!���0H5B�<�W�'C$��� >ul��T21N�T	z䔷d�����V�'��[9%3�pҜ�E7$���+ˇ:J�����6�:#��SN������r�.X���m2?��j�Fi0wO1�F}:�Ɉ�h�G���78bM��0>Έ�l7~�VMJ��mCYk���>D0�e<q&XpOp'���K�?9F0���ݵ���Jd}O�u#���!�C�7�J�E3��Z�e�h]�&!�[��cw,訾W��N*Т]5i6�W�z�U�J_�h�K�-������c��d�kǴ1����|̙������*�+*��M5�ge�U�)O���3�����d�VT�_�-��T�g��o����,y���"�Kܰ��W/�T�*���ώ��<�6	R:#@H�����H��!iɥZ��.0C��]�o;F�?�jh��yߥ��h��<X��t�?z��֔��?������e�<dcCmV3K&�'yLԘУ������zA�tmi�|t`���$D��e�\�� 4�b���Kq�ȋ'���w<�H�"`�Oظ���oAO�3���B.� �֒���1�[؎��U7�݀e_$x1��)/����Ga���Ш��fL�܌&����p)��>,R� ?r=�vp���	 �M���	Vd]bs�?(�s��Vd�B(K&U�[	<��p�N�_˥Z�60���Y�%�gH�����@�7u��Hy�����R]׵�Z@ǒJ:{c�S��F�� Z��H���,�x������F���*����ڀ 4X�$'��֪�Ik������o�0�k���o�����T�A���ƦcOD�b���<�~�Y�I�����T����=��g>�1o:��[ĵ�O�]��M��!7d�X��C@i;���I?�f��S�oِ/<v���f�3���~�h�G>�$<]>�P�(䎂�kg)'Ԁ�hW`��r�J��10T��H���#�f�)�R.oa^���t�'���2�c�M���l�-a�D�T��x꽜5��C��_ʨ���m��j��>�V�'�~q�1����X�V=q{,��/^}��B������\�^|x�)�L��Tm2�p�w��3�˖���x��ɦ� V�}�M�2;� �6ٟ�;�G�HoALt�pb����o#����z���m�#��p%��8��K"�xo2�LJ�i�u�N-��D����y9mN�80sp�@,�5��C��^F���P�ܨv�ŧ&лP,hl@��Bg3���VZW����>��X�t\.vg�Yl�˟ș��qQ�|���juR\T(U�_$$�&V�ϤpKu!E�^��C�H�\�X?槟C ���k���$��7F��%.x�U]�?�-��k�#G�z��U^��Q�����`(�nze>Z����&_��=0�wXS;|����֗�� R�c���'��f5M��!/�*0ԩt+/�o� TXh��6���.ސ�(5�>��d�ӥqD7���0�tzMn�����w͉��{�6��ε}NxI�d�')hR x�v��q 79�% `Ơ���S)�/ZY�1IJQ�?%R!HI8Y:�����y�g�n�V��F(�j�ح	�m5�8��	�xdU�z���5��Z�sTFn�
�y��n �$�%��ƍ5�݊kɧ���ت8l�8�&����T2�p��V�������ΤZj-�;Y�w��)�0��nd���X�����f���iob�6�,����������c)��g~�Uh������v�_D���@�N��搔2�j���=e��^�e"�T��Zv���$���>����`�<$�$J��1�^���?ZS���U)*�������������6���>����j�KE�!��`�D3��u����Eh�%T�|d�G���h��e�~���icE�����RX��,��O:{��!T��J��, K� ��I�s�����|�5��%L�Jj�1������EJ&a�}����,������U�)[��+}ݳ,K�$Vb�e2Iҽ�Rn�Yp���un���9A?�t^'hau L��S�&)�Yh������5ο�蝗^�{fr+Zs+_"Hkm�s�k?_O;�"i&$gv���F���k&/�b���"�71Q�i|Ń���3%�~j�Tʾ��Z����q^�C�,|bI������C�RO�¡�HŞ����
�M|8�'�߅�?ƿ1&bRv܆��e:�~+𑖄�ª̈́�TXʌ0��rx+И�ԩ�zb�n�8�����e�%{�W&� 1�0�������(38�ڷ��<NnG5%��e��cH�c���δ�*|n�D�4,vi�3!��m짨@���:��~��]�*m����$n0a�W*C��N(�C6}����OkE5�2��\],L��=/���V�Nd����WY��m:)Z�:t���a�Lj\COe$C�;_@j��ؔא�9OΓ,����se<��z �;��ۿV�&R��h���D�%]OI�3wŁ���M��9{���碇	ע����Rc�`���
[󔈮'5|P:�����d���7�P+!��?��jj���"�eo��č�`�@����e4�����`��Q1կ��Ǳ(�;�o�+b���jG�w�c�A鉩&.�Qv>f��1�(���!՝�0�5:�$*odh]�S��4��E8���hn�
@9�]-P�v �<�H픰�PN���|d|��d��O�O$�d���2wR�a��!Ԍov�N�s�xw09�n��"d�R&�$j8�H�oK|<�����u��e�΢̒�;��K!�
)M�� �ia>X&���J%w�=�����)�F|oJ��(5itD��ߑV�|OjI�� <�͖�h��*y�����o%O�G��Y���q�r�Q-ˇ�
���4��3\�9?ҡ�Ǌ���rX�b�}��[_;o�����L��A�}�¥�D����u!�!�.�%O���b��{��!hZ641�r����^�1���ʿ�s��%�i�%|�m"�"%��<�;鼶�'{�
�}潕+�R�0�7ik�Ǧ
]�ЙW�~��,e�rK�GK�����|���@���[Gi����'8e���S{�f�k
V���V`�;��!d������wX�|����oY��Oi��*.P�wW�����E�2��Mo��9GcA������R�!j�ş_���a5�D/V�<g�?�c��g!��(Ax:ã��e�XX���T��J+��Q*L�:�	Xy�ħ�M�Nm�`౔�O!��VK�s/%���M�y�i�F�Վ���c7ײ ��]lLj��Θ�Vq#���(c��x�s{�y-�ڂ%c��]��{�n5���uYp��d�y�s��f��ز�P!\B8�H'��+J����h��I�@L!U�}��J�ˬ�#��J��\��W���?���y�g��>ؖ�G��������9L��y���?>�N�I�>���ř�R�]��l��쮌	�)Q�4���o�s��۶,dM�Hߩ9m��)�<�)���}��u��p.�|(�)��8w�,�#��pͳʋ���yQ-�oҁ,���k�>\ǰZ����Sʭ�J�Dg�\3�-��g|V��f8���y���7uT�j��E�vN,2��[o� ��1^Q�-�A��?�\��]{ ��kAE	�B��2y��)m�� ��M�{��3�XUK��e8�Y�6��&/s0��gX�x��g4 ꢌI|wM�7������}�t�����C�������n.*�I��f��G��u��΍?��}^�@���?������5pT�]Z�K�/̀/�]��,����V�xp�F��3�\� a��z�1�QF�PF�;u�Јx-7����d�.��!K�{p�^��I'��g˲_Uer�#����<���:M��K� ����e�b�e]��	�#��d�g��5-�M��p)L��������[H�H�:O�_�举/)$D�8��]H��!,7@��D��L�~|����{W�( Ѐk}a�1�%3�	j/"���#����Mڅ�>M�A�HX�k�Ú�tT�]*�.4hk.�]o):�2Ѐ�q0���Ы$��ͥ}]�+��m�Ȟ�|G�R:�6	\���%���>�-�8e��O�G��O�/���M%\f��b)/�ʿf�HfsY�;许���w�*Z�!>��չ{�(��.)ƮXƧAeؾ��FZ}��d��vEP��6�R���n�At�'�%����rᚅ�:�9��q�D�^�������������{�Z�/Bj/��e�R���e�;(ä��¡�ݿ�oƕp��X,�ӡs}��q\Y{�&h�_�~($�
H(�i4�o�~%a8����pd��Te�#��M }�W�#��K�d{s9#�Vո��
f%���p��Wo�w,$O��k��DB%ԅ��[�^j.��}��ζ$3tuEƗ�ǣf�|�ox!� r���$��F,�>6��)�0��1w�
��_��G
���LE��������`��B��urj(�X��#��*��ŝ"�\�K���:����W����	�3�\Q1�sSM��E�6�����	��l����}*":c����5�(��}��u��sz�.� �Xܙ�"���t\U�d�\Ga����|渟D
��L21������&ղ���
�Kӗ
�TW{��@���蘃�{
XE�=s33xim4{G���-����YC�|��F}���� �ŀ	�L��}���k���	�ct,g&{���E����{�&9pH���3I��d�ew9��M�)���4��o����n73��vXv��>�)|�^:�9�[].��f).��+��3�u��髯�:f�=T\�8�&��+�(n:�I|�sOT����x�ŗ$Ǜ+S�/�.����7o6V���N��i���L�^!H�刿��CL�a3�	8�O	�'�D3��t�&�� Vz̩f1�Y���k1�݉G��ijTT���>��2" ��ݏ��^�����Wg Sď,�x����hNn����vFz7j|���ZH�������WD-~<;�׊��G8�]��+�o���6+'�(�O���Fr3%OQ�L�}Р�9�<u��Ũ9�����rn�`4#�!�C�Y��}�����[�[��7���KWX�D�h�Q��w�m�����u���)��=}��e�+�����	k�0��褘5ְז�X��q�]S��;잝��3�Z���P�T�uݠp������1(�<f�'%��k��{֨R���^2u����p�m��R�� k��&���a(�+�"="��~Xn����H�� �g�6�'4T���$���Sˎ��h;��G�5�CU�J����G�Β;�B)��B��7f%m�p��z��4cH�1ʲ#�'9�s��4ي�Q��(����9L"1k_tb��gŖ�_c��;Ey��Ʌ)\��9{,�2L����ϽXĻ�QBE�Pɓ؝ ��&�U\F�L"��E�u�&=aS�����m����V(���#;ʹ���=�� �
u�W�S�qfJ�j����Z�?5�_��� Z�����M��\K���}�Q �Q�M
%���y��b��U8u"=)";Nn}B��4��h��KZI.!�@]�s6LߨD~��9ۋ�˓Ye,�����g.ga����6u�(��B"?���)�֐Jd���+I˰�o[�� T^�G�i0u�;*P��_ �Z��
�L:z�n�M��"D����u[�����QQ��&ֆw?]) K�d#SC��H��C;�n�t� �ЌA7�^��>�=����6�p�5p/��s����cCI.�ra��&�
#bɎ:5�־G������z��XswX�b�J�$~/]:_X��uS71{�s\IZGo:W����%�iv�u>�b�RT0��2�1$i����)�Y,#��Aه�du#%e2	EW�R'���kJ�7�T���*�#k$�fYX�i4U��5$ѣ\<��gg\�� ��5�M���C/�r?����%��:�����o��}���O���l�֯�L�X��R[��?�z�%��x�ʗ����M@j�"r�������L��x"���:��������_j�l�yg�3��h�C��3#<�ҲCR[��t��2Xd-�M��n>�ԋf
�3g�e'"\�f6�����X^�7��6HM�W�r�y&��-~�؋��fՅ?9���K*���
��t�v6�W��%~�� <�C���MyX�^�oB��.�'�#w�x�0r�vj�ȧ�7F@@�<z���?U!PR�hΉL�X�����v=�m�L�	`:��ygu��M�����C�5���|Ŕ8���Շ��ޚ:dt�x��X�]?�P8���-%v�ԡV�p�z�u����	^y��1���!j�Z�V�$�s]�Vip�7kB��}���oT�/�7a/�.�sY;\�Yl���@�!)���P�¯~3��S.�����Rw�R��y=��氚�s�,�ُ�1��I05	E!ʪڹ��YĤ���"���f��kƸg��r���+$ӱ぀�q��b�O�p�*W��mw���`�,�5��۹���ۘ����=�l�_���%5���f��S�,ӊZ�U�����v,�{2ϗs�W�TX�M ��̳_���ӝ0?�c�&k(���J'81{!�z���ԧ����<�0Fa�Llx	�v��s(_�(<H!�k��k|���I��);3Q�R9���Ѹv�c�̎�a \����f ԟ�0�t����t�Ss�b��$�������6�ϼ�S���Z� �;~����	�S�,��^9�\���>�Y����=8�6�U��@�m�2����N�]�zOg�ؕ	Ӧ�i�ޓ�|�F;�YkT��$�D
H� l�f^��] �����=oNHd��K��\���y���(g��*TV��Î���5V��74,�G�%�S����BL��m�Dz����^�LIwڨ��$I�!�S��D�O�?E�jW���u��X5���֍0w���Bh�*�7�/���97 ���!ַ:x��C�@�xk8Z�4`ܶ0� 犓��Usz��B����=vZ��D��<y�O����!�;�AZ4]7Bb����٪8�E�.����<�x�@��f��r�9.]��S�b��� ��j􆇉�t+q����3�O���ƽ1���i�o���~���M+ԋ��d����E�y���i��H?Q2 �p���}.����bY^E��@ѰD<#��:���a���,%"[�im͆��l�R�����ֹ9�U/S�Y¢I�Z:��Q��!B;��� ��L��M��ֆ�aI�	q���z�>��<y�XK���oL� P�׉g�·X��J+��P�7�>f�x\�o�ݾ�	�e�]!1� %��� "3í-U��������P��8�������"C��Y��0Fc��+l=j����)�#Vk~�b4x�+�}��@9Ļ	�h��Ǆ�y[(b��Mgb���a�����v�#���~�Iv�=Fr�,/��������O1!s|5��U	�.*Ş�f8��}�}[J�nq#�+̇�yW�
r����p��񔒥[N�ÐݎYΖ�Ez�$�NP���ʚ�Sp��'=|N��lZL��e%��U:��[$郪Q���۶i�o��u[��	`�$ l�u�,�4B����>���%��]c_�y1G��U�iJ!}SEf�֘[m�ǃ�-��Y�Y��򉔙c���\���&=�>����Q���)��G�`�$����`q�J��|�e��3�*f�y�f��L������Vei�t�ƹ98�;���{B�վ v�Yk�*2��q�Ԯw���%a��-�����&Ah����T�@-5���I'!d#�`C�.��xI
y��A�A�A��A��˻�pYvy۾�'+��'3ڪ�ҡ�Ɛ��!}�jUD�ָ^
ѓ��}L~i��w� ΐ����?�Ld{�H�_˨,LU�J�>t�q��٥؏[iC۹�_JDնºb�vy�����"!"wj~҂�<��/�0�F[_�d�S�ͫÛ�1��r|x�x��!���t�-�hb�׾� ���� З��D��P)����4�OJ[���s�h~Ib�}�n�f���b��kV��5��F<�Jס��H�#��)ە�h/�>$���i��.=P4��Hb+���N���t�S���9����ag�`ԞS4X^/�x��-<U���U�g�ޯD���L��|eB�]Iù�C¹�n{�Q5�x��'1��+�E`R��Θ������dj:���V�z�~��݌���<�@}�����)%��lg ��`:K&@*Z�M��'	#"�3>$��?��lX�����3yR.C�����_'%��D~��On��U��ﾚç�?�Q2�I������$!|~��i��,I?ĽMu
���=w�uldT�p��! X|���v� �<� {��:���d�h�G��f3�t��b�~�Tm��~�c(��v�C����pm�l�J��A��=�W1�6�^�
R���s,xto��s�O��h�׿��6��Bdi����6am_�T��ņ9�կ�lٳ�3�J�kq/�q�Q22C�v�@���r�g��,{�Qy���S�����@�L���Rk�tc���~��D!�P���
C�Z`Z��$N�AR����J���p�P]�M�υG�|���ZJM  �_{�S���>A#
ݝF(S���|�;��*]����i
��JGQ�v�}[a��cD !j&ݒK'6V�uV�q�"�>J>�d�k*�E�'F�%�ﯳ�,6=���4�u��t�h%\B|7kh�tY�xO�`7<0q�gW�QU�|3�2�������:�/�G�B��O:�D��6��ly�ZJ��׺�H	tɣ������d�QSK�9�<�����y;XI<��_r$m��e"1��P��6��G1���M�'u't5�GY����f�9 �-�
!�h���b��}xCb�Ă���W�L�:��74��}NH�dD�o'�C�5h�HE���~GC��C��ށa2:S�PV5�o�����pC�ӱ���W��cvG	�����R^xo������W��&���	�;P�(�8/B��"r:v��*H	��	�Ϊ�|&-tG�'��0n&�k�D��#;��"s�%&Kg0?|���Q�3C	���[6�=l��>�xz��p�ʭ���e����Ň�Iٻ>��U!o ����1fbTǧ�#h��NEO��-�c��DK`��p�qr[��(�q�j�8�bI2Q#J��'�Ε��w"�\�qad3%�[�5TF����z��[��+Jf%*)>8����kͶY=S��́T������Y�Ϙ�iC��V,�Y�8�l����=<∱��8��Y���y�D��X�#��3ͩޡ? 8@����U�[o%H��~��b�'BN�v�ސw�$~*����wÀ-�G7`T)��*k*�i����=��K[�9v��ZM�T~�u�S�ǭI��9�jY��� (9@#h�_����i�2nn�������	o=���S��Z�0���������q�Ռ�|��Q4$�h�Щd�=D>��r�LfӲ�,@���m�|��;,(�C�N�����Pd(��:��d8u�� �t4����Z�[{�Uu�,v��r
�>��h�9�cL�{~�X��wc�U��9��'��!�'=��	M��;��YХ��Җҫ�\� s>@rCā��.E �����E�_��*:�#��+yc����?�b(���.B8��2�wg���_!�D�*��H$=㹗������^��͸	g3>O�l�WL��k�F@g�>�f�Y�,V��}9JW�	eP�~��}�3���'��p�y�{�gyvK�>�����!��Bk�%uVcG�_F!Oz�M���E�웵%�p�(Y�RBJ�X��S�m�\>��ۿ���J�"�B͗�ч��U��� ��D���~����&u_�-3��z�����s����q�K�/��+�&�lg}7�-�;|/��HO�-�>ҧ��jbh���`�<%�!3#����� IbV���ׯ����oO���X��B0�ci�ͦ��x��o7
P���� �tBU��!Vw���pX3d�	QQ���?��t]f���-{ �����MF�֐�����-����,�k����0古�k���;�t�E���Z���A��.��.�)썞�L���������`@8'g�K�1:�8�*X�Ѳ"�)�H��<�"�9H=۪��Yu��Ǥ�SfQ#��G�H��&S"�"𣫜��~K|�+~h`�ሕ=�H���,���}"N����j��0TG�8k����U�%t�r�	��z���y��Љ6��eO�́  ���)hN����w��񶂴-�H�5x�j�V��	x}x2�l��T�{J�C����f!n�o�Hgr����oF���R�9O��C2�ŝC:�JU��%K9�'u�����|{Z?�>���[ �?^x,���x�Ɛ,d���S<2ޑ��7y��*�Y�i��;&:A)��c��3��������$�~8�x��?O�w���Ԏ��?� ��8at㫜H��X>���C���T9jR~��¿¬��.N�4ĜoXcd�lv�Eꉍ�	���i{SO�����yĘxx1��􀬊L��E/y[V G����+�`M�؜U����iHf��7��B�$�8��[Q���0u~����eC�fL|=0]kcX2M~Clnk�W���Rs�}eagY�T��uԈ�*\�8����6�p�]ft��6��3���ua�Q�2�"#�4�e���@�M�m;g�diX�OF������ރ�8Oq�iH%�Z�?��K�8��`Ȗ[ex����yJ�j���~t��;�M� ��S�������}��O,&sG�sx� �/W�f"��rn���<(3!���3զ��q[���X��l
��5*8l��r,�N	���A�m]\��ggJ��h���Z���Z����Øg��(����{��"9Ķ�ļ',A��kk<b�g6���N�da����uy52S(�h����-�B�us��.�m��
8��e3���`��Af�>ڥ'n�c�����*I�#=.�H���$����d˘T�A�,X��5r��<,k Sss1�(���[fx��A$�$�j���'�Im��LWm�q�
p�	tŒ����^�|�Ha�;�Τx��ೈړu̹yY���w��3[��`mǟ���z��+g���;�-J�I���\��#o��*�=WFr��l�7c,9D��)M<=�� �=
sۙ�gP�D�xv���N]xk�b5���d���``c����bz�[F���	�L�}<-K���#�=#��K���|L�e�C�H�5�P��D��S��XX�����u�%��ƻv�����[kK�k�㰆qb�δ�bRL�xy�;0����Qx���6����<
k�t��:{>���hi8�9J�D�DY��8�4�.q9�*�V��Ż�%��B�`����1R��Kj�j��v��_[�ҽ�����om�'�iߧ?4dmZ���s9c\dL��Jv9Q�Gl �_�
�e���e�e��5xkO����i2��{r:ٔ�!�n/3�+��!z�Q{�F�4!��)��"�Mw���j���vi��������z���B����[���R$�3.�Ҳ?�O�Ro��юC�1��S�z'J�g���� G��-��H���E�fK��Ojk�ߙ������c�_=JK�@
Eׯ?�[B�I�Mi��J�����<+ Y��6vRu��/�6@g2yL��I�|ȨMiH�oB�VF���q~�8�o	�C���h6�A�u��{��tJ�t�t\�]��w��-��痒��1�̸;s��Y�a��� "�3��q���d���B�}���7��r�1
�ѿ���[���U
M/���l���_������X�I�?d���?��̼�����Q8�i����T��r�<��u�X��H՝�/��3��U�&�8�ם�E���Z�*�{����0*�'��K�,��'��;(Y<6�H�䘳�"ƿ�ǔH�j����?�<d�[:�٩���
�{���
H�u}����떄�Z����U-~�}@񎱫xh�;q��3>y��{|r8��VU��}4����E�\�0��
�^.�{�N��gm�>ɵ�%:�ũ�f��"�\b������y�$H�!GN�kl	ϤA&5י�+�e��>id j�I����ÉƐ�RG�/�gXd��55m�	T^SɼG8�v����J�fp §�t/FW'��A�q��4���6��5��;�_cn���RF5�D�$����G��qb]��?�rf���R�p����j�7����#O���AJvq�_K��5�y�7�����)r��*M}`IB1����烃ڂ�q#o+z���q����Vi���N˃r�<Z��jMy�Z����VÂ�tk1�B����"N���0�T�h�L�
��~��в Ufږ��$XZ�&��� $Jx�ל{|�hW5�w|L��~L����I-(G�5���0)ل%ܩ6�Xz��PN������ޞ*q6�F���#_��pII�V-�e����r�F����y1q��s�m"��`~B��[*��k1�$�3�G���4E�O�h�K
��4Y�q��B�҂�5����x��7aw�P��1�Ax�� f1G��Qf�_�Cd֤� y�1��E����ݼ`�9�i�Ǩ�o�W��Zb�&v+3�|�N������^��Q ��HH��������ZN�4�b7 ;�	��ŮuQEae�>Ʊ�+���LG<���1�7u��?H'G/XE�P;�'o�>�,@V۰������2�d��[� d˕����6���D)&�MV��CM[�n��\j��VI�f���-����
����HƬ��W�E<��[��4�?�lk�9_@	��q�a�E��eZ7�XjLsWΘr�/w���vt����WNu����b$����C���mE��^��4�b�~%M�0��u����NnicK?��G�j��N���܊�k�!L^D�{,��M<ǁe�xi�Jj�"*YԦ�7��?_s��ĳ�|��#8�ؾ��]o�Q���k�g��d�ɴ9���Y����W�u��y��5(󥳿��ru����7�2��p_������K�ռ��9[_���[zے�_Kޣ'�x������rܲ�q5aN=�dX��z��݉O).M0�^KkCd��,������>�e�&ΰN����]w�y�=]}�����x*��]Z��l=)��D�뱾��;{�l�D�t��6�����+�i�x���9��t��&v��D�%�U)F�����i�S�B��hR@ܹ��i�\�1WS1�I^I�*`?�G���-C��,��Q���F��^��ԟ�s0b`L!eG����"���f�����2�Z�K
;���Xl}���bV�S
_�L��yΫ��0�g,�7�� ܹ��C0D"%��I8)-;�6[l��I�p8NT�)~U��Kh��1�QOV���J�ۢtpy��H���H�Vw&a~$y�Ew����)�r�z���aƘ�k5��L<��:�:�, 7�Ը	��WF!�e� lxP�jul���^"l�<�m��B	��Լp��] ���c�ݐL,��e����0��ؠ��Gݦ1�#�Q4��0���tՠ�����"HxM��y�j�	=�k|�aE-"��^�W��g��OH�i���/�A�O�ޏ�c־�Je���D�,"9wU�y��kC7��Šf�SܾTSU)��4OBq?n["Xj�J�C��|V��R���ƉQ���~JZ ��씋-�K@��{�l;�I��%�YI{���P����=ۈ�z��]���~�/ET~�;߾��넯���64c5��쑍�/M��ߑ��`�1�Oa�.u��O�ǳ����(5�_3�L� ���	���B�]`%W�>��D��QH���^~7��w0��;D�:�Ǻ��b�+��n��D�Jj %.cR��D����Z�}���݀�c�M=���xD��J��o�%�ڂl_
�҃/��6���̾hdl�|fSن.�]�gk"�Д�7	{��Ԟ[д��;�R����/0P��,;+�ml�P��d�M(�ݦF��6>�ʒ�?�k��{y�81��olx��4�o�`�Ec̕ۇ�(�[t�O����ڨO����~������	I����ԕl��'�t���֣=���l���Ni�c���	��ܪ�%�� ׳�u=儜��d��dIn��w��1�s߂l>G��l�i����{�y��_w��b���/+zh�����P9�|����vO��q�A��U�t8�A*szX*:�v�����:�G�=�ð��Ξ[��G����CL�Y�(��K�ˊ�e�����G� ��B��w�:KfF�(������g ERQlQ���Y��I�
����ߴ������ﱳ1��{�K����z�=�U(�$�(��:��s,N�	+Z�L%b8R�P�!y�g�X��f�JNU����SƊ�k�3���sl��ngC¡�W��$fA�;cg�:����k���<���C���ӗ?�L�YdL����&WS芫`'E^��!��"V���z"h������;���2QÔ!���#�AD��\6>0�ϻ�l�//��DaUPcC�*ֹ��4<;�&�6z���݋F6V���"�f�w���6�-c��`씽N�]�Ϭ�c�6.ͫ�)�!S�t��,,��\���+��r��0��.��Ʀ^����^��g�ṽ�7�����U���Y�{�R�[��m�?���Ɠ�~���Dͅ����hM|!�$����CJ��7%�QdH%E[6)7g)^W�21PS�A7|�?����7'Z��`�т�$�H|�c��R7�%z"2e�<�?A�m�Mw�\�r�$&�7��M� =?PDN�����M��G(�ǅJ������+�7�q�9���E8V��AV0)cbT�ט���ï�R����fY]�z����}���]����Zo�D�P�T�M9�48�y�FV#٧�l���|})F�/���+���6iMA8�
�2�V�$���,d�0Ů�����մ+MuЂ�T�#��;�#D�����Q>�5�\[���ZŌQ��I7	�JI�"N��'D�;���%6^�j�3�T�=�HR��<�� �{YRA��C�P�%��х߼;���0��RTE�J��P֊���Q����fd�_��M��'z�8���9{�e���I�Z��e��*��S��v�i
%���ڑǼ}��l�z�>>�����j{WY��U���/cԩ��k�D��<iN�^n#X;�)�����eM�d�d��x���Y���x� �4��Mr(��Z���N��a��,w	�t'!佲�nF{M�?�`�A����Z8n$m`����n�-�ɨ\�2�V��D�m��:�$W�V0��G�R�
^�M�ͳ�Bۊ�z���6��1�1�c^�@�� �/�7\̑{N���:�<<�����$N����%�<B� ��I`*#Ih`��۔ ��9W �Lՠ<j����=�l}}�j"���u���~��1�"��6��3�r��ƙ���%�30Sܝ�aF�"������n����(uB�4&�Ey9�w�aU��|��~���y4'T?�svof��	R�����L$�qS�|C}�wV�>"gI��4�{�7f�r+���RՊ>ܳx����;N_
G[�B|ҹ�����Dt��tV��i)4_��_Y8�?;�"�`��	���+8r��H�p��Vz��8E���=���_Q��#<Zk@�_e�"�1��y��O��@v����A�k G\XJ����`��d0��yI&�|j��Q�7���ҋ+��� �bN�uh��X0����@�mmn�MЙ�o��W��+�-S�R�4���_#�F�FE?�����6K�*R�AAi)}�#���k�m���Mk��9���=+����h���*�@������N��:u'S�i��IL�Ԏ7��U�2!H�m���4EUغ�����깷�D� ��
�Q@�s�'g���0��� �6��4��h�<$��'$0�L�iJl�`f�~1Z'��d }<�O�>�����1�����L�7�LPU�X���ؽ������0"<Cţ�y������S��F ��؂F�a�ߎ(bʝ�}a������� l[~�!ŋ�&�=
�ؚ�Bo,�dm���@S����>�r&�)��-A> �y��\�"M��zԤ�Cd����$?sT�a#$���o����g�+�j���=�o_	�s+E��>>li�0�t>-3m��j3��c�
� \a�o䄡	R�(B�vj�9A\��ւ�Ѐz1i�7�h@:�{�����F��7�����0�-|ـ�N�rR:���(��Ym�,]��7k��HB�ql8�����/;���H��>�7�,�A� t^���S̪���f6;<zx�(���!�~ok\��y���/p��h�l�¾ t�8��ɍ,�"�=9va1�N�Aw��'�s�j+/�#�0�UX,�r#����T`�����c�$,w���As�7j� �^�arơW���Щ��r����n��!�"V��,�.!�T����`����F�l�tz�^�]�>�݅faCl�Q�H�Δ�ڸP�)<�r��'�	�w�����! ��Ƭo_��#��w���1��{�N-r����v��]4�#�� �����*�A����"�-��%�	2�]PC��r�^����^�Rs{y8��\k��>I�$B�n?w������5��oB4��o*c���D|j��J��H֏Nհi�T%�S��mЁ�ݕ��T^�Q���:�u�����M��4Բ��iJO����p�3QsJ��mW��e�#S��u&�0�8c����}�����J���:�C�K��:��ݔ}J�E�'< ˩!+����-�?]��ԖK��ʇӘ�hm=��#'�es��g!�SRr���:�w���@坙�:p���fq��Ö�B�����4waP�fkT˼RzF~���T�CW'?����n��4�&�j�h�nl��;�IUӠ��y���S^��1�H6q��'�#�
:��sDq�4I��z|�X	D�jZ�m�"6���b3R�6�+�8����d�s>:#k@�N��	��9��}��4u74���� ��y*.�oj�$T�o;ȏ֦$��'IM�7��r_k�Ds��C�D��� =�����Sձ��f#*}�N���>�cHI�!��ǯ�j�\G�Á�rz�"s��l-m�_�>���-�U��$��Cuw����I�*t����=;>,fN����H�A�1t([%���Ow���s��э�����E7�* ���-��G\�������p2F��<��(��h]B����a�������}��9.'_��%�"./��q<��=�
'3�Y�3ʁ+�G����ʺ� �H:�AQ����;"Pg�(Jn�	>�A�q�gW�pyv$#Ⱦn�|��x!����猲�8E�AD,u����˽�/��K�3���l�gz��&M��A��s�es�r�~�
=�7t��IzZ�̯�= W��`�+�k��Z��Yo�k�{.�'��|��*q�6>�v=u�V�����}����-W!�jyjc��':$�ل�[��&eup�96��ֆ��n�+hk�n0��zJzdN�g�E�n���F�~I���י,�~�� )w�T�K鴋t[C�>�G��Ĝέ��OI�:rh��]{�@���X"	�g,}��ۼ��h�_ǖ}
�^ܐ]�~}mAk�Z��V@鯧Y�{W���a�TE�R6_pI��8�f��mZq��c҆��0�"���̐r&+U�)�y���F�͞��lvHe��p�<(]|~�M�M1��G ��y��鶤S�u��⅝SS�KGߔ�WO|E�1���׌o8>�{L�0kۜ�~�ɍ��9�O�����`�Vm��NGܤ8��������F�ҕ��, O<��|	]�ܑ�G�Aߋ�R`Wfw�q��7p|��{��tx[��F��[�Q^��7��f\C�BV�kW�\z�:$oU��$��� ��0�Fa[�k�)h�2Ǩc�|	���_��Q����djc��ks�o"��!���_����Y"�j�k�'����c�hH&��8%l�V��*LH ]��}���H��
�B������fO�M��~�D�9H����xj����K������Ĭ_�Y9��{L4M�$��ҸEL	*tP-�7�������Z��lu�7ͪ׳�^��͔�6l�$��U3�H ���>�q����#�����K.������@jr3��k�x�a�W�(�$y��ܮ"��f;2����ON��8��� �0y@�ww½�\
,[C�Թ.b��Bn@�K�}����`�� mѬ�{-���Pe� Y�l(�"�:RV��~��\�;#i�%N�r4�?aZ�*�n�(�]�tQ���jSx8"�=�H��eZRIQ(z�픯kZ�����ݿ�c3����楹��
���N�K�ګD��	�����8\ǲ�����5�~ơ5~gIlN%�]�|�S�1��yI����[��L��]�.8V�wS'M�ę��|����
���n�xO�"��+#�P���2�թ�~%���F2���'������5�=)�n�]��-�p��Қv��V$K�ͮo�S�P���87h�_aD-	ە���4�_i���N�O����Z�#m�/���}���&�69�oE�Z�$��G�e4��؁�?�"�ﶇŞ�R�ܺ�6�� W��sk�����YQ����%Eh	�n��TWBSۀ�M
�_$p�1�N���E?���,�]w��'���}�c'�{�J��!]�++��b�t5� z@�`�U[cK��x4aY�]�ˮ��or��?��N]�5A���V4n	�}|g5�F�z<د��\�Q�� t��)4vv���8q���vcw����K�����)���萐 �?ē=���Z~�L�1WLZ�M�92I�!Cn�ir`��Lo'��;������y5"�>=�S�3tH�	
x��ӑ�Y� ��}V�߆�#��v_�>:������i{���[0��H���4a�� KB�x ���8HH�`���\�5!���S���k� *�@+g�1�v�����"럅����h�&��d��~ũ>�U��.J���}�"�R:��?9��q��S7�d�kKk�Ө	F�Z��g�֖��n6
3�P^�w�
HɎ���4�t�c���ʾ��qp 1)���!�G �4ue1�g������&���c�ʲ��q9�C䎓7d�"f3��)�Lb�D���
+�2<8_�tr���5�X:�j�����B#H^=�|���:jH����+�w�0e�T[��~z/��d�s���1�H�LT>nMŮ8��|�W7�-`���,i��N�r)��)�n�Jq#��؊p�����w@����c�z��Cz���h���:�@諾"b�2�{ޅ��������!ׅH;um�F��~�|��G�����錽�OķÓ=��9�j�;.�XH���K(����k��b%W�_��*\��������I���~Yx&g����!$����T�#�ڑ̊@����ϩ -u���V`�7	]��KQ�&}5�7f�?���v۷	B��:v���R�g�df̨X��3,C�O���>1���T{Ēۭw=3��{��N D����1!|�Vp���:��ӏ�4��@�gٲt�3@i]gE�EZ>���4�X�d�M���U�O���9���m�����s�z]�F���mG:�X����%,P`�s��i�fJ�_��^�T�wE.�D|V2��R�N���5!�FX��V��V�%����Ǹ��a$aV՘h4/��!�d�z\3��C�%�@�Y�>�u����h�t��tG��m�n%k�`H�"��������Ö��$��՜E�b��:{i`:�A�R4Oe�cxs�����ʾݤ��R��r��0��{�_֜i��7��5�+[N�\i8�q"hOPhy�J�6u���Ӿ��b�Ϥ�0U���:�;�	���=�����V�����oeA����$��F���Tk}�0]Z�3Tp�c�8b���W�����X�>��f�av��%�F�!������J3��p�i�e��{�s����v6ǣ�'����	�i��C�=$q��uG��~�͉����o�M��7$�㬪p�:@�`��ɵc2ם.��dt�֌�y��O����}��Zk՜�����������D.���h�L��&غ�N��������g���J&�Φ�����S+ �aв��"7X(����Ǩ(�:`,��mܺ�c��FU�4��]p�[�	[��w�$�tcL{������?�y<�RQ`�Hc��)�"�(���|��e�c� ��t|E���{�wV�B���j`�Y���7������2sBg"C�+�/��� �ƽD���+7�Ć}��8U����y�Nmd<�.�3�D
'*5Z����Ci��0Xė&�'`�@Mm�oQv���V��[���O���}^���S��k*�竍|A�w�x����T3�t��no8�#ͱ��Ҿ�f�	m+�]c�j���mn�@�ɗ!:�݊�����tye�x�X?��y����H8/7R���L.r��r��t�jmǋN��}g�v�gPÀ�%%���j3R��׳��S�<b��Π��;w#݃�
�Y�R��
��=ڤ3�6��I�.j������_�Th/�.mHe�y�ˊےk�ޫ������5���N�}wP�}��T����H�)�?;�i�1��7`Ȇb{Y���kC	$��\�]����m]K�/�U���#��g,?��RE��}N�!�����!�;!�`ak颪���0�-ѧ[�Ƕ�q!0�k�����xA{�����<��Kt�f>m�R	{�w�WA��,���z٘���|�/���5�ً����?���\�
e�����n\�5�?L\���_\[G1
��i�Lه5:�R!�L5H0�O4�8/�Z�h�@\,\
!����e,exlK'/e�d�/w6@�+�)p���W�K,�>�|�u;6�3D�>fy�PVK�dj�3�������Q��=I�D'ň�G�Q\��Yk�*���1C��D�j[�i�"ޢ�}�Q���@���;h�rh�,C�5-4in@������	�UE"$��R�'�*z
zZJ0�q��BA�vZ�y��<Bl����üp5�(��H<+���q�~J$���*�T��B]�����v+�Iݑ�^8�Ap�*�ƍ��Y�i�����I
O�(&�������*��k'�mD(��1y����DL8���sP����Z�d)�$&����*6
��U���f��<B����*�^E��-�f�� gd���pB�����&k#i���a�����t�����0� }���:$W�Qo�rY�����kRB%�Y��A L�'�ԟTwd6��op���i��	/�ޣ������L��A�Wd��K�w/�V����_�a��?-�)��Dug�"�j����=
��}RQM7��.#@��;p�#�"���W~T[���������_�;���D&�i9�������8�u��(V�{����8�7��������2���#%�����T'��X�N{�k���̆���1�Ose�dE�ĕ������,�0s,�Ί"������1|�P$u���� B�,��e��'ֲ0گ��f�ic���igv,��L�^7ہ�,V�a�!��~T�����U�5�m�a�_�>�'��>�sH���bH�C!5P2#f�$j�c�41;��T�����E �e���@���r;���Ϙj����7��,FYW�/ْe�{�����Kb[:�cW�3@C�s�=+!딭�&Ǿ��0��0�����:�M��o�ൖ 3oy���?� *�n@ւ�QH��������JW(���N�Yv���>�������n�U;/|���	�/�̱�n��=uǗU5�j�ɗ�<�[P�u�#N��{C�l434ol�Z*�/�=>���Csp�]7�tU�*vI8�E�������^��P��C��	��Gk�.��_U��D���F����{>�\5�L��?����j�V�-���
��X��v�Ta��?P|�]v�߸+@�L�?��mEP�D	s�����3�=2Ë�{�m,ק��VBV��0i�<� &ӀEZ ��"��љ�Ҹ��ً��j�h��_\Y��4>��'�I�dIb��|�,��p9�5'Ѡ���Q��+��k�`L�% Ǫ�n����S()���k铕ɘ�S�x��K�������.ʢ��_2[��%�e���v(���"���29Y�� ҊC���@�ax]o6S`ƁևG�)iVv���$ԟ,Z�����4Y�*�C���@F�����.So2�P���)@n!�M��" .B�f����2���#��)Q�e�/6_�_�H7���5���t5�n�u�oo�����H -QA��,�&�X��/tW؞����-� l�fI��n�F�=��;�9�X�&;�'^��I�[F����~��z!T�=��]���
��k�Xr�ٱ;��x����ð�`�R�;�A��~���j0���=B�2˞K���^�ߖ�N�5��H�6Q�� ]��=����أ����$)�Cϧ붦S����u��vf*<����'��/��r����5���_z���Y-q�a6�}��"�'�6��ͼ���쿞��(ƒ� VW���B�[hZ2MzU��$�K�W�{
{tX"�u2���f�4�5�/t,��f����Q;�\�$�],)�$�w��>�FM����W�	1����O�	7�ʿW(ucw|#���kE�sNV�{ģ"����Y0KٔJXC`ŉ|��55]}���ϱ8zP��0W
Y�0	���of����L��:�w���A��T�'�7=y�JB����z&�;�����ַ��{(*a"���Q2d9�i�9�s�{8���@�
8��o�<���ڮķb���,���'�}�����U�#
�Q��{���� ��U,�'��JBΪ�Q��V�#�0'�r��j�}%n������B����`&�LE�<��i.1����)�|���_�������r�/�9�� ���5IN[+��6	�q�PJ1ׄd�ϯ��h�_�X� W�F[J\��n��J3��)[��(�|��>6�U�^Cb�
�B��W�Rw���S�N�&�)~��k�I�̂��)����E��8��ٍ����h�χ�C��Lg�������?<�f�R�.6Ư����N�\ֈ+��2�I��"Xy'���7�~��9���A��s{��,����T���AY9��NU��(&+���o<��n`���΋(�4 ��%=�����+�Z�8�v�'����8���4��a�"�tWNBw�H�n�RO�U�x����1w�z��N;'6�WE�]W�s�ua?��@0�2>5hu���?�oJp�N#�p�T.8Ѻ5��9L&`�)F1<�䙡U�� a�gqz���F��k�'t��/��[���@�;zRm���+ŒƘ`~S�~��_ز�p�r�1�m��_^^��Q+��,lFe<�0�9�ݡq�����9h��.����_l[�VU,�6�`F ���M�B&��\[���u�����{�>A-�B��D���n��eٷ+-�%Ψ�/��"�5Ѣ�b�v6'E�Wy�o���� ��ঀ����诼�ĩ��;Y�b�%/�
4�� ����2x!:a��%�&=��<��x��v��J��_�l8w�p�h|�dR�`��p��ɝ�U�б��F��5�^�'f�W��6�3��l�iۺȷmU����.�生�5|i�M{WJo���'�g���<�x��"1X}���8c���y�ɷ0Ƌ�$�y `��B5&݉���j�Ƀ/c��q(�5���W�:|U�Uz��x�[�1��
��fD�jcV��h��h@vʒ��c��c�LΌ�}�])�Y�lRu�fw��Jj�#�L��	�\�C(����[�����vԅ���>/3�x�]��$��Ԗ	ZB�)0ǖbI>1��Տd�V����T`OzV��`�X�aH���6sr�M�8������"�@9c�Խ�w�?J�m&�-rM>�z��ͽ�u}��%��E��,���_��9�~:��fR����Z�_�n���{H�e<ma��u?��Lg�c�+w� ����'iHj�mN	��y�rt/�gx�'�O�R��d}Ri��7�=��S�+���xц�����H�����
����>Y��wt'��M}ϕL�C�~�n��������d���9��-Yy��3���^����&�5 ����'�P&��\��r�J�M�``l�+��=΄l�)N���"���K�"�����	)ȱ=p���&�BE�C�͘!�5�6!n����u�W���U뢰��/И+wp��:O�{�N��~�Z�{t�M;���n'��y�0��Y�v(C% �'��	��)o�pw�D�ۊ�=��k[äP��MJ0��B�_�r8 �yϦ��s�3� �	�U���>�¥�"��u�f-�8�~�N���\O�K�F�����MT�����n�xO�l�S��G�Q�?���Џ�Mv�����(M���5� ��c��4lL6Н�Zxi�N��4�
�\pJ���#�hA�g��:����$T.{�?����OY<?��Pu�q
��!<��<�,��N�ӓ�I���F�j4L[9R����(�3��\���">��6R\��t����{;I���T�k��қ]��0���Wy�4K֘;�QőRq	��w�;���4��/���T��7vE��6�,�Y5��.�X?���	���ߦ��[��.<�U.��e���/iE�@��K��L����E��� >�Pc���4��H�WY<��29�������M0���G����?�ù�"fՇ-C@��hɏ����q7�ڱ�f�!��EW�4VS[�"�$���+��,�S2�!�ڂ�����;�c~}u.��n�G*��
������"�)a!�]`�tN��&^�p��t|ų�Vv|(k��hS�1��,���k�l�q@�N�Uy�~}��@�;�?c������F�
���dl�|Z)��{��J�vS]�|����6$�ኂ?'�Gʉ�l&D�w~)�+���͖d.�Hd���We�$��h�,�MuP�PnP\MQ�.��}��9]�v�4xQ'�@l�5g�c1h��6�`��'�
�k�Y�^,;�Q�e��ԝmm��A�˜�'����:!y��-u��u���s�?����P
D&�6�yH�{z��+�ښ#jz8Ͳ��߻��k|��9�h�=�(:%��,E� �B�#�������ezN������}k��֠�为u�����/�;>s��zV!��:��-��S|��Z�N3�hWy+�V�޿C�k��|u����X����UV��?��M�|��jϏ?*�mP�F������R�I���-��D
!*��|]3�6(�:��U��r�^On5 
�K+�y9`�Nf/>f�d4�B��?�.իFN����3Ag�'(������X����z�G�#��cA6���.��r��u�^>�7y�fm�k`YcIPj����,�+��7����,�8�v�u\$O���b�ľ-z�K��{�o4��-g��ׇ�=��$�4�����Lߍ(/���A-�����gt�Er��٧9e�ѩ pe ��Ѵ}pN�<����CT?+?��Pבw���}ʬY�g^��q-\����%�j<��m���EߪR�}
�b���"���~\������(�
I�
t�9NΎ��?>�Р��F��n��������$C/d�Y���q�WR+T���<���-�8�E�cA�:άk����Ki�	������߻�mA����n�H{����i?�b�L���GZY��t�\T}EӠ'��B�Β˶"�V~����]�1hˇ��G'/����u�$-+])Pn�@!�<�T��A���(�Mx7�OiI�f�1;5F_�d"_�J��Ȅ��K|E8���!~V8	샮@��oHW�%�C�i���Ҵ��?P����2В�|�=u�Zj�O��o�|��m7�rZ�53>�c񖉑{�H���hM�����,�%�u����I����O�=�5W��ݪ���,TUY2j��̚4��/N%��kZi3�>Aa>Ɯӡ�I�IߺV��~����׽L;+�����q`�!Hc�O-b)*S����w���g��?>G��z����B��lڜz�OT�Y7 �߽�����MӪ����;��w�E���<�r��?b�� �O���p�JEm:�r[������XS�I�Wr1�b��E_
ݐLe���a�ھ�G3���@��Z�!�	j�_''��1$qa
�v�RI�&�C����R�?�����é��Q#���X(K��`u�3"�E��T�їS7������&�q̝*��󖠖����>5�ip"�G��0�,J�0��+/��b&e����),�ЁԊ^�<=?L*%ɐQM��툜s�?L-�${M���ңV�2���� �blI�'�<H�B��.ŇEfp1PS�t29]�v���3�*�i��gR�k��3�Bx�s�����p�h�̙�!�WC	�{�65�5�<K�Z��t&���CS'BZ�:�ۥ���@P��$]����,�mV�\J��]8�w�!5�䢱�}&�}��H��P�ڻJV�ؕV�����	�숗�����o�׈�+�[�ǀG.�y��%�����䪬�1t������%K�O���f�O,�����
�3���($��F���Wb�W��S�S��S�RG*爺G��H�f��~Yȅ��$�	�ƿWE���oOq��@�aB�g�u����[E���e�fH�ſ�l�ll̃":X#�*C���w��`[�މ�Y�e��#�^�l;�� p&r���R*J��)�6���(b�v��Y-�3�^�^��?�7���Z�g�g����Ѐ�,j�1+���9}��}/5"ؗ����qT"Q�q(�&�:���՚(x���挋JF��5���'�����wV&Ju�}ӘE�1ÝF�9GAbK�y9����i���5ص�C�UsDK|�ah���Nn��Dg�fp��d
*�(�P/O�Xu���2��e��D���O��!x���:�����_@�,����9���CO�ٍ'?4�T�Vz$�����PlE&�h%�;?>h�<�a�Q�ҩ��[{J�Ywp&�cv��Wʈ��y ���@�(�p~ɠ�">A �g�n�d}k��e�-�4k?N�ݹNQ��Q��MH��~�xfϖ��!��=$q�;�
�8Lѹ�m&��`߇6�m��r�ۉ�gebq:��:^��z��«�.�/TiD���u���)���N2�Ξ�G����)ؼ*@�5�H	����]+m�!!<�\Q���ۭ�_7e����ض�5흴B͟0�Cԡ���T���_|B�6S��֛���n�z��hYo:��xv��S��'��� �d�"_i0�X{�dݮx1��c�?�F�Z�.�ߚ��ٙ�e��A�c�?v���璌5�30���KHz�}����8��?oj�U�G��؍7�za��3��C�3KX0�"�4�9�X��u�`��bD���|���6t]�B�y��"<b���<j����Z0@�����q�=�$R���Ӱ!�{I�p�(�l!�vP���<��k�*�d���N'�K%.���>���K��h�uPGt|���Q¹��ӇV�	6�EWD��gNE���.������o%��鹚��`�� �H�On�,�~�3�H;,j_��}8�V4C�C	�B�E����~ ;u?aq=�d,�DKUE�J�������Fc75���`,G@�B��ŋ(I�tɒ4hK�Ŷ��)>&x .0����\K�����㐈�9�sIqÊAh���EJ�� Ә�
�N�?���M���ض�u����؉�$��&�ql	��Q�F� vF�r��0�Y�X~�b�q=�G���١���Ec
�Ѽ�-��ȼJ��^�-Y�k=��0'�r)��y��Z7�ЁW�fkzabQ����*Y�0�D��lǪ�Pb}'cj`�Iuɋ�D�Cwq|066pӗ��7�H�L��aO��:u�31���&�ň�_�7\ք���Z����I�3<����Ǐc�N(�s|$ؿ��Y��β̠�K�S~�ye ��8q����y�ڕ+�w�O�Eo�x	��^�@c�1���#+��������J�=G6d:٤A����4�WM+����#�'&F���3�?��V.>���;�r�����*o'�U�d�%X#߶��j��D�},���c�ha �u�!"7n���J�6Sa`k�T����?vΗ#;�V�b�=1� �72�B�n��ڴ~C�|B��	�>����Z�d���'���9r:6~?�z,*kD�1`9Y>�[��Z8��w��,hƆ9��C�Kd+!&��"�z�0��f^3�U���Uߞ*��h�ė�ht�P�t�
o0]/�{�̩z^�lv1V���n�F`�2*(������V@:m�-�a� �C�XgKˊ�Y1�E��תm\9����:�*�ֈ7H�aH�����ٝ9�.{�
Û��~ȱ�^����0�\��~ ;��F�?�,��+�K���|*��\� �p2$D�q�!>�YVy��=܋�=ۓC��s�(3���t�&/��S��K��4����5K���}���֗97�'�{|	u�/�~.0�>, 
� �|��T(�6�:Dk1D�XVz:嗎�H��!�!$�����6����+��R=��ɾ"}N`��sDU>�~�YI�q�2���(-�w9�#u	�702�$�#>jLL�.cg&�S+Gpq(7u�d�qC�ޅ�b�=i�]J}�~hF�6��>L����m�<b(��f��P���"W�sr�տ��B;z��>�����?�-˃E]J�����@��Z�	V�C�B,d�k߈�e���=��L���T�����DeTM _�n�S��4Δa��ևh� �r�2ۨ�/���J�t>��5ӏ��q�/�Y����%��.�j�݉W6���w#����MDy�HxL�"ח�7�T���x,<Ht�d�)������?#�4�V��X-�S�J��K�{�l�����m�L���(�a�����Z�sK62 ������T��q;;2���Y�%*�7�N%'Ipy�G���;��sL���0N)�L����X$��P�yޱ�9	h�K���j��& ̒�A%�*|�=�ϊ[6����~1=��Kh���Y�zS{��HG�K�7�2��A��q�&��f�Tyb�&q��Zķ��oнB����:�sF�K�ZL^��=62ʁ�s�����e�#��ʉ���c��� �;��!��is�y�>f��i�t�z2-	��B�lL����2s��{)4w{�J��h٨NG��P@�}$oQ*�<1�tC`�L��3�A>g ��0"�8Eκ�4���6��p"��|X3�$Q�'�+���
 ���P�6�7�'�0A9,��m�W��"A%�y{o&<��}���p��3r��*�����M�foa���OE\(�u�������&���aQe��m��usB���c`g ���9:��s�c�����8&	8���	�����Hz��ya>0����F�ֶ��
cmĚ%��4=�V1Q[=F�Jz��Q!���:���G�2�У,3�!��O`c�\�q�W�A�U�XX��;��� "�Z�0�
�8��r�� gj���i ��)���תq���J��u���0� Ξ�(�"<��Ҁv�P�C᜗7b�q�a͉�5ib�btF*U-��(�+������-Z�ZY+�(+C���#��e�����{�к�"wid�S�ٿl3�u�f6*�	�L�Zo���\���5׍v��A�b��m,E��kh7~�L�3d������!V�,�bI5ܝ���OMPXe��5]��#,���y��q�3P��*��U�9ŷ�S���4��%�k;GR����nM°���I�������E����y$�R�D�u&�MSz!?_�y�h�s��K&Fr�)v�q4��Cx��[�����3�Rh>�A��������C��D�õƭ�w#;l4�p��I1�+�����){,��#�z���?�U�g�3��JV��?�\���&zju��!"���7p�Vg���R";��)���j!*��^��;�/�w�-��yYK�>Ĩ��{ú���C?���
%�婖�����C��I侦){�HK߿\Z>�G�w�L����Rٸ�.֗}s3��w)+��qbN)PR��х�X�"}���M����{s��6��f��j��$�Q���d�A�7O�K����ɂe�@j�ƠK�2K��Hwh�/�3Z���(��������W�p��S�������g&)ؠ�P.\�e�{��2�j	C�ޣ�[<m"�Z4T9��4o>����K��gz�z���!c�r�w�5f���:��	�#���7�������%�b�cro�|s����_��1"S���ѣ��m��t;�m�𭏴��h�:�(%����s��4����Z+���0�S7bQ-'�&I�8��O�8ZՃ��/�SӾ�Դ����R��S��O1!^+H�8�/��kZ{�*���  )���b���n�Q���x��.fS0qF8t�	�%L A[��]�)��L�.D������L�z�,���O�Dk�m0���'�[�����8�o�BH�_s<^k�.�O���>��.6������A��B@*.o
טD����6��W�Zɸ�m ULC�5Ee�F@=�C�M :�`�q-�ɸ5��c�>b��*�B�j�M����7@,�2Q�p��PEL_��H 	Yn[$��#z��IA��,�*��5���o���P�-������k,gi�>���;��Ƈcy�� wS�C� @7��W�e�DY)t�|-�H��F�`i����
N����ۮ���섡;%�mB���ؽ	�b'�<bc��Y�7�d-�;� �o0�>qz�H�-CZܧM�T/^5X���mg�d��²Ak�z�o� ������0tyJm���<�5s ��+�k�)�BBC^�[@B��l���6�)��GIa������^�JA�Ge�X��m6�7�q�(�$�9�̴ �ө� JO�&�T�`�H�+�z��R�3[�LX����C�FIj?F�[{�a��~��7�Ԩ�;
�0� og���	 ��\��xu��r��|�TvT�L{��%�-�C��4G?��)����E
2��`k����(�X.ՙ���Y��Ӥ����a��еM�I��mr������	�Kࠬ^i��Cnط{Yq*���(*K���U�
Z3;�gJ~uCpVu;�FY�d���f��'1QHx�N��b������+�@��`��IAt_�<cSJ�қбP0��S@]���N�Eg]z���B�G*�_>$���Т[7���,�|��M5S3��gu��-
h�9:������B%�р��e,a�Pd�P��A|Xc��%�
���fA,V���3\0������?3[S�oNۆW%C~ ����W�lYJăb	��N����W����,D�p��������MI���
����=��R�����z�¢��m]_�}�Z��-�9N?�����Mg{�}���������ԇ����$҅�.`R달���}f�)�N��I���х2M{IՌ �j���k�|�kV�!�r��|_������E�<���O�f�3�²f���B��y��k{���d�zW��nm"'�T�l���?�8&"��r��BF@G�#������9Y��j5O�'x̄�<Ƃ�~S_�
׆��.PE��ɤ�ž�ۖ�{��;[#iE#ư���Ń��x=�$&D���kHj�k��jx����X�p������{�W>����fkw��g�P���tfz������hRt��Ss~�ѕ��.l�B�0a2�����D���b�]�%�J��zƩ�Ok�(}��3G@�'�Ï��BK�Ŝ�"U���8�������c�k��X"���ّ��r��?KԌ��qvG��`���N�>���v��j
zg�lm�X%g�) � �S��	�[{-�6�.�mS>@vz��B�X?���G�5�!��o�e��ԷQt���)OU]85�ҊG�Gc�E�['M�c�R�r5�E�*����lݗ"�8��l��8>�0G_���T��R��9b/
��R�['7ZĈP	�9��
�����W�Y]��Vo&���%2��]F���  �{1��6��{U��؞1��hxU��F�;'����ꪦ��~�g�|�_��Pٲc5R�:F���H�_&$_�� U�)N��o�dx��a(V�z���`7�l��y���Y�t���͓�FQ|�Q&��gb�)���N�0�ҭL�K���;�-D] 4$�m?X֕���ca��ذ׸gR{j
VD�H�b��LJ�˯R�/�E(�^��욤�G^R�"yS����V�|����ܷ���A��M��R���������c��$��U����|���<oi�$�"���F�-�F��.������e�Z:�M>�.�s=�ӹ���&TWm\�5N�D�\�K8A}����y�f�!�ρ�q��%�QtMݩ����e�;!��^���»Ǚ����v.Ĉ*'��a��dڡZd"z7����ŝ{�Ae"J�=���:��Aؔb iYQ�><i����2E4��l�_���J&Cl�d!����`*�J/p|��5,���Y���t�;--@g᳽�����.��H����$B���k ��\��U���K0�׈6����3�0Q�gI��}n����I����
d��φ��+���J���VV��y?��a�o��~�M�h
�8��Ito%ߵ����%$~�A� �hT�j[��<>����䬽:U8��C�8L�TA�s?�L^�����݉���
jwQF�\+�9�7�\I4^���C���U�9�F01zY�r?N�],n�*�UB�,�x�0��i}�o�)���n�M]����Q�i�+Fo���I�yt��Nn�1*>�M�?��D���_��Z�\ ���
�|�^W#�p+~��R~��g�ߙ"��XG�M�,�v}[N4��"�`�J�,8�fN�F]�nST(��FN��8��GH� 
}�V=��5|V���-��]�I1���\������pN��cK��q��_@"��� '��3�Ds$tE��x���H�|��r�bw�d7V'���ﮇ[J�"mo
[�\�m�؆�z;��g���|h3����d�/���S�0NZ��۰��S�7?��R�F�G(2��~~��	k�����z�؅����5 � �0�O,Z��0��dS�(��j��R�B�(�g��w�jo;�6�f2���,*x�#�.�Ss�<��<f�������_���B�Q�4o��$�fx%L�b�VsR��
���1��{1��أ]��h����� P�/a5��_����ʈB�:���Y��wi�B����2�c��_�qT/uQ~F�g�8��fU�ߡ˲�G�;Z�JZg����klk1�� �ҏb��xp��|�|�]�LŃm��}�+&ޚs%a�����I�o�r /s�1v��b�ɯ��g��"�W��0�1��tu���p�1��C�}��zA^��F���S#����N����K�d���l��02�+�0����I�
+w�C��4��1щ�"��~�dټi�����ُ�]}�>8pL� %�+1��n�{H/`�W�f��X��9+֡A�kZ��:�B�j�
���1|W�	�+��Z�b�aq"yV�91�P�B����T ��k4�h�F*���v��yVi6�:&}�����8��RO��2��gV�覫N�V�U���H�d�ؗ��8����ə��x�sJ.�i��rWU2]�Ŗ{�Qi�)[�4t�:�u+�	d��I��'6�"�C_	úZ�0�~� n�F0����.n����v�m�b��2R�a�W�w�8-�;��{ߎ��͕�-�T���$��p�z���'�A*�Q�e����@Yw9ߋ܉G��>r��{1+���j'U9�"4�'+��f�c>�j�1�j�O�A�tQi�q��q�V��lV}��Z�F���c�3���B�$�� �ke*�oA9^0_p��`��%m�5��Mo�I�P���usY�Dv�����ۛYM��
r�1��9����]c
�#;B���a~2��Rz��[	*,�!s �}�����Gd����<p.���#��\����6���dcj(�no�����Dv�E����HM}��D��ޜ�L�mI�=�X�B�l*%�_{5�^��t�V�K�̖�X�DZm�y�m��!� $U��P�� �CO}��\Ws���u�ֈ����Gc�+�$~C^H��79,Vڎϙ_Y%ec�_��Sz��~��y�X��W%� �;fS�}(�^z�K�矵��c���왲<�̧VIi�U�����u�}+���Zh��N�V;;cwW�P;a�=E����TS�B�*�~�u����t�͞j����{�Oqv��&�V���BE�d#֨x�E������	�Pa�����20ڤ�n����S�Jx*B/�3�(ja ���8a�r���\B�rxS��`l���z��F/��w�� �S���Ũ*�B�o�\��.�M"$L�`|(3&�X<+B��h���#��n���Q��;��@�{B��h�+Jb`R��.l�E<�7�=\?�@C H������`��V���\�V��p�x�sfk4�\;?�ap��o��5�Ǧ�t<�*�c(����$���M�������Suj�W�J5�V�E������Ƽd�(��Z��i+!UOU]-��x����I�>G���S�������[�/��5o�I.�ƏŌ� o�48&Ӷʬq���(eØ��~�^?�t6�ܟ�)~�����o��������'Ɗ���0�_�D�]Ҷy�Y#'\���9l�*{�^2�A�q�t�'�;��6|bK�p&��29^��w���l����<RZE:NL�ծ��L��M.ٽ��B��|5��N�B7�Q0Y^�����4��P��N��l������_�kO�
N�|�I��J�D�RP9Zq&4�0���&�ǰ�i���k���+�'�>��(>�py��F�k�ک5�����̚���U��J��;UBe~�]�|:AL"�q���0���\� ���~3���BǏ�;���,���_4p4B2����W2 ��s)��uǒ�ճ�+��\S����n��}��+>�A��.�����B�PHR�r0Q�� �[�� ��Y��E��Jp���Z���,�����n�(��I�n�U�1�)i�ǫ>d�ۀac��t�ʢ耪����F�>���7��ӧ:���߽��t�bxS�J�����}޿Ȗ��7$J���b����l2�D�t�h�"k?����J������a����r�7.X�0�.,�K�9��M~�({��^qR�u��S{�����N��_(���lsj��_����"Ƚ��pܰ@n!�@�D��������5�2�h�&Y�
��E)]����G&g/��Wh��܆��7uć�︩S�p�5�Zk�U�"��� �b��J!��U�o�Z�f�v��+Zx���h���>dz�����g�̗��F�Q�
JN�̰����V�{_\���(�8:�葐@[�r��O?){=��]G���E��X��^yR��� шu�\�����	V|�O�J`8 �.<�T2���J%	�sꉔ�,��8n��-�X��3�NLF\5	��NGt����(
���~�.�v>bi��I쥯��\��H�:��'q�"_�.&��R��Pm��<)��M�fy(������P\pF�]� b���(Ѫ��;)���-�S�0��sQK�O��B�#1��w��A¤?��$�
��c&Q����.C�wH�q��d��id�DқFM}�@��y;ܜ����CY�2(g�R.��}54נ�0�y�L��N>�*_$�o�[f�X2�x����Ѓ��)g���=[cȒF�4�Pq�e��k�b8yEHN�����1�����{�VFg��}L�]���O��̡d~�<���vt>����D{�ץ��ά�H!&"p(�G��34�rQ�Х�j�h��;$]��p.zJ	��ޒϔ�U�(�⬕x�^�U͌���n��I
}P�'�:�bY���f`M�z,:"r��k�dN��C� `�72}��u0����u��$��]�Lx��i��*Q�oUeDf����n��t�T=eC�m4�H�;(�P`��nQ}".~NF�kD|����V��{�5m�-�X����ˋ�� (Lf�'c�|0�lI��\ă@&:7J5}A����T����÷����%��͸i��[C:�S��[`˷�1�/2�s��\���ˑ%v�(\��
Ųx�y���@+iH`��(ğ_�V�:��-�{�u-q����^��֒��]��3;K4���Q�D�Q��^�	��$�.1@��n��������x�TVK^�.���R���鈦���ߥ{s����M0:��a����i���!�j�Wc
���q���1e�+�'�A=#z�%�A}�m��Y���*ˡꛑK�^|�#*�w�V��׬�ك�b�6@b�Y�&�g��BT�x.��;�dNQ� ��E:QJ�m�q�cf&l���x��m\q�DBE����\��m���E��Tg���V��$�aI�U}H��|�P�P8�������V���'�(�[�UW^6zmΖoj=QG��F<�Clp�p�D�ռ���%?�|��Q��5ZZ\�E�g�{fƍ{+A��F���N00�qcS�q�������*$�#)�����T�`�	��d���*�*�a�
=5�l�t0�Ȇ����@�۵3�#8�-�{�z�U=:��#�uꢉ�Io`#���	Tۓ�C�yx�y2C7�E�ZWY+��*�zy�Y����N|q	��i�t������楁�cͪ<1&0�{Ns���"�����e�G2�N!|S��(����N&��̫F>C`+�C�{�!pi�4�dTG
J��G�I�V�b�w^��8tUY��Ԣ5�����1h��ԙ}���W/0��e3L-�	hb����x�-q�����m�c�\��X�J��v�+���/�8n�3��������ۯ�ȷ�w�9[�{������β����;$I'�
x���I͈���t��{U�<i)+�Ԓ��r4�1��Y�py�咑T�F�X]+%�͝�a{{�8����6��~qh�\M)�%� $�h(�(}ˤ5�m���MK"���J�s���d�u䥚@"M.�����	U^ h�H�����'��>�َ%��ũJ���]����x�Kf~��i
��qK%-����U��JW�*�Nh�}�ȍ����"�y�����ԍ�s�r٥phԶ��l�������xvbFeM?=���'p�Q-�3v�[��W�=��@��Q�&"�������9A��a����\�xܗ�4��>D<�jB^u��X�d�(�!�yf��������u��%�v<UcPP*SrJndH;$w��>��#g;u�y�WJ��klAsCш�rЬ�/ZZ��R�h�aԗk��ħ%�Ϧ.�2��fR�HB���X���-fio�bj�y�q�����IW�ה �$+�[���Ə��Md~��b�(:��z&��t6E��[��3n��S��:kI��n
����>��������眚[��5D�N+��^3x>��~�����#�6�xgIR�	F�}��B�>�c���н��|,*�������l�!B��!�3A1C���Q!����2��'Ő��z_�K�L)�O-�-�:/۽i�z�����-�D-�9u���ܓ����>��$�#�L��x��}_hcDO��h�#���.�'A�̊\ޮS��)��Aޮ� ������WtM��e�-%8�L.~�UV�Ö�J����bc�k��$�����\��ۜL0�
�4QXz������<�b�@alI�L	lҞZ�y-޼M�Jb'�L:?��P
S#Q�[��M	�}�<�L�N
�?z�;i������@Oㅴ�UyŠ}FY�Gҳ���݌�6�eq8�����$
<�ry���p�;I�Fx���|����z��r�mR"�j#9�:����z�\�>0��b4���G��|pb�u�2G�&2�B�mX\?��93�����Fjq3�[�-�\���ï�&v�-?#�k�!�h�&�'��F�tՒ�l����;VM�dK`}��X�6�1F/b�
�u ��'��p���X���G2
���r�P���o?���SN\ݪ���H��� 䤍$P�y�Ɍo�T'�^1Z}�~�Uƪ ��f7�!�p��og7�P�v�5�(Q�D���C�b2P&(��v����)�GE��rx�9��U�l{����× �$?"g�;�FL�S��R�!*�`�(�U��"#uY�#�~X�X#��O��(�LQŉ'�9:�^U�F4�-����~�|�Э�/�Q��x���n9�C%VDx�D��?��)�++�b�V�^��7dp#���h�RRo.R.�Zu3@�v��4<g��%��?�⓼fC��Q�>��r{{���O���@6�ݶ |U�o�-2��ibٗԨ9�n_Qĺ�+�#+�b�`@q;UӲ۩��H��۸��W^ݙl�Ѿ&@¼V�]�۪	5,~ݢ&���T��/��s���yt,�v�l��L=��/awKCn��ts�x��uQߋE����D$�@�,H����'R��K=�����`��%%J�e��8�su*�4|�}����-��=Ę�$�B��4U$v�����+�{rm I��B�"tG"2�~�͡�Q�޺�2Sp���k�zPe%�V��o@�ɝp�kv���Ω���a�D����rgar����]=6�= ��WD�;��X8S ��9v@sU��l��mC����BI�e��%����K|f��?a⻭��6��at�#��l��"�
���`4���jE8�g����h�� ���&E���c��ͮq�W�̌$G8���.؜��!�����lױ�����qdӫޫ
	��<:�/\jM*�Բ�姇��X/�:�5�q%�*�kֈNL�sXKX(�e��C��lU��>��Bd���ڙR�u�MM���*�͝Ƚ���ɈI�f+O	zF},��[3�¡��H��ٖo�?��y�JqQ�lTli��PHB$ nf�)�go��g�p�D�����7Y�A��T��/t�k]�k'<4H�����swd;@FE�!�#�G��m-1#�f�j���]�����-�uT���2T�./7f������"�b��,h��H��\�9ȑ
�bs���j���4M�x��!BO�:ɰ�Ϧ]4\��E2�#J,��rv��(�V C�j��h�HL���N΂�QB�Ad�}_�\8�Է�{�Um�K%\����:�������E1��0�Qq1:��z�V���.S9�`]i�°t��!�;�%? �)S��TPJ5Y=w���Py��)�k�h.I�7�q9b�v���]6o��`����u��eI�~�z�#��d=����Х0�M��ji3��?,X(
�:K�s����b�0MB��S�O��g����Ls���E���;e|q�^'�
OI[f/u5N��Z-���ett��̌~�fh�=�߷�}G9�b_� ǁ�iŧl��o1:�4����
+�t��z^��φ6ΚR�50�:��.�G�S'R��0&��_3��DwZv�jsuX�ⶄc6]�h�2k�,�洩^����5���6ԧ�;���j�8U�DQ~��"B}��\E��Q�Rv�����ٻO�*Cl�n��fRo;����G��"l |Q���f�E�s��?�d|�]x�~(�ܗ�g�{ퟒ�j�2���_��Ԍ(��*�W�)X�PI�BA� j���N�h�.s�&h&W&��*\�s*[�g��GI�����@�įH�5L�
��g[�5�W��(� $������W���?��
�3cx����L��̿����[�1��|��D�aS�
�p(�a'tA@O��$�E��D#�	��xvA~��@��#��f���WW'��U q��*=�-:�ʜèP�������N����4�nWĖ�{��[ff�o�J:���d��kL\�cv.���~5k��1�(�O�դ��4+�89�l&�t�9�ЪC���ww�Bڊt3M����<Wf��j�?"2�cE�`�g�����Q\�m�v������u���o��X��S4��w�$�{ʨbkIN�/x�ؒ
T����&���π(�X?�A����tª�<Y��b+��R]�m�I�����Y�YF���1��5��t;�"�F�LE`���� ֿ�������1e#9'�J�-1�ɑ��� �.ZV�?$�n�v�O ��R���c1C��$	m�o����%$���+)���äluN�́�ۺ�3��=g���{u��iDa���6�sc�����$���h�t���F嚨PPT�H���7�x��K�O�H`���p��8�������u�fbܱJ��	���"�xʟ��!��4%��腐��ψ�+�GB�y�-�8�������y֑g���Q�${�C-��򼌏�d���tg�ϱ��"S��U�f9d+�ŵy[�uw��S4��¨��Y��R�r�Ppv�*#q\��n咔��nAE�ƚ5W��Q�x��&���P�T�gD��������\E�wf���b
3XU���ŉ���;��uڢb}�����M��|TA��!���]�Hǧ,T���5 �븿�Rx�s�Lȶk(�+xD�9�	�[�NrhO	e�`�Z�����U'��B��;pƔ��"\�'��A5֤]����u]����� ���&0���	�e�k���ƍ��o/{8�A���1��!�*�萿��A���&���=�?��\���L3�\_��q补���
Bsk}V���v�����6�*C0x�x�9W�T�4}b4iPU�J�K.�|�*��'~�s;����u�"��!������0ueU|܋LCX��KJ��* ����&�����hCH�B�Q��eOW��Of�}f�TN���5���!����:p��J��7S����{<?a�P(�;c���#rd�G5	�ph����	q��j�q��߯�BcrP���1��;-���
�޴�� �Gi����:��v� ⴊs�#���s�,��&8��2�o�٧��J��v���c�n�~��ֵ��%{��wy�d�˟r=��൶�����?����1��㧗Nes+��aU��E���a^�ڪ��+hȧ��~�$��òB(�_��V���/젨p�����U}��7�^p���(#w���x���@ӧ-�=�=�㇫��"ZԷ��aд�!�|{�����wm���M�3�0�gl��\1���_RT�E��THVDX�j�Sa-�j�#�'ަ��TWj,Gm1�%�V��r)i��M���X��џa�m�m ��$o�S�ѐ�A9�u5kY|�զt�'�GCh<d���)E%ޢA'|�@�͈:u����(SK�+x�fy�{��h���s��^��TWiyjߗt�r~��+�NE.bZ�8M��@��n��3�dTB?��*�4�'��m�3M**��F?
̔��D��3>�,0��_�o5�p?e��}Jf�4�����g��Q�}���U�޾��|����+�
=�6�C���P��$�lPr�+��9[\�������:w�=Z#�P�{qd�&�D�l^A���&�%*GR��UY7�8?e2�lQ�f�@Z	��eurj`�,J�MM�W�O���/"��B��P�c��u�{��a�Z���q,��P̟������&�P_�C��s�0��w�l$�� ��g�"�.��m�ս�@{<B���tx�"��z>��y,��o��Cs/���RT���xȣ�-��mm�ҹAy��oW+Aw�ϋ�w����d98@��.��W%�������6C-�N1�k+�i̬n�E���'�p����0�pA.<��%��[�v�j;H���$�w�iFtB�3�'��b|�N� 5}���2o��$�H ���bKh��e��È��q���IFQa�Zpox]���!{�FZ�bD�������H��������x��y��;�����3����FFR�i�����7
�9;�<9ͅ4�}`�?���Q'#���I�1��'��fO9
М�C�����.������\H܃�n�x��R�@�l"[ֳ�J���#	_D�u�Ib��䘷��G��{f�?�,��f_1P� ���nSVfm%�<&�f��;J�SA!S:�%u�N��ӹ<���C�.�4��7��� �1G�����6�q٬�� Q@~�>Ý�C��~\>cA�|2Lᭉ�JPU裣s��c�����P�9�:���<��d�XRBT�����A�6��=�x扠���8��P�Ǌ4�J�	ؙc5��a��b��uC/VB%���%9.|�s�����]{=���� �᜵y������|��LMs���ZO�Q���51A6<~��˿�y:,�(�*�2�Ԟq�뷴�R�vɏ�ױs/U��5��4:0������o�;+���.'�]b�'2�H�~k�j�g� 2�UB^*#�7��w{�	�!F�S����Bm��r��G���ۨ?E�6�hK^h
��bk�!XEoQ��Cg��������qK��w��s��ES�Q�t��'��m�N'm����
�kǹ=*�C��6LQ���w�AiT��~��!��<���9ǣ���|7��n�҆|Źs�i�f+Z�yE5m�MUt��n��;D)SY��{;.Շ a)�m^�R�p�W:}�U��k�=L��	bY���`A�$���.��c�%/����DudO^1�G��g0B�k*��n�q������t/�q�u�ۈ%ҫ��=��H�5���|�ןzW%�w�d�'d~��''6:PZ��B]dOR�8�։��� �zH6/�V����S �8GX}T}�W~{�L�������;���t��D�^�.��j����;����
׼���_�����abO�K/w����	�p�ך	N��ɬ.q-A�?�`�D_�o0�*�}�ȝ�EҴ�V�?��Ǘ�� ��/y��O�^P�uuU�=M���M2d7�FT��h	�G����g;�T��Ӈ$A"�Xs�����-&.2�������[]F�[V�g�ѥ�i�?�c��Kꉫ��;�㖍�)�m����x���(���z�Xt��?�l��-Gv��"x'n���ʩ}h��\�ia�"?3�79�`Og��atr:�E5��w�8D���և8Z�B|�
h!��i�b ���m�����r��IʱA�Ji�Q���x�N�Ņ{�����\j�Ҿ�)�A�~V�R��bdfiH7�E���ˤ�����9-�X�l��zS���`&1!Vk��=Jo��AG�!�	��"��2!�?�{7o���>(=���0�Ժ��v�X���j7��:�Dd��1!ZQE1ӡ!(R)�G×^#���AC"��V���F=OϨ8�&��p�@i�.�bqHH�
�>�[���$5���v�a�3� �����Q~d�����_^�Q��Q��Xq�V_�X4��E���)0�����0w��X�S����P���b9��kYBN��6���xr����d!�Vf���#{֛(\V$�D����N�GQRI_FvA'J*<�,X�0f���b�j�^�Q�%T����F+�2* ���eS\o޴Y)�C	L��v �����|����D#��˻�u����;�i������&gjǱ��ĺ���$j)+���y9&x�.�-W���6����4VF��������X���H�~�;l?_S�OxE�8�2�Y��W҈����Z�ftG]7�W̿���n�]�����,r<FS��`J����QY�aT��|�a��Ż�k/�UKKtK�F~_Lm�qM�|����\g�+�x�❿Umy3c_��qEts�)%��YJ3��ĩ!s,���24�0������Q`64�bE|$���Q�2�F��*�i�\�gǸD�_ƫ,_@:�L��loR!w��Z�8�[���:=�z�Z��=��@��j��	��&����/$�]N ���D�mk��;��r$ݮx5�9��������M]ti������tR�t�~h<;H�Rʿ �q_��_��N�R���F��,�y;������;!D�<XւC(�]WJ��,j�o����'"R��6DP�	��t�=x�p�3�
=ԙ'}�@�Һ#l�i��$@��i�]�t<���߾��ĦC��`��f&�mX�z�,�4t����.�y��K�MG\�a��Џ��5�����E�
~3!�&m�a�1����g���np�wH��q2�����<9���5t�\�ZDO0Y,1Z����l	(������S�ud�薏���Щ��ݠz� /���(��/�z��@��?��u	�.�=������c�\��b��[�'"ã3��.�FuM�t����?��U���
b��wb{��v���O��2� F�s�"weF��9��Qg����ҵb*�Gh�74X� m�җk�_ʣ8�!�ёP�w��q�VWc�&�� cM[QӾ�g�Sj��{ee�>�0�I����JC���"�=�~��&A@�K��f2�oi�����@Ǣ�TQ�W�>�X1���<�T��l~��6 ..A��b=��'�d�l\ꌪͿ�����X-W��>�p������f�=�����%�'yt�� y�Ix�OJ����>���<m�ql�	W~\�;�n�	�y�Y���&��s�Ϸ��\e��G��^������7�F�XO�Wa�!�T�����Xec�7{r���E�/��A���+�R�}Q�J03�@�̱�.-Ċ�dݪ���+Ho�m����������vP�\���K��@�v��3h>4(��$�|��<ul�4�
���ad�ڱF�y���q���d];�p�<s�ÓO�+د:��e2���ޓP���&���t��n���K��c�u����;%�Y�ɺ�ϭ~�!3��[�2��c�ӂį�[�5�VΟ���U��`��x.J��L}EE�7U��G��
���KL7�0��{{���*��(e^�=��JXbp-k���7�F��7ĉ�&�E_H�
�RH'M��Tw�,w��f6�Z,Ε��s��˘���A=���H�=�$)zi��7�K?p����Xĸ��"{<kW��{��u�N\5bd�ɴG�p���iL��Z1#��*"V��[u�B!�m����/c���h�Q�_w����8ג�E����	[/afJ_	8���!�r�r����z�̗ͥ�M�w�mZ���آ��f<ZS	olL����,�iV�BG5��]	3#�>��-��,��E�t�!�z��N��S�|�X`J�u�R1�id�uZ:Sk-��,��O=�6�T��w�;(�iȖ��G�)c  �KM.��uI�Ī�OT�����=�����']!ѐT�O�l|%S�:�K���9�Q�'��/���x�3��i�u���u��^C?�r~����âͅq�\3���֨gu ڻXK%7�i�!�LFO��/���Ǐc�e@B�[��}�����~��|���1=�Q��y�N�����w�\ �+F&�Z~���ـ���c�$m#ŕu��ֿ�9,"tI��i��2Q'�ћg���N�����e�s��'�rY/�g��衜���O�[Z /��z��.���^�$nܭ�Pl��ƕs�����^@$S������Xhy�a8{��h0��⬼��j.@�8Q_'\�fBs^͛�.�@�^�J�m�^�b	��1�g�P[Ʉy:��͂�0�Vsic��d�bJ�U�B�f�y��^l��n\�T�m�O���N���-tcN�?�a�"��d��r��y����w:�ȋ���!^M�i�e���\�jC|�b�]ݖ�ZA�rd�<����d|�^��b����U"$!�M0�|�o�[2G��;M��NK�����yÛRE��C�\�E��4_"I�^\�B�2�Q����X/W��R>!��R�ˏ�:4����N����P�]���J�}$�|�U_-,� �n����A:-��fĹ� u>Ӷ�e2����;���,�*X�Z���kr��,w����.9�Qfz)E<�V43ԑ��VQz^����-c_�@�囒|�r��<�*��,ɩw�n�,��]�ܭ��������b �̳�����$$�V�0������4��G�CK�'
��j�n�%ϭ��W��1S�P~م����]�u������=& 	�c����DO�}}�GP�:�#��o"'���Q�Q�6���g��w+'��e�F���9wBr'�S1��#�,�}q�(�4�D �X�,@w�'5P%6x۳oF$	��4ϫ�]�Ӧ۳���'�̐���V� �;�ÿ��� ��!��7�tl��PC�y)vo!�[�X¿���V�Cz-��i�%���4<�.�)���ڇ�HƯj܇m��u��);Q��]�Y$��7���P�a�[�.����8���q��t�a������2����LPϱ�����3�7�
 ��rR�J�Q�tw��@4P�>�x�`�R(�g�����m�n�u�+`�u����z�Y%�����v�Z�pIRC��O�P��3���?6^m=��>�WnО?�~�rp�rͪ����~�/+�"1�]v1�?@�\�;%κm�"&
��MF��)���&o��|��ʸ��>oSR�.�����V�4c�8'f;�k�yp��\��(9�ދ�Q��gf���bx�3��U��0��>H�I��ktt �v�*��p�΀�gf����q<4�3o�{_*-�(!����Y�pX���}mm�N��r\s��|V��������:e�Sղ��BL��1^H�0�ZB�Ĵ�c�߽o~@~��{Q�0�����+���Z݃��ɂ�m/��Q�қ?ިX\��nRX����w|p��z��g� /�I����clj�U���?�.�y��.6*�c,����N<��n��������������Ox��`��KEsװ��}�� 	6)�p�o�%�S�#��a�=l*
M�,�T�^�\y� iдc#��}��4��u��N5u3e�y��	3�ˤz\M�*��rDdp��T����C'K�1�8y��ٞ�/5>�$%�~���32d]<v3.��-��S�Mz�Fظ�f�#Cl���z��p�	Ćw'¥z]�9P�aწF��Y�s��P+"B�����l�/���N˙*���Zcn4�H��Wѐ��Lu=
'j3AZ�]u�6R��:i�{0���(f8����C��`�cW�7q^�*���Y�kN��P�S�V�/���A�Q�[.%N|;R�Bb�o	���K�8�������3Q����˒Q*�1-�]͌��̝�ƼBZ,RhVt��w7��teV����W��\�F>ԶP9)N2��߷T�;�i��m�����0�Nr�3�e�e/f]!e��#�y���(�
)@��EJ"`��kQ�9����s��o������W*�;����%`FP1#�̓��-\��\��܍�Q��V��{� ���v�Ǣ@�Ԕ�-r���w���Y*ؽ¦`Uf2�aN�1�a/'�TkZt�B�jiZ��4�'Y u�Np��>� $�*��<:^�S��]b�>�k���f�>&ç0������S:Бl������ �Brv-G����"J04�)+s�kҁ.;>�Ǒ�=�=�-� 
�a�+�z�����"���<����:���o�Jz�AO�X
:<�M�Zq��7\��;O��l�|��K$�A��Nx� �K���M��薉!�X�r�@?���œD���[��tpF�����:��ϫt��:H�<���@�5aT#Po���܇m�hV!O?�!�̸�0��F~�v��n[C]TL�N�1���A�:n1����z؛�qI�>,��_�>�8}��O��^/Y���jS.Gi&���8�Zm�9����5V�nu����4�_�߻�%h��q���:�?P�@%�؉�T-�4d�%���!�J����_���|R��I V�f�p��ꛆ�y���:�z�
��OU�oa��V�Xs�M�9�G�z����I��:/`������Bm6�6.8�t���	�<WkY�ZD�U�2�N5b�z�L��6a���r &
��̊}����U�u��j��&�x�z����Q�{�gJg%�ת!Km�c.e4r��Y�2�C(q���t�q�0ny`�g�����[7�s�E2���&W�ˆb�Up*D*�%W

��FS�\�����$C�Ȑ�t�2,��>��^ߚ��_����Gſ5G��{L;��\B�e��f�"�3��(3S���ܣ9 d��"Ul�W���r��S�]T� d��G+� �tS��9qCEe�Qu�Mg>�tP��h��#����E1.�Ha��F�]�؍rÌ�����J[�砋�3D�|CI�q6�l4��A����?N�z�\rsdmB�(g&��݅)����gBc�@����qͰ1��D����YP������p�'�.4�%��X�S_�ڞs.�E;a��T�	���:�+�o~�����0c%�C��>@n�����^�& ��������w9gL�ʻ��W�����v���	%�@��o�䏝ń�4)���C��܋�a��B����c�
ٷ�W&���s	��H�vYdДR^0ly�Ɋ�"��T�� bU��`���+m�t�o��z#�7�:BduP�v+v�R���]1��U�V9����Y�Wz'f�0��HZpw��f=���A�4b{��>c�6�>u�)�z_�lDcsI��S���c��G˗f��֛��H�*��N��<��8#qe��m��� �|=,R,/� �H����-@zLg�j�%�����фb�Y���3�9,�A�YLu�b=�>��>5GP;���/�D1�k��֖ ���\�E�V��v��z�#��7@[�+����]���0Ɠ!JTu�?v�պU��w����4��˯���*ú,��H:Uї�d�zI'��s�����xv��7T�����G]����z��7����?.euWR�Ԍ�p�f��6F܂Q!����V����׮��K|��?��k�|�[4��0�t�����S-uJ����go/�����v��3T���_@�]�ecOE�E/��p7�j����`�P"s����\�1��>cp���MOS-F���^��Ɩ��,�u<�E���W�Y���P�~?��m���P9�>�`�p~�Z�bC�'j�)XΛ^k��2���b���>�x��߾L�q����J�y��L�B2���� ���Ќc�a�d���
��a�v�DKȱذ�	�������P�Êawh�/����AH�O��<�E�hB�g�ǵ�*֪pO6y�'�������9�ʫ�����dY�O��gs���;]������yXAۉ�����l�5�$k��A�b-�R>�8��Q��-82�;���/��z�\XTZq�.�%�a�Q9�� G����Do��k��稸7����)y2� ��{��G�,NK3�Y�P��𶪁CM߆.f�'��g�ͫ��́}��x19>c6����������s��5���ޛ9�bj��N���o���}���vO�lA�_Ʋ���p�Q���<nX�\�˦E�K����Of�녂7�����\�Y�2{܅�PӂkQM��-l�/�]���.p���G��ƪ�~� �#��wE��i�� �g��~(�:����l*�s��l��������L��ֵ���G��������c]�oH���:?�Y���6&�cC��
T8���]}���8ٸVkJޚ�s7aj�g���q� `jx��*dga��,���V����ؐ�c;���a4�d �#���-�h��?;R+M��d�su�*%���v��s�x��0H�n2P�T=��jj=f(-����EQ��]�z��&0���Tz�C�0���|��C����>��K������x��j�/8"������
�N����Y	A��� �*�!%��qƻb1z"J]kĞ���\wW�u��ci���K���J#DfSb?N����'n���SX[�9��e��ы �kC�
@���_*������B#ץO��r���nܞ�
����,i�ZZ��2I����$GY{���T�ާ9�b7%É�YW��(U=
����B�C�.bZ;�=v����f��A����?��k��5�R�t��yȕS ��Um׎�v��y:X�V���p ����	��]m���e�뜽#p-=rn���vv˥>���M|mfZ���Ei�}�pf��w�&��i��u8k�Y}��[u7�GA��'f�-K�ovUk3"�G��+n��y.��]'*G�Qd����<f�n���&ؖ�xQ���b��<�иD�+9������{��5ZY~��~�<��!}PL���)G
�h��w�&>��8*�� ������0���C��}"Z��Y�ެ5�����ף������oÂ�yk5D������C.cb s�#�+��䎏���������h�;�]����$o�Z��E�3?L��9L��M���w#���8�Qe�J��O�U�MwyD�e}����M��n_`��{&�V��WF���Lz�}nV�|��Wb����02�\�����7����BNn'�ow�Bm��k�"x*��6H�:}���w� ���;��\�/&h�N<`��d��S������}��ZQ� PSP�}�8�{�C)&�1�]/q#�4-oN&�*D��s�L误v�q0����� ���Z�&)�H�) ����(CW��z˞�?�έ���)��3k�n
��3��qUH�������ܫ�c0�DZ��t=�������<�d����i�6��%���od�jz*!�z��`��p�Z� ��?�в��y��B2^��탓菭���*��$����R��t��Tn݋@�$cJ(���~;x������RŌ�r��Ab}�\O��+c�s�BT��~��mj���l"�:V��#D����/�M�k�y�}F�j����M�� wL/��R���jŌ:ȋ�n-)����f%�3�»|7l6��x�����S�}Ǯ<^}�f9������ђ$��N������z���l(��o���	��QT�O���õ�g�φQ�=�t;��I��[+]3�Ȉ�j�%�yUi0���`R�S��=s�I�ҰtsjR��2��-]�Ҕ��Q�I|�爧d�>R��Z����+�t��6�@�$©-Y6��J_i~� 3��Q:d_G�$w�x5*�پ��J
�r �O����EM�XQ�+���� 7.s=��s�e;���R� �3�4�-nK-��K(��*�ܯ�.��]��Y(��4�V)��>��%����"{���K%|�Y�;��T]܊�������)⺆dM�(&v4�ps�W]
{b��:�|��yCĶa����X�Td�擝}t�㺐/cf��mM��f
�Tu1�V�Ёᇮ�v�t(hiu�]��y��v�߿��,�
"�֩�
�m�/d��P���������ݜJ ��G��,���O�~)��*A�򺺡P+�E-�UW�k�A� L-4�,>CD;�­C��=���x�����eKx�L�l[�7O�G�� �4(6�	G�m�^��o��%z��՟���v���� Nŋ3*_���������Z��:�P���r�&OmO�����J���
Q���X
��������O���+1Š��+ڎ��v~���`τ�0t�5 !�|"8�<�k2D��	L��Ƒƞ]Ip��-#��=� �V_���ī����(Acap����Ś�	j%��T�I*���eͶDr���	���=���V{�{��0c�X�j���E��Z/��I�MB�G�*(,�Wh~�Q��#V���3��Z���*�
`F!�[�s��:ƣ4��t+ф���{��tM�� A#�e�#�맯��<���/���{w�子�h{=��D+�M�\�6O>�Hh*�����q���pL�~�iT׃�� ��nΤE����n�
�P�sRN��z��ˑ�*&L��Pk�+�;X�o��,VT�m�#w�>�q�&u�k��ʹ�/?*�|R6�����|�p�H�����)�h��$�Z�aZB��|&�걧���T͞(��K.��m8d�E8��Jp��'�1�_Yz�[�W��H]����M�7t1|$+)��	P?���q�R�+&��\��,U�v�d/�.p���e��g:e�z$C���V�uB5�����N<]�I�N�C�D��4S�C*���ɽ�ҟ�V��8�\��c�h�i�.����f�_����:�Sa�C�
�t�l�X�!wkB	䑣�8��M�9�R�oC���=�[��?��n�n��ν�ҽN]\_j�˞�DC`��:�Jc�䴳�(z��)G��zj|	�r����_*����,~g�I�6��w��]G��)��&����H刨%�&��w\b������k^V�"�x�T��KAE^�(i��u������de�j�^�rձԨ����z5�>�"Z+�7����vA������'=����R?��`�1��ӧ��[n@�����[��k���g�N��� E�3�"c T$<����4�.6X�ۓ#c���d(�a�����dd������:~�4��[���;���,�wȉ�A�
�Q����~�4�Q7:4�{�gJ:"����L6��Y�+�K:�r%��6~Z7�������W���y�F)�E������r��>�7��.'��� 8oѡ{��0�C�W�`֖"�MG�H���E?���|x9�����,/��eoM{�:v��������[)[ |�X�=�$���[��M�x�{3��
�-(9m�6�m��'D��W�w7���lweNH�i%C��H�F��+�V��$	1ң�>��_�3uZ�pJ�U(x�����+����+^^�RZ���C_Y��OL|�J�
�3�_bj�7��E�Ea0w���Le��������DM��-�K.ՍuT�՛BF��4Z�f���]�ϖ��ϵ�Y�]\�I|���]Gb���,�)gSʳ�ז�g�}{��f]<��/��l�܎�����]���(�h�KSp��B��f��<[�}�����wc�_/���r��fy�1����_#/��u׍��kt0O���
S�\�1�e#�$��~ ��%[��7��>��F����v�^.ݳ�3u,���ԺW�q}��^�=I��rQ�Aۂ�n�@I=�g��h`�]��9]2vUi��R]^,���#�3H�?�-��3�H�ir!�J����>u�����74�v��敻=N�"�Y�yG��[D`�r�(by�)83}�w<���%� �E�w*���L�����:?QR�f�'w�L��%m�a��r#��7-nɏ�΃�!ʴs)�{6[>r��jj��"!�M�gO[�#f�v������m�D�丌 	"�#�o��ĞNE[��-���8=�
1b���<�o�~蠞���|Xo��y�Q���G�k�nS�S)�X�n�+nA�*[>�ﵳ�3Q+�
dU&_Vŀ��]�W����u���������slσ|y5���[sl5�Z��=�#iq��7M�?�ۻ@�m.���h���>�p�x��F�Ĭ�a�n&|U�������n
1�נ�X����=P��M�;5��X0�b7���Y>�L�[����Wc�-���.m]�{>�}����$�l7�TCQ�:�΢*��x���������(TQG-���;V��N{�F��>H��sn�	'��):y�qy�9/���/xL���?��R�E��[�΄/1�s�?����t2ۖ����|~��(�Fs'�_����Õ�XW������鰠=���coi���bh՛��{x�i�Tмj|�n ;(1�IO{�
ϳ�#v����ܔ��ӝY���I�tLM��y����pz���KU�^T��r�f#�݀���nW�.Y/^��s	������6�&��B��$'��fi�y	�9%�H��|�}V�ֲ&n��ĥ�(��A0���)��xR��rd��e9It�^$�{L$}���_� ܋ޓ����l�"���N���1�m���j%����<N�m]"x�S%�J@����n�2w	�<S�Q!�P��T<w(@(C�dob3ׁ�(@��ȥ�� �n�_�]҆��%hǢ����~ӗ��<�	*MXu3�;[���',u2��k��a�˧N�5�e�і�s��:s�2���}h$\���;�+C��,�{X!�}\�Я�n4������	�H��PV?�̲�f��Cv'rr�O+�\���\8O&�MD�V~Z8ڞ��H��3�s��� t���Өo�c���^�n�G@�����5Hm�r#��Y�V	��k��;�1:�ܻS\��}W)�MðG����+�lBP��y�^̴͞�16~z�5�&�\�ѝ�}�֖?M��k��;�t�� ��QYv�R;� �q��틾,��ͭT�]{�S�䈜O�%���������<j&{�{�b$��ΥAz�9�]��:�K��r���CJgHDQ��W�=��}�x/fJ����qĉ�c=���)�ח���v%;V@aؤ�F7"����9��r�͹�iO<@�O�h�!�K[���P�/����.7B�;g��V��}���74xO�"�E�F{��f(Pb�7#��`7&��p����q�؂��_���x������1��˥��^		)�@�KºP���Ywl�����*��$���(��b�#��P��X���q/��,�%����/�Ӄb�knd'��I�l����p^n�rG�BF� ��x~w�$��Ag��R^{�zv����,�����\2Mֹ�,��e�\r���w�`,��q%\Ϟφ��ʐ����~.�~=9�]�����֘;�~�������ц�U��7km���/#Vԓ}��1���!CH2�q�k���灇;댢n�&^*t���1t��W��	���0�/̉���<6*y�}�YM�Q��o�.��d ����Ԇ���4��ʅi������e!�ї1���Jo����/&�Z�
&�]Y~Aw@�0�|]{B�hЯ��{,�(�E�
y(�<�H����^u�����9��	f��lǿҰ�L���N������RC8J�b��k�|
�u���V ��tf�C[U8�B�T�!{j����8
W)�.S7U���+�ʱ\��r��Yp���t<=m$F�� ���jGM���;���=��6����(7�����h�M�m��$�q��ʝ�(��{�5+2&�����ڒ@]Q+�`#���ڳ����!-�MA�o@�b���Lѳ�6a63�
�����VRH�˦�<�[�-5#�)��f��ζ��<7���(r,��?�.)=�M��69d�(X3aЌ�q\��g<�8bT$��Τ����~� ��1&z�3s�៙ӊӘ�l�(��?j�2��;��O��X����3|9��hA��	n�^#	��Pw�C�A�l\8z-�������#.�mDU:���.�|ߏk��ܲ=S�,>�/��?�H��K���rd�A{L�v��@�Wn*�L}���eR��z��%������Gw���X�Q�,����Nz1�&�|sD]9�D"�Hذ����b6����A"
ښS�^�6Շ&l"z�%�fԒ%�/�1g=S���S)`ԑ_edR'
27��Cal1�����d������4�|״��1s��(x���m)��]�0�NU�A��˧o_͋r\8��xT+����{wr'�2d�!z5�l2쒗s�����gӐ��<n��a5K�	ĉBV�����?����7#��o���5�좮^ۃ�7��3�s�������좺tve�ccW̐�u�G+�m���@F��[�֫[)CJ�ް�(�q�<rA�Y
Ǌnp&I����"�j�@��+�ޓ��z�}�S�zO��'�E?)�d�q�`h��*��4S���D�R��0�~�!ˬUax�2"���@�K������.M�bR[H�����Ժ?��bF$��J�Į�!w-���^y�
��Wu�Ѝyy0�_J���ޡuY4�0�CoL��U�t�y`Q^���Uo���!6�(+\u`�@ga�|A�Rq�Jzu�a�~�}эΐ�yFh�Z�44ܹ�B4^oZЂ��,�7����Ū���y	a>{H�z����<�>��E�A���>����~�圣��qIm],{����*8˔�o����U:�.PﾐEY�UO4�⏸X���������*���m���Z��|�0��=��i'ȐWO Կ�t��c�<܍����U�>��Cu���CL�̻
精�B�1"b5$�2ͬYLi6ĝ7�g1���j�ɞ�c"˿t�OV�@�М���wz�tw5�0���ȜF֫�Nq�H��������6��*�4J���a�;���`��7��� 0^�Z.���%z��an��j�٫�{>�6Kj�PQ.��]��Bx=�%�z�V��6D��J؇T`���M*���!�f���,EZ�g�荘�f�=�6!t��l�l?	,�n���Ȧ�:�,~��������H8yc%/��Ҕ�E��
"��O&����)/��%�[͢�ZR^p��a��FvN]϶<��='����	�u�i�����9�|��%޲ȹ��[B���b�R�׀Q��r��i����OJ�##A��w��ɺu��L�bl����P�D��\���N�#�2
�0�^��P����r��e���oR�t�tR�����;/�g���_���X��Ym)���PA�5i�9���2BJh�?g��k��Y�BP�i� �a��_@ѯ�H�)?�`Y��������3�8�Z��K�8�P_o,�R.G-t�#����D�w܌X���cǌ��ܖZ�ۭ7/+C�o�I���s��5!���r�U�'�,�7ܥ��]w\�XY�C��wloa�,�?f������P��v�vaw��z2��!��ؙ�'��󖡶 ��ȟ�"��
�����>�8�IgU�H)9=Oz�wq��݃�b�Bt?�� �/���)��RK�8:��Q�̦N{!�}]�K��5��٥p���9�a�N�� ���w�-��Z���կ.@�wV}��S�[ �G!�3���\\���(�J�4hUZ���p��xH@��O��b>��.���a��r�$r�tW�7�eN�"��>nr[%u���4�헦���<�{��V�����n�,:_�$dHH��s����7��J-5����҈���.�>����<_B�1 &ι�x��=5y"��C�w\r�%�7�r���9V�����O���Ѳ2�J�GO\X����N�c�R�!i��[w�O O�v:|K�g`v��~nu5bQ��#���;��ꁒ�s�h���s �2-�p�7�k�I��fD��cE�'���smY~��Oa} ��Csk��p�p��S3�[[Jn�Yk=��7n��8B�d�'�N�^²l���Ѯ?�po��p��������׆Y|̺��5/#ٴ>�%�e��z�+b��%�`8�	 tOc��HM�Ȝ��7�}�n�m};�@��g������
0f~R���=p���z���|�v*��ۏVƭ_�b��js���ɝ�(NG��c%�B�ty��m������v�X�<�Ưj����R�D3sl��<�C��B�TMȿ�晝��^K�lq�SV��j�04�e��,a�1��0���j"e��2��
l��������i���Q�d�0������Ył����4�B!<�x/;�kM�Uڮ�I���Ʈl���*Nh��W��/��i	C�)��2�
�-`p�#�/���̜�gA՝=x�*-�Ѕ�"��(Kb3�=Sv�z	4�o�Q=⛋�gm���;�2�L�r]�����AP��z?�o_��KK�phg���6�r��yʘ�}�}��_�?��uo�߼xQ����I�U+���W�q�,z�bw���a�>�n�pz���[?�̝m��o�R#q�u�1g�7�0�()=5Y� ���%Tk���遊A�Qn#���h�Ѽ�~m��#���t�xU�r��5@�!��4�!ĄpyCoեZ=��;(d� {��Ǐv�4�$g9J�b �\Suʄ%�Ò6�t5��ø�	��m�1���/�F�Ψ+"������h,�b|/Ӈ:�9�U��y�J��w#
K�ƥ! TB���h�I�`}��\�E� L���J����F���]�M�>�63rUڎ?A$��A���	q��s��r��@��Y)ð����7��Bze�p��+h�.>��$Q�)�I�]���|�Q����5��+��a��a�b��x�� �2�D��݀�e����#|��w���ܘ��w}��b��۪T����R{;z�l#A��*�,3���F���uP~!ϖS�xM��K�V,��	�������ǰF^O\	#q�I5<�4o�a%���ONG����z�%0�"��D[�X�W�����"��RNj� �M�0�����΃�t�"��9�
Ιo���_#�.RIߒ!�/�cџ��gŹ��� %&څ?sb�ŃTYxУ�C+�[��-�/o!�G,r���G�(��:�"GP�n�������=���s��%6q���0搬8�ޗ��q8�M�����j>pR�J�J��ǯQ�����
��W�&�n}0�V�VC�iu%H��R�w���aD�!��?�H�����T�ꇬ{o*9�7%�3��j���Vt��]�L���c!=�e)��-�e�Y�_ʃ8=!�ٓe �n��L����P�Vdؑ�J�ډ�ؠ>�r��Xn�W�^��O�Α��CF��Ԧ��g��3t��J|cG���P�/ I�
)��g��DI��1���d� ^�u5G��vw����o�+�W�X��ak��Ƕ�.>�U�Z�d*U�����t-3c��AP��N���������r�bÝ�s
����vi�l�CXT,�f�ݭj>��F5�]_���N�x�,X��`V�$���"aA��K
�Ќ�9'
\[�0��E[�x�g���-�C�/i� ��6��R݂0��ܴ(k�����U�����FG��z���BI��R^}��.�hhUVk �M����VM9�j[e���s��6\<�G��/��k�R��<�`u����ř��!�Y�A&ބ�@;	C���x(,��&[rM��lY��>n�=|�Mמ���v2G�/m �w�yG����})��G�JlØ����#�hd��+SUw�F�'��E�c�K2���A�O��q��m�j��a^q�ޅ��]�$�
�����q8� ��l��� ?�����a�ªD�+�7��>��a�e�8�q����a0R��ΏkgO:�E�R�Q%w>\��V�~�O�z�wn��ot��(E����~A"_�]M�9Q�=+YT�֝��ઁg=�E�)�#%oF�" �sk�OB��+�L��/�]�I�j
��Q��*NR���'�N$g@H��W1O�= B�I"�� ����c�I�9���_�&��ѓ(�H�Ɣ!I��-Z��`��4Hl~%J����P�EH��$�b7I��v�G���;i�!z�R��"0�t9|F^�\kB?�.K���+m� �w�1���UbT��9hӇ!���C=~����HkƪQ��ր<r��E1�b���&Cܛ.�����"�D���Z�\�2,։3ɑ�%[�+n/�.��T ��b� ���fA;]�g����ߵ���}U��v�d 1Բ/��p{¥��b��!A��wL��胑P��6㿐~���a�'�E��rzhk'`��F83_����ӷ�g.�� f�wcԟ=����l@�����9zмu��>2iNT�	�Ɍ�S���É����V�)d�HLj�Dņg\8s��;��n�V�"2A_,�dG*)w�~�:�	a�v�1��N��?���F��9�\�(�E��|������`�,5S0Ŝ��n�!��Jx��-rFp�̨Ѓh�kJkֶ��Cg{�JC�'��N9�T�3��� t'�<V3� ƿ##�i���j�]�0F��oO�bE�M�J=�H��Ԭz�<���p5���E?�2TZlr�{�u�Σ�nق�1��JFD�W^X~^�7��U�l�3Cw�!d���Ѡ�Pns7���rxq�#�<b7�.Uҳ�)rL4�+/�S���`�ɑhp�2[၌����f|���9f>�r
��W�̧\��5$�A�aU�ӡ���!v<8������3w����ץ��珱���r0+��[��F��������!���B5��(�;O��u�;ފm����@�I��jU�B?D�w�w�<�Җ����y��5���н&9�,t(ٖWe� �0���p5�t@�#4�����>��1g���gS�a�B�#<Z�Ah��'�8`�7�)���4;\��TU�~sӼ
pQ+���f׸m�D�v(aaVV�ō��PM��Z������x�þ��,V'�G?Τ�t;d�?z�s��<�(�'�ZuƜ.L݆���g���
) M�}=a;/:��~4'�D�t`��Vd~�T���߂�<G}3��\~5}b>����:��I�Sr�l��X8tA�I#ь����L��׃�U�
�[�m�����u`�xO��г���Ώ��e��!^֦�L|:A�@J$���!�"�-���$v��T{�R��@�OďMs%^#~Ԯ���z`0T>o��#Z�GA<�"�,.�?DBl�~u7�0�h�������� :(7��O�C��n`�4M��ZsI"��O�H�\j��nB\�P�����I��m	W�<�
:�
�,�t�8E�,P��E  F�����1JMz�>�Ch�$�&�=ہ��A>�0��i�k�;Nk?�Yҽ
	@\m LKy�Up˪C@�.(ⓜ�#~R����7��ٲ��+e�
�DtJ�L�A&�-y�q�>: '�l3��4uȴu$h~@=L�D�I@Bq>�ԅn͇����.JE��H�q��P�9i6���?��n%�������#Ō�m����D_7c"蝫ƣnR�,/I�����&�'N�E'rEG�S�j�;Q�oI�%ʦ"5ǚ1mI�&+��&bЧ��������2���C��:�ʅX;N������h�3�.�`�����E�5��P/cą:p�#�;�H8,����NqQ	��	�,su~�ʀ *��G&����X;I8Khg��
k��$(Ռ�}<%��^;؍犀��c��Fj�G�$����~f�-�Ko\�����y}�5�W�	ٕ�Y���6HY���}}g���Dʃ�{��l�g���~��MI�Q�w�}c�k$��f�MBBV:��2�p�?���I-E�@�R�D�B
�e"褳��e#�x�ÊK�K����G�ED�����P�t�Z:�2��9�6�����a��SPɡ-u���`�Z쏳_�GO+����x�C��Ѵ�r�|����ĝh��OAN��d9ZY�	�Bl���kـ/�,!�k4�K[�Uv$�:A�Gr]A�E�Ŋ)+<u�4�Rψ<�j)�=YLkْ��h@5Y�-�m����&d�>UP��Q��c��C-�#�vC��Z,��@YA��$�G�Ie22���~9~�DʉJ����P��O�{ߪjum:��-\�o5҃#7��w�^9��@B^$Z��ǘ%�Oc���V~��K�%�nOl����U&�i+����w��@�B񦟾�����TD�=h��3|s����-V�,� cC۫M��x��
D1��jhG��(ߢD�ɮ[x��1�֓/B'ŷ��=��&ǥ��M�No����o�a1�Q�o����=7� �g#Ȼ+IE�:���^����や"7��4-	��8��V5"Z���K��h���x�o{���9X��:QJ�����vL���I�/a�l���g���/�����������fu0W���w�5)�%���uDȿ�7���9���>ܪͅ�S��OQ�f]i��!�H�GQA��H��:�\�tPhWrn.�r���}�!������}��̩VE&�����a.�b�L�y��t����D�lWh����{Fmo�5`W�}�ky#�9C���������uN��P��8�Z�Pg�߳?23[rƤ���y1i��h�����z�.���hS�H�뒁]@V���v�f&�� �f@>��#��dH�N|<[��y��lc#Ő�ܙ ����/ �qF4�$.50t���ƌ�B0K%�4��*9��h��Tjfj�I��� H����z�2&��U��C8UMq�-luM������(NR�nϽ��AIof���^�[EdM����{g(0R����ϴEe�����S�6�Ʊf���E;Xȅ������f��-HӰ����K%��;�. =�?���s�����%��nп�1p!�w������3�"J�x;Z�L������끠��p�T;k��z�A����[��g=��.3�Y%�p��c�Ҥ�R:^�T��I�3>�t&�\Y� }��
���v�k�v���^8���� �X�%E���+���!ڎ}#�6�}#N�ɠ���>U0#���C��Y��[��ጞ=����g'�� Al֮׉"Ji�u�34mՂ<��x��n�	%�@䫘:
Z�9��K��I���Ȱ,ku��_���&QaV�!����ns�nӿ��KF��{�z���:��X$PH� h�9~Iv���2�K����82u������Ƽ��XV�ss�~
���iI�3q,
f��*/,oa;���ٴkF��z|��4>�Z��-�W�'���6�}��c�1Sf4��d7V�ȕTay�}^9�Y��"գ�Vt���|'#�K8�wh����ZM��c�$�M����+�;����K8�:j�%��_m��: �OuI��5p�����%���� �2ODz�I�>i���5��i!�Y.吡�������ݱr�=�}�i2�,m*�}i�1�����8�Jupپ�Ї`a�����:��d�-����Qa����0�u��l���!|K8��w�=N�PΘ��<\-�C*)W�M��	�9���]��A���P�Z���r� qBE�p��$��+N,��=�w��<�<���{������g���9���!���A�:�>a�t����JIyv<��g���!՛��p�'ф���&�8���� �������j�ߍ�?�r@�����z�-�g���~�{P7)��ds��j��6_�P���� �P�|�O��-�����,����	��J,N��/>���A��d.$��2[3y?y�G�@5d�VH�W-3�C~�����'��*؍��_���eN��6���ZܐƗ&䂤�=��f��(5|�Qm�9���͟v��cF8�P�)�ī�H5���M�/�6�H��) �Vؘ���F(���,�א��G/�{R����Ԯ���!�~Z��n4��	���Z�c��	����,?[ۋ;�eX�:�o1�э�.)Xn?!�vF��Pg!LFN�[V�}�ᰙ�{�Tߢ����iK@���4g��̂�����ڮ��SD�^O ʫ�8����������7$+����e�W��`��%�P�/0�@dNv��!��$����8����V07�������[�-V_<�����E�ihȋ�n���Bo���p�k$�>8:gu���X�g��J8�Ƚ������W�MeF��a�3c�4��Zs�U�Y�#�Bk��N\�y��o<,"��Η�̥�03@�jI��.|�xg����\�s�7�T�Agh�vjz$\.m^{�O4�Ȋ]��"�ޙqR���}�:J�!g�н��c���o�=d��yv;�fPM��@�mﺐ��o��G���D��Y�J fg3��)�a8�;(?ϭ�z����$oK����O�	V6x�i@����Ap;�,���@��2�����q*x��^�"g�������d�-T�qS֡Ĉ�2MkI�X��NB��*y1+�~���צ ����P��8�;�Le Q��`�T�.���0&�~𹡍��;�$չ��x
#������x2hG���)�"����L����� {��A�0rK]�&�	}�tĞ騅n 1�{g� �*� �R��B�Y���/�|d�L�Wa�*4ka���b�r߈�m��Q���l��&�γ�Yӯ��w�'$�Z��\�8Æ�O�?��<ӕ�^y���)�y]L���A�Z�d�H�&���HW�*w��'o�q'�J;�ª�S�Kϯ�M�z����KfJsv�1�N=9�P��p�Aad�^~85�%��>�[�u1�lЩzk��;��Ů��4j��qپ�aG�&���0^#�'y~'�����-x뾜�p����2;?7����l�
����c!��_ٻņ�?�p�~����I1�]<<F���/����s�]��\���xo����q2����AV�\׈ ��fn]��x�%��9��n���=U,����'n\�	&r��x����Fh@0�R�HT�+����l��¨��䘴x"գ�겖�5����~�ߟ��H�=��h�2hX�Z��V�Ne��:ӭECKj|��2n*�H�Q?P��}�rZ�5K!S������\|�m�}h��ޮ6�� ��-6����ɫ��Esu���C�|����E�_ɯ���Ni�z@b��%vA��P�l�&?2'0:J�8ؽ�o��Yh�q��w"%�S1/�Z�R7L��@�ˇ���*�[t�fSi̡�/�$2�Bq9���g��C��;��ܤ����I"��8P���׺�����@t�M�����H��Q�c�*�ԥLc�s�0�U�}2�W�0?Cv�� ���I� ʓ|~B?�?��o�]�ItL7�z`�1��Y#+�덓���B���x^���W� �Ko� �q6�.�y��j��F���U�p1�4�)��n����xh�%���ѭf�e�nb�*��_� �LX������H7*�=X�5 �O�� �����$�'�����lq�����p��۠�PU�H��ϥ�-�sN���j��6,
��H>���i��;����#^?"a��h�ۛ.�(ٍ!�UHF`r2�۸����Τ��T�N
fY��H��B*�v�1�W+S�&K��'�����;)v�p�Æ��<��.Ao�\��	��:��.�$ۇE5���cm��z=�h�����Ո=%\צdI����N�cB�k�5<��)[%�U_��:���[�����r�P���2��WBW��l%Un�&K��Nl�;�%�x�Y��}���8qfC���]�̉�U�Y��Efb�2x�JV���g�ՁT���rp~e�<-�Mܚ��cτ�"x�&w3�-�#�bC�Q'��V��z���o��hD�G���H�^�(�4	@�0^$���GV�j�ESTֶ�^ �w�(N0U�>x���n�,#�{�i�CSg��l��P%��|ՙ��^ �>�6��ɨf���&���`l�b��\T�[�
�{�Ԃ0&��N�ǻ�<=�;ϳtR��hY��A�?-e'��Mܣ��'{��?�^ډgg��F�g�R�����zܘ�'c���ԁ+'�܎�LJ03��s�9����չ.��	o�M�I+�ǰGT-�;�m�Q�������nH��e�,P�F�.�L򵸻�9�?����6�*2N�8f�)�T�?Q{�ޘ���8[��#8��٥��IS�SYP|u�dk\^����0[w�J*]��ZE��*� �~�C�)�	$��J\k�<,��AJމ����J�� L��i�Č����^�G}���m���+"D�j-�rV�F.]��~R\�S�*�Gc�,���#�*���E^�-H�R�H���sh�<D��^vZ�	5q������$\D��^'��	�����O)�ܟ�ҹ�)�hY�h(�ѱ�\T�1��sqF~*!�H��Cq(��iF��V�A�x����e��PIЧNw0[7��
���(�gyns��m)�eE�|'!t�9�%�m*V�l��7�T�F)���4Z��������>ع�[*ץ[kR
��ٔxЀ;��H�	R�XD�����I�B+�$�g�բ~�ѫ+z!��'L���&�F�⧊�_�l3��M�].��w֣�19">&m��L�#L^�3Х5���ͷ��n���b�?
Ͷ9���@}~�#��5�;�-|�{z3�������\M�t����$���͖�ٹ�h?�=�y���\�*[��Q���>t�
&j�p�|�i����W3!n9�s����HI�t��a.�X�� �4�����\{liN.M7�^T�{�	��F�3[Ш�X5�=�o������q ���EYi���>>����fs��CF��Ԧxq=a!��#+dgO	���H���n1Z��l��x��	�kq'�5/�q��ON1�=�������+���ǎӗ��4U~���m��rw������S��V>��%��D�~y�c���9;�(���F��Q�P�Y2�wl��Żx�{JL�F��Рo2���v%$�4��/��:D]�q&{�A��c�Pջ*�ͤ�����9��%
���>p�$"�,��� K<=y��m�=��x���j�rS�]Y_'�;'j�WP���$���5�GeCF��odlR���ST�OS��Uf��!x�	�=�
ʰ�M�@H��[K�oS����E��߂���YŪ�,�R㖭Z��Ǿ���\�%l��qb��:�}V0ʇcl,��eJ��R�/�Ѵ^�F�<�/#�ϒ1���O���n�쐼.�VCui_ѣ�v|����ӳ�x=���F@�9�j����,�z >���t��4Ǘmt�q{��A�.Ց>-9���cu`S�A9���}��*�n�SDR̬7�L�*�.���?iϚP�L~�]���V
PңN�����4���V�(�"nh�Y�n��mԯ��Uj�����a�$"UѦ�+8�Zu�6�Y�.%�6e!��V�)���Bik�\�/���Hn^ܡ�_���XmC�� HN��H�8Vb/?��(타}E�u�H���Z2��(e ��h��� ��� �^�Ѕ�Xfa"���<�`�ƾ)�9G�Y��3���{������g����.�4rWG�����˕�<����m�(G�&���E�u�_W۩�șv4��3&�T�a�5��K0gC�z�fʹ��ٻh���i�M*f�$����,`*�"�W)���$H�t5��F�5�je\������LZ=W� �� _�߂u���R����w�a0�V�=p6!`d���=��Bk�'�v�1��ֱ��f�K")��#��.̌1��4Z��M��26�r�>�w�������?3��/@Uo�9��𲈹��7
s8Et�Z@�թ�P��z"]��3��&7�s�f9@�������e���8���:�vh7-*�e���n�9�8�n���O��0E�$R��՝|��Y����S"yZ�آ!�D.;Wϸ�5^㵿|�s;%����p��A{1Nc��KJv�w~{��7.��ؙ�0���i�k�a�$Ґ��y�4��߷�鍁�LeV�8f�-=��В+a��E���o^��cWK9�#0?L�⃭�M�#��/�xcz�J�=�+!a��B�y[_e�8M�h�b�h�'����9���-��XN�7)���� T��Z���Ԁ���b	sG:��̈́�(}�4׫��Kh�v]��T��s`�uV��Gz�mk�ŵ���fY�%so�\Wƴ6{��A|ɓu�:����<;�ꁖ�jzgMр���H/�� �#S�`�eDb����p��.`W��)e�y�>�:-/�$~ҠmcnH������'�&�PR���
�	�É�-7�����*���ӊ�mHc.���hm������Jz��bȝΏP�I,&c+DW�w!;�'[)B��AgPy='P�Q�ʡ��|�	sO0��~>�m'7���6�;��>T�!(��o1x^���2$�����F`G�Xf@nr]<���u6�;�9�|`��#j�2�yk�sR,��:8T�s{D�2mD�ڪnåI"����ʌ��#/F"/�G+f�)0�j*�vB�g�� 3H[̖�H�����
��oxj*���#�Ts�eʪ&�x��ge߬$
>��.���%��]�]@�gd��:d
+���s��(g�������;K���9�J}�ܣ���Dz�ŉ��xs��t��sPf�Wۆ1���j��`� .���n]3����S|�0�kvǙ<�;��U|�G.ʅ��i��Z+�|z2��;j#+�~;�����1Ǣv#�Yx����4Y�,>�Re5�Y�VF�U��QG����zå�	|�� �ލ�Wo���
�6{Q�俵;D�'�;��
�P�,0x8�&]�|��a9����d�G<+,/�J�]W���/�e���*-�����T ��8�	�=_���J�wG*p̉1��R[?IIk������m8����K�����=랒�+���
<Pl �䍠���w b�]н7���'��$'Tī�D����,L� �I¾������@s.t�����gS�8�v�{�C�L!.���f�Y�w9'�2�����
�7F����{"�a��m"y�����sU������G���9c�i�E��|D_�`�]�F��.��3�_#�qsh7}��5�Ud����0�RAi�hg�h�t?�;4̝���Z�y������NA�1n��d!ъl\�3�A��Ġk�«�W�X?��8���B	d`Jc�w�i�k��� 1�}LO��ŜJ��c�7���4�m�բ`��Yf�|���YE�4�EIޅ��.�m���5Xև�ǌ��ޣ��\y���9g���˪I톨�8��2X��^p��i��3��J�ꎿ�Jkֿ������.��#�
���Y#�~�e��!݊͡����T�)������\B���Շ��;��=e��6��i-�%an��eOLw�q[���su�d��â�Fj����y��$U����`�mY-OcXQ�^�"�"�if	o�cwL�C֊X�c֋x�\�M�+ <W�d�n`��Pכ�/��+C�<������jx�R2����	�d_F-� wQ��|,���)E�B,��\6�ՀpH ���TxF���dd�;֐��<���qAE����p�$۸r�9�.���Y<��� X�4Dñ�9.f4�l������?�huwÕ`�[�=l�HwY�5��t�`�0�R�y�����t%7��P͜��t��+�	Q�N`tZ��|��zEX�*>/�_��l����!t_���t:��_����U�-޳�\��ݒo�����
JG�]5$���êؤe�:E��J��àj�͵�CX�'�m��%S+�e���f��i��T��>u�X�*��J��u�̉�k����,����E- h<���"�0s#����b�-R�ٹ3�E�m�����qL ��9q��CiOVi A��O-&�b'���s8J����vڝ���D+���+�0�}Ja,�ts���Cԛ	�M<���ЬzXzc�^i��:���n��JK%���F�.w���J�,�!qiVY���*
��� ��F��y�m�L�x��L�Fv}cs��/(WR��ѻɨ��񷁆�x��o���'&���Z;�1�]���*��=K�@�i�W���}`a�K���B���	驪�D"�A�VB�((����O��˧h�ȉ��Q0���}�n�^��zପ�O�yu=i2�y�0*Vq6��aqW�dU<�eJ\nq��6J!3EE���'�Zl���o`:ե�9��g=OG��4�봵�p~�����YKA����M�V�pe���{5��6��
f���
/?|�IZW���c�X���'�jlA���JX�t��������&v���̠��j'�xi�~cw�������!��+{�6s�nc�?7��/]��'(������:��$1y����V�@��:ʿc'�����'ӹ����q�{��F��y�����"�GDP]�L�3¶wʭ�����\F���6�,�Qt.�����S���M��%�DM��S�ڇ뤧�2�)��K@�E?^ŋ�&�w����P-Hu��d�з��KFů~�V	1x�N%���VȊ��e��:�6u2��⌆�D'^t0l,3v�_��Z
0�8�>vn�{3U��{Q�L�o'C��+� ~�cwQa%�Op>S�c����V�O�@$_��Ӿ������'ː��/}���΄�#�L�	1��[
��+#8}s3��zJ�^�~%I[>����|���כ�^��侹�y�(�6�����TOc�&p��G�V�� ʆ�)��[�q����:�!��\£Ƽ��V�JQ��V�c�Q���$ZAf`��3�fT�lR�;-�}�a�T;p���غ����	�0�>�7/P�\{H��+���'���yp�W�P��	�p6�t9ٵ��m�02���k�9]RJ�z�� }���-��<v�A�%mx�Hm@�{�t���-ˑ������ ��j&{��Z@�8YQ0W_\�� ]�<�	�4�)��Ƒ���V����S�%iE�հL����j��$��~�R�k4/Tr��dG=�ʥx�,m�Fә*��6��Ц7tL}&�t��c�8�獂x��t����(ɁAoX7x���c�-�7p�,���,	!,���Ox�lu5�B~U,]��H]x���׍e2��v�mZPH�(e2�̴�K�����$D���IO��b������$0�(�%����;�/[yȴn<��2��Է���C�HK�T��N�{B"YU���R/�F��칮�R�F���)����
_�_9z�x|�q���q�i�������B�b�N���RϷ�|���[�؟�C�Mby��{ߤ"ľ��>�Ȝ���P�>��q��ɏ�F�[u���q��-�W%!�b ̕@�snj���*69~����e�18~꽍��c[��ل�k-��4�͒oJ�������օ�Y����x4��p&�*�VKA�[�������;D� Ձ�Ћ��2/���<q�HL%��l�	���y��x>��0uZ��	����6�pf�^�g�O������Hg�Xn�k���%yV,�I��qH��d���YyB��&0A'�d��Ӝ���T��eץ�2hxs`����J�K����'4$ȩ��� �xo���+#� ��Q��$Җ�be,,ӃO��{��V'�C����" �i'��{�e m��ډ�]�g-լ  ׄ_*;bC+��/����憛�|��J*۳|��`�n("�ʟ�a�ζE��l�j��;�7A TK��Q)dN�{N�e�И��)�8+O4��)��É%�7ׁ��08��m��&ceXe(]q8f�3�@6 �_0 ��-,��w(�S?+{=OU7�`Jz���fU�2GK�\c]��\F/+�����d4wCv��Z�-:�s���Q��G-�l2	�A�@(8��g���B����.�fYʅ�����[&_�i8�I<���}��?R���ű9�����FN�A�X̙J��ﵝI\�3$�r/ڙI���f]��e�b)W٫ǿ��'ح� ց���p�Y�q�n�#��T��i����V��#K����w���$B$޵v�V�wɔ�.a��@Y�me�����f=����v 4����s���21�#�Z��(#��@�.8h��u�m4S�� �V/$ 4ԁ�ُbm���>U�G�z9@��1
tث�n�(S�'^�t�.lfw8���?��G0g�?��ED訄�_�-�͇��H�-W(��A&d�dx�[�ױ�9���]C����OI����R��[����nP�vA�.<�'Ghe��xX�{�0Bv >�˭B︓�<]9�5~N�(�u>~��sp���E:t^��	oݧ�8���Ϗ��X~�Z�nD)���A~�'c�UW�|iN��*ãG[[#K#�����Ox�8K%��h�Q�J�_}�G�֧�j�u^7���X�QS}��.������y1��i�\�a�a��oR���.z������o�$�t�;�+�~�' 
{�G��'�@E�A����\E/���d��s=���Вç�}�nV3PZ 4����^���ce=�E��u�Z�.x_��Qn*�D3EL3}� @�圮S&�F�0��KI-����}9��Zg��ax�h�t����8��Z�����m~r�"��~̩̍������ZKh�P�=�+��&��g#��:}�E7�U��R��\���S�>� z�MTKQ;��ǆ0�u4�����1w���Z�|��"����0�T��4:�j�o/��~����?0�hOy�=e���A�5'���XC&��5�M����6%�uv��\CUE��!�f���� Φ�렮7��"�<�*�Vr�"��2L�f�N���Q�o�1�EDe$sL���(�u֩�{����<�3���[�Ul����M-(KZ�K�'����f�Q�[7z�\B��.Pħ�u�@w������J2�C�hDi�9�7�� 4�UA�	�;܆�j0���yr���w�����˪*���ٰ4���h�;����aʮ����^������w�v^L�6��D�,��:��`m����'�����"e&tӆ���
2(��J�)g��g������n�,R`)<�[?��o�bD�2�Ͷ��$>0�����֭�M������n����\���F�9�^�Ӓg�@.kZ�
Q��Qe#-ǂ�������Nԣ��fV}1pZ,��d�Ty����8f$�
�"y�,�+#$l>_R\�#	g{��� �;�*�G���[q�?����V+�bkzLw��e�7��V�3P�AжTA�P>x^ti��ڷ a�
��-��K;��]�9�����<��{n��F�*0A_k�C�l���������8A�:W ]���6��,��o�@X1�hY�n3�r�T��Nc�1�4�� ĸq�v��)K�Ty5�]N;�n.M�2�b�����+Ծn����}�,k�D�<�*��aC�}��:���eb	��d��S�H�3��YGU<F9Ԃ�s������^�H{RR�,ӷzR?(�`�U��
�@ނ��E�[\e�9��߉2"X)�o����!5��Z�g#�;�s�>�i�H�Mh�fy�?2_;m�)	H����1�� Q�;m��N'�`�i�Z��bx���\
�JI��o�F!֤��`tE������#?���ؖsJ�S�YH�ݺE\����l� w3���s쮲���G;�l*GC]�>����w����8|��+�6[^�{2n����Ro�˦���X�"����c?3�c.Y5�x��6	���=T{-j;\ ��s�b�*�W��9�K�Y� )4�����u��[._.�l4�X�x�H�n\����Ql����`K��*�Xx�[ ω�5�aa����Լ�����^8&�뚧z#�|#�'m�S�Y&:�#yrI�,k2T�ڃx�F�J?�� �I{��1�B�J�0O�Ԫ���i��_��O�	Ł��x���Z����=�}�E1sV�������N-��
$�]�흙�}����6�@�E5�;Y+�07�v����I�E8��v���F�4��,ʤshY�H����m[���-��\[2ɍȬ�7�.Fy &^��g_�<��Q����b-C
:��(��VE��������9�@.x�=�e҃EY\�=���0S�IA��BI�
V;��	*)r�P���
�!��%�hYT���KO]�	�3U��RS~�&_���f�xP�J�˗��{��r	���Ǽ�l��t݆}5BjϿbf6�ľA����é�lA�Dm�Z��lA��\�-�E��z?�Z��n�e�N�a�0��o�A�0DXr�������#�`J'Q�)���N�I~+�C�����/KC��8�BեÕ�;] �v�F(/�?=��Y�?�[L�hLq�Z�ۺ�ɨR=��� �o9^�\s����0%���V�{&���hn-}��z�3e�j�����3Ѣ�̈́�_P���m�kE<�u�q�����dP��e��@�@���7\9T�?j/3Zo�MT[�ԚZcf#�Jcx	�t�JN�����y��BiPbh؆	U�\gk��2-��3m�KtQ�|p�,��v���̻(��ۗ��2���_��`6#�,��F�Mtd���ۊ��w/@���$��}.N�T���H�e�j��S�o�|��|��ᅭ���d�b��I��l��Ń���5��������z��Pw�4����iG�~���^�p͑��۬�
�n�E8^"*�n:���)���VS"����<���6X���z�ϔ]�l�a2u|4Б.cdUƷ�����{����s#����W5��T%RF�$ba�a8��� R�1�?��5$� �Bk��<�,+16�+����*����C���(�܀��{U��K;�s-�T�)� '�\ ���;UP��3������Ŏe�r����J����̣�Tq���HIG)��~�����rx�mU@�冶Bi��{��7�����Jʐ��@�#��G�L�4�[E�'�B�Pw{�eR�Иk8D'��eU��K�-��2?uD9 �t�����S��Z���ȥ��;�i���ph;[_���,-������n��,��8�;�/�g)
��Η6���q���5�⻉�x���z�R9�|Le7OO�Cɐ��W���$�:�u&�^n릅����"޳�r��?� ��;�Y�ui�)�%��7W2a g��w \fr-UDI��0�䮿o���ޣ2������*��%�k	$Ft��P��2Z��9�R)���nE���v��p�[����ÑJt�P�����C7%F'�n�]5l@���y2czj�4��"V$���ixlدm��Mp	y�!0�Y�g �ѹV����v�E�'>g�����U�I��{�÷�� �~4( �>�v������H;��0�M8�c�a�`T,X(.J��dk;T�.o��I�d�	r������_	�t[M�^�l�Q2��C�?�����]��p(�>d"��w���|Q�ZQc�;�\}�s�(B�/���Q��*�g��_C�ey�bs��@w��-�᣺�f��f�1.o8?�hH���ָ��[g`��]��HE>�MAa�h�`uu�`}� QqO�G8�H�}�lSv�%,�u�qP<��cB��(���OQ�)��r���ꩨ�$G�%h
2�6{<�jc>4?��R)^r��4��$j�`�~#L?j���-u'�ӣQ,�clel&P_]�z�E�Ӫ�Y��n�:�e}8�OeaU@>^�g�*J�#�e��%� 7�FHraQ*\>bN��M��3~�:��TTv�%F�5J�2~_0�'8e�||h�/�u��?��V/ ���_�����=���]*�UZv���ϋ��(Ep���Y�mP��L���5�q�*յ)T֋�%�On�4cAN&�c?��J1K�F�ƅ2����sp��W�٤�i�y�h\��E7�����p�Q�.�by6�qD����GB�#���T��0sW��5���\�.j����QLn\\�Ge�:�9�k��՟���xc���x��Q�!�K�,-!h��@��}�p;�/J�П��Z��2a�l��#~�/~��g&q<�(��z�5-��Q$Ǽ��������:ݭ���_h���-{���dj����l�w`7����D�a�\�j�����o_�;��m����Faޟ�g,�0$p�c ?���A��	��{j�K��j���5�"�4n�:!�_{Ż�Z�FP���6��D�2@�)Vz�X���'�r��HI-�:�V����� Sm��ۺ�
DڥD���1G<�e�b[q�c\�>����!E����_�q�鱌��LW;R&l6ӥwHM%Y�W%}j>xy�Q�yR� ������������TwAQ�������%T��:@Xqk�6a\��ʞ�\�D]�c��\x.n:��v��Bq[�5�(_���[<q�A�Y��R]�0������Ha��U���{�"���?|P/n[����I��%\zV�}��g
ܰ��*�����PH9Q5�斎b���}���G))I���e��h/�#D����P����Q�*X���>�A�u�Kc1�g�BG0�Zr��gz��9�K�D��$eޥ�~�W�-\.��Uy�f[UW�[X�U~ӊ:��0�����U�[��E�l`��H[k!���i0�7C`�,��c�����LG��9�^a��� ��f֝���#����0��/Ye6�{�XuY��2�^����9�N�������yJMG���b���ȈN���p*g��-t�׈$g���@��aot����6�����xe�I�4��6*�I2M�ȡ�
���v�3*���gy4�Ȏ�sNҾ줥�)n/XkC�;�Z��rB}%������ҞTc� �-���G�M��ʦ�C�:>��P�fށ��nw?�uFDl�C�WL��oMר&1�]�\��d��7�)�5Ԉ�>"r�|?QE�5ܥ݇���ǻ�?��g�����P��<���Q�����IQ�2��Az��؇>J��H��^G��z$�U�C�}bSN�^��sړ�����5=��Jϣhj�S�W�r'���6�Z��Rƣc)S㚅��q��2��P<�̴�9���e�Ԓ��e8����sV�0��,=wᴶ�`�hW��<�tf�]7�����F��"*�*�!������O�P�<��0>���A���y��?��ۤ�4���B{�RN��8MQ2��y9%C9�:�$�sb�����ڶ&g^ ��-Ы�wS��c"nFl�n��w7ǎ�j�ٓ�2=A|�T�9lQ�72�R:d����̈�3��r[_&��'����LJ{��pP��c�s旰^�r�EO��p�Ｕ�5���T�ԄQǿ��ZGN/�7̠V?�5��P��غm�0�����8�S� �����3�q�o��F���jl�z��vNaT�h��
����*���,EL~��P�6��Ӊ��� 1X�(UJt�)�.5���i�f�xG�ylX�8''�g���2q��sǽ��S$��IUZr�n�2g���mE Q\�ؿ�[j���Z�S�H�����c���_��YA�`��$䡂<Sb�3�^<�z(��:����+u\kgvZ��k�9���vC(j%����P��)�,��vFU�m����eeH%���l��=�Dh�ޱ&�=�l���,?޸�Q �4�E�����W]��,�;=�VD�e�tCݲ�k������ M�DQ�ʐ��s1E8i���tR�;ssP�&�����M�G���Y-ˎk���ǽ 4��o��:v0�l$���ٟ��^�[~+÷6�ڽ��n�لΟ��^i�%��3��5��p"�gO����r�C,_��:pG{2�@Ok}DɇV,BU�h��y\0�6�Vl����&2ȹAHo�v�H�KX�ҴzŖ�V��t�i��BycY��޲>�(�H���db�8lf_�/$��y����]M �c�f載\	]z�R@�A���NK=(W��ق�w����:�>��ŵs�3�\ͳXc�G�G��S3N~O��ff(w;����aV�)v��_3���b۾�]É!��i��+a�t�*vYš�i!�7�����d����ĿO~��۶�'f�i��������-�9�:�ݐa�ѻ�V\a�kg����,�I���E�'�����k���Pʙ\gb��lj���j�d��m��otjT����M�/�:P�X�b��&2���Ս�,�Nu��"7މ�.giS�Ak�0�o��EP$Ǫ��x,�$�L�N��ۥ�CQ�Sx�G*���ЗG?u�[�PxJvx������c�b��6	��ް�����$�Th<`�.p��ʉ"n'�m���y�3(�YkrnX�:���W,��5���_d��>����ҟ@�b~sE����=����q4����G%v��}%�+L�!"h$g�*9����:9�
y����/+��X��UѾ�9�NL��<v�����-\��S����A"(�L��U��z�bM�����<熦��he��!��P���J�G�P�����H�o4K&�X"g��q��]S&�>��2�W�F;�)�Z1��	玜8d�F�4�� E�H��k�=��W*n���	@wa�K����� ���ko߈4� ka���[���<���a˛j��ǭ+�^������e�S����@#��9S�2R����h��Q���隣��.dzL�\���Tm��rZ"�+��i�����W6���f��(g��&Q4eftuo��	��RkUՃ�뽢	雂[���
�H��
���щ��J.l��=����+xu���t��b^����+�a�D�5�!�C�dg�}�A�������Ш�M���c�/�4���?܂To�����MZ�ZN��
��P���ֹ6���g�S���g����n��F#���T5�@T3�j�|@����v>��NU�&�^��s�D�k��$HpiHPM���~ԍ��S���z�J̒:8�Eצx�2,:���/��v�a�V�M�������x�7ȏ��:䊄A�W�H�]��.@�����y�*)[�Me�]�0���������gZrI ��h /7����Q{�%����&�^+L	��W���h6&�}�ಭHh�N�G	Ϸ��\��%�ʥ{
�(�*�ǺB�
%�á���ה~��*�w��3;p�5��;]�aE5e	wt�3i�F���;����'�MN睏�/�h$v�O^�'��&�o}�%]]�����2��,bEg�^q��
�����Еƪ�g�#"�9�ڮ��J�v��(��ڬ�����АT���f�>����<}R?E(�.+��`���s�¼�D�l�����|�ڊ?��dn@�e�\��/��L��6Mv�l��Ѵ��\D�}>�׿���%�T'.b����yφ�y�q����PL���|v�n~�#a�C�ЌUr��,^�wh��4��Y���>�ǥq^֊�U���!��for��ϕe}�[ �zq2I� l��:.��w�	w<pĈF���d֬��6�g�S[�Bأ�\"�r��`;�p���.���+�M�!����>Q;ߞϕ;f�䭌0�<�SR����j��c%R�^Ϝ�cp�Y��}~y�-þ����	{lXlnB��o��X�����n灟іT��1�H���Ȳ�-췝� /����:�i,�(���%��Vds������mw$��%
b��� �H9��i�J%!1���ݸ�)���XVt���eEu����9��� ��жY�"�^��8�"��*�?�r]��4P�s%#.wSe/�ԯְ��ݿ�؆ȏC"V�69�}Я��ˏ~En��X�Q>4��'�� �I駅_�����ʶi�-ɠf��	�+(�
�x��^W�~hFqߖ%iަ�n6|b�}�2/ Up>�60�H��h3R�^���[�i�_���g ��3X0Chw ��Z����"c�v	��272Vq>�Qm�m�x�v��NX���� ߫O� �u�	�L����+,M�����Ol�ԛ:ƌ_Ew�����2��5��V-Fr�
�OE�⾌\\=S\��Z�Y:���;���mp���t����"}��S�����_���r#Iol۞��ߨÂNm4���y\�a2vǮ���-��X�,H"��"8�2G��ڤ�+vhtT����!g�Jm����C�Ǔ��1���|B.�8}�4���G�z�IA���^E�̱���D���V̳ rWz
����4�8���{Ě����[9����4��A����Gl&�v���n��=���*C��0�����3��V���h�>X�)Tݧ����jDU�|��[�F��?���E�2Zm�2u��3M ��k(���|<7�8'����xi�*�&1O�vμ!uw� ��f���g{�+D{"��2/T�-��R'��Qqf�!	֋9�K)����s]�~rԁ�;|@> ʤ�	�c�-9l�x{HO^��WG#��$�1�bZ���;���[�H}c �j]_`�J搔�v���m�(*N�N�����]EK[�>���Sj�^+��sDG[þx���ݎlPO�`oz�h��]^�^5����t���WfjxT�t�ʻi���3����W�M��Ie���[�*E���59����n%���}OI���#�)�ַI|V�B���qV��g�<͆EK��]��q�b��hpG�I�}x�ݚ��Pr ӽK,�r�O�:�^�!�0E|Tz�({C��;�m�n ���@2��dB37��rj��K�����S��V�T/ڭ|J��\���W�o ��>��W1���D�����R�=s�������;2$��F&��ӂ"!���Ţ4>zC8��/������.�W
4�i!	V%�A�O�1�P`(��)�n�{���Bd�t6��>6t\EH��h�Fml��h���YJ�qj��(�nxOGp���r2@W�@�(W�Qz�:z�%���{r$�y��\(x��q*��%�} _ o���Ɖ�/K�G��v/3�5�FW�P�k����������e���=�^�_��5_d�UO����`J�jJIS2���ʹ�z�x�C�Fl�M(v���G��O�< �u�aFp�����s�7 ީ.�u���*o���%D$Su�e�5��ۍ�TT��ZumP��;�-��y�y��vy���_��g���&+Ȳ���E��tz�|.38�������a��P���$(�iٮ�'H�}�,P�:<�s���kQD`e^���/jK�mA�jѴ�ʍHI�'���j���ATޙ�����8��}���+��҃]���-wL:�%�~�Ks��EW]Zz���?���^:���ܒ�OA�H싣g��3������.hȻ4?�(Z�*�cS�w�.���rg���Rh�A�d��&����Ox�����LKW0��ː�0������4��YC3�&g�`EO����T�����J��>�;ů���=��A�_�(K�-��0�'��$h�p0�e���ӿ�#4�q�3n�~��|��Ӌ��dh�t>�c�ޭ���_Xr�~X���	�Ġ�/v��Q�F��K��!\y(�A�DV���;�Ѫ�+��ⲯ�;�в����,�L���"��YΔ�3' �WT��m�����k;��I2_�Aa�U58��æ��~�tʟ�-�?4:.�؋BPu	s��rm�Ծq�M�N�b�U��%D�Ӟj g��j	�ۂ��G����=����D����@+x�Zvt`����%1�1��$��8ʼ��r�)b������$�\m/�P+ l)'M��UI�i�����b�Q���!����_+�f������z�qE��z֮�JV���yƎ�k\?]C�S*�ӎ][m���@?=����G{���OV;F��M���W/e�&����S8Z�ö��Wij�7��:Y�f��ٯ��R�

,�<u��+�̷~���̚'��*���w�h�i�4��v7*by� ��(D�tz�vNC#��k9�Gk���,H1�A��X������	�V���E�u�2S���N�O�8��|O�.T���.]�1�m��/`��6_���w.�޴���;J���U*�:�ۗm���<���N�/���N--UXIbÎъ \vd=h�+�����4�Ê��#�@S�������R�ʑP�^1�s��&	�w�&d��S�t��bR���M�o=�'��'�$m=�"�.�/4t��#&�`F� ���0/^�&�[.m\�P�BC���F����
̐�PGH�F�X�����G�f�`�ƽ��[,$c�v���Љͺ�Q�o2����Š�v���P�����=s^6mǫ�|g�w*�L1���)�K9�Qx'BU*��ઍ�|��\[ߦŃ��ɛq!NV�kn9w��̕01~�o{'�1��;;r*��<Ԣ���f}�\`J�����&�"�o���_�a���M���d<�H�I[�?�~Ǯ��PS;�.!:�D���&}�J�sA���<��W&�����o
�~��|�=׶"9vE���'C�>��"��p/2��/��I��1�)����`V��m�v��A����o��.MO��Q�9�+����T��׸fjO���5�-jc=:�j���D��se�q%�v�Υ:b"�ܫ���$�j�֝�ZF�qHR���x�Jwʜ�I������@;�<2�w�3jR�Nx�(9k ��~s�������B+�f*w�( �۝��:m��X�a���x&��6�*3;x��M�0�A���?4e�AȰՌ����+�¿�����_�ʒ�/���)6�xy.#�R.����I���d_S�Vi�9�� ��,5�����7^׋�}��I���U	�-��%4�\*	��]���q�[��g�'/�-�ndY�������#G�+ٻ�j��-���A�\��s�.�H�4��,�1.�1"�}&GҒ�/}l���\E��(��Ź���������h~�&�5T�X���s˘(P1���"�g�0����L5���[v�� H@��J+��cH�Gv��:z�7�z���/��P-����r��*�}b�\�����.d0�n�ݓ���6!�z�mJ'�)�1T��I��d�g7��&�	���e� �|T=��%��?���N�&yD��)X�CJ<�F���`��׬�	�s{I d�f���y�c�tYL7.�E#s��^��j
`0�1��+�`����t����6J8^sĳ�6q�{�%\A��(p��,�x;y�d2��vd�H}��n����e�3c��i�L;��0�_�)��������G~�;�,��r���u��$�J�����ɌS��>"&�"��ك��=�����QC���E��x֣1���nq�D4q�ӹ���!��(��&X6���Kȯ�}�i�Az#�jإ��sF��s�ӵ��n]þk��F��q0]��@$��p��]�}�D0=:�����hX��䁻�B���x%غ��9W�+�z��/-����]4J�e���>�n�V.����H���R �_�۰|�~�s���%�:g�Ƀw�O�T�� �	�KR�I���{5ٛ1f�݄��OJ��Y2�E�koȅӾzc�j	Vt[�;��Ñ�Pz����]��β1��)��)�u���t����2��Ǔo���0�6n�HQf6�<�����R��R�y�����]�T�Wd��ź�}v�(N/8���x,DB��`b��̫S�i�\�ަ9��K�X��k�i��XVg�T�3i7&k"�wv�D�F%���� �{��Y[��.� ˟x���J�-b4��M�ڔ����Vj��D���G��玛uC�`<��a��P|[��A�6G�ˡWu�Q'����r��[���%Cʰ[rwv�l��='��@RH�;=����6z�J�4��F0���KM-�~Y���p^b���ց`���C��ƻ�㗘�r�gT�� ��gt�J���;�K
8,(Tf�Z���&X�n*��')���̉� ���~,͞6�3���-��X� L�ݼ����Q�W}b�,�b�>�lK��p���F����GKڨ��s�y)Y�7( �8�d�k�r�p���(����! �_�ק&;/���:Y�;�}ʽ��"����XZ����O����S1�S�_��&~����6�7����K�)"��[P�f�0��e�+����F릶{��Ot���u��oH��ϟ͚�L� �u����G쾙l��(T�Q����<3����TGwna-��v� �s�cz�F�v��ܱt�{+���n�5�i]�_*x��GC#��^q��b>
�$�V!��*�$^:iZ^��)�{��VI���o��,�my"��>�d��A��&�����=��UG|G��,�i%*O����э���yi�����p�Ywi04�9i;ַ�k!�ǳG�����O1uYz�sI�Db)��|�$�+�c�|֭�x!h�ɨQ����P�)�Q� ��v�Q��<���/����m���]����5����\Q�J�}�ZB	��_�2;�߈��6���]л���O��]%�O�c�����g��X�k��E�P�­����8�	%�]�{�߈�9��i]�Lc��i���&Xq]���9WY������xۍK	��|�Q��4�tzL-�q�Yx2	�[�W���%�#��+�~rA��~�j<{� �z�5���I2��X.����4� ar1���ےR�ݠ��kbH8:�E�F��Vd&u�TVRou��h�����lt���_f F�M��y��b��a*!�*��'2�c�eRߖ�\c���r�y��>Y噳Zd~v��2��9!��	C ��c�j AKz���K��"��t8��B��1�`�OX�%�V��Q]��{���&���LBD��p��	����JD�Z�S��ً�EP���S���Tv̤�DX�T�*�B2B���B�P����!��UKܲ��z�v�蓪.��%����Dm*/�8�y��D�h���a�t� �����XT�͋���|C��@N|*���'{��p�Y�v{I�_���_	�A$O�����?���zڳ7|�e�C�*��a���lQ.\��rTq��fVh�_)��V�(���|����<����8�M��y<��9�.Ӡ�V:��s��%���޻�b�Ƅ� �S��.��S�yɦZ�SK��'�W:cOu�g/����[p����U^�u�@o.j�x�4�W��%-�����n�Fuպ:��v�@�ޔ� �V,3�����)!L>�Ef̄�>2�����D�� ���%}�g�B7�+ǣ���R-��.~)�)g G�V���r�r�z��S�>ٴ���Oᔣv��xe��΅�#"�y�TIbka�+ge7��!�H�4G��+��L��1p�m�n��VJ�\������7����X����\G��sNy��+`�Ը��4��҃���?. }�#��Y\������(6�+o������_*y���l�#ʷ�\��ӝܻ4���<{wR�4����5���3jD$IXI���90�����8L�ň߈�A*q�V<���z&�&��XQ�lzH/�9�_]`,��.@bE�D"��N��M_$��@{�hِ(�4榚O�R�\��z�IOF@ɮ =��iّ
�.�a.�j�G��gv�9<Ca��I��`` ؃�yI� �N����*��yM�i��%5D�7�8�do��=�y��W�=XŰ0�W=��.�g<1s�ı�"�� �D���а���S�ATlsܧ�]mww*p�$5F�}�o���kRK�4��M�0)��6��_�17^�D���RP��1S�%au�IDk�P׭�Q8���I��+�?I��W��<פ�����w�'�h�g��L(YUh=�*���AT��pgt�uL(��!E�����$γ^�k�9G�h; )>k%b�ei���9b�#�~��]��!T�tr���׀�SɭQ?2X�32Qx��.T������y�h���sV���S"¢�B����e�����B~$'⠕�y��yt8W�c��q�����ų��2�������A�%L�y�s�\�����	�GN���&4X�_(��%*�?�x���A��o-Ez�z)K�J�����D_P���h�Z��1lY��&.�SN��W�f���+�"�T�J��s֚��k�D��o�%����e����3�7R/ob�<"�⎮��ig�.��9�3#rEvv�
��]C������=j�=��|X%�,-.�̒�����҂'�8����/Ue�!>,�]�2���j����x/c�������m�"�V�v�%����K���
�	�����?����j&:����5�a|�c���ɗ1B�S̲"��m[8�I��^~�A00������XD9�n�c��7��m��+����Y�]hېh�.3�XX�~e�\\����k�+�˼tb�1m�P\
Ѥ�p����f�˺�z(Z����g��DT�7�!q��*=����)b�qX�˜������s����WO7N�����}���$��ա��"1[&6<���"�|n���5�g�
S?�����{ۥs��"Ѯܛ�����<r�����ճkDy��m_��9;�l�᠝K�����n�l[Q*ҍ�g�]�q4�w�:���x~&wCS��Y�0��g�2i^�����m���?"]���ޯ���b�w�H�20��]�>�*�]�����Y�L7�Fn���5�8���
=u-�Y�o#"ҏ�8��R��1C�
����V��>}�CƆ�k����Մ ��Z�e~��ֺl��Bދ� 3��L��C/�
ǎ@���~}�������u�^����+�>�2��j�bųT� �����S��ƍ�w���"��'�*�Z�<zZ�ш_KJ��G7ʫ���Ec���F*�v�v��@%� \�~�\6��R�{�7�Y���^x��0�i���I��BզKI��Lm�f��:��Jo�Ϯ �
�&�r����Z��WT	�_��i��BG�~��63Q���N�y�	�d]D��Hڪ��I��Ha [�� 0�%o�ӽ�$]�J�6}�A*���v�뷎fś��o�T�G}n/��	:���S�Vz�����p����>��
�SZ����Gwy�;a62*�Yv��$�|�`�H�����=��jK�|<^�Ͼ��fQJ9�#���".��@_��(^�7�J��GR`�1?Mx�Q�G�C��ל:����Ӭ���Q?j�H�i��-�P1?�X��eC.mp?z�U5��3U]�OX��R� ��ȭ�@Q;H��+�D�=��r1��nG4��*�kB�����5��v�iȷ��²��x6�i ���;���k�EZ�=�M4�з��}5A��e6>
7*q�fI���d��3�7�k��OV�?"o1V8��}\����{2�y��-��^�3��."%�s/D��vwrӃ@L��"�?��o_��L��:õ%�I���\�]ѐR�ғ�\�����ʖ�p�U���'B��鑢3<��βV՝��Uh\����=勏Ѩ���gNYa�i�O�)��yVm2����%]�Q{b�>���w{�X5�T��]Ӧt����\�2!��!�_�����F���s:GT���ϛ/T�>`�\t`ed���ә�<ʉ6�0r-҅A�{	_:��CJ� V�m �B̘ιn���Rf��k3[:��73;-4!�U����(s�zϒK^׮���/��WXL�0���\ZH2"����,qD��%C��;,�|ˣ�ý�B0ꎪTA���r�n�s�H>��&���pj�L��\(Ӥ��]���[E�VX�h���B�����Eܪ��
翹ب�=r�&$~��9�=
��۸5�d��ݗ��|b��nK�-�<� �ґ ����fe~^���\ӧ;��uq�m���Qu�+��	S3���G$�_��Yz�T�cԿ�RS��7���yD<&@�o�\A1g��p;����d09W-��s��ӓ����4k�۰#]�3��M�ۑ;���.��2�C{�E����2U@V����z`�=��A�Xii�ζ�'	�&v�^�]g`%����Uw�i�Gr$n|Ls�gJ�J7n��T��u��qU%2w����8�m|��
K2SP���\$l!Maby3F�8eXJ�����[H-����PBAs��K��i�u��WJ'�7��W�]�����X�m����S��_v��#��%@O��b3�����Z6��-l�±���z�>���R�i>�ϖѠ=)�4> �kxp�����}�z�O���~���D�ܣ,�q�=�A�{P��e�r���[�ٶ7��m���b��l�����.^�k�6�e�	��d�\�qoyE��b���u���B��rK��1D��m�9Aݍ�m�t���0����1&C�SM4���f�t<�eS�C,���1�"�k���� O�?���^��=��?�t*�Y��"8�WW����1U�x�� �^���rNK�~K*�I&?c���au	_5�.R���sX��s��F�n�N��8��#��J��_hb�4�͝v���ݶ),1n��)I���{��]���T�{���
�ߔ��U��3�Gv4�7`]�=��8m|�[	�����M�\6�l�b��@�	3*�giZ�/���qB�!�ħ������g+�3u��y���qV��aU0�Z0C�5���3���@�rb�J��?�!�Q����:W����g�+���b�a�7F݇�Pc�I���S��o��	�3��fB�ӣ��K-�נs���>�ߵ>#�̭M�U�zp����{��4J�ه5-�k�xxbx�LL��,Oc�$��5ɮ+�6Eg��D!��Z���۹\�HO��m��_�l��¨!��8���Y?��aG﯆Cnj���f�@C�K6:$� [�c��YHm�|�0jTP��-�/�0!SQ
t���)��QH�},x,��P�"��-*{�??m�� `2!s[��zl�"����������`�?��hM[q������@��炌Q�iܥz��]^�����%R�0��p�FGE!*�E���9����&�c]�SDϥ�Y$}�( �p�oIh�&��b�����c�a7��I8<lx�[Qs�.�EӋ�3��zʽo66�/-����o`T2���^�s�U�h�g(���N�Ag4��'l$���@��.n|���.�Rc_��J4���eU�Ϥ���j�H4̐a"�}4<k����
��D���1��� _(h91ԅ	w-}b���s��]0epݼC8Dg,��bsJ��E�ӻ�*T,���1�_K׳�����G�4���S�`��Ꮎ�g�R�
Xq��N�:!%`����~��9�PDC+�++v�p�_f�
��i�����N0\�2�;�!�R��z��Z>�ϮÁ��y�@��aă �ǿ�tEk�ũ��4��D7o��cE�y�1��|�i2T*��j{�C�$�H��qӬ����E$�+;��|{xӿB��@�ȯ�(�.]���)�g\��ǌ��k�*.�k銌�O4���r����e���3w����mJy�,������l%W���R��e0�~��R#���)����9�#��� �4r�$�^���)��K����T�BRۈ׽m�U�r ;}��	Cz�����}��MՈᚓ�W�#���_�W;�G�эUO~%t*�#g��ni}^<p�L,���?�[�K[� OBK�E��j�f���S��l��j��8*\�԰]k����>���PFS�.�{��b�J�_�{�~�h��1E��4ѭ����!a�'�c`�~s�O��?�Ѕ�E2q�b����#��u�ZX�<K[�d��m`��} ������?>7�8�
�s�2���F���D�`睂�"d?�S���ꯙ��4à��pI�\}J4���q��W\Q-�zj���}'��c���^�8j�K���S�M��J�7h��G/��rQ��UH-��/ hN�����\?�GEȡ�/+V��o93*�>U�n��ۖh���ò�_1���
�q>� J�[$&s�����<1e!�b�ۼ��
����&-z4���k����"/=|���i�gL��#��}#~1�Ko�c%����qэ��������5����= ȁDk�W��1k#�D�V�o2�;�+^�$K�:,�ʄ�&����ز�yb��.��)���Ͷ��ADgiG�4�������]�/#�.w�[��/[�7/��C
髣!�	 ���B�
q$���7�z[{���M!�d(iyJD�뱀.s.�����=y��|H����҇��t�U��[���F4�5V�؊��ɪj:����X���#�j�/�����~�ᖄ��X�b��W)͑2H�/�0���u	����W�ȟ��D��-�uӪ���\�}*�/��[?zl-�Qd���c*C0�D���j�qr�N�����  �DRɅ���Y}3��K>��e�oǸ�������G�_�P�R�hFV��ik5��ͤ�?��JM���D+Q>H�&[��*�~{vݟ�,��(p���qیn ����k�k@=�rU�J�3�E-� 6��k0P;�R�4�Aؖ=��N\�HkrWM�9	���E35o�"�y2Cq=w�����HE0��9�yf��G����U˹[�c�N����z�(B��HЊ�T"�Gxp�W��;6�n�� �gg���+0:P�zd.�~
�*k���+f��	����=?��%��I��k��N��5�V*�\���ސ3�1l��(W�N��e�t/�8��V8V��y�*��n�<s>��r1/wh)�%pD�5�k��"}�ڦ}��cF٘k\u*v���\E]��y����^��~|�N�%�Ҥ���V�ex v��xm��1�;�\i�Ic���f��1�Τt������UI7h@u�}T.Ɯk��ȏp�'ڥ�ٗ��2*Ԉ���#I���]�	S��"R�;��9#����⍲����>PD�QL�#�Miʙ2�OR��}�S�Q�Ǥ�l� ���Њ]�D:��MZ�{��#4HƋτv��F�P������� �\�%S+c�ӄ�*8���a|�l?�S���
��`6u�������5\עi�S&��S@�h������:lF �Ŀ��38�4�}h]���猒�u��xBs��b`bf��ES�"B��
T��q�W���I
��ux�y�n&L���=a�=��	[f�JC�U�Z�`̜Ϗ[�D�	Z��bZ,)���>�箒�EC�}��
&:-Qy����o|�w�{3ylԿ{d��L?=�zI���� y\(��a
�7n��[ ��zݤ����ހ�����C�_�M-�~��G�� G�������{A�[�]tTUh�t��e�ť��6�KO�X�䁀!,�Dk��C��²0��X��Z��oL<�:�_4'*V���A���}��
��1=
���\	��4t�!��J�F��Fj������B_lj�_���6]yg�4�7:�ktf�F���y�O��U�*y�+qZ�$��y��3:~;M_�W����:��:�H|�/�R��Vڿ��K��5ae�������Ɏ�1cI8�/,�(}�w�]^�R.�dT�"�}\R��<Jp�9ld�t7b���@b��!��LbC�s��t�/��N�������CDUZ��g�SИ�� Y�-t�R4e� ���i��K��$O�IZ�D����c{�[YX
a�%TPug�o�J�fA�a{q�n !�����"K��V��H��ȏ�j2,� bp���y�%|x�2�����	�q���A~�[P�M8f3&�'fo�OSɹ�1LGt��G�~#�ޭ�{$!k����D�;��9Nc20 ��ZO�p���kn4�������p3���@��+�=5ʭ�a��i��%�fր��W�6Qr�\�X�c�{5���^�쁟i?r�b[һAb_�"��C��k�eF�<���*�7��P��!�\u3b�&�z��m�b�U^F̉P���I�y*���=
CY.��{'�x�))�j������/n�Y[� Zey�(>XF��A��6)H���N��s�����|5�$cq�N�����},`x��A1O� $^�	|��Du6[!���[m�z:]�r_�����3[����S��~�YN��*�ل˨���N�qd�Y"z���~JgK��?O���%[b��]�E���>c��73?���AfMf
�E@���]+�I#��m{�=�.���ǚ�\C1�Z�"`������.�A��&�&�
-�_��H��(r��%�Bb��x��<Xe�vh�n��}���Y��Do�RX�+�CA�Ӄ.�ʁ�	W�2oh���1�kr�|#�K!Lp ���A�$]��@��o�RJM+�op���T[�K��P�MH�.�r��[��;��p��^ܓ�٩10�i:�JB�<�.e��A�>Y
�|*і>�m�>�1�� 2��h�G:��с��v�9b�#�Co�~C�1�kq� M[?�aq�B�9Ylc��G�1H��TN�5 �GG1�Һut^��0��+Z!�3���rg���	
�i���������c7a��AB:9r���u��ns���jp��%�w�tOr�>�O.��4�ުDE��YjG���%�X�*�(ݳ�sl�h
CmRŏ;��Yx�m\�˔Vv$�<���$G��e�P[�	���S�����R���
�!T!xf��fvK���e�,�gNG��1�A��h2��]�0���~�2��&W9����
Rq���+SNFC`�ykS ��T����� =���������J����5#9oV�y�
��_�3K�e���LG���-\'2�\}m��V�����yj_�oڛ��m�E����-�J�ؙ��'�
"~B��tQ�i�Q� ��J�Y�
��HD���e<3J|�1"�Bw�A��aF��t�S4���B�v��z�8]6��+�Xh� �
h�*�AFE�D��[c��a�'��kY���$�b3.⊳*�]���?���u�_�,4+"�8�eM�Gj�n����{+!�����'�
�wf��>5���q����
�v�"�E���)��o�ýX�n�y%jʊÇ$�涸UFr����Bi�x�sܽ�a�g�4�^���/:��)�>�ʔ���?1��]�}KA��w��]��'��:ο�t�X��w.$�P���J�r�wE�N譹���N:,]J�h���lؤJR�G�fd�C�`����a���HV�O<QΆv�����rg��~�U�(H �:ݖ��o��8I����Y�����p��U�ʵJ��<����F#Fi�c��|���N��Hc]y�POϏ摪���j�R➆�1���M^vf�>E�B&�s�@(��<�M\9)�7-��2ws����4�]���8=�6��9z-�rS*�7�q��;;E�M�hZV��� Ax��Z9Bؽ�ɧ܍��c�y�\A�Y�o�k<UM� �:4�S��ف@����glӚ�tK���㥆b-a�}YI|�I��?��{Z�ċ���>o�G����w���� �u
�h7��L��L{���zH/sڮk�s