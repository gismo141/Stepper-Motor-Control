// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
ThZVLm3zm61drQA3ctQeCJdS0S8iNSEsQgtaMa6DFNRnRPBuOzPSYXb3vq+sKMkT1+lGLuAI/LAG
qX5DreOZOAuBRD28MzxkU8h4kL38LuAaeia56kt4/N5bQ1QGlLsZ4xQXMirWgJOkclBz/UQ6AJlM
MVnaxoZN8DAo2CoFneeAiwde/IKK2EzWnzJ8T/a20q1wOJhCFWpXVov9LUNW2c/78l8zvP9anGXe
eVbL6pC3aClgY6slp6z5WUY4S0KyIORBRcN/hF/ch5hZ4wWxq/PiwcnXMqfJzkQpfzcM3Snzdk9p
GtAdpcNVOH3IXP25HlwomNMiqe7NrpgeRefQdg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
XIffv87RfC1kYCeZ189HpX7CFtSYtUvon2zDHupHDx5+rW2AYGvpejBwViblrPCKkOVbAc59QJuu
MvT10i24rcbYjsjwu4cvy7qFDz+XiMT5oM/CZJY0Mu8lwVwwD8fBnzglVn0r6bqUL845DZHANJ9K
bTD+Fdyb20u03pkGT7RwRMzqH70TLwPt+0+AsDArdzrnlu1qKu7mW676MCN3IMcqHSzin2Sg8+Hr
3R5dgv8b1SpWqmcwo0uNTHNwtA6qoZXKhTfdXSIpNNY1xd7ZMr4rxVAy79XyehlzNXWUg+FsQOHF
8cr6vi+FKDpELDf/qcsfLcXIwu3gxiAhGmr3w8BoVDcrpWtUygQhd4cJLcj5Q955bzAOd/efpPiK
/w0NFNmUhwUcnPYoK08jMeRXSZH9xR+3jm2x0kho1TxrhJNoLI1qbhzuawDC6ZOvIFOZKDjcerkM
fR5dIFjGPxB5IQ22frBRAQ5qrXjYe0F6jWnOh9NCpw+DBlW/1Oux97kcLEDe5iUXnPgDsm5Uzlat
nV4x8PeKn3Cii9clEFDtjb0CFOnWuQ9761v2XjNHzvhwpS8dYxjCXFCg+gyKUQrGX2kgGgkEZKMW
lAhkxbULbTru0le3zs3FWtHcxHIa/Fn6NvjEJCulzim3rgGBd+FYD7NbWZ4rDtjNPNkvclVmOzKF
Bm0ksWdjpPt+mgD3fFfjBkyQRN9ogEg0pVxMUvzHavJTEaZAaIWn3JuZZ2OuXYLus+9dA1MqpK/+
OqZmB7reT7jlPoU577gkf/3ZQfEepqPdBOxNm3yaWawky3w2EjxdjTariGqTvoXGGK5hmBloeo3q
FfGBK/xOOX3SvY7r5YVPpeGLgWhYQLOtyapxUjbuVWP6tLjql2VEZpJQA+HgzmGHIjlkUQ88Y+PF
Mi8pZ0LEDukAql9oV7KhVKLdVZO2aZC23ww2JWuQbagMYPKuT+UWNt2GcfeStpMA7TCQVLEbfC3s
i0SUEZIM/3Y5uc+hLb9rtYhaCT05cLTaQtKTtWMh1DdMu19yVF+ozmQPWsIYtKM/hPZSX7QA6mFx
wPKgV0BwwHU40dMjXaKTKgrCLV0TjJQ9Z7Q50S6UlQl23omr+q1RwESrNw1awCwYpbf8O9efVCG4
U136q4Gdsy7Fhh4AG3+HqJJuBY6ASDhBqhpeMAO9j2sqoR/Barurl1mGM/wcx8gsA/zuLgIxKY2K
HTccK9Y80CPgczPKjePJEW6Y2wUZkHY9iex8Zbyua6zVMyVdvbHENZyYQ/cWNaMIVEm2l/HyJSpl
Quiqhxh4Yi+8UtSUpOllBHCm9fZbsqzkN26kkP75SBpw4WQow2Cm0qoG5J5oy1VN2ujvPxLpZha3
WRRdlvAU637MqMH18uhNzu/g8hJUdaUGTjMO1LT/9xlgss4/mju3M57iwuzrL+VFsf70Z/+O8612
pCfJK4XsgCrUjEEfLfQSzEAxUpIQtzFSitUAin4P9k65L90izum/rG/Exm7GHkQw660qZT89BqV/
xBIwZVDRSf0xen+vV1fIhhwTnScse8KoXql0cWEkmrDhQA9yHzG5S3oI+WP64O+rPjdYyIsRuXPe
rAlnMecOXkN8Evfo3S/Qemp37lPRPtJ2UFOyOq5oJGqK0A1ZlCc9Y6d4yI7pbg9TknRXih6KHDSs
BTx/jEH4JMziCt6HtFo/tJg8HNG4iiiMYEa0I6wHmezw58wSRfhjp5jFay1cv/23IUMBrZ5DYwOl
HR25RHcfA7fsDcQ7e0bFYcA50VzOQmrlrVFjrA0SpBiupLZ+RGY/il0qFgX/FSggSAUvg56sD6s1
8b2hMHJSIhgeJ+kHursPaN4lAzAOO72WucbwGwkvsBWasiGTlg2o7uZw/LpWzSCzNlUP+rT/bTYD
Hwsk3/veUHIzCUNV+fubTe6WuS0hKjzSvA1x7wuoKWuWAReZ1bsyXhNNSS8VPShju/ZfwNSBuSDd
fQviiGMsgAbv5t3fAGUPikdMNyLZV6jDadTsiiPfcJbWAAJMlcx85vgmGuW7n9neE+UDm2NEfeJL
85r5lUE8+zbSCjmovbq/kIu+ddxpOJrNGeoNB+aY/yOjcAEihbW6fNQbSDtexmIn+GVBwkjl2CaI
jtIdUmHnIW+ZjxrPUNnMNQvzQn+1CE01I6HPc00EPqsPm90P4Q3k8+KyXbnHhx/VVlkB0zljsP8f
CoUWU5NUwp8WDHrgTqcunQjJFa+LF3n5Pc+RacSkviZriH0iJNa7tOcbQ/wOmZ38O5cmC++xu/Nz
HT+mQWllb57PqCJGr8QsUnQe0FM8/0fyPC6XWyiunooSbxltycJchuKalq4oA4Cy5ITGIq76qrgG
VG98qF00xZI1fouCbzflTV0ArLNlK4TjsIl8QGjO28iUzLcRrvSckyQyAU4g+C2QJfkMuZ/A36HX
csdl2J8/CqOHLj1ZqHqHZaf7+K5fXIIWPkA4GiUYoDIxLfUAQDEKW6sNvQKG9zIJ3VttpU9dmAkV
/H1oLPnoozGzy5V5tYTVyJQTQjVrLjlCvir/4ycc38YoEm5l3LfHzoZlRY99RfG8oNq4qIdF27mA
jXkKeKPKIg5Ix2r5sw8MSV9j8iaw1O5eig9oBw+7sUZxWa+imSSp1bfLewS6hY3Lbx/duhbQ68c1
Esb91s1TkJOHFDMqOi5/ir8XYdarSR25EpnUbBEA8vnPQgBRpT94Q25nhJa8sffBfvMBV6Auu5yJ
1K5L2AdAlTIXZA4cSnaHiywwdeIBlRO6O5Vizk/a9PJdpz9UWN5P7I+mhN0itAGeczX4xfcvXR1J
2Ean5TEzBWkQlBGF/H0ThgOvIpc+AB1FWrp0mW/l6UiUBQySTOWIjcHHWYjW3GVaHxNWrSZsd5DR
zFejQvKHN3qYxuRS80euN4To2N/RFoUD07g83HSk5jdZQtC4euqlTQncPojHQRPb3IZaTsOMT0TP
Y01wF0sLYPgnewbw+ewcGpo02CfRqHV/QmZOE1TH0BVSQkEBOjyNoVMzJT+CxnR5z8C2g42S//6z
V4q7/U2mtzaLqu8TtdFyM6lEXrIYRXDWHNQ72Rwjgd6XBraGFZXilGTJ4onn0gX0Y9+9oy7M0TDT
GnkDrVt9dFynGqPuARB45NgVVnGIOqAAZ7DgHUOgbbLH6iz2YMAtVXVmqwqpVXuzgqgVJ1XmEhzi
yE5G9JBUJ54QklRgsQcOxOKjuyeYsWIwb8LpFXQIf55BZ5V4+FTPNYiSVowB6NcVv0lz5y79aAON
gpDIXAJNBigVrALA5A1jpQrW+cduCTpGJ8w4N2h2YCx6tKy9SkPO4rFqke827jzdIzoT1XrINDkJ
QP/S4tWV4hW5ztjjm0q7tLVMPuxLSqbVOgT8roYJYZzBG6kinyN1SIRWf4XmEWyV+fhqWWmbukLc
23GLpPb4r/lmtAbg4TGI8/BhZcWS5S+StajLvbE05VOLf8CtTnUCuG1SQGQ3/Mo7KMA8mvBu3Abc
JTfvCRRevYwTVJx5PVpykH/H0/6NfiBMOFs3bWK1FE04jBG9tVsB/du1tHuGNvsh4HYluvLw9DiI
yla73SOPaN1wP3SWRKaflJviHmsYYkktBt7TodNtCDRsZlASvlXEq6IPW/Yojg/K0tNaVpks0yvw
26Ecy3vXZ6tk8OgxwZM6FjIYL7tcuR3fkl/oqH2EkeFryZxYS2B0ngfYz/1CobbL9h4GQ4fxQQs1
EVM6pkb96uZahs7C3K3XYTk8urD3Tjdi3SAG7wl+O80+sh4jA11QIlWaQ4zIxo3U0ns6YFrL5i0a
zDrh/Oi+j97h/rWJ0/vFaowGnrRIBHqDvoK/ZqbgJF7ScE8VV31cLUrn+DFsqerVq18RVyOJbQOn
HhvT4JLydyLeEirxNRRxNWeW76vmPw2o+berkAmOKyb63nlgDFtX5h9NzUYzxi5wbO1Oxjsz+FJD
64ByOVfqxPovzBOKN6ZDsPGCkw0aZoU30DqGF0vodeHh9lrEo9MZP/a/sH36fnvh3f1IO/VJ2LaL
1XuCBn7puP3NAoHZqbaIJiWp53NiW3+mLoJQ1v719lSMXkqeqFrs+zqjzRp3sdFXW/+nYbJxfAh1
40PHpx8c2rhnZYyHeWv6KNIuuCjfG8KbPUP7McGQRyKO4ws2ITPeYS6O9hrYHMNKCo7fvuMC09xI
YAusoSW1jxpgQFRjEb2BUQ4DNEcgAVKNvIgjol52D8pRsJQnPx1aZ0zt3aKl5/Knt5EzrSvxAc+1
ix12nBzi6HHKkhcrQcLVW6SPkaZATyF796K6hO+Jfj628RfbIGgCWflKtjHccwPCh80TXUsjBeL3
aR7v81va/GZe+ylL6sqbP96t1IqbXWisnx9vzTRxETHiUsK67Se32W5GMzhvYalHoRyyeRDkdLw2
vnZhIsMDQUpNTGKhTGgPQU0QYGpq3SqpAhPx6HHDzf3/wKBAWTLLml7GusqbabpLZXQLe7IzU1D7
gUrbwOs4KZdwTWv62x7Uy7qlvvvtzBl2ao3n0MWOwGW34xg35lpWeiPlotjjE8jcWJ5tRIJ8ei71
Qt7l16O3IpnpyrHkze6qG5dFLQv+iWM47Xv2wep3UfcbhiQAej894TI9EVXQl7qMsL8gzGOpkH69
ciG2H8zecSQOeAsyFDtwiy7jfvgKiaSyY7xbFYMyilqG/vs5PCq5uWuDkUCjnIjCDKcfdJeUr6XE
BM6ub8flRjtgQeWJdT6UFRu6VpjbFdDXRuhfwGIN6BBrC0XjWFLehGmyYzeoBKgkoMQHVuCMkUZy
EwMbrU41aCJBDUIQSra+TVu/U1EQflvd6AycOugu7P2sLEr2m7it1DLAI/YpuNZI3RJD2SfuJvoZ
Z+DC6eLGuox2tO14gGYdis2nsdEMagTk9N3Tkpkd6X2Xao2r0elDxvxy4daf10pjezuKJJJvMw3L
0GuqZsWxNPt2reE8JN+y4IGtk+cljGGD98EPEsgcqU12t+VrveD79TqcsAmNTqVs+81xe+EGWLvX
3IU+K/B7PjiPRmqMvG+yRqfCxiPaWg1PBJsfuzLHAI8+UfT7DxxEGWEbohC+dQiM+Pkj/pp8ajNU
f7CuUDGKKM21jIwgAlg4tWf0+WFjZMAAY4++QuoTEk2EsmS8+oV1TO/zolX2ePbDY8s8ls9+62y8
XlEBFDumlaCJr2TJ9qMl+lzB1V5GcDpJyFoiozdnLpfAfYs+854kaGDFCSuNcEkja6MWy7QaSJtB
GiDQ7QmwAYNKLi1eP/jNk1Lkgr0t9tni/dVldEDZ+1SKEGypByyX7xO0gNm1qfxsoci2Ph1fT77t
531IgzciWbVWkiOFHJaGH0hqpfTVnM6kuOZiGzNFPBV79XZ14QpQKTqJ0wyy2ADQIwtoun0hJCiQ
hp9fp3RUCWQJItvPIlefz38mavdXT3Wi/2mjtziB1m6TUcDzlq/X3dY0DxeCfhkcJlLgbvZGi0mb
MDjdZ4WUOevB3mfaWZedBbiO1HQhCEJ6TiKThYkm/0Vv9DRCVO235KSREs7avwthFFGUIvmM/3rz
anvCzTtUiaQ+hpf20G8kAlfeGDKNR81jQq+z5bkN/4kr8SUII1XFyQu5xQ2fimT1P7aUiMh2LDQ1
mWy+Z7WH6iWkr+KnXBxFGKFYebD4/7gyn0BOxhz7HfIDcHO2T6yZ8UAPEFiR+idU0tRMA5LkVflL
pQXk9dInD3Ar//FLTBUhjvXnU+I7PzELnQ1HysolpHqHAivuaWTYeCi9sCHOCQ/hCOYKbf00R1Mj
CFEXOJnaYi2faqMIgEbwRYqnKmN7LULLz/yhIZvcIzeZrMIcevfaAY0jIYql6hToI2MmSxFTA8B9
S1SiBFwVR5z/1GDNbZgIXdKPM+oX/5zY2GDccu3iBNlMgSVMz4m4gQ/h07xcO8sQ7x6Kuj5FGc2V
sjczd3LW3HWsbHZdCZS0Db/6V+NoHthipCliYU2uWYbrEDfM6caqJU2NbQf1nRyMJa47JYiyrtXx
1AYvJI3uuXV3k4b+wzR66fLrKokn3fLPHXQCVBcpT3SB1/rb4CjU64kO6v7aBpMjB3KVjCsw7faJ
ors26y9eWPn2SU6/lAuAZWi5lcrsHMdP//8RKE865bCLlEVcB/vbiAUwYBmm8jHcsZoqJX6Gi9e3
hYAdvapc+dEOc8013vjb55z8xO3tC66cWYrSfbA3lGfBVg2080VpSZyjLVlTHYMsdvIXm8jNYTyp
BLa/9VQ1CwvjuQWAc/IuMJdlKjWLcJYPn+bSjXEh/xZHQiitPS4xp+UtZA+tmnVCDTC1kCgGzmXS
EfgjgbLPpkH2OJ3CyYKnUC62BS51ZAml7lfJidacNRRVgSYFCUcMjJTYNMlthg0H+krJ/laaG2ql
GsZUHOLbYHhr5BV/H0ZPxbk17Xc/W9TpeqSZAQo8K2bTjFOcyV3N+h7zYb61NNXVUQYgdAhaXrOI
c9KyDnvo5eS/14w/iVZL1KfNpR9pQ7sm/30kIVqTbsIPoFmAYitl0bCrh2E3mIab5XtRbrYnl7oY
hzar1ECzckh/3iRgQ7wJWAQiiaI0/Gam1RuooIqipequvRYs3mvyUDF3z48WWAkcjM8ogTGz6bcs
gtnYnTahJEGRfkYuBAJoCyOpnBkOCgZ/a22FyoimQsqa3DNwtBfGpw0QfSUGD7TQ9yg6Z19WDwm9
1DJZexrZGGaZsvZ51y33rYTLklSSPCo0kK9ogOX1qWgzRDFo/sq6p57JUADY/1TIKTSZ+e8R7iyj
HWFeEC140qJxt2oujQDLVdSoCznx7N6amtAfUAv9VXUFwe8zRyYfGbBf69F8goNxN2cW7fT2u2Mr
8TBzvLfcOuzqj/yds+PMZqPShEYwOE3+5zNKhSWpzqjHeLoIi7jHRVQrNx0PAubekkCBtmoIAObS
L1NT5KdUVM0bIafxUcV5I4pguuO7TuRg1dfqOZO61SEPd8jdsUNaLCBFV25Lna5xBQ+WHYEjFpFT
2maYKpMzz2qK6Uu/TUXAhBHApe8HL4W4z6+YGWKUfMaQlgil5OJd521hlnjFIMWGGiPH0GzLILDd
dEw99jztcQmFIu2KLnpc/ksCG5rRuuaSM34AGI9MlpUsXiMlfA/DR2XOc68ix/R3s8wj602T7fxH
jF+G9SMv97SgiM22Z00q/mVtKGSf4WOyvuTac7UbPmrLLuzJgYY+j/eobxn7m+o+M78o30H2w6YZ
e/3O5Xs484FFfcYt+5N2VvScXKYJwdwvaSHcXuvXMllbJA35ZDW6yGK5i8UM5PztCkiySgGXGio/
OI7Uqyv/LZBjUekozR7NDw==
`pragma protect end_protected
