// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:48 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
k0MIyRHbq2bwrOAHl4pfFCVWokxevGzSVLb/Hc4e71UguJp4wIAwAkNtMvzTlsEb
uV3ozK+8KEX/2X77/A3cXBaFryFrz2qD2KCTNIwN1w3+dl8LGcqOjdfXY+waUWhs
RCuRCW6zTRlc6s/cXOw0zE2DAuSG/qPEnIYpvm+awZM=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12064)
xtZTkA5lJvVGFJ21qu6ez267T5jBqgnW6ERU7OLUKbX6sVVTVJ2M1ZJCPuAmDzWQ
dIUF8LCMyWFGKB3XPSZoo+mDkplq3jSAIhQNVvmrx1vdyhLgkdBLxkHJmTo5eGYJ
gfmV51+97MuM1RipD+zF9eR9qSwF928UczQ1R08otDdriP5HB7Qg8e6eKRc7DSBz
pKB5Y2BlBYUmXlCpj+KnvtKi+be+zJANMS1I57Z+cGgplAwzzZxL2Hq5uKGEElYE
MwGLwlg/+3mTlzdPp4MKnug213hSZC1W90TbkvWrblAVkiiDduSq/h8ij6HZI/UB
cuBsYJTDIm9GRCaYqnxrvEIQdLzk9s3x/OJwr8LuUKMi6Ma2+aSY6g4RfkbqXHwM
r8Gzi4bledUghKBBB5WfyA4ogtq8vCwGwMkfRgjkKlXhuykeL3GBLa0CNyuHOs+5
yrx5h1Vx85CJv2HgEpRc9JaIqRQhkERRxSJVsZP2+oCARk84lJH+wwSJTppXuyGl
PxbzEiIgLm3UqkdBOqCkXZEx8AFBD8zW3746FSokwnlGlgcIonfKmlmxm534WuQ/
m94/TF0L87HBIl1tPgaD3mwnmeQ/yvdoB9dFGD0RFy0OIQ9v5xQL4hDvLS9780fW
nPGvF3X+8vpMF4s5gqMugknaeqjgQ3+tbL/F5m+FsJljPSdJ+v+3d+N5NdfAFV5F
RjeWwLUyiRQWIJX+0++kHfoJg23CmzumRc7AkQXew0WLFCzkAqIRt+RrSfcxjj5b
jXIRsp0NyuCQ/5TzGk/AE71P44JkPGBxY7I5sStJmXIwFWRim4SpC+BjGDVY4HfP
ncAQ0tiBAC2CdEM7KJFUUtROUTt3J26aV3ZMpWbNHWy/WsxX/ym/na1vH34sfmkV
tkWY70Sdw40UscEDyosneKnlhxzQPUu5ygSPTxYu+ZAaF9mLKmNyeDePEa4a8lxF
i8owY6qxkpMB/59Pt1PU3oNoUpbMlQi7kXEM6k8ylwAYdqRh0B4i/jjl453skJ3c
uDZFXopCWiq0YO58VdIMrM/CNzfmXb4h+QI+BNuC3cmceMXhkPkv5KjWiU08NfLh
6zS0LIeHKhKZFtsWtXUH+MMdjq7ot2aDhO6LlPWzP4qBScYCFpSC6g7WaTV7EBZA
PdlOjmLpTqItCe3g6n4Ebzq8BDZDtQeMwNuQel6RWvktwtMhkkUMrsfuroz17dZC
dnC4J9yTZ+XZEzvCCwmLWeO0C/FDl/9eZRiwzDBBHja3NLtOoyPihpNXg94HjjUb
0KSF+fDQsPon4rGzU7/Fx0Ab4AvAz5AEiXgTRgGUejJMvoAqkamy3L/2EjetrX3H
FE0bgXVdvFkLXpS8k7ksWohPX5EELm5sMLV1qJ4gRhoGtHPXrOgkEc4HA+W7ECs9
KIHryzTNcdtOdZn/j87GsktD57I7VWzgFRSJMcRSk8qX0CpqLzil7lGo9Z73ehC+
Abywe7Kyt62Sglltbw+7v9Sw+MiJ+H48bbTbblAuipw6DWdcc+XEsYl41sod7wNh
pobBGjVY/wLLG0cfn26pJ771LpVhC5PYhpUoj/nWKSyjnJjJbBPaWrWQ3+vh7E4q
/+zR5WF92OaNk1co0Nlnx1vmIuc5JxIGvnt5TL7w2kdQ9FTF0NGBUnDpuq0ptYv7
wfMH11u+DPqjMAbBIQxqMdZJ6ptYnreyGSdJRXe1AWzr2VQQCPKBZzh+bRXEr5Y4
Y5g5M9X27oZMjKaZXQDidbPreGpwNuTI4XoHYQuwuA/2eP330BuIPl002hTaReT7
mQ4nwlD1FoaT+vwQQ5X6gU/gFn2TgTdf191mPNXxyy7M61qNtBlINrBCZbaO0apf
P56MsUv93UwxEGLBJkjn/afxJA5Kppl6J4jfcqU4TiudxTeyfLRdcjqZ6yCay0+X
3c9TWawC2s12IFSLldixfF/kpo5bJWzyKk/zmmJ9p2tkAOReH+riFZVkOurhWp4h
eQzDUIPk6tbx+To9eRGFUt7jQTj46tSt9rLkA5BLmvKJSgjTjjXOgcl4x75gnps+
scF58dtLueZxpV+4WW7DQApaq5HW89+XMcjRx+Vtrec4L0F3c+ed8R4AyXUv3ZBQ
UtnrICK6TaB4Wf9WXoHsIdd9PCzZzD9LS7nYtzcljIhowc6TWHbFwbtUSecHqb7B
VsE/soxNn2ROw2cmVaEkF7Cysvx4liWrW/e1r8b5tk+5QNr6//y2sR70CRIlKcVN
0gDJlh/6za03yPWJXvmEFNJ03REE8I73K0PW4QvAkqoN+iGyLApdTNbwgZxztV9n
B3XsBwqZtPA0nca8Jr4NRAn0mGB6jZ2P1mA4YuKcS7QqlyQ5YvR9dtytg4ZzOKHU
fAXvh3BDzvVt22giE+bfYP3E2QGaddF5geRP8ntHdzpJALWWrhXbCHAUhKKDxl/1
gefXn+Uko6/4YhvkKDYZOz+ejCZp/IgJ/K5kcujIISWVdgR3vN3KBcRxmdEMddIB
AqfXL7nf2leApoq5a1iAWlVWk+wA/VrnVcbD0zOOzCDYxQN0/RPNtDxKcCn2DhdQ
7yEbpyg7/YrF/jiBFO2gAiBwPTTJRD5OjolLv7JlvBtAP/zhxCcwZYutioVJA86N
rX63p7FUZfCMKFyD/psey7khTMleRsWgch3r+Wi2WZsO629sRVO9eNX0pCqw4wB5
eKNlawvesj7NCn6HXy6bpseBfcwVLDQgGrXtCE8UrCz7Fio4K4iH+ZdZ2w68J6o2
kQhd23lTSKZni8qFOqbUFdfhH10vR40fROJrrVG7Pqs9eMqsFAyTOBlL3RZJuny0
FNMJWrVJkweqXjTSAQ8X4XVJTaxp58bpBv3224BGy3gcZHzUhKVFycA/d1r9WDKc
zDYRo3lFiYGN5VN5/p0TM/LRra1jFZiaoeAeON9Ah6LNc/BE/k2e0gD6llsOdOCx
Cm3eQagy60Ph32yf/XzDDY5sw0b3SbaoVpq56yRadqaDnGftU/zXY/kSk9I1Ssdl
pM/mlooAEU/+x1rvVkO3563+HA9whylMEIDg+lPHPYHYEZL1rv85drR+9/ZGYJ13
V+A5Z6sw+iAbtSDcsDdISQvZsYI9bGCgym2z/7drbIM34lIE417WrQn/87K5Pemn
JSRj1P5mb3rSXHFjVyKevfs1+KIoeIzflpQpj3h6vcDKURayKfMWf/VgWCiioKXP
AY53Eu/o7X4pLUTG1Xngy3rtR6RLH/nYf09aZ+TFjxUKdjyy1OVuoBDtUiKO/63B
WKgZp8T89sx5juR0RqCIcI6CnTqGgSeTRb4OxaTyANM+yQ1Zpg8CqD4Y8wxmfSk6
Qu69YcN0hyagCkqyr1xTWmWVTzcMD0IsU17i5BbOXVVXXZP3BY9zvchf4kbE+5ym
HXcpXQwgNDKnFtAFLXGtz0FURem9Qi9hK4VGb9gejgW8sa6glGx/QC5FRQbkkWf1
KXSL/9D0a5KjDic9hrX8HYJEsqgnokq91yxuz9YlQFI8Zs8jIXMRJ28cKZsFG2Da
fKrPEH3N738gwstSmeGn08Unye6Vd1NM5V+O5113ARuYFL2lwMArzUqVOzf4O8tJ
cMl1malsr2sJTaksyEzqTYOUkSN5cidwF2dFYo3tDfaIqvOPy1xKPVZ/+ETP3at9
by6Qb3K51AZUPDi2ErmG6O+tfM3KaTWpH70eIjb8twwalNjslvJqG/HkoTCotGqs
UX6yJxUIU8jFPP6LfKlKC7+kJX8aiikF0sKBBtbEiY/HZhaBBbqcSNmsscvS/s//
kmp1pyiXNXGfQZ39D7hfychtOS1nvPEoeaNMbv1QHxlNGWGnDjoBIp4lFnr/5l+K
ZPdnznrr4QFpeRgDQRRI2he6b45IQsWT0V+HihH2nMTlu6g9MexZvm5ltE3CzD6t
4MVD0/MXlsKa/tGcStGg8Sx+aTTn2R6trr7/aS1U6eTcg9vfrVrDJPzejFMUcWWY
TX422+8rsMwvC0lIXpWxCNcIZT0GfpCMnMXMDGliNoJ1k9YdNhzqJ+bpdop7aTm1
eshE9L21jKVmafsDFHsw3dzpIyzP99Xw8IuiVBv0UMGZ3gQyTwUnXvfndkgww9+H
4p0bkK8VqHF2KrAR1BzN/8jFLu6eb2gv9gC5/MtSbs3CnrOIfpkoyJQbj4AKJ7aY
tx8fnEZ+xhTcJfyBDULei0Vsi+kYoUxH56VlBDqnQsBReEOxX8jdUEYKvyWdK5B6
ZdHoUr9mpe5P5VGYAXW3dUI//xHJThvU3yVTby0BMNjzGtYT6EK8uRrvowhJCrOl
gkhtaBk7l4FgxvvQgJ6YYgEn0A2DMg77+brVgU3cn4PMZT1/mYYA6VMvDTnuPovO
nWRbjUcxl40K94i1Jh1192ppfOuJosCsvY91jWE2nJ/CY+7wH1Gpri37MPJD7hL9
5Trjrv+tUMsTP5O3wtGSoV+okBtATaP/UZ2URsX/km5bHOv3BT7dFjRMr+RkKLjC
bPEoI1qou4GWHVMj4ROgI0Mqap/ExQGqOSBJu1C2juPAfeoAEWbpqd+dn4o+AJn0
W5p63Fp7D6z5sAyrGfbZORwLkTlR2qp1pOiqm/b01LjI27RbbfQ+fNZyWsfRA2d9
ZEIbvfNp/E6ZZNzt8ga9mxAxkwotvqEvZKoK9169d15fiMRLJKfhXEwyvNFR2iew
efizNoKB2wcakAt+l0ccct/PonHIJH1dAn01kinu57Z4j7JK/5PqOaGkJNoEQ1cs
e/3uuVkfS30UEh6pnTanEsNLETGf/1nMOqd3TmAs4uwIh/6xeeJFG4JXPKao5/6W
OP7b9d7Ro0JG/+qIKhoKbaInuQK6wxhui0msZ6fnbAvENIcJyqYUNAJMjeHkMAm4
y/60bRAAgB8ddyaw7XIDCVLu1/PKUg9yT9dBJ/0bssdO/MMAdXdUSaOcGSanu6B4
pnRi8LtU5CUIgP6AqFnNlLm/7pbgY28l8udaO0VJz7qg/mGQgc0NAfs/iYJbI2lb
06WKbD6TReaNFMgn7q7l6upCADVV+zblN3ukuSxbdawafbRdyfEW2gEgp3NLX90m
iHe2hMJAqDrjbsSp4LDMlIA9oMg7P5+fxph+V3a+5rxqe3lT59UdRwM9ZOv4VH3r
a3I/NScLoycWOxMQgf3YQ4KSW2FAEZvmCwsLms2Dzl+eFkA1D4rRwPxhqdudcQc8
LHUB28OxNDTGezgNzczAjIdn8HXdvm6bI9cMXazv6JInrgNyxoQu8q11NlxZd1lw
xghvlsxevVg7BePe4G28wJb/0ucxVQ8sjty/mHMwdThH8xvmGDFslk6eSf7AiQz7
JGna91+Fc4KkZg+SqYaJNKiNHUd9nYmwcvGpMNfQ7ktiOv0JS31iN2e+tEbrXHt4
SZqHQaehdhJV3tEMSy27ODKTU18sHAkm4Ya/mWsz2yF5zH9fHk8DXHJ9P9GWNvk+
j8Jt1HguStS94Y4UleMNtt5gNfVEl1xShGr8BI9FyQOP8I1/jxOjKdgb0HkhVnOI
TePzJiq4lcKkjewG4A4V89Zxp3m19iWquZg4NFqahk9QBLdB9n1Vnrlz43kSs0iL
ydh1UsiEHcAMDsZcgqcRGxUSK1MdzYdvARE5Z5j2wEAYnvn/RdL/lTexGQujdufq
8TEvnkLzvkKNT/F7CSwfJ2ePdWEAy9rFwV0IfEDPc6aS/CGiAvRLTP9e6UuFtuGg
L32wvB32VCFznSmp+TEq+nE2Uvv55dk1gXqCjdF//uKnll0p+AyHH/zthDtUrXI4
AODHDLsytzxabKCDDqqEqtfZp68I5YHyCzu5gX17L4qbgGZqnndS8nPjuZ9x35XF
dnterRBfsIiWd3ypx08UjrTazCY5hkjevHIhg6R9eSjR2JEJY+EuySPplSoCcE19
L0dj8rnwxitrv/bPm76+W9JtoCWkYKKxi6b2Zd1Jsa450TJ9DBU5SVsg+VdAKJ/u
AHe221htR35kCcRcw0AZeWqTrbs4JLzKuVm1BOq4qOEGYLqFjvQnH0fNAOJCbCXN
MNFI6E4qqc9UjZI3ycxD6IZpOJXgCzkNiZgVyA5W7uNEjkCLjhclDtmVJNRQHDSp
TmeM5B0N7jQVgj1ozynk8v8b+qd6a06jXCaoNyzl+TR5lLpLNCfo3Vn/eA8hAylT
U7pXQwno6DN2VMpx/oW5It22cNbtk9KkSPQhMzWP0vO1HIWcH/BV8jvQrqmAj8bH
AUlK7Eq67XLZ6xmTaz+GtOR9bzPf86zNVBqSBbVLGhnzJHL+qfNeH5+ZMUoLf7bv
oHkN3r5YcKURzaGxa5r/7JuefqJcdrmex06PJlTqupv2RuD9vVlc33HLv6nxe/ek
2kUyONhbUuhRaj50K8fHfKS26A2o0kpo2+yWu6RkNhqIRMiMHJmlxian3PcpHjkp
tJGPLqxEv93w9yHx4gtqliZehvWXJ+SEfgJmCSmCCiS8WQHSpz13GnwbMn73ZQGF
m/LE8j7OA7T7app+ge7o1jckafOBGbsZTkM7YecqcD2vRx+Y+JyqCbyLHoaY+nKr
AHbo/dw0ts7qd2sz+y3/ilwPDlxQZQSWsnAeWucao0AsjTdzW3smZqvNX6oGoZow
Czr9t855lYMae77FYS6c7aAGjYd1rEzmlHeKaxpQui/MpdITUGN32VK6sAUXL+Ol
9OTWtX0ulbgP7ZYbt1QT2nQ0ZKaXpl6Viun/DuMS3NyyVWI5tArcqJfptj7oD7Z0
jms8wfww2Bxza72bZfQ8CHdX/iPiNGqEuG23O8ALzmS0dACss+7TVBlkJe1VgVlU
T3+rejGJQUYFAKSeS6yIYh2LxLM04Zjp89Dpxb3uvRVqmGOqAe6KX8Uw1efmXgWi
kGsAZYWJVQiodn/LloBqYeNRXl6tebysxyRSp3UbcauGzd7Y5sM9SCDovrVWnYcO
AF78LMnJZv2bPgPUoBFeizHetPtIZq6DyWVljJLf4GWZgf9+Tq8Io6tbb4kF/dqp
ksayokWDM4+8+5tuov5IN8F7XFefFXIL4DXM5wWt05lSa2qi2c+ERFagXGTqfSA5
lnyLJNvmVFqcPDci8/3L3jVIbar+04SKJ5dFyrj2MApWp5MhOkZaZ0Gaad4e6cGx
BaziKw8AD+nVK82BvLTNnDBdxyS4GgQdelz06IwWG3BVWLrxaua9IvX0/gex7RIC
5xpM7EymZ8WM/Z+5SL/1wbPeRIifiJybY7BKbk+YO9CkgUefeuojXmeCekttkBWa
o38VZhdLK4WRSnpAUdgFx299wrfRsPrxrcpfT0ajphFu6M/s4WtNMYG1Tob8lOli
/dZz51tbtMTbvmCTpLdBwskr8HMet4/LFTAOiSGxPGrHjrROLSH316gLpAjYf4sL
zxjFiaGRv+21++7smNqaynQG5fui+aWloQLLsNjHpeznvEDmMwasdICMEd+Osc47
MeLusk/h4Ycp0LVwO5aO4FrrtOvOJctQy399rI83YyUnixkEjnQ16YBhSUPgQ2aB
7R2uKFkTEKSqxbWUUlfL0hqHBOAcJM2R6Y9ViQpxfwdl8y3M6ABTjP3qeYOrkYte
Q0dTTGyBGyu55LLm6DQ8f+Lt3hp0bO4sOCfxqjkLmoGH0UFUJrOEWnnmIjbgVOm8
lKI/1EbN8YlSIME1IZZWPNmJHSmPn3NaRNmEYVuLUjd0/3UExCy/HOMExk3wgHX6
TLHifqzjj6vlC4sOWMRQjL1BvlBdK6FPi6dBGjhr4FoVY7prxmqZJBww/IZnhWcb
ece22OTCZjR3MLKxHereSCr1970440DP+oHx/ZBCl3nxel6uGff5besNApnuQNDL
Z/4Uaub+Y9En9J+DuBzQ5tkrJf4Q1LU7UvpFsvbK9qyQpHTVXWtCoVRQGAgougiH
ImqiLTwLAxoXdgdZM8QIWHd3qznTwY4F+FjP59XtJL/mNhm5c6rqDxmWuExQPIsf
IG50isdYZwDEZDIfr0U9A0ufgYmu+/12zhRkMCqMACvnxF5/ltXlPQS4yq21GP3a
YlXRk/nJroeM2ROpCFnJB32ajPfA3waiaI0/fxSaVE/+6LL9P8DXo8fURc4HD+Ow
AVf098m2ZiJjv/0W8ADEIAU72YaKAQjepIjHmbbDHOw50Q9ghbcyiRjlP4usrEi+
Rx3ZKAhfW4jJzBwM+uLof4o0oFKgHB8bKLmhOSUaOxpp4m63/+coHA1oWgaMMIcz
XDUbWwF2jdZ3Miy47a9iUCw1Ll2M/BMeA7Qp+rVSN4ChVpFwI78pkd1qPzyUflaD
A8HT63/SiAvMpx2oJkLc0zh1WkSK79xBwNhyUMjTVtuIaAXfilj37xyvmImX+dB9
zBTb6YsK/lV+3xH8K/53A21RGopobfCUTYy0XvG9eda76xWTHPOwIIJNoWE30QZe
Fy6WHlby6F/p8ZqsTpxXeABURd1xNb1M/IwhMda8b6D8uNqUJ0muMnuOkCR8JqS9
FBn0KwRZG070NZhUafQpvto8P25Eq7YwujS33CCzcYad1WwYqHcc5SvHN48hQ4nB
3PFHLWPf6UIiVEVHdHdfLom3T8hicweDCSnUIgkK6BiKIVIL2PBI5naVBfilwnH6
sr/9I76TCtM7enRWPI6Zs73rhFqV0L9RW4funbSF0D2vGV+dZRYeMcx/m+O1wbBl
z3MedosymGoyUet0Yauz2R7zOZoYI1rxJWfOIAkr2qJ5Ahx8cndU8+cjvb0lx7WZ
fF83j3sSmUOYhD6hNzyTYG7Q3vLl01BmvxTIEPaGM+vLkcSyPE9qpWniCfVLsNlZ
ySdtFlxlqFUayfT0jppZlqP3YFEcvMXQHEU7ABCQsURZ/+UCQkB3KEcybcoJwjem
qzFuQnYTvoMKuAkezbtNf1GlU7BqgxUUX5RFVXTvtL7ed12P67Uukp5QNAG1RRlJ
v/dtgIpyBFE8rcqVOsUKErTC/qgDOGyRCd9D1mTX3ZrSZEY6uVmKHVzRoBMhX3UH
Ikfz8cY3kzRrfGVUSIr/dwLc/+mU42DEjA27IfKiKQLcbCYIrBlLciDL1k5oSfTq
oZZFlDFzUBxxSTuVJRgA/iqgRlWk58On4OtLE8c81BhlSqq+bPWlPw6/a5jVMX5o
93tjy4s2uDMKPkZzmblgMgLorjeFpzpczHo9vMEp0KftghojjnpuqSUolfHCWnFO
nxYzSWLwh1z63Eh26qEII0WW5mRdJMZaXsCrpJJKFBzm6Il0IwC7k4nxc3mb3cmI
j+uCSWMogQ9loqYZe7xUsnvzSLLZXfc87h7ccpUwdOOueVHnpEgujuDMKuL3sVyl
B0wSAt1GZiKmJgX+Dp30qhK1VavemY4Qo7ZW0hQKyGQhckLfOBZ8XteYOTMaDB1A
cVlQqNQd4SH0qr7EfCoEhqtD+thoBVliyf10WTw2zD0XiOLJ18AH8k9rFJnpao5s
LJa9utMASE02+A3z/zjzeMSASOZ6ZCcdm7HmbMQpiQT+nJr53ryGr9tXLBGE/+ab
MQOizemZ+mB88c7sVqtUwWmG1gunYIsjqPnibE3CJ/JfrI/cWVEs7tRiEvhcITjL
rcT7CBLBQXun6dtz/anDvP4CP0MVx7J4Y4OC6/fo/68aOlbIlzNeDOybZ4TH8TdO
/FbPmUfPv0sehT5/hdeDYTja2xYRTAZYkwoGrqVXYAIBCp0Znz+RlZHLvpbba0Fb
ioRr5GszyELCS30fhyY3CL2cZKDlIXlyIX55uapIAHlJC/CD0MKVq832Jltfi/xW
IkOIj6Q2uwxxBMkdA5Bfvbf+ClwAF3TI8MYU30680f2xn7QKK9jimo1PuVBTckuU
5CKe6Hu7d51L4WqT4fO5nI459EwWdYVTRj8U/6Ac7M8Y3csRf2jLHLuvUxOzfyv3
+b8qrtP+P/vdrC0xITw7P9LOKz49Nn74W/w9mOR8cx8b40Tk0HpmggEyiiqisWCv
7vRSfsMq7W0L3PcIi4NEvDu3E7ANe/JKUfxDvnxXYg4O9klRRD7GKVAuLAH0TIdR
zb2DQ/WZGBcUx60e4k0YgdC7ITUEUf/M1O5ZMc2Bs1o0ok1CSAPtRMadfH0rhsd/
7WlGe/wr8TNry8BBqkoemWh1oyt+Oq1fhyhZGAomFxEsJYGvVDMTPfo7bADaaFv+
VRxvTrOz17WEHmhmOc5S+urXeOcWIvyfq3AN409wV15mfsNFB4Rc9Q7tUdY05n95
EdBGZmM5Mj7c4YWVRVv6GbiKTY3Z9OUuDXuLXjphiYuFV4vIdXNMYlK49o3TM+ZB
8Kk/0Q9c/pDsqIqi4q/M15qdVvw2tRlXUODYZSf7ULTMv4sHAmwMkCdc1yb+pV0M
sZ/hqN8SAwmMwxCgJoya4UXTnbPBBYZ//o5/1p/+UN1vnjmFfgBzXLh45F+fS82k
tOxMYGZu9LA6jmzmVFn1nG95xCRzEk+mEngNixUiek5kSHzLlM9Jqjk8mTmCMLGd
pIXn9KEVn2QIF1GraBb3z2HhoonXiN4jIa6XRIaInK6QCJC0NrsTp/ElLukQqFaU
nO0u4dhqYGqdcSe2bLAcP+p0ovBdICmGwH+DqIQ+gBtYVU/BjNBvBPsNtIu9M4Vb
AXGz347B5/oZUAJx+14CAfNb6Dbe7iODVOMtz8Bw1DCX9pwdyvxzIURzVfOQSNhN
QGpxLEaZ8tzMOrK8XSZ9TSqsK9dxZHjWwEha4v9cozEXCnWyLxQY1qy22NZmL+Id
8af4MJPCvqyXTcJNGgcbcyCd7trMAW3o6UhW0mQP36tbLe8qV6b4ZYepqTEcTzaI
iX+/jwqhFXlYtpKGnfOVG28oYesoYerEsymLNJEsYQZg4KheiAr7rZdZ6ZlE0ltR
62hgPv+XaQav9x6R42y/Dl4lqpSl7/PXX00msB1P+RrfeLHTViJ9FsrN1oZeTY9Z
5xt7GvkoO7ZpyGq0PgfJtcRjSUv3YvXjL+tAJdD9fHuqD5/JZO4Rg/5bGJoze1yg
xGaMFbEC3BfX8Gq2RoIhWDOgUCoZgx27kdxBdJS5zHzivVG2JkxZ2Sig676+pQwX
lu0XPEgvHSgPxlHgmGDi/QJYOpF4XWfIfSOM8sP6d8v2ciZlUigdNT9Ek1MUdkH5
wZrbVwKsmVAFxkTSjRiDR72CaFOGJcuhn1mb5LzMuCf9o4EN4almRNZrFQU1AQbc
POz7pOaaMr03wxoCbNoN2LQqFbkj6u2IiXVUw2SWyt0UItiISx39/tbhejO/8reC
FjSAotIbBwrbdq8eBT9AlaU7my2E2l/mR2Rpbyr9KdPkIRRKDD4JRhG8Ahyqg4DS
JA0x+hD3y5GvZnhoVcMSvLPR/fenShrWJsOxpKOijLevF/ItqQbJBLKffELUpP1/
/wBytm1IlCIVXv7+d/k/jgxS3t9neO8922019CCghtNnPSmGk1JGA61ovGlx3pTn
YVTaMq4/hKNX/RPYq0uPcriyhHEbAdy8sssA7cJJMkfsz6TV0d7ELVlKwtF4IXx8
5jZjmv4sPad0O+Q/VhibHOVQky+zWOiCX/YsF3S2ZvYDk0J9cCZOWnlek0MDZHfF
3LpJ1gVGySXNOjXdgcvtyGnKljI6xR8uD+zOriPuphdvRyNkZjwaZuPYbaLR2fcX
ydbyW/q2gdnSxvF+0DuKK19XbIchvP6MsxGfjJQrl2ezz8D0a//UNoXxSeeWFI9C
6kQBcIKeTWghhnc9eoTaRjHNEJklvw1RVxfvgIxIEZR/B2kXufa/jMqveXDqKatj
Ul2Z9SLviuwu23j6u9xJZS9zRNkVd/LY0G2JLcJE9hPCt6Do0uJcvTK5loAnI8Bf
fH2T1Bh7T53GaQzeozICNWE1030zMR3mX7LpBvsBZBBYPymJM5ux523UxoJoxnBJ
0Vy8AuwvZZU76AbI+Q+T95xVx9kemOsttU/S6WP7pcmmB84DkwSmXv/r6TTxau+8
02uBhEbshanXEmUYUObav68WaQ2rkY3PHvKdYFcWd2N+PNTmdwS+eZfTTxBRkBD6
SFIserdDWu3/ID0i1zuEXrcd+4c5LGiPizLxhMpFnzpatiBrbwWNnlZlodiJNET7
15j6SoN4+tlkDFd5+ircKQmuJLHomlw7KTLknrRe5qUQ1TL7cBMGgN3urN8s6m7w
HkR6VU+DlL9jts1UUJoyEXkuROXq3NsqyEIH9jyE5Z0bSw/4BBmknRW22+CypXeR
eYJZiMs+AcwzkBU+gouKiCK3UvykqI+kmO2bMWkpIweZXTzKLH3SWH3sLThAfNUX
QWJvM5/XbqULEe7c3WIKt/G5q40cYmQpGq/vPigVB9B1RLRO9rnDV09OA5ZEcaw9
31LkzFQj4RXCAcZV+YHWk3vQkOeexyLrGGTOUaF6FHmrYTaEYMCOBRaOYwBRfW+a
9DfkL4+AgXkMPhyNlNoQHedpY56nCthhKWUJ+VEN/6D6wgIhvYUN/M45QbOVwsmd
Plxc+W0r4dxjznhNuQpu9I9n11uo8bVh+NdkJHnbNW/59zfc2vWl3O6VuYTn0ycT
Rds6p2CHRZVvQUzjPLAmgPuTnvfa4TV18WrDQ/Ow1ZkiFE9irj9IXUCipBAjN4Tj
JeA7TcLH38gisMamLitBVyn6qH/3YSrEG7RVvs/fEdSKmLcHjf2Q1Sv8UgGB09rt
6pPyP6viJMO45SrVYEQj0VL1H/6VOOPg4dDYLGGaxdeb44/KLUPmVxrPtU9g6pw+
EpbVs0+UPf8UjeIL1ucUhxlkoiAbWm0p5CBRUcUlmOjTMAUifdZcoqPxtz6y//02
afh3lnB3XJkOp0qNTxgiDDG33J6doqqmPdxSE4h+OHSjImo4hP9PdJWlZPmZLLqo
rmgX6JNS+e4DKJ0U4eSr1abKL57EGrA+PwH5P+qV9FfjroOYbYkoXqsJ8oOsjCJF
QhaXW8RjqKb8Bqi3pn0gtpPfwaQleIDLV5x3/20JQXY8ycsmu22LVKw85z1v5hLB
JlARVysJQdTo9TodlEcsarUFH/NGtTA/v52JJhE4AxlPB3pL9yEF7TbVDLNFZBjf
zFVoB6X4J6s5+M2MH6OybMCHA3Zqog9djY/K5pLFpJ+EmUlUpr0kX8jqovrOT2nS
wC/l3qoxy3aj6lzq8yvLOVevPPVXK4eeezkif1k9pBLPcQpvtpjJNebV7DJE0iBG
JWYVWYFIKhoApgS0uWPp4PhsPkgYKUkyJ80IcPIJGzU6tACbnrEUBEE4GYp0klTB
bKkM7pPbSbOZso57zGgE7TUFLbw2ZZXUOkeKOoYBIr+vuGQU/V4cm/ePOQ8fBgYn
5syYFY1DQkjIaw4ABNFMC5fY+aw24JA3PSzbxNTiIgKIKiVH2XUJGUS90LH5CQOq
bGPi7WD+ZnL98UXnXamYgQHjH+j6LMp8ak4UcgkWVBkHyg+6LeBifUI79hkRPET2
iusA1GZl6mATP5+shQD9lWSNBATO7afe4F+by3O6lS4lKpXutytLMi0WHROiczZD
cdE9Q0Pbwkood8VxSF/dgNt5/akRDFpXgP8/u0WO44kobIt2t0tLhCwYTbyHPiA3
CvjKE2kD8mNqQkn4CEHw6WdS1gAgpMINpH+KYXhBLYXy6uFXk6tl5Ea0R0XbGKIK
oxpa6j3OvrU8yklJyD7TDF5cVAPbL9STbY5U/lDss9bNG/OZ3Rb7zrSHb1F+gSsb
G2OBmnrDXY2Jde20//3lgQ1F85u/DcDFHW4HkeyLNBFmaCfWn4MXhgd+lHoL6Md2
OfvFwqJevdMP38OqvwI18yWIdtk8FZpekEUCNA3bZJ+k8O1+Ym3Pv8fnlkhhIr/B
k6N6u1/2hq8woS9m3TjwnQBX6NI1yaeMJxJ7a3yGQqaO2TEzqSh47je5DXxYZBCr
U5furaIMU2cLoPygDFGQoIrXA60pMiJc0DwR1n6Gisw8TBGofEvK6ifJ8pj6EtL3
/G7TxvLcfTRkCyFQJX2A3HAIeGaLVttofd7cgtvArWBRbaYeKPDXC8u2x6afdOBN
/Uggsz0LCHtwwnhLqymTBOwMaWcj3cbMWtzr6OnKX2n1up1IW6HeMnXCwGrfM7rm
RFn2mFpCbBcwgz8XNXtiS+HPiPzOQSZ5c8LyOIXyXJwr0i5flRFc85AgbCxBnsz9
vF3tA91D73zuta7gGMSmXId9yg5OdL0cHWXDmANnZznV6eN18Fexxr6MRYeVB5Y3
AWBKlEPF5HCtnPRf4zjHCzpzdamzLqHGbhQxzeKpBIhqjv2VluMOBBlg6BxgxHWB
hILQMnm8zVcehzpkIKeUPvPuCOekUrl8rfl4KCJ+FB8BjahIvtdXLQics/o7NLP1
ixtAoymNSL8OkwVrNR/k2t4SALrgBiyBpB+8sIeU5xJ8/pJZcJv2JLubvLJISFay
uu/HYC7OupHyZHc9V4OE3cVao+iXqclGFjBfWP6iju8W5cybjLEcdGGdp4KLPppw
A1PUmdDTirGEUlJaC9BYKbHo0Hkvvx2eUllrIUs5oEYJJn6UrvN1XQeAtU5eLcyz
rgFTY8TzovDqy0wkf8lsJqEIYQuqbTiP5uEEh6jsIgQr4G9jSPglGd1nsixigDH0
VS9YrB/ecegB9EZWNVqLYL6GUlsyzh2HdHe19v8m3b3GIINFJylEUcGgHJT78PDy
DBUVmZkct7LVf0YJnJp/82fjbI4XZx2U6fDsbfipZEDQxyEi24/9timaYhm8pnuu
Z27nsCRrr2enGDJltylhiCjhYp7bnSW6quSNiOrgWiYnp76MgbbTFFim1zg13j3+
iQG8jmNGr+s11CknNbONz31jyV8OBNQLasF36vtzejjLIAUlAOEKBq/Qvn3uUvil
tnjHAqkrNLCUDIXsYFP3rQGbLM1EIIctO44DXLinktA7/WEZvXlfl9hfS7vl4RhN
QB6KDsSIXp2uTb9K0XpyT1lQPi/haiUaycpS0mGDglh2ZxVoufWE1Ldxc8WsSikk
nm+sG4iRtUauRNqCMd2qEXB6ewMsik9nNrztDIT/HBoHIsy4qrDXRPXjo0P00Elh
Oi0mu0d3dOjyfY3br/80cvSFCulInv3xiTEcct8rObWpY75orm/wVJd1n3tL7BKe
OmsjtCvKpWf71oGaY3dovm4cQUOaa6G/9xoQxQ230uXVE6wUfWi9EeHrHTOTy8ip
c1dhrQ1ER0E/sGq/+Wfi17V8Qr4LOywApzgg2NEZymzWVxqG3iRvNKILUzzmu33J
dXq7+pbbBKbvks9W/IQoXJe9184ySBuICVHM8/Il0fg6SaIBOqBzNoS8uSWn/RVm
tiWVr6qR6BebodJ4elg4uOnIOcsSqWNz7UOpsc05NpvuyqwNNnD6gi2HrQGNp5pJ
rXxiAeyNJl+u0Z2mOB2YfPQFKDy54t4HIokoQ4LBy0BHtLXPSBtKYKmO5Uv+LI68
ryu6xwf3ccjEdfMKMzIyXu1vazQA3g4VvTPsjK53vWxmfrfoIpjNWto2RHB210QL
geUrQ0JDQqlpN9mVf7kqXdxrKnbBYW+OWKhc9XMd0gC35t/xXEAwZ0Kyj8MZJrq8
JdkvR7VwYByWqQyhIrT+K4F4QEK6Dl0q/Q1cgwgMsDH3wRgrb8TITv7b+jY0kLy7
LHYT+RBHmtAPWZgD8Ja9eozA09snx/z7qZbxwdgs++6VFAQQZnplgtw0stwzfzDZ
ANpQqX3h+pAlLpoSR3cKvNXDBkpIcn3dUtNXTLtd/S8qnuSxpA7EsKCpT9aWzYjE
fcNIyhzdBc88JI3wjPiMWiDczdW3OAiT/4j4BsWDISc4IRiUdo+GH5YXVSaOAjFD
OddomCWuTt7M0ovfOtNzVWBz7PgB40Q5k9los5ogiUlg15XQhQk6rmvhpUe99tcJ
3e76V9WghH3eDtAwLn0G74mi/WeJ9hcp7JOZN6JnJ/m+edfuQNJcxdLYMg2RaXUh
Y/3MRjl62VofiM9yQ0lYvsgSPS78yFqz8TCIHtPLROkh0Wn/D58FLVhCq8MdKWYx
LHEQOVeglBOdNmMuWjQwiwIiw89NXJORVk98qZkNjVVrUzlmsZ+aeEnz7+Eg1f7C
qsXQl1CIH1/es5UYWrk+WRue8gMYAHr7rzLoRtDHknyACzfNJaSyvdog5s64pt/l
5pbLUlgzrqVpbXY37gEnng==
`pragma protect end_protected
