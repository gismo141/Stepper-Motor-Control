// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
be0B7Y0Vah9xrsV1maslARDesjebWhak+z1eGnx7TzHyUu5riBWtNuSN0Bre0CHy
xgcraIx0thobYlCAdialJ5NnwEYj5tLeLke1OqH+2gsbCB27uIoa9rulkw6j7uNB
tUgwEoRjyTnMwgrCzgARH6GUkiP5K5W3CYOC/0Bk0J4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 131808)
lWeAMXRUg9369UbASMcO2k1fzk5FeQilvYBlNsQdXJ5ao8b8QRAWPArdwkMi9/Yo
/oBhuU1bMbN5YXAhPiWw5Iz/CGyKLXBUiIyTuO/MQ4csvMzzzhCMfQJOKbI+Lc1R
J20TqfuaOGlGzlV575DoIJjIFjrmyH/kp55azNekuTn3g4IQrIsNWUhgZvnmi4s8
qfk1yO44uV2IC5YrlHmIN/yw9BnCE5Nhua3y2KZhL9lCfAOjPpERCakY/ai3Ljlr
gITxGGB09LpFlPn4Ydp0ZSbcDr2+9gjLKFwGlwta4CRSc8iQCgSfksq/gVioTiy1
ewkaOQPzgZ/Rfnz3cRDme74bV+Zz6kMTAeKWePcBXOruwB6ZsFcwu/S0UZQsuiR2
gihWoGo6kVG62La3qgbC+u73hf8mXdtsUaiK6ThRZSV8GM6Rakg+uxwE5ufkkhaz
KoOveD1KJWL+9S7icQuYXHGtvrpfZi5iQI7KajSMaXAbqwVohvSeYosZ5ZnnkYmP
tDgpMZ3IOBbwLQb09iUFYzWkDElOpAq8a53C4dU8qyJedVdDppC+JRuugKYggSaW
cTdCeC9Z11mKcO1SoqYULb6+domzT/JGNXPuy1WBx1LV76GK72CC5jz1O2u+usxe
G5EBZwgEMnYGD4hdQUD8DavchEJXyRgEsr6anrIoRx7/Kn7Rrwv86vEOvlNvOGU3
UUJa82F0u4d/xuIQRUqpl6NHsWs/LP2k8AVM24CZO3BS4uYvtCnwWMtBYImethXI
taaUidscPPFb74QPTFhVw3s/9m+rXJ6UjgaLD8Xo3QXgcefiJHkcACxiRUliCJbH
QClkGIUdyM6Z5Yu5n7/1cxUJTQef71e39BDd/NFwZMD1Modff5WsR2qsp6pXhwe3
CCTY0Ymvqa1V/tmCfssgexPveQTs8PdguUPSavn35dSQdM5Cm4kzMLDTV5oQVidR
tATRbRYYt+zqJLaF1mEo7GevufRoJ97UTCvLwP8Kt5PAwPQK/ipoQsf7Roe27qZu
3L7h0ZGdfHPcwH9KylEQfwfmkPi8unAGDE652cZqNIRv5IpADtNuVxjRPqlzZF7H
YqYkRTCWI1wjS/oLhPmUKzocGF1GyI9V4K0UeNw1UOGFrwsQHeTc6b7vVxK/pyU5
ZlCj1mE40nwrchpgESyYmTTk40MmeUwdDOmjlM5QAsCrp/hVm99gDdyARTYda0H0
8f+MKYPVtpGLtDVjS3iue3J9Mfxsk0B8HggcNdIziRsXxKtDYwqFhceBrfW8+/f1
1tjdjwfrSyCaZ4DV5DmzTdfxu9Gi/8flCM9Jxmwn5x5qzPzua3WzqDZFNSkt/oH0
ygdS3Kx1YQrggZGSfyKffpZOhnRQBERxZ2Sk64JqfHvGsKbbSndk6yLtdsdvR1Kz
bGuDKro7JpWtBaX8TgOYa+FQhdCyQnrKwmCqcq+xFQNvLi4vB6GRcHfalW2/xX6T
blmFk+LCK7fVjzkzwBt1gGBm13wJmyrE8fr737xEIY/wkfJVO90T/yZ6KfulnqDK
KM6IL1q58bSK4D3YIeum3J3vCQdV7lnwgvEEq20vdWBAlCqMbXmsg5mBw6xCEx/5
QfRgI6IQ0HKxdPo791rz7dRJCG7uUOcYp8DtFtclBp9ohd+P1GvUG5VdWxnIoCuq
Lw1M9hWHkRZKqVjioxIQjgH8VlLSm9RJiM8qN/cCb5G5SWOo1qxx3kSF1SCJ4+r7
pfIF9ZakDo9jFRUVfQfZD69Yqtmx6wyCnidxcZhZqRwK+GHpjrIKU3pFlFwppZH+
LhWd49IXxrWqWxlXGPJpvcld+K9hLNXH7I6Pyu6AudzkdE65ZjNXFVgIW3bNoylG
N8kEXeVrfG1QaCC58GEDzPTaCmcwYpz6sNztytCO+wdMiYK7Y5zOTK2IFTa+IwW0
Lwld256DRMJTL0yP8ojAG6F/zHlloGsC2TsFWZ6McfQaRj3fCNUcPLk2ZHQ/IKHR
yn1XYE+/l1ftTuywycCRNv34zsoh01wy4M3LEFUYXWxcxuqoLIk4Yf75ydQAOtBd
3Tz8WRZfh8hxhYXIoeeChWZlqNXBTAvF8f+RFOavcJrMBmqVIYfJFo1J7XcV4/jr
D1dEa1pmhon319c8ROxIEzI+mmKOh2CMtmukl+jEzyU6h4qUNscDRl5WkcVssB6+
OhAV4bLGfsna0Rir/N7/n4GQcQurToIFkRx0jHxSSd98gjVdrb9XgEFo3yFRWfGv
e+Wv0gbfD3zAV3nvXs2i8Rd9ONkldjVd7hBZ8/2rJ9H8seUK+uPurUPJlIoKuBcq
9QH+Kw079SJAEArI9IhR7GzwicbMJrKWm0VbJy0lUhVxWlwx8/JvyeHz6iszHUMO
p0eWgjz/PyBkFu/Yu96+PQF0XT2wvo1Qsj1Sdx7+J0ByZEllkywqPQgDeDeu2owt
OuZ3CBRC5pHauZcQuyVwtIcW9uh7Cjg9vDnVuI29zgW9LbMH/6aclCef69f9Pr3g
+AuPvqKDXI6YKQ9JnTykjvPmjRoVZ+U4MmBHNDtLj49IRpuK4CofjlAhSre0Bq/l
XCJU6mUvf6JC6okFunSBHNFfmJIAlhJaMeM30PuXgsPHgooRgooX3JibN/cuA3a1
HtSW9CExaSWwsB7VLfeE+j58HCWoNcf5xhhoOeO5ue0os/vI4mMjgWT+r4LeDCLv
LkRIoPU8sNGHblE4PyzSBEp731KIYF/bLXGIOMwQrUpi1hU4la9jzIyQm/v86S6N
4KouTrCt3rH3qwJ6AxqUfqYiHQhExlJFmm7xVfbkB8nCxohsAfZmFi8tVnIZuzvX
gw0mLbkZmom5tENFqhU43h8DZxWSptxw71SrvAlHmV3jPYJkQB2HV5YwQsTF8hVm
BGwd7IohJ+RSo3/WHY93GgaARMlv1RMo5kGNMl4dQpxFnhIsTkroXMDhWJK+nw10
+K592ocCpUEGloCF9Noas5OtNQxuMlnMareM4X29qdqJuotzHpuIFvd21iDtYVaF
T+85h/xXRw+f/qCgeSI/AbDPkUdJVq/+a7s6Fqj0XVnPTbKG3Di91DZ5PiXAPQGF
JEMWhGsTTfBZtqHKgYm+h4Q2EClcQHevjgR2323qNrqGKjxaljAkF12MnqF5xWNL
eI0pkKW6lH7aPg0at9MMI2IF+0O8GCzfGETzIhAOmGDAnVDzB7IAvIwIum8u8oDy
HWcLY8f4ak4xa+vmlMdBAKfTVXsi3rm1coIn1MyQAEBVk+vjuPnOVvnB9NKbOjUH
F3tT2IulLw6U6AlatBtNgknWlNDOX6wS3TCU/GVl27lSbKcyUHLiVjaGAGkq02sw
pP3fdUFBYV/iSjiGYfFuepRACVmH0iBfAJJaE0fFhdUYim82M1LXJhJzSom26mMN
Zig7zXVdx7LLy4SgEzRQ522gQKRlj17IAGsfTBOtPx3qVoERsMIiVhobDNEqWtLR
HOZNztAa3MAw8FHqKexr+Y1X6N14bTNgDAezGqcAf1EGuU1YhQVjBtBwlpAXqkKi
WPjqD40Rtd30sNILZ6/KmfqvqNCNmkarxDkA9E1Vqw96sC00E3wNT+dJOe/lgLvm
amE6a2sKjLKALl1Xihi55kZMfv1WuD9uc/QFKCHugLOv4mNNWR8Ul4bVRZrB47Tf
9/nxacYA3+a8UknA5AFCMefVNdeXOM2fMmeOphpdxdZdJ2Sl8UzpRE3agomi6ZC+
0uxqpF9gkFRPABRuRoMYlBKq5FraSAbeqO3jzuVzyIUzhWHxcphpTdLk+v4+HH34
0+hWaQ0reasNFgWtR+PtDPafWwRXivMaH+gd4cko6NgUjTzMB4cuNutXyDZns57X
iHS0BgfastqQGETL0HwEZ/X/eI6D9ltPpeM6z47L613YoQi2jQsVHKxydPjzdMSt
xuXtzwlwB7Q8hVojuwHLVmB7t9NiKZiIJVupAcCAM4ZQQ8qXgPDfBsV5uvrOAXRW
nNmeNuGnP6Cj7bVvY+4IA7qcIohG1eO2XWKyeQnOcj+nMdE5RTyRaB51rwU9EZkF
BM6iW30BOWlGW81qSMz6JWPzZHYsGH474qK7QCwS7jxudMgzbqz8wuYXlGKH4xxh
GFMSkYKljEDmmiXHQzi6dfhFgQtBK4hJPVr4d2Hd++iWkaQ2i1qXDm7qbYQWcHwr
VGGRbpzBK5Lk2c+Pe1CNnmqFnE7cFJIX1t9Ipdk43QbRv2dRe54kUa5LLJnCu8CI
zej8u2m3Tnv/4mCdHOHOsOwrx6X33e8SLWao/Qo7JdxOz5fsoo+czriwYwbkVxnb
PMXafQsqn+IZCtXJGQ/h2Cj3lalvJlEF1FWnFKQMqep1QvhrPG+3yae0gdta6i60
zFol0xOidPknPUA4wu8p/aC/p4fwq5eFCl7nYVHhnjZEll43vXtgctR1N9WAcMmW
fAcXn+fjItDjyPozG/qAxNgYAlTl2hNP8QCqqjiAhEDGgodcjl9GvWj0jnVvWFoC
NtF4Q0ikImKBVdM8+sk++Ls9YrpHSESEYzTO7Ti9mlePk5SWW8be2oDP80F/JD38
i0pMYT0pursg091jGdSo02UvhwI/8c1vALwvO3TX7KOFkOBu7CvPU+d1j81GstZ6
kG5l77wNvHgNrn61QmERkjWE5pUS8+pAXGz24nMIChj60sg8Z7cTwkfyrdp5DbaU
zoPwzwrWOugllqzFM2wvVAx0xMn1nTICUHeGrVgttMMtKXVlht6ZT5p3s4I5TQec
uPLwDePPnZym7MxjCap8up3YVpLEAOVrMt/n3DZQ0lA0x6KpcePUpSUu3KqCR3XR
TI8od+olSFmzh4fN45wFScb2/cvwWxzhVS9WfVvzCEi+vSTApadXXMwzOwVMilQL
yu7H3hgf3OMCj/yOGyDsuMVYXgdls7p4KHnotMnsY+ZxvK/rcR1UQ07GWyoy3hLh
NclHvwxBJasYEcfDBr0wha+QPILX45LbNGUZpsbJ0yPYp9SKQFtTPNUsd9Ib5pbr
vKKWEHkaTXSf33Q08XysI6IEJI0Eil4FicEJiBI5xmxWQrIqB1lhNzds+eKWZtqK
1q+/VY+9b9IdcPI56DNVjmRxGIVPgN1xdegnx6kEXGrrRPw7N9XcwpFTzKSFnMgF
1J1Rhjw7OOtq7cbiRabeQWXJtW9Qve9EKStbWxBEuL7qB9rUTcX5YIIfxxxPDIiP
b7IwHyrHaO0dX4q7MyRH8rPIKlw4SVLn2lGqWahADCTzOlMpV0czZ6GnLSHgqW9p
nrIBx6jSMnlS0TU8JymfGWrixznZBR2MoNpRQn8PrHURoC+vDx2DhS87rIhC3p9e
gTerPRfqqFyREw2VYO0jwftpVkxvlcCZBvKy6f/T3sDZ47tiPFx9M0Tf/vpdhZm6
2xCUXhe8LhbfQUZLse5KXqa6Df47aYXhUhXu8Xl1LC4MTqDBJ2PvQAYlVZRpm+6Y
q+AAbmcb9Q4aMqN6vNItLUhA2ichvEOyWxAOjrrLUkCfD506hwqbhYM5B6YPZaWk
hydjk2AxqxR6lNK/qy26lr2qECUtGXqD7Wtu/DqfukukK900O/ZPtF8D440mI89Q
waNFanEvyXMQNqNYXB5el/c/VqxmGws/th5Q88MDdqw9c4sRZxiJiHg/7jP51XBF
c06Hw2XB5uUb3rQptf+jZ4A/L86baS4qgHrpeFjxPTwOcWq4LIV9XHy9wQWyJvLf
G7T/G+yLhOKmCBJa8hY+DsHwADk8UHyXAlPz2pq8Tcpo/rV/97GlKmoJjk7hFoXB
3ib+8irCNw2elQo4rG4jRpG7p/64YPh+c7tVwdC0Aup+qDabpCKeay4XGdIXF3Bx
9uhgGN3IIF9+hejvsv9Kyd0wnw3DKff4c3Y8z8pgggLSdjbWmG1EUEyNTfBNW/MZ
kQui8SJm39sACLQxdoa8dVXz4r18WyMHwC3I3b/kwhRv/yxvfrmSmimrv8xfAZ5x
FVlGGRCJpkoX+Fik6o/oXnQas3mdKxeQhN49dlt4Fl4XXHR8Sp2qXw+4M4t1Tp/4
xbD+XqDDTVgPmMDoM2+dSbXAig4WOSlqBL+z0wtgs4jneMQU5hIt2KQJPdH9LGBA
odurUver1trboLW0QCmZNS36G+MLAyUlO3qYJ/+YaQ8ek/qvgBjZ0YpBKHPSCYgf
oXHX76FVF4qj1Wn1JUXk01Q4WR7Lp5NyVsNzkpIz0yaOlSX3vIJl+g8lcL7Whiic
TumU4t5UaHhatQXkfWEadpNoJVvNWL+jgk/RKmzT8JRojS1NBk2yfKh3pbQQG+iG
UvtRyHSGHozg+qK0AQzu/KW9atgFELX1SDIM+sunfhwgh1C7B+FFb8W8j0Ec2iMa
xhe+zV01joQSo1m4EffoWDuX62dm25ixt/gUTrpuVQBdMGlLEO+OYyZqqM6DKQhq
1AVnPXMNwHpqIey/hcEFQ1JIwVZGumzI+Ex86L6tbt9EMeV1fkNbEuu650YYpVnh
2HrZmecXiOHB2zPIbAGYQbOkKxtMRLv9fYvrrlrCmsN00TlFO3koVHGJOIUqLqd+
VtI1uqgxKJst1iwJHFOv11kEPxFQb+SX0ahUFegtVGG1a0w4U0m7fvFV+ve1gBKL
f0HnUNpVQpPy4gsK8Ct3+I2aVNK0v8V4IyREEudZP5wpLkmVAsVKo5ZbJDG3cVJ7
tjlhz6UoMxpPXE2SFmrV03mhOwScxhQgmuldwd5+HS1NgZkXzGi7AITcMZxbsFtY
4Y8bRe+Yim/M/LzUomPA3hv8xnIpNLW1N32bFmfTXLkq1K6F/zo6zrjtqwafrLVT
IDcIPBG2x8nMy2uqFJRpdjhBgDNgHMbRM5I20q9ZzWeD8ee0hr1WK7kkpIBPhp0/
OyB3lpHrR5UyfF4PuJ7kUTOTmxUzhEj5+GZfbv9NyRJ8E1TZzIBNY4N7a9t/G29a
f2h7MWQTflMkSROKFHzbxZXF3tMj1pLHFNb5R7SKyp2dwiFdeNhn7/pDuraITM5K
G+VuJoJ4O4iWk3RgcmFPtizrgYOZAJP+sgQzxjqEgsMrp5+qzFnetvct5jk+ZdbC
yIievCazJoQ79aGWi68NZbJEmyCDztmHt2UfVTZsAcU0ecGqPDlUrlT+lJNgKAhr
sy0aROZszR3+C1dkR9zBYLsV2MoYxq7Xe98FF9qUNFsLGobZ1DWZLjQr60fPh/br
Yhr0HmgbJgtf3/xbU2e4DSGS9UUMQRJpdRDfqLCKH4SvbnaaB21ykaGKNG+anbTT
eFJ+FOhd1ziPGv92WRU2u0QmasNgPxpNcV+wZEjy/GjIbniiY2g5VhHCz9YKKq6t
bHfh8eIPmNaD5yptUh0emb0FAhpN0n/4AaMZOi8u7f5T9vuL12o51m1QXiGa2PEa
B1o7zqE1ijsIInwJ2WsvnFO0hj6IQpCJRmBWsWaTMBaAYvRSM8plumVVksklcDZq
jeJmqfKCMZersDZ+g41Ivxtrvfra4R8+YFfR/0ejsgSesw2O0hbXfOMcaihF34JS
4SPwHK4cgvTFe7PYpaKgWcLq8ABGsGAGAlA1glRlyTHpBWdjItjr/pApb8BgesL+
fRzlevTx+bS5UkBax7p2xiwofBdOww7SVvonoB4S5FVsFznHd6VUxGu01UhfPTQX
/vOREbT33PyMGHi8zJkMRnAi6AmeXOhXNvSCnuZTXPdI1c89Yt9KaWe0saZJI5H0
q88+YCVs6VHObiLKFlO1InVjlt6LClNs56+UNQoAJA+6UIrPwKDrgiMhk94Phui5
mihMwewlDXDk7b8YKoYZENpwsQ1WGP+ANn/QI2LVAwS4k/v2AoZkf6/K0RdbVAbR
GIS8ZyytJlRZNh1kjo1xe9tgvYmKwiZaqNEegqzCiIEj6Aj7NOIRQRbXSiF7+j1P
Tj01RyO+fFdsYUnAXQTXrXFZFFEJdIY1qV1b3TioMDft/RXMWJGKH700agt2HKng
bFjENhIRNlzelKcwI1hmn0V57wsJ4WmiDwobZPHffw1/svz4kJNAXBlfE4cFDsrU
depULoLfsjMWOrvca9au6iU+NFYrUC0R5n7eo78sbZX8ZKSKyR89dMIVwe4ysZBq
WljZ1+f83Lu6bFouuDPdiKoMB2/SNck6DeQ31DDkI1uKyP01CXccQ0u3YRvwYMb7
I9dBCsIrwgGMCKNGBsk8tOiiZZ7j+gw61Zmz8NYcTjNUprsfv1TdUWCCw7nd32ev
3yqmLSmSgHrDVlUwXc+of7WjQtQPRp+ertSPUaqmT8RKVsVEnH6pMFBeRKfaWFRy
BZ6r/+rlthC4mY7jDQjTXwGxWX2rVip4kEzJt8XgFooYhS/LAH7mrTUKnsOcXaHx
LmKS3j4O6TkKbVkSfJ40U0KMuvmTwd42+15RTpydqsegObBoWZ42tsLjWG+OrzAm
Qc9IvagSytJZ0Iv1Sj3yM+n47ALQoqXk5y7s7Z8GOe1PxlURL1UC8jUmTZSsPd6h
GzFtrU/yDE5SD4rZCRxqIjjvQKkcIpQPqNBb1o9LfXrSuD4G/x8EYHapN6dw1K3q
2ivFOHfbC44102td62udLroC0D2WrfCt3zLmEj3zO1qyge549N4mo/TZIFr+bc5t
AAATgoRRhgb2WettkuoLRi0R55EVZQUlibM2lARgXHT2iM7T6jLG3LgTJGyQNMCU
oLrz6g5SyeSsDt4+P/Q+ug+pnrEdcHpNvrBBmjIDe0ofIBH31AEbj9jOUwYz6ORW
ApHGtRCJ3km1cltu5+O0cp1HMZpiWah2fDPqhpeeWELBCGlhgkR2xTPEBwEWqfIo
3o8+aiP0wHFGvxDoiEkPAtA0BXGPx6V7cgL1yysFWaBWKSLKuH1utRzZhNRM7dpl
QUMScnGUlp4g9A6ta7DCvpMN0usZimP/g2KXSvKOa9EMy6QaOARDMe+DIJHAjsYz
pK7cIiPlI0OG7S+aJdTLQwGpcp1KooFjVO2vu83tfjO4MosxUk4JsSdWGuJ8fDhk
j8plXf+Ad7VEasXxG2mHfoijG485zy/nUIbupIzhk2hafQzLQcKUBsYEuY79A05y
0Q1eJbBNJd0sCntqldRAlAH4/CxoYOxcprrWCf+LJvKSCANoEJTKlty6P1uqO8hh
DgeZaqKDQWuIjZgr66XRp4SWyYCMOWiw8wapCeAzKgM6dg1GfgGMsCecZhNW4cSc
V/XIsdJfe0J40+JGK8lw/1iSxHDLf+TGkb1PftxRtD+2yXEawjdXeyo5wKMfSFBl
PBMENueJ7XozYwNjfMjkR2iocZmQ5m4KoygAjds6rhgwuqWHuSUV9dwvQvv+y6Pa
6jEB86kCE7tsx86S8FYVUt7t2DX0uSghGhRHMqEJYUTvCWEhmk1QKGJ/v999qAHR
lfwLihCmXsE1eMGrTAT+nvXOBr6to6koLfuvHbjVVKUn1QceKk+pyhiek/lIwNPM
fEB+CiFggFdfW7wHNIpQ+61MWLYIDMa0+pI74V5md5lONB9EY9GRgPFAKa8uMwJM
bGakz/4Gp9Z8rSM0GM+0wCqRAQ7j1gcXzBmwvYqAq0OkrKwCgIPxzQvfwsqFOqwY
O8dB4HWok4emZInVP7lbmYyo2IAcJZ79BQ06derm1LJWBUAqOv8hCcdtH1do8tvR
PJOHwCMfj95HQ/kjgJlm/2zLOJMCpSNu63YseTWLvwSI838vbYG8q0KxxnkByh+K
0ClPiRU8iWO1GQT8LHYSHSoWJOKafOiQlHALeTQ2JmP4qnWL0mxXX+vhOtAv2FPf
AQRGD+YOlysmzXFsnuOTCLqxPmQUKaxsfpkfGSJ+7Ln8StfFdh6qOS/vUjaU0dSY
7diMNI7hsBazyv2Zd1PgUgccP5YvGtu8Y0jJeIyymAC7Tijpfkswsrn6lOZ1Ubgj
g2MGDh6cIND4XMqPzN7UH2Q2Q9ON9H6MA8t/X5JwdfA61KNLmi5RaoYmorgMhUXN
5tHC1lidVZLJ9UBNk2vXTLvGQlAsJtqmmzEo/RrsNMDNRthCkM+t8weauDqf4gin
k3QXhfB24mY3KTiTxWWmuXpHSvlQl7645Ptfs48kcnIk8IBhjo6mP+Fdnh5CPCDg
ERQHNqx32j8YasZojloKhmYiBo+uedrCk58d0+GSN+ZYw3eggDfhCAke0dmRr7Bb
zCzZqAT/Wv+MFuSvBqKQJsFqstL0Yflns76TvlmK4vzSL7QSTrPoFGd7vBH8bih5
dA7Nh58OtTbLZovFB6r19937GsIAqeCb6iiYiuVE8wZ+29zLEi1Ql5EH4dwXGnid
wMTuPp3whpN2PJ63y+MarHUBk+7EFPPD+mTxKx/+WeWdFyzo3nL4Rt0N7a/USjer
lMF5ZQk5UT+uZowAmFl156Q9iWcV1vWzywIlXfFvIpw/uYhIc268A93I8N1BZx8Q
AJ4zOUsb4JXzlzU/+T5m16luEQojRxOtqYG6cmbrnHWGCQy0PeD575h4mVyzRq0e
FpamUK1uXjKUMxNDD0WB7kJIVsJrlcqAboz163E60M8l2iJaZ+s3Yn6ISMfpEcs/
GF6Kf7pFFDansEXhArtvVl4cEc5aXNwfn5oLwrfg2ZJ7Z0Zn9A7BTJ5yVRvk6zP+
aPTtoHEOBwqU4DKdJwEmoZQwm5mS2391UL/E3DDwi19qTWyVsbhp7I5C++WZ+v4E
GxNsjhE7QzElPkJKj2GbdPgSbilzSHRlq911dNcPKocUIwqUxYazpSB7saogsMIe
pmcNxT2j112p7EcQNKMHk3NOLZAT2Afomd7K8ch+voHRBDW2Tvj02sYY4NnMyJfF
/KB0LV+RHQhUWhM8mzVgc3E1A+JEQ9CWZq6N9nTYfF4Lbi2XJaOHIqqWDEVwH2gR
YlI4zuehEKIp9xQH5jZZhBwqT8CMQaX6WpyXiZpixlm73I8TaEmpepQEGz8XmTxf
K73Mk/RH/BXcTudobRUjnweyVhrUh3UHRhOS/GSCFD3bMxwkf1K/4//KdPBjZrjB
x47houfG5KXDc4Ej1MBWy0c0jvRjZwndoBdd03nPRKjZdoEEbiffmpUHK8PJ7v8V
nHMVtPAz9Wqm+PxoHZgsos+FSvPLb0DZxsNIXyB8TVRIOzl2AKRuHc4EHVlvKiPH
7DBUeiXApSXOTBoCRmRHD/O65fOvJ+8F4jN5e5p0jzsw6hdBvJ+R2ddN0ixeB32B
24u2HdYOcKAB04JEqB5CylIfKX+NHjPibS1AzFYALtwj9Oh0tbpVKDhGz03bHm1Y
aPPB5/R8Um6OoJ+rTza80vOCKqzESvlKglS+7Pg5tYb+qJ9EGokupgHhOCK+BfRB
WsvkBw3QYPtjoX8u4JZRIayyHn60tWaP0Ioc/+nlUW6W2NmQ/3hxymdwmCX+kSHH
/RzbRemMSveKJ6ZdTMQDlJFH93tPqzs8Ru2HaJ8v9zLbWR5bupZSpXbBVdGV5FtX
OvCR1KHiOO6jjk/RW7tTcfO3L4OSv8MUGC+TtKyjJ2UWk+/03yHynlexFQt/btGk
SLtuWwI6NQeGz48z3xKULwxrBwNQ1IZFp7HZYm2Mz0vWgr8h4w/A2tXhPTtyVhez
Ak10rImzD/BrAUkh7+aT+wn+4t7pGp6AuTX+79CPctrc5C+dkB5wxTNxAx0VEqT0
XgI6Dzk/AvHAIwJwqy9Z5s1wvN+AfSNlPrbGL3R+q0hAAnlkqwVqWYLzLElh+Qfp
TneAAI8KmNVofBNQylhSc6kwpe7G0/TXaYTron6aPP++1K3BduOYMcHYUre23gOx
TpRV6EBhJDvLcIQYDzSAnsoaF3WFnRzhiGTCOaB4kgUoSKdFSr1YqyKty8lJ86Ee
sjNWaYccKX/e8Jv/9I4zo6RaUVxB93sxXM/wr75zSam+BcTB6rY4IDbVYwBUO0Kc
bzFX5UmVj6eiZP4+bqSMZ+IElco2poxy5ZyI8EFtLRFVV4Rkp/+nUgLOG4qbsmHY
sFa/TfsyA8ytAwrqNgC5W4tST1zCZWPC/rEB9MFbQ6qhyFLPiYFNljf6EW3CQxcU
h2PSi2tfEhPv4EHcUUNGy8YMr5fbjqIsaQLXo2eE2GAmdFVerjGY5gdwg0yCkfYb
QB5ScmyouxYRUi+o1dCGJYY9SMnWlVNjDaA2HV3ro9r17y6D1Wg4AST4wKcl+xw5
zLxtdk3X6k/lxKn9zW2M2+DirWTKdIYZZoSBW5vEc8/ZJMimLrKxpq68DfznOjUA
0VFJZ6phOAzZrPVzWc7eiVFi6SUx4NMiOZc+/RFzQPTFKCIfDspo3HxLTI4NeUbB
eyfNc03VHjWkPbboW0rqibOMx829AEw4SkLg+MD3LAkSv6hShulx988bvqpfRLAR
jmsBxwx0b/gTWD9otvmYZrpjROyjV1r+r2MV4RBuYSzJ+0Jh5AE5gs6chjOdhO1n
aQYW0+IOo7pqvnjkSJz1OCyrpr0sMPK0kwCmeNnRwvPexl+F8DcYCOt0fUxOW8/a
qlarZhUxWGAIL1n/Tx5Xs84TCaMYtEyQSDZP665+iNWigeWxksUoE5Ofa5DcU7Iv
PljyyFLjWC7mKubfJtBfkRxTWdQZ3xmdpD2qiScMIkeDq/egAtfQNiOAVuW5bC4j
3H5OiIAj3lEXdCuS/XHplaGNK5YSl84qqd4q4PzjYbGlpNHM8uHmdhNmAr/v0EVw
0N6j2wFEjuFwkKeG4+38m9VIo6fN3pUeM8EkcK7v1QdZjLG6FqAoYclz6oWz2aPr
VLZ+KWJb+F446OwzLW2DTRu/AgnszQiuiY5JY0NnJSjAeAnhMmsV2BVZW06UrhdT
b1vU7r8xzb+2tAvDEY0aHpXIp5/2NaGE/F6cu2dj155eQrW5G7QGK5Hwh80H/tKK
fqWgC4by41zJwVwS+2uwJDimeM1NbZMXywqW9zVE4fPhVwXu5Urg/381eI12CgIO
SPOq4zY3nZnxWQTVdwE8QzxLnyxbroP6Hi9RrJGKLtKsZQMLnhTJuLxrF5Nm0afY
yyvpUk2+/dCUrgVyoHMP6o4lhGQF2MUKUR/TMMYHexLSPWIRfCjENpxk3sp9d8ML
bCr16tuUviaAqM5OIRTZuYofVg/mSB2xraiyVEDJ1AEmBKO8p54NmsoFaV3D8uFo
aa9SrvyaBe35u5vFaO0xXrayi3TC2FvPtkxO94xX5V7aX486CZK5S99nwJNYWvvk
4pn41EYQUfoYw2o10g54uYkCb4qYzQ3bOw4gU7SFitl4/PwbFd+DbfwJT44VJHSV
JvuGw72nu2LJgOTMsIjx9lttWarhHFoFhvdKAOcaEQo6heRBBc8+5ukxa7IA7jjq
tyIPKAC16mStc3GPGUm3B5dsWXSeutKiYLB5BBE6jdfy/eM6Xb1HvxFdeSYeEiNF
9vlEwQulGUFQ1cfboe759lUbSs4Lf86dqYhW6f6H2jKz3758Nv4MishK9Ynp4XK4
J1WcabxTojXxHXFqdcS/+Q4aDsp6o6j8RNRljD4FftC+Lk3UdguNNGhZMuMJkvIH
YqK+H0yPjmpUTsRHXSMsrBzdIn2uPzVG8WFdRWgMnVdy0BUyfU6bpX48kUxA4UX9
Rdr0g2YPgw1hh0mu7WCSqCLAgWsGtKVSoNM9v6/VCAEytALBtf36HcB+ukzSgwVl
cQQOWJSXGQEQruUg/49c1UGHDBo/8aOuQ5PefLw+Yh00b9aRUOqwH6SRYEM0uMpd
3z+PJe5/YTw4/bP9kz1lmFHC0bKPW6GIvj2l4MrO9Mo/9PH4/nH8qhmVpDQMdHvS
e01F9VNoFGcUDBw2/HQ0Z8nTVHNXXEAv0bJ9uZ2ca/XItPba00aTKYs0Js5HLJhO
9wa4PX0FEyKBWEljzsXr0cgAQwoBvxiHKf1JCY3IARfnvw5MG9KZqluEGJOo5gI8
lyr81yj9ZzeIn5gXHV0UlasKyhZHd9XV8UjGHAqe57zD9Oi8hJmcm+tb14tFg10M
6g5HqSyDepBvKssl1Ky8zkeRZiG8UrFONkS6CQx1+kNhsvL2/SeorgYWAeoJ8d4Y
Dou8SlBHrxAMdMxfBrGo5xGsN14kEBO4W4BKTYe/v76H6VptVxRmscYTFqp6Zmz7
UvxIT+BXAgD9UX7paB+oNYlzoocl5g/N/V9hjttPonW3bdsIGCvkW7sM2iWgwkyR
tgm1xzu6VvlAQ2ttFMhrvhc3tY3dnupHsG6Pqx0aJ3sP/omIXIn02lTwLIN+4hV6
F/n/Ixjyfckfo8fVTZD5CXMLcHkwFugUkS83DAn8lf+9i3gdxgu0nU63ZbgG/Urh
IAuj5OEqZ65sGAgNJ/mOc9CIMx8hgRLEW7Aa8vhbFKl55ySx5WanFaIyCQbiQqTc
B414ENYLpvaywLHo2FFH4SIE9nzyLTLAe0OJ8dWcV2BftPEn8TAn4ebLQEb3xTnc
03WPFFnf2p953dDAb8HVFmc8NZ9MrOuAfVvUhudnChuo3gcHwP3ci97BuOTWmaGu
m77gnQ9Sp8XDbghxpkdtQv8A4N9ujawIgmM+vNCt6FVLvEfYGFL6mmGWlB9/czq0
nxtUDo5npBDoYpLoCojSzsOnphPB4NZ97mqR12mC01mCW+yPpt6RRSLkh4vMxGZC
S9oHeYYTmkVQlQTzDtDB6yFojKewsKDZzBlWbwfo5ULcgIfA17paARfoG+DJ8Ss/
TwUt2w1fwLs5eelzm2x9AzaCE67Wzh9GJiVWaIclsmnzYKLa6jNIT3MgV9BqSA1M
sre349zwyR/OK49knATykaVYWuuhX6z9yzJVHcDksrSDN8MaYkBTFLJmqVdwUkza
DJ6DKUq3fsJqRRx7A8FKjL/lUCp5zJZYGeNfBvSbcZ8JIjJQ5gpwEUZRuCvnIXB9
KP1Fz9EvmE49SaBUPYszg8JSWhZFKELEbhe+5jA3dDk+e8c52YfXz7dVAPTIYHe1
XHNzlgp8tQrRu234ykwloFz7BI+bgGmhtELI6iBtBq2PVyxcqAIQ/8CKPnEb8NDg
Bh85a1JqM+8Ngb5srI/XpTaUQy6F//XMdAxUdcx3l+oN4+vlwmGUkxDTfzokWVbf
d9BCF225lnngdg/IXpDxiBV5gMTvhcQ1+cGMgsKm/8oZGC9Tuk1nlc7G5RsyumHL
Ku4bxOcHBkjFcI1qoeMX/32UisX7008QYzjPVwTmTNxnhYwWdRd8LeC6zxol7NuO
HVBvWY5P1B1yLdI6VBki4g2XzZB9O70+CwWfxedjA8VtdK+X6WdsHt+FD9oyqIsN
YZ7Y1+/x/5R7N8xf3m5cQxlgwCy+scW2NOQqyag+SRLCHbxmvaP0MkNEFVqhDN7X
ikfCq2PilRPHBd0CzzF5rep/Jc1ZPaILqp3891UAvl9zJKmYHGqmL/TKMUV0XC10
aCYSHkXYWbCufS0BBtGLu6Sf3TQ+uzMX5Kiqqb5eozxY6QXZbhx8YutfpkRn1OhP
D/kh5FYoiDVE6+0eMpLBHAbA1U0Sc67xx8RTs4qQLqxro2RGESJHthtu0fKEUam8
hpb413gk2xRCfuEM9iv/P6AsyRczJ2SLCdMeBsr98PC01udxTFt8cRdCMrItwowR
81krqTDEqE1tdCarZe4EOBRqQqwfLvDWnUqp4tTXLccmUXPeTIc7ZaX4t7b7R+Vn
axGXgsPwPUFuHe6jUhJjhK2p6fHuTPc4IuSAWyS8aio0LMj+F2ykKrP+rXF25RNg
wnWUlkWuEkuHT4OPsTyxdclAqfCfV8m8weh2oBBc90WR4W5OTSAAbRj2bZglJK3R
1uKSeClPd3LX+EoP8kQg+6CU+8HburXGy3IgWdAx8xORl9pJXuE9pK5+QS3v3Vrk
epKkZ2+N2rVQ3q0ITcJoAD6IG93NSCddXDEptSn5O7K8LKNpXTs+UBxd7p0AxWO+
70NB7Nr9Bpy1NFd7y3VRl5LinUsBvH3UWq7HuRg6sQokb2W2qg8CAbW1ZDnzP0rv
YshYH4cg9YYtiB1K7hLmtZwfNBMoyoDJsYDxF0N8h29hwEEOLXloJZJEkF3j0dFi
2Yus4i1tqn8VHyLEQ2ZrB0JusQxiPNM99ut3usbAU37ypFHM7OnIuDh82cPvJpA9
VkM3k4qTAMcZ4s4wQtnBUK0w9gt4HoMTryT6njWYXhKXgVMAjLFRfh4KhMMdadgo
8nY/wBTM8AePkbBXKwrRrj0U63uBfSpLYlLL+uORCQC1+pag0rbuurLLS/CQw3xq
Az9rdvIVAvk3WW5tvAlrZdDNlde/b/8c0XGAb+I6+I590LQIma7hO8oAWjSm+cBZ
rWHOkuXebnti+8gydiLtxMpABxkLT6sTi9WTqv4AO3pERqQguyXPZbxXsk4FcY2t
Qa1k513qEfBNK6775kEy261C8+6zdSKfcyrjNudtLnimn8PiMUQH9AQ/RpbY+MdX
3Z/AY6dafiJQMt6Uu66ywZGGhIeXRcB/Jq/BsQ1/JYH/zPDbpbEfvIaYlBGy70Bd
2vFyooY0XFxxCtMVpTS3hK9X8D3wDEDhe/UOAbEAh33CXbprmdq856/67PeVjqEi
e4+CU0FX9xhJ6l72ywn1AJ6PqadCNfaYbO9Qfdnnm//bvNKuQKWHOkjGv99jD2lw
yfCHjOxPC21Oc+ONsW4p0bMAgpVbiFsyCylygIQp/95OKLMousO15UvomQ59h0YF
QUN5/UoqFjNCQaE9hpENDStNgWFP+aYEviuVyVFoolk0bODwoWVB6MAq8uRZE5YZ
d744m2Y0V+0D/O35Zc/IIjVDvECELcBqXGeW5UEVANm7m4VFBLLsbMJ54jzAEEbK
hlHasAgU4vnhQT6h+LBex7+tMOywCAVUYx7mGOWstvCmJna2PfpFmY36mvDdOARd
9O8ZrQidb/ma2I5U9srvDSA0nvXeht/cy58mF1rAOLWle4pbL0q81A4zRTT578jj
1NSjsHfjqTA7Tag7HqXTGyfZ7V1TpNgqVUosSLj/N3B8kiDiKDinuBKzPXJFZ2mN
YyJbc3AB7ANS0kLpbWYxZoLhWGrHDfvhP47d/YVV+kkWL+hp98jUBgEd8O44mUy0
gAg38DxhForrcdJQHRDrh9zvGoC/hkmvKI3RxfDp6aKJ2rXLtDfzvHa5FkY1a6ZN
g9Ev9NH2QdsEq+bZ0djvIqvRjm4eYzwYpmA8AT9fK/4FYgav9+E7KYpr6H0NRctd
zFmsmaHCIvXSpyUWZctyK37PqwyrysIcNUS0RzL/7USNCCh6sMwbzHCnM1jq1BGc
AbYk1Z8B9wLHP4WWhupplENVpvvOfoaME/8IYuds7U9w40xJ6YYkTYWLIwx5tcy/
vnS2TE3MuexffOvSgyuFLMyXaJlepr+ZPTDY0IQ0b1Alkjongqd6s/yHUjTFPRnz
23A/XDhYgWdomSsCAiQO/sGuh2+SEH8uUFujAJVp8vKaqeDQ4qSsZ4GZ2V5s8SPR
+BqPRAdnocd4xCM3W/FWgkTG4qhtduPfugpKLmE2jZPDtWToThuZgPYJ7O1n1W8p
7Otp37QUm3oPAckthZYIEHVhdbwPytWEX+MQFMP1uevdqYCguRtj7DyUoKOEtEQz
+FjFc7tnPO8LT/QFYx1awRzxHB2i1Hze68hVq8nOXcSMxC/2p66560DqUxOAYyyE
rZpYdsj3mzs1P75eijnaYiVIoBNbgT/pFyx+4uGm4qi5KD1AuOlYwH2zxfOtZRfY
qAducfWWH7es22aULf07L44UA2ro+AGUi0HtSxi0O6sWXSchjnhn1iSg9nw9MQSU
XGA5InW+AW8pvZWq6k+75/4Knn2VNeAhFMjetIZqmq9F6IeBFNIVzSyvEdWM8S0m
kVJqZU6LKj8DAUTHKlO/6r2bas8opunp/imHKafsumbZHeirgzc4GrRMcNsHQ8A/
ANAcgwSGaFw5Tkhl3Def0SnvDg5Ac6A+fwzgPySPFfDJO+nkIPGNqf6gAc7EJii0
Lq2xvBwf2Zx7oYnpjmK+L3D5pjchuSdhOVXZUFmVu6j86gmnvUsXavtgkDdnZNqB
3tqTUJB5VaItq7miiG4F2xx9S4Lq2wOEiR8A1gJqZKb/nc2kmTo1qYRGqlzfIrFU
3jdVGy4J7pdswdEzLs/Dq8vxtR5SOBUgv/k0CL0KTad/NnPLyZ96KZuESwMK5Fli
zzwdNqQHyEk5uDnm5qEo98oaMBG5+rUuFjml05Dj07Ii35NVD3NHE4GlX4Dpdn+0
FIE8WI1hzgapqrLkd52cOsfvUI/8M/9RdTHowXEUaZ5cDkn8hdMaa2QPLWIQGC8C
HPJg5wICMuKz1M6vZC6e80wCHjgE0JbeRunApC6X97bjDfZZpaxAbRqR/KM0d1gg
f+p9FLmekK15MqqOB8UX84lrfbD5T0bDvIW9M731XMROd+CpoIXLIVKB75d1w085
rKQI4KIAdR8sy3uc7Thhg0QP8zWKusN+pPTQvFvLaorbslWQcVKWE5ScaVw1hSZw
k9/3leE/3IhrhN+sUrDOxpnys5T3rjgN+zq+8Mh8UnZ6MT5mxbsbBnpqaQDIW+jD
i53zu0xDp0E4ZIJ2MRwhs6Y2TnxNs6q5xvDogckGX6c4XlDJ4Zt6lyyqzXEheYiF
7bB0Y4Eu3BRNoGINAHVkzeO9Wk6U/7k6ECJg3COflTCOLjMLIo+dYBluAyRrKACn
0TBMzdyIg6M+wsRJhJB+MDApbKcU18vOZpa0qn5+S0E5a8sTnXVCpjkjfWvHT9ju
AKuUIcf+Urvv+zHc75FBkAr4BLWvKIpgWZesFdQSagwtUL/059H0HqIALMWjjcJV
tgHLqTom8NlVxfmaKwQOk45zezCLV/cXuWS8gBkbyXn3QewbGa7CVC9LZLt30WLz
CC3ZWCt5CZgP4csRBWbHtPexMXR94fLQlNIkXsF3xLdtuVmMErpQR1rob/vGGYeB
yow4bDjy5S6LNZU5sSb2I7t/hnvV833g9uvNVrgHx/zPkYeAleXHzCCt0/X2Gqrn
owzm5I4PIqOwwqQlZXF3TttCRM99GlgbKS3agI4nkaGGD8wKXDdksbdB1Mja+Zu/
qMYlml60J/b9cKb3ECOo8kRsaUXblwFMh587aYau+pEtDl6qa3VIb5/ELrHLOSl7
/tEwp3cQT4ws4SNpdlVq1eyxMtsx3UJSFXatdE8l1RwCt3MDpc8TTPR+0BfwsKX1
JrYAlH9F3OpF+DdFHVxHpJJRO7f3ozGNPM4unNdXBQUmxD4CM7b6RjYSSb2IY03Y
A8Eq+Qp2ZWAgz+stk5+S0LLmN151lVXx6YBbQulvYwxuirNAb3FcD9zJ+fwHKpgk
nXqc+1mRk9WhRZdurjMrdqcvm5Ith5hfqclIUjkHlUMAeHdX4Gd6GCdKDFLRVZ1L
AJRKpdtQAOOpulv87OPpscYHSUJ+JjsothzJT8TIvxcw1X8qjgM8yarFHXC8IVLr
FqU6xW0eNwlsYkQ4IBOu7pP0i6TnniaIhmAKrhpZc7i58w6TV248cHif7jkbQRjT
12d6iLcCser5UA8LxcYQwFA0km75l7Rh/GpzCGY7YR2U8aQr7XNpOph1s81bh1gM
qlHVzyIdFL1/ueroUy1pRn6dWvJwnje9/dwJn96HhdPaUQg7wg3S4+JcumEfrgCy
xuAgpFCeZtBi4JBtwCcShGY6qXsCDSuHTTJFW1Yllt/3ZwfId/tv12j8j/7uiW6+
MIBmsgdXCR9f0WbSxRPxvM2/XpMQQYA01uaZaNaEb070J95BRQc+DlAWssAv6UpC
JzEs2Q4+S5ak0UJuX+etdn6XhrFsX0uZ6DjDGJbUtfcx5UvYtP6ziOzKpn4NZNOi
zjULxKVXnMW32eo1XBmD+Kr8YlRjDxmBg3Jec50npmVUq/WrPV66j6bHMQ1ME0Fn
Mi+YZqtuWV+QlffAvumDcYLhz0CptTvEkuMmBMHd6kJKAoYA5ovwsOGczbijvlpF
wNwbhFe0zQHOrsRYi4hPIdTvW9C1Su+aLyBqWi2iRlDWZPsnVxAZCej6JoHW2F3d
m7cHQ2TSCafb9rpp9+nnSarMzfmEPvbFeD+8myoe9CEUChg0NVnjo12SPIIM43qr
uR1JYmoUrHV8py4asTKlFaZpzjXhy9MR2MEE05FGIC3crA+/AqYonstTsYGY/Byh
w1IMBIyfKDq7PaCC3ay/AAO71VxRdEuhw6XTYp836SxdPnbfWXG0ZwOQulEpg02D
PG1mDGM34TgH3TaAtJGx8XmQswgTKzaCLs/3gpHEdQsZd/fGzb019WBKu3i3Dfbl
0yMEooJ3J/MgZ9UL2E2ZiJTSCf6SVDbBnwtM7UU+Gqe5P6XqxmwoEZmhAM8mnd1h
EOucUHNochuP059gDCTznDfBBhqkX7gI/tamds4kKjuN9WEaloUuffu2xMnaWVFC
9mNfqLjLoiiG51XuN13M6terF+mpL3QGwzK84qP8C3mQcpYkWCTT8CLcLIttBmfV
NqsXlH/SDspvYbpR4JKnTaPzrMHbEwpGbd7ZpTmDt7hufUdDFhQAIiQGDurLNjFn
p1HbwVfR0xVXZvT5jlYXalP708qpS5iaLEndwxfaJqIhfeTkUHGvqGSyo5iOz5uB
x/dBju81+WTOZLuKAGTCNk4GfdGDI26RYikRrkYEEQ3jPWX2u8/+ML4Mf1fRBd5l
RSFsOhUXqdkw4INjSWisLC0XCT2twawY77bsfhjHOxJYxPnDYnVEbxrJ1fc6qRQW
eL/xQzlZbhIR9Xn71UFDm1MVlfmEvOHEJPsgIzIVte6opbYhcK7SU07FDIQqIzvO
tkCAt9c+H5ybB54MQ+7Cei/tPIolU/jAk7fWoLvHdlYh+qGDh7NAtGAZAN4/5vCf
5TsrY/J9go+5AnJxcmKy3FEmT340jNb+V5T6tJK3D0Fz82CpG2lwLucfCh63Huma
SfZrMZ4H/ir5r8ZtwpIY8VeIeV3LBG0jcmy/uEQWrvApqVKaukhyhEMvlScVXg8A
IsZPs3kGW35ubGs80HgiiZ9KL+JRGx0X/YWf8J+2UfQ+F86U5g42wiDJr1GP56nX
bjT/a6nAK5hH3cDTFaNvSz4WObZHkNFurq6KR99o//RNsSmjdUSmd5p5nj5ZIVfF
/EyZDJcUGKIs4WOJvjcFiGs3xbH+lAQS2W/DiDY//21u4j3CqknGDP6IZf4xAn5i
Q8O08v2G8z8h/CAHmt/FZoJFjpXhP4FrKFuDhVV6KS4+U/uKUBiRzu1Jg/awIUMh
UPN48WLtEht/5c4E7SUD0sI+BhZzZ2+oBTUrfLTduoqGXXECQLM9pNzqC7Ols+Re
w9lc5A3Q3b7gDreF3TzDA5anjj5bGDnjbOy1k+u+B64Iyp7VhCCku8k4JcwAqXcs
f1ioIOZ5xt6+aNomNhuriH3/IK7AgPU4Qlnibjtau9friy27dBk49aJ4YMGsTVKP
UpsZyVuo24+xW5e5rzfpboztbyx4NHQj5THsAhuswgb85KEi4BBsFSI/5nUDc4dE
GoPUpmmfB8tr0YFcrf16AKj4F3rjPyU8j6l4T1f/ObEm0LjJSGx+QCOFkiC7z2Dv
LElaaV14+NIybFpiiVuTDcCwuAh+jUtpJ5RlBbXsOcF5qFR753NfJ1i+tuCn63wK
KETGqtHid/NjiACEHUoEWzvHuhSSVEPFT3wqDeAb6/tN7ywqFM3xBgAqoY8IzAUc
7qWlHhZc6iam3fAzYPkQhIvSMGiDod58NIAxPy1HyWqhL2gF1c72G03iUcTTrymP
JgT0NxdlU24KXNcK5TzjZrHzbOjpiFgj3cmfWolYBVYS87uA7hBw67F+yvIuYhM9
Qo1BRdMlyLfDvKYug6MwzV6gkwpWhlN/Tjl2MTGkYbf+f45kNHycOuH6yxMZ8lIc
3QC0d39aqQ0nxWubbUss+EqhQl4+BiaUvjnDqWVzV2pnbKxZmLjgTEDIdyDRE4k+
NRtRdekmsET7qsjlK6y+EysFginbwyzVF3EOiN65Vw8H2kY0Ss5QRIcOPJYDapo1
Wr7/9dYRzIqiJMibzSyEuCvx+Wh84xJ2rGKqNKXpH7IAReSIMKhS+dPcnFdyD8jF
anH01a6JW0Th6d/44geA1/0k1VJSOTPmYPj8+aL8zun6L3pRmSVMoAsI2Jifshq8
dqKLCtl7wdUU/aloHd/uImFlAaXBCiOs2/0+FV4uBd0wvulE+L1LTMcIJJGsMPV+
RbR1YJO1mYT+Q6uEODIXk2ZzuMlqZYGgkS85P52qHnVHMvsUPER1C8nlMspn4jsx
4GvUCy5nnEX+8mWugNBDNvu58Jx0r962TJtn5xAnBPVz2xSN9G9CM2hD3mO8YuFC
SCJ26V9RLuMhlk3mNPRtiDeBP5Gi4FU3/tMXQ5hP0xSxFkS7gBWjpvUrrCIbww+Y
Cn3lALFqumyHefg26qVHaOBlVs80MeV9a6xba761D6TjP/N/yfGuxosxWyJD0HZc
5JJWsiIpDRTpe/8dOsSRpxTYIECKECLMtHiiSTEEnUDiKeXbsp1AUV3bmbyR20Jj
382f+gVrJvAiyrt0v3P50aB6fFfy3O6rr/9yOcnAUlQdGa8eJqO11ajixz9mmJHj
Rek1r2VDl1tbZgDRpe0lH8HgJbkaXjtDu7xAZ4esbWLBuRABwhRc/sjyc6Rakrmx
R9QBqmR0pt0KVxZD5De3B/kwyiSkcg6W1M/7eY8hQmPw7C7uAK7Ry31OmuearSYe
o+EJIfYZOMykHUbAT/VPw24tCL0ho/VeOL/QezajqC08PIDbeYTjSmsp5ESg5jYH
TQCRAQgVw2qu3ZZm6kB0MZjZOx+39+iwMwTPYhMY0U8k/OyMM9uBI2OoH82t5FXY
on+hKQo7wsORvNdHEhKNPMC88utTziGoHH51/iImsmm5R1iTkp3yIcVfjUdaCpvJ
1fPVVFt8FyNtaNoU+niT3kfbi0TcSiEbKtWAZPUKgxYi5vgNlqpfFG9AmuZgymdY
xPZfR285wDE5I8XdUJ89l66TxObA5nXjsaO2ohi5XI8VI/kbgnuheYvsMaCFtU9k
XIgAO5SC4KOJO9UY6vCLRXGN3OpkCIpXMWkXXvo9m4IAg1MJNEPgLUL3e/QNtbBL
YR+JHLJXMFCLex6AA9Gj+G/lIXl8s3ipYnXH2foS/s9h04nQ7Jec4krkQAMX9oVg
24nrqLndoa/tsupMkyE+f1B2cKCQ9OCSZ08JFAVd9hWXTK8kMNs/mMEEoPxdRf1r
wkvGQMTDdX00cIot5/MN1/xS5A85uL0bKO34MusGpGqT/Iho/nv4QxCxGgw18KVf
4UJQhni38+knQioBep/YKGpfWBsJDPVz8ilXEiJ0+d2TYXyK8SViuiwYojxzOmGi
kfAN4GoOgF548wBqg2WWDO0oGftDgyGjcsi0gZa4ZuMaT6O2flgzGpyFusbDHGCz
YKmJaMdc9BHm0Nmc0z/tjDZTT3peLZwuKVXZFt/As3yVZuUTzmlKltfNx7s0nX2E
3ELLzZWhEVMSiyvRB2HhUKX38+AESj8lzizjp0xyhpOhJfd+u5fNP19OjVlpi4j0
3AXZeXjY+gF0Sen42epSrhC3htwRZwcPdbjJpfIhsxJB/AcpYZ1q4Qs71nOFtdHH
J5Rceu6OlOAM5darOVWILkdgU3zEfoFt0g360xA++RZtK2kxS+fyuXLcFdWCpIzm
eVzYwTyiCSQFDxcuUb+Nia7qbcZg5gKadRbYNlJEs0JgXzFSwU1GIYo94Pio0kMl
VdJ6IEtap+ytnGwjtfi9Yn4t7kddo11r4lWOGAqcVvknuT1B9amrsGkYXpOTyi26
yHvCrczZZJ96aG7poTeQTD/rcR2iXYFqm0IGi5YAR80/UQQnW1YXVzxPWvxSFXKB
ZuwkYKb41ALgWWYprLHKUAZsxbhZZMlqHkxrXj2omrAcL6ODA+/IYoJsbUU3048s
wkQg5UaRJa0YGRhSVs1s+Zl7Lsc26IaCeu4AWJUqQvdEiWVSJfpnFCcV6Q0bcHBC
Tt8hsDO95ntUAKtuOhQ0vXmgLhXKqHl4KWxpfNsjZyMirYD5Qm/hBebX+qBeTGRO
HfqErw3ps2P99H53hYjcbR/mnep5GNossTlFE0NoQQPfvd+Qml3qK8+9AKo2MDV5
iOJoMbjLxX2AdivnOwZ7+TRh0TvZK4bd+JQ06NhVQHG97iVYiFBB271rndt/lbZ7
/JMrX0Sl68+Ki8il9EOtSrB2r/SV8pJAam2VO0eWA1Jw1Snl3DbI1HzOqER1kwPt
N7YP4XkAl3yYI+F0GRaBeKYaRoPapsSD2f8xR7Uk/lwxUgi6ew3zqEFOyulEfco8
DVHigY/J+F6+UeMxEDi4TCczYcCQlra1F07TsZirzJj30roqZ/LqGrFp9ORLZLyJ
tj2xxOGS8w9gcFGeps7jEt0NPZAcC3Z5XorqqYbNbPZ8JWFUmxgeWE5uN1e9Zmfa
HTdFNJA2NwslbH4vwxqornFZ/0KGi+qz9CvU76Gi1QvEwallDhgg5w0uzWwI8le0
YoaSnnfWX5ZiZrsUhB5uAYPEatb2OifcHXcrS0wZftpE7N/uU1uD6wJMnQ0Vep/6
XfSsifqUQB/69m1NogSbh3IvdAZo89D1AP3+sEaT3vXyRJh8Z6JNUNmKB3ODFM6j
8THiuyX/m7WFwOQ6YBiZ2SobmF2F2lk62BPbNWLu7aHT4VuDkZSCNS1nNFdyWPur
GbD5oyhvB3GHwpbCZ3CoKJuNRfMPwgdguC1EdMNkkGy5V6cQYyZtZ/WNGy/4twcX
/pGKglg6z4DNT4CXSotOiq9PDFxKLQDT5GKjlnZGBosGSl8e8PrgsHKRe3y1b8ZL
UjMr4IcE7ggdZBLjlNtoXfM0Ogvc01pGwQuZ8axvcJF1CXBhZUE58RzGyjhXrZGE
zk8nsneDQ5ApAC4AOjTYLXFIKqyH8unN9gM3sO6rOPd2kjOFHL+qZE+fSgjnUx6v
/ZyVU1VmmQ2+6FFtuAEf4bFSdrNlheZWz5ljqTX8k+DZaR7OHS3I/rsid/w3VR44
ZQxnfIXxr5d6wXjdmRrfK0vQpfCD5x4NKAGOCBVYjJzt1+lgDrazYBfXp5iXZr8b
ybADH8IZeWz8JUdX0npW+2lZ9g4pLDh7WNnH8eCL1mcqNYwKytIPwYh4VnV2NcJY
4ikXmz8XHOP8qSEeqlBOyF3H1e4f81tIGCy5KpTYwA4vcY3+raalXZexOPrkGpkE
wWg0oqtqkm4iQUkRKPXoYxZ7Tc6iCjb1hTkiBrRvZF404LTjS6OmJ8PCAJxaLwjY
mdSCzGdpD+kXvbD94L0u0wAYWQ5Inmy945Py1/l7gI0lZPLNKg6jXHKaBanxPzx1
TnvFreVFHu9+DARB6HHT6VKtDftzubQRmgKfXpPbFhtCspVWvAXxDFZafPWi+W41
z2yWzK9p/20GFEn3Gn344wwAEhBPSh2VfXwGlgrSdgtsLx9k+dIk6+MPLF+4DYWz
7Ej50OA2YAKaVOMBEN4I/Ku6AWW9j4r/5qyQFGAb1n7H1tMf2u7BuHkJfVmc5q6n
FD0eTrFuR7Iyvtapz8/GxKa/VHYCkqEqRKEwqthrDzJdd6hZgosst3sK6o17Ijoh
G5aBr3jL0CRTanYMQsCSVx0YzkO+5FLfr5Y5M2zpId22eKwg/AzjFDqsg9J6usWG
kibJGw/+NcTEP2ZDtSFo6PvGUhD6HI8G7gRe0xaq+kmETLGST8a7sInlQo9LDhZl
Dr/QHkROOlMK8vUzFPynrbWrUIUkVuFKQBd5l86Utba2bouIn3/KGvpa2WAakYNv
Gh7wT1lH/TEIPqsCszhyyQQGvFcZAdJ0pEgxuTPas1QN22/Ovk8o+Th/W9xfPZdN
2nFAO96N5EwRfliBJ1QEndc/p0AzCNUDFQ0PVSFplE2Yx+8PlgTMXNPQJYfA0e42
QJOroyzbJKGj/DiRFNRYfyeEDrDzkIvjXpiEWjACrMVaKINvzJ0nWRPgG9lPK5db
j+e0JAdQqkO4uzIBPWZsf6E0RyvYsm68x+Blr4NQ+Udodr6cQXhZrI9mjW7Rs1X2
lTi1lk4UeEgz0x5KzXcfLg0j46Un30qSR/Z8vjMKT08RDDL1zTWpNOuF14870kiV
cZud8tJPR0keAhKpUj4P/JfFx6T6MNKin6wHm8fwJfD9zXalae6DOnQ3TXxem5G+
XsXEjtI/KH7R5BFNm5o/OFWZ6zap+kJs8IZ5kc4jDHXxQfSJNuMlR8jUAKhwvZWV
CcojHr4fbvGoAmTiYNi4IcW0rUZgrlYUJWdG6gJRX16oONLetgIXEhkULCsgR1ge
27gpwiB3kN97H+Op7zoXZEGevl5VazclageKsGAmvh7FpbUhsBwiOv0DV0c6CPmD
CYvBYlnY9IAUSGKwiR91fNCqolS/by6coW6rttsPm4+Iz6uo7A3MnPYBVG2fATEG
15FZEpR2kKJ6YPnOJaCl3L0AU4p+mkaIAlJ16X/EmgM89yf/wpW7kK/ChwmpVdfL
8+i8gVpgl2J/7Zik0iBCt7ag0aMAzpj31YGfnFEz/ZGvtpWHi/gReId7dB+pisKw
9zMpApqt9hcd6Imx6veZMavcUJdu8Sf1yH17ZboCXSSY5i/hbt5pLxDjCqW2JFep
7IIKxrY8XcBA7hm7Kr7tvCCR9Paq1JTc1Fbc/GU/1NlrnQK16bGRBqlQ8/N3/QGq
8IjG3v1H33cwk5DJ3V9XS74HAieE5Y3uRU1vRc0uSwnTdYRgNt1nch4bhfxRXSBi
m9Vqa4CBGeR2UubxbvP6yTpjEpVM92LsUdrA5EW9LUVc939VIKQaKnPqaWjCOJ1Y
lWpmD0AqAeeRFTZWyRg/GkGnazkaIjg+nM6ZhBKwhQdpM36m4FrCa9Dmuk/EdI7K
CL2RuBZfFduVkA1VyrO1nvN+gIJEvN6r5Bhf9f8aRV/SuTU9LpIsE//MoTd4cW/0
frzkPJ5nOrQVKz7IkMBYeK1FZOUFxyIjoj+DC3X52UaO/yCtCKw2RcqcpFgSxJcC
qNBI003NaQOhc21pkqXUMjzL7TD4JaveuZII4NHMHPQH8WTD7MPAPqD+0wc5kUwG
n3ToK9cdNOB2yQrwzNMgTJ/Ga3U9YevBgoOp1DflAg0VAqm9IVHXOTa4JTSRSnOU
pQErQ7TfXyyvD8JS5IHdjBMncGzXkeRB+7qkdQtvIKqDPTdoAHgAgI+k/V67aGgF
2jjQaY0SC/AEeZzSA/Vjrviy/h8pyXhHVHaQyqhLq+HzDbkdP4D8Y3V9vZZCkNI8
xWQaZmJr/oavIGxym8zRcVVNHKasOQDYfy4L36Em/KtZOtUOIUJX35DueOy6QQpc
BqP7f5PUHAWPeyGvaZp2OQcom1xkxDWF6B4g1B8LBKW3mhKS1lNJ6V+88wvglaYD
vIFRFSFj7ZKWsb/a/FkCZOHf9WlwKTXXK5YqS91e5g0weDhC8Fsdfcy9SOtTEHYr
WPkXSyC55APwF7Dj/fuGVRuuJOJPDWcgQnHmZI/8VZP3Fs0+7AiRfjXYo8W3cZcP
7lpSjTl11Cl9t0fz0wW2ZJnMq2xG1BUDg+t3RQTrTl3Ywm98oaVQoXPrhQFOvWVg
wpOvvCyzS5mYSSbrm13ncth9LPVFK7fmXg6NbP/kUX2EQ9eGYFvO8gOc+BdEnx4m
s/tUDH4ZZBghXd2/vmG/VyyVQMIjzLVmfXYrHoZJu07QIjJvzQbfZuEudZzswprS
Fy/RDAxYw0X0nEl3JpjRzjFNL9zrUqjY7cO5DAw+6nGAvABO95tOLaTTmrf6cmCI
ilNGbZRiMehps3N9XE9bw7ms8CoSrXuxU3p3MaePiPBvWrKfvlMrYQg7yQuR7x7I
qNN5bxZKP5lsXarLWZk5ip+ZTLh5RTYmexqWSey33E+IlNwMxro33bYkQu/fYIKO
T9ZtRW9gT5LCGyGnu1RHDu/mNOtF1Ak0npIhBAYaPhNFl98AIgfqraWK6IzFdN1P
t5JXZfysjbGZlegYxPXAk4Y5C+/Cq8q66c98H8uqrlHTU5kod5yzo0pQHc9GE/0L
IEJENpK20MMWX3/oVQ7M3lbpRKkEDzJMV+Zl/45VMrU7knITCv+n8hQNENWKI1uY
UI93c5OYPmD0BNo9NT8OS6smO8iH7Dsq3o3foieJAOuFwVekjNto5iX4JFejUfHr
ctxHZifH6iGMBi39U7bP/S2w12G8uz4d+jRPFQvzhVrid9iD7jTYu37mD9oL9ueC
kydzv0SB82PCj1t694FenLM2XvUd4pbzP5v1GrMDU5b+Dg7jpvWGG3JSPGT5g/w0
lqGPKwRgc6ePadLwkrIvq+VJoKO4BNKKOKwK93OPVSG9rFMzM9rsHPxPLbUDy4uT
fwR0CWPxIteGTUxFsifByadcLnVtCDVirCX0dq2fc5J+48io35B3+RA24LXnVr8P
SxCW2WiOaIuQJpI1Ffh9dm0omygkBB5An/Nd7HsDe4fQKz3wKFeC5k3Fc547+++O
3s0Imr0yTYV3nHP370LSYLolqv8uLblgCnC+6v0Rw2Tuxn5lukmZBjRVK6Luzubu
2I0b6G/KufT+CuDi1yemDi0xPrybHCpYEQ4jqsJokPaq6V/Teq1ZHS1GUnEojdMk
tMkZVUV9jIjMvg9WnvFIT5uddd7vXBPEnxW6XFzpOoK9TQAmHd77RJ039UCxdgJP
cThmBhjj9bRq6lKNTBXQAXX4NsktPjshAoo4uze/7L6PDqGFHcJhHoi6DJDhGxi5
ruZMB3wj3j/ng4D0ZpCvbBTZD9dPjl8fiHaG30z6CrfGvIiOpmUO7ofle722m8qZ
hprFc0HUL/QmzjPgUOl0SELmwH9bfjAYNRW6s7IHbJ9nGLahGP807GAOAiL27s9M
6I/+JCsVD+nWuz8SNNFzEWgt0SA+fFv4krnMtJG1cM/LUdqsbjLu48FbDDivBR/6
QmANNMnBmftBnZzLa+bhA5OVtESBkCIDmYkpjMx94wh5dawdMTalcSxgm7b3K26+
4QoK9I+UobX1nS7wvG2/Va0KShlPn6gjttnG7M68T1ziVEInTFvkj2HYuWXMWE+n
iQDsiwF224MFt1OA0ppBPsmx4wbppz7B1OwPq4FmiB6RAo6rTLjnBBb8jZHk1P22
/DBMpRz8ll3V4ZsN1OJnA7841ZQyEyeAHwfml08JV4PCvilonbmLlOie+TDI+gl2
DOzE0NLK7miX22+rwW9SQ7nsoc5CLUfczTYFrFS2Kn7XjK4cTj1qJEfSfgPLeiCI
hqd48Wqq4f3dak4UYGekiQyYod8OrJx8CuIsbT53CohW7LXnvLeZGrUYOQ/gmjsg
MPoePKkemofZpKGjBrdxEdfA7nZsH0Yp9gw7qlg+6EGezBW4oLhTFxcsyNiRVOKe
QwLgD/70c9NpGNqpEPWopNQjm+DLEKdoUcJxsIPLFgI75vGltoUJvrNAAp1gyGbE
hCq2pmCIe2M5sRKaSoC4Hek6UtJcxukQS375pZ2NiME831nkQd3Gc30/0Z8OKnmB
6+Ta02ugDxwpPcWA870NmpE+ypDSAZA3mu5twzedBsxQPBGebyI76/beBwPwo1gb
05jDnAAkNdAHtq3TXW//P+yeT/qF7AXnqLSdQKAmFbn/icM+P46gXm1q0JAIowcj
aLaaakqIs2Kc5kOSnxOFiXxLeYRb2pYvpA1+FDRVo270XBzHo5cEppl1U315dFLq
vOxD+1epYIK/LcdxQWBIlN0+e07GSnjFzIdN4uO5iQLkc9r7cbn1j9jkyxmoQLyq
l6y8W2vWh0nmiJKPgisvXd+0hzetXVUul/28boVMpaEpMHvJofyCgeTiFHTBRXwR
226a0vp9ZNj5YpiyxDrqF1EUANGMpFsSddb2GVGIr3dcn2uDvS1pq/WLCwDme9PE
MNBrvciGP9AuNa5MeT+yOmSEPpafwai6bOAAFYgj2IkTxrgHdXj0Y+AeRQ/Ma1bA
nepIXgDuu9xOfftncDTHBKhmJ+RIYUFoMIITGZorbT7kiL4hbOIYo8gG4EVd6Pym
OyYjUjwlheuwCjW14J3RUYp+fC1vXZgnkiq40mluBdy3GacC8bJEajDeFaDxuKJt
5B57AOppsz9CgBmmTxmkvlEzxNaAZQiMn15+fxqOlGS5y0b7deVn5JZcnOHg35Ke
giXPjnW6H+5ufARxCp5swpJSEtSx8HRJ5SfFFItzqbrHrgQSluM8wAyDRnZSqn1I
uI88542049Xlr8/j/GPpr0WBEwFWiF92EGu+mrJpU+8WN3AS55woXqrGMWuoBaA6
iKDQEfJzC09XtrB5seFSLX0jCrOshymPeYHvVpRFcfsmcddMtT4UUcDVkoDEkteV
dsxWcG3ddB3XvFnU4OpI4KM3uvQ2Nylym3mnGZXZlfMmr0L2EYh3ENMXNl8u2dAG
j3wleoG4YKOYDWzqfLEPGgn4MYTfnKQpl7p00ZEG/J6Ydx1rNZaiCG4kNi0Vaugl
9nFToyfQ7p5tsHRMCSjy3suxNHx6SIgh3bWVhHb3aNx4yiqKoktKxqVUlmRmYdjv
7IAKKLEyWx/TnYZtqpSv0Iv1lkiCqQ7oo1pU5qFKpfUkHCmgwF7gGe7lYhAYMYMB
dusor9w6tTUSDQCiSNYsNJJvtnBQeHq0xCe32994VnZGTb45P3GcD2qKlDY70A8N
ZIihPNoOh2q6/uTsye1LeOrGnut7XBb33PLyitnGe2tHRvbbGQJzzr8gUDiqaAHi
qh5Z/AUaOSU6DGudL1L6m/EUSoswrdqWZvx5G6l199A7bAK+0PJpr/7mQslEi6yt
01MEPK4ZaN5bw/u17GkPsPHDZaQdtxogfgkdDCRxhT+QXC83LnXlr1PEsjCBXLQK
R8oJYkeUCx2DrAoqyrNDQ0z3CWm2CYvh6UckzasQLCsd5ZDxookLhSF9aIqh+Sky
kF52XxbN1cRJrr/Sna7ZyYBUDQo20vc1bcWEyUghmBNf+Z2ixZauVJPEUQu5DkDv
oVu31J+pksqeKGNiAETnTY4hxTaE4QyvoXAgnsXTPPNnCSWC/4wsOVM0v/2y+CJ9
56hKxiXo7u58YAvzXUxJBJ05EjDlNhQVJwiPcxffGxC5IHT93r4mZ38yG3SGisd9
eeCJ/qqYBmwjql0bzPEZgcC4SZ4vk2iiL+B4yMua6zkpCkx5rQ6D54C3GUJJNInj
WMt75jTvvM1D8R6yTxdK5BIIdphkoG+VncmN+RF8SFTp1DLeU439TsiUC8wfA8Nh
PwMN2cy0GsWz/+ImDr6NzlI/ip7IQCCezQ976hVlw2jUSWrBhcjj4PC4NkVojvrD
ijAMwSZEjpsymMhsrTgKguICdlcwTrQtq/kW7XoBcZmwhqEIYSckc3kdFAJgy9Mp
Bw8xGhPTI+0ZtjW+82CVBkDOfAbJCiPaOwBlLmIMYQPfaaQP19cv0vcOmiPMChKE
jgmoAqTbecNThQ9YZWYMCSjgIdmbdeB83wrdZkvEAOFpr0rNVozwSrdSJOLf5SVn
xPs2TXZQLlVoILfK3CevkluDGWfI1Mx5uvEvzhvzXyuoePflDjQNUbIUUupOJi63
M+9CbX3mKDu2LHbwY/Dz6jGzzY/pdt2Xgyrbh+vh9S/LoOtZvdIkHi3xQTR1nfzI
MXC+mCxtwlg+HqXljNHDgGFGKmfELxnKF2FioDevKNkTh+6qEVy/XJJrT/MUVzJU
7CV+mJ8AeAaJXlVwrC/Um+i/EuVKklJLfDpRpMlZ71P8c0aqKXoTQVdehc31OL0/
ZPjkE01LmpQe/qmTtQrEzyQodPsWUbeyH57Zqzk5/GDh9JuFywaQpUuJxvEpP0BC
HkWneY+8BAXGC8xwVyLMcpG7TIkCr98VWU+vBNlcbfMRssSEylPtQnYPivffYNKL
PPypIGhArbthrH9GZ5oziYdBH1JMxVS37xRBZFI3gQPeTSNc8u5pnx7B7RN2YB0e
rwQ+x9V2xI2dFQ0aaAv4iBEHgUwtmzd7rSMLLaBRo0ev9MEjOyVKh/ZMK6DuA2Aj
pzoGAnS7VQrNXhMKn5mfUP1anS/9gRQko2bYE77k2QZ+EaXKrtfBa/XT3MYRR4Pu
vtcBaUqAQjgm1ZvGLbCiavRFR0y9un0wHuuHzfOsNlzXuIM2OuliIBPwMD6sqOdh
FCkpAKfal9hiuU7WsFCEPcqmAVJ9MnO9e3rGNeQihPEjM2L4GiTOhQn++hmyqF63
VDeJ5aKpyidCX2dy9F4iy72vLhf08NC10TOXWS3rff7uwHTr05QiSJdvmQAW1TMV
8lcZXxkhtCLuAPJ9u92ZZeDhFsrZp8Nb8mBw5egbB8/FrS76SXBHuWg3nV+d9Xj/
PN3XhCtwNF4a/Ggd4ZNcXdlBujNwoKmw4hWiN4gw19DAphPNLuPvNptvVexGlq/W
Yyj1RxlQO1OUQMeA69nz7wjInOt9P+oZlu8p64OIrw8Mr1EHTOgAhX6Pm6ITMtPI
bPdwKJU4ITAd76ie5/WjDRl/S1zP8VldaUjoH73R18TL16/oGiDgLBh08jdnLN3B
WWiZtw7z905o7idzLnyQNjqnG6QimAJWWD+x9MH/SwwA3R2kMgYXiRXqVOHbAJ1b
I4Drzrr3wBLZRvZ0jE6u5mu/zsN6YDPPyOrawTA7qDnuSls7zzY9LzDYFCqlE5lF
810idiNHcAw7I7YoqXU6NnWWEzwQgdPcY7H4ZYCxitXaRF141+QKn/YIRqnlKwXM
imLc3+EFmJCxsaOmtp/8MmpSpoDLs+KznuzOcNpW2jW4674LFNYhWM5/B4+wj/hS
iOiS5nKZ7otPSl3gqWHpVGWMHlY7e7OroTUQxA7IlhqhjzyKz0OGrUnywiiiLr3s
+DuC3t4ES4hexi1NEl9YnOi8hwMsmDWUSCPl7nqD1L3TFqUUc2rENjC+ctFUHs1f
xGz2VhUD0IT8yneQhr7d7ARwa9OW2ZBfPJcBStIkV+NxmNaBv5FyHudJ4dHTJ6Zg
gJk/E0N5Tb6cUOk/DZhrSG4kzyDIxW2YfkYDs/7HsbBFjjq+gCvWtXKaamsrVVx8
jIE0LwRhbwSHDYS+4lkoSKa/u2P3iObQI9GIBTSZsKV7N3m61A204KL/qRU2Hn90
YeI6sj10XbttMmWVOhE05uZabAyVlrKi+lpuBgRDndYqspZ/jSe/wUtLIer40l7S
RT9v9tZWNbNhFzHUyW5UStb0lqQIw6eekkqBljkCdwcigQj0fq1wTd3SSvt/ZmbL
E8MsHKDNLTvCBycP2A7mNyAUDl6K4zORPr0sirV+KkDyPnppTCHgxsrU5SGh4xGk
tMFmJCaZkb1BTP8vcbkffBVnaOyus6J8ZoEhiOTh/zy9yJSIJR1wkxF9dVcOaRgw
ZhGfU6lRiW+sNp2n9WteIqCanERJqLkMDX/iiOsumO2Gulh7PM8iNgLEvxNMF+/T
CXZReDjh5jwnW+9E9uYdMJYJFdNyufCDS+k/MmVvFPtzerSBvbUNZRQWsVbT8pdR
7nvhC0uYnzVIeF+OuF7UUFMk1KsuB67uVCUAsTYd6Tw/BJxKCOLQAgSEj0PEbnvg
minHdsMMTRkhFxHjTVVtBIx5Iod5kc5Ot4tchNldYJvfxs6XuOd27n2m06XWWQ/a
8Ca69SdWQ5i3LN9aKol23W9CEdvbITqUHOzr2mh4Dkl0pCnyJi1Nj+RvbOwQxrc1
nH1hulnaqQ2nShmr+LRzsrZFcFydHHDMisGP7fZZcfxfRLCxkYakwbhRJmT8sUNZ
iTVA70bOFpxTbbfnFkEKwsM4acOgvUkYbz5QMNEy5wIvL0e5w3qNzHe/D0W7HiSg
jCbwvr5L5Ngd6Lqvh/dTTWCsNlhbuRhmCgFolloim9c5HN1lfNyjGqLjjqMpDJeK
YGBQx+BR8nyyTFQ+xTWrI4+XwtTdYc3DiM4JoqOKfbfRqv/zIRfuBBocwDiLEfB1
7HM6rBdV+RNAyBHxiQw6n3x50aO5Uhv2h/F+NeR0uCG/Q+joDnYg1Hst06fGF9eR
DNAZ7Ue+pF8Wp5iO/gRGXHDGcYOaeXd4OEzObySGTPjz1qiSme66sh3NPFN2nDCb
MFsVl2sFbJodMpH4fIOuspO9DwarLzx75Kp5LKLCeUCQan9nAcnxvuqquSjow5zU
NPFFQLh0e1fCVl7loZWlF2LsVUzdt99UsKDE8Y88KzUbKmH5y5BO5mCkvZsgvuDR
IoG6sIJy/bQLZd+inbi3bvWc9qg9wnfO6Qjk4HSuq3VrxbP1ARiBtuLW/f7HnAvk
f63gjQ2TURgQZkMisz3D+QT2E9GWOhjXG6wueJF9Iew6SXerW7k8vV7D4UcfhZTB
ofiOnHkYXwxbrroK7afG6X0x++vaZJiPl57QRNRcCtfnotpA19YcWgXeFom2UGLv
02KdGb1NsVPQN3OHTYsmz2gXi6ev9sAqMvrejlo6+LfZzraZ+aYdMrw4nroj/yqK
+utgzJqNYP23yXpuQE0P8l7z9a3buzw6+Qp/ywMdpjR88JlHMndVJ1joNodgqv/V
4AJ0FW9M37tE46vrpoYPqvLyeNp5oY2ryk5F3Blkfb7pBvyVtAFKBIt1mTU1JpB7
xfdnXxAj7hcZgEUiBxxGmg+47DkqDnIJxxIE0FhICR53a0Kbi0KOg5+N+/fCddlP
jggT43GfaIQHCwyy5t9EJCy2pK4qtswo5Ga+Zpe1T0/WAYuShqYh1vEvzt/d1xvv
3Nft7PGPj9/HwCcOJSNm/FbwA4icYm+ElJXopyeodkaBmVfRH43B5GnULpY5nYhm
88SQxb3nfdyP91icUPuGfP3crJubiYsPsjJzbtchTh7S6nlNQnbnN59Qri+Qb3b0
scRfm8oJzi4HqPl5ByN9Ad5weY7zwEqieLx7q6fjBz50wORIP4KMoGcm7TmSM3hm
lTlKaP0QH8EuSuSWRdaZOYqabRKA4h+w/R7TqcRFi0LBJHKTBftI6CBhvgJEmMyP
6QMXuK569JqQ4lXyP1QabRtQemNpuA0lexxhZoGDz5R3BP70v/JPl0B2w2joWAAc
vBWDtR6P2kAyJHlDVOTTeAXkYwiq+PS4yr6nGZrTjm72xFFeSz5JDxcPWkTfjf4F
TDlYBicxDR/JV41wF7tkmfEfnLYemx5aOec4VbQq0Zvs9p0ukO7bLkXlpJT/9whu
Fg5EHoM6/yJg2UJ4FTFddZx7xv8rwVSUOfiuqjrw5gblfQJE/8m/c7w4923SF6Ev
1NTKEhNkvjnoifFbQN4SCWjGdIUmFp08VMPWx7CS/06isRyLo77NQ7BUyY3leLZT
Wad84eEX7hRhF21R3EyO/2B64VMaf3AjjU+GbB7ehNOZv3N0scmDP6LyakYhupNQ
eZHHtsvXxdfpG4aybYDjx68igPcc7g9xkiwWLdxyD0V7+x1iPXWJzjxkQqD3vyr1
Ei7HW7Ea7Fr9RtDCB4j+NERHjX8C04QZc5xbX4y+7b74ihXyXZ31waBvnKIMnaCp
rDk9sHWre4rtcEBNEGAgepaOk/wPyaYZDIzf8ZvhVBhsdauC9FrYAaOl/pX7QFy/
M0Ixtuyb1B9e0S33RcdtrkrC2Kkw5w5qHW+Pa/uS3QXnW0uVqSHtsh5fcI9xLlDS
UIa3xZue7sLhcotaqdj+dFOXBy+7AeIr+F8g2f0KnlCvGvcF/ENsH9R89gIZvldX
u+xENqCYVTLSCozFlKpO4PCVC1IWE0JBpE/naAdWLBgAgu4pTbF7xv0dAnMOhIwb
UwMduL0afpnT4wnkXK2ApUwRpM/2zvKLMuGaos6hgT8+E1leIyqohjP9psNyP5go
Gdjz3sggOTJMOaEDNdW8W6NUx8ew65ACNtOK5m2FFRwuAmFYpflF76s/bI/fsFUs
1PQIY4yweXGh+tNBve3wh6XwLpnpYB5fS0jL2ay5eE5/yj51YvlRT3X1ByfQ1oE0
v0g0LCz1sGPYS5o9bGNTtp/pTvT0rUXhTsLty8EA7vKpsUI4DfHKkyNfZyZimQmZ
d31CGZ4/fRa2jggmclfqiHSvgVNzuUeFWdHL8eTnn+lLLfkb74f2joPgbnKLBEfi
TLsEfBc8INIxaI/XxdXRxgl/J1RtIS7z6QqcC1UOmdDjC0ze/pjKpDhnjouxLuRb
2BXBBHL9Muj2ZnOGy88ad+oBMBbknVu4e75cETDrb/ZEjaxmsjpfEZMFVDQb2eWL
w4L42e9DP3+7p5AArO8kqxotQPqv15dGsecNLXQ08MaMewDfuSQZ+VY0wmdkWsoh
ndHXthjAugkIPsJQlmbD7J7FJ6r1pLki6MkbTX/BNSXn6lBi5a/QeaK0mTyKQjsg
Zt7SdqyZwES2FwTCdKLiUZucN7hWZZRB5wIqiNXZsZb4dXtEqZZIRdyA54e6fTIs
1euz+3i6ifBG1Mu6LiDRwDT2xf7FoKHpKT9M36XuoynO44+6Hv3Z/sFuUsU7FHka
7TITEYMm4pJgxMt7pg3K/jBJmWd0nAsiAJE8VALtwfrCCiIoViMDveGmxhhNGk7h
xHkr9JSkS8ehofLbG5vdkybVE5CvXaD8qMSInRv1dJ7CJIgdUc2pnaQmXRrGHDpV
PnGHlTB9PnIxgaM+sqaUZYTP9VhA5cwHVZphZJAgWOB/GWcSbq9ZqrGvhzDfYB2o
su7e5fck/+vFGgZfyHgMsX+BhrKJq73aEdviiAeEB3gvJrPamyl7xFq6aTlfg2t/
MH5f1ha3Lf6hkjAFovUWddJ4pjNEAtlo0RKjP2EmBJcVRHxH0MBwtuU5BmQG9Z/C
wcTgRtBtLuDkk81RGrL9tXLpjGTigqoN4XHbZsjEQqr9ETr8xGOs/c0wp+pktwmk
jw7MF8DD+LfZ1eNaVWOBKs/pPfyUQ+FQXATCASc/4oGnSzICkEU4bc8JxEXX2HNg
8sLB8h4LwoHIC67JzM9jM39J889Lmih7jDYGAsu84bMD5gRte0IYtJV/pfi3hv1v
0Ue2ezzoo9CHw2oHNveKSebCQLuSewb3swlxFdxspqhIw7VvfXelSJz1Z08bjKxo
BieYlUCjBYGRTg3nR2MqdId9WWcexbX8YSJtds1WMGevY40YMRwx7Aq3pp0Jz+X+
rI5MUuuPchGG8yb0d9lX+t28Rezj9mgFx3viL8l3zeUUOLNTf69lBFSTo0UAKQHQ
4DCV8+iyUOWDCE1KbeyvutHYMHgFgUsepKdOjG7z0pxWQbpjaGHwVmLGr4J34nRU
NBWtCZWIf0NGg1LuPlt/dQ+B/3ASiy+XvMxssbclD2ija6mlnyzfMTAXPl3MM+Qe
IcVhcddN6ifI2Y5N6LNJW0Wcetay2z/Rk7D3d8QA4R3nse4yUzEqu5iFo76624/o
TOUjzik52e48x7t1V9+oXCiA1jvcmfh84PtKK11w2riuugsyWkwY5NIzuCxqbO2L
Jf6cm/u4hw9FvaIwSfEf7IjFnnQ5OsSQg24ptNfAfrONdT3Zijq0BDu7ppDJsKYA
OxJmt2LJLP3Mf5skr4On/w+sndNPONNI/rE0P50gCSvSrShDesf2LMvhAnJZxNz0
cUojFnDdWaPmWYhHem0gj9r/zYS+GFMpKrM0KWDCw4MK4COP56Zh0CXL2C67EbLT
p4d8MY92x2Gvc1wScOUKfoXK0XeJ3yfSeYG79oRp/fa+oT1HzHzTEKj3Axj0FvBd
V7oNeTSxQTl+duB7miZHJeZEn1fB+T4bYQQGErTLNFKsOyJms3ltcA/3CKYkTzMG
ReJqJdZkrc1PFTnhNyW4wxwr1J9MTPXtZ/mn+4bjLIS02QAI5V3vARbZQJgY/f4f
uM+XhA2dIO5NnsXnUH1O2h3TzBvY6ll8t/O2kashd5qCHqURRjStJ7xmJhjVJCZX
FolS+6L/vDvB1axVKOiK57L/zqoug6jAogdxGBLXDYhZswFKooFD9xemDCXZvp/Q
jnCk8lhAUMz15qsfBHotKFO4nmKyMD9WSBCK4T+dDja7lhqenj5hb3YM2b0VVfl1
lCzZvaHOe8FcVDCD5jur5HVpq6zxD1vEl5RFzUIOwKD/KdyMTuChYV28No1LeKlX
8GrNmrCoP9o0sAxS4sWcQL9SuVlVw1/EEQZCUtldidauskZT4M9fKTiUNgM4j/gu
HAvPTloIwch2K4xYN7UIrUEEo/f8yrT6zAyWw6IUdcOn4tTiDhYBnRW89p5iOVNt
3+QwBHPoF/38AvrXnFZpCV0vPi8LQ5tSoccCAmsh7imEaH+8cOhExYvneu/qY1Es
aZ9Yzw/0qfV82SNNGB5lHcc2ap1+1FgWlwWbXbztRCi8ViJPVf4jLAHLbS//lz5d
Mq6tKEpHvd3zUM3cS0G/3W5glppKVHcdt5xpNwp7xLGMufAA7TXvQD1mPDm9ce/y
pi7+fdOL8mqR6VkhwUDsjVu/ALTovJh/ndWZuiQvc9kKEZUE8X7MqAB7RMjU6tEH
HqOeWShTyz5HAB+xaUkVFgZcwERoudylcBKwYAF2fqog8CKpgfhNt5Gh9Sy1vbA6
xImAhI4uoy+WonukdRck8glaib/Y93YyynJyM0NbVqShltelrVdVJaPP2La/dTg2
hmLL/37n6Zj7AjCwKMNpKtXrvow4+DOrQPdZJM6GrmUzWMt3Vvu2LNJ2BuEGEZNs
GQa+Y/Tsa1SZurBaoiymR3cCNW6AyASSoeNKS0joX2eosHdXtAwXj6xeTMH0lvUB
qKFSAL56zh3OPz4zYAM+eBnq2afNHp1srPNVyFhjNd2+TtDhtjdu7mIgEf617byb
r2Y+SLCPwlbX/zuAQejRjmj/+FOQhL1TSm/coKldGQU3JrFXLLCSab8V3UgzZTEG
0GAmYvIF2l362FjSPCOLX0G2Jqitkglmhv0TM5wQcqbNJbUuWH5Pk2A990F3Rt2C
hz2K3VFjW6Q16uB880LHYRQISzc5WwvhGy2PmOaqC3f2ous+xmBwN/aj7AMgAFTl
8J+rg7QP8TZT3/34KsILXnSI+0ZKnSvpYmWKa2LU7twsk66S+jeV6Z29NOT/Ehy1
ZP/0QZWh2I7qcZyJK8g0GYT+TYiDwrSSjeQ891oNJTp20HCVaNFlv1fZkAR7G71Z
LT8D4AxQCF1yJW7UP68wIV/s4EyZbIvSIDSy2FQbVFfqTGentAcp8JP0V6w427JK
ECVO0Fj2bPTF7lJ2ao+3LUN1FHSY9KLwgSRJTRtfPeqkNYF5WVKUl2a0HeepV5Ll
2S7p2xggGYN1RPXiPi5BW8jp5Z8oNUgJ93kE28aCIXLTrTvRc9dNbfF3qjSwjWxn
5V24a6DaiZWiOzg519k35wJYHLv6FpYwkpKZFXqrAO5w8GEVMH8oliw1lBwYoNob
z9EGx8b+IOE0UJq5f/7Ob37qzT518dxJkHMolBoaExnXpORMOCKsDF0R1JIKkDDP
FRR2OvN4r1JwAxbc3sTRda6m2HG74lhOUZKQRphCmL0lF6+d2VXqACyS04XpBjoP
DBDLBZfQglqcOTjwBlHej49jGwowv/GJs3/yLog7r9tJdqvkmUk3G9hjhpcUErSe
YuYYDEpod3jWnFYNI+AemUhjzKW37t8sj0M714YKbTbpj7faVNp5/azAKS/xUqFL
xKSqKPpIZucLWdkE+c88pRO1WxleBLiHoIotaZZtM8tA7Xy3C2qjunf/3hjh3bmm
KuI1DLqnt9Ggir5xe++DlpRF87q/1oQ3aTdtm31wsH8JwX6vdylepBrkmkqmr8y9
ylB3JmxZKJQvelDXRwVz5HyKGCUdhPOCJACtBofnp88pD5RuwIESpCP+xnU3PzQE
Qr/oj5bOzznBGdwaxdGy/ausLwpZx/DDhqQsgLmSb3V9LQqi/Ov8A13/C/JaWs8F
PQRC9PQtbSlxK8Cyu/owh9nHIwNLdjt0UtxosW0WK3xhVd3/eEmMdI2VZ7vOt3xU
lmTmuEf51xuVQjRFSxFmavZ2M10dKlkCCliYk/hOI471uq9xkvfvHSU8dC75cLhZ
DYrYT192dzzVZxw2cJX8TgXECVTgcpJ1PcBENCMf/lUy+l82c/d5WSh8pnEHISbK
RRw1GZ60a8Sc42vLux4g8ZQM79L/ytSkoGOaZ1aoB/zW7kvwIMc+bxN79J9e9bzp
JeVpYDGnRkNE1Etqc82Y1hoOMZlvfvhv4P+BnZ74fjE+vaxoidW9rkOLzT+HjRLX
Vm/jOz15NFeayaMTocGBgPXzJXavUXd2tAxhKO3lmXV3JDqPyG6onMI+bhIXBwDg
qKlfeFYii4VS9i8sUUJNHhrXifMc4zMU6MiLA1VsAcCRC6aEGks/3fMIQrnqowyV
4q83jplHqrXf7BkFaPRyonCTBrkT/50rRyOg+phqIOYVmRQVCTNC5GqgAXIKB9Pi
OqENgUMJJq8gfThAgBZYOEYgsVvXvg4O3qSsJg/wQ0aaNoR11NSf0weJ5A8dHZrn
Qh7SkX6POZVKFbXsLPgKDdTI7MRqaXE3p36NlvHggj0s9Yh2tst22uWl1JRgUdLv
jNk+KTn8Dq69+wdY4iQrrKytCc3R1u8tnbGBW13eZQpf+muX0fhU+FNmIK2UHFjo
WUVj5mtjyat/5AJPmbqOcF7bU9B3M2FI5gubTHub3CS6F6vMExexpmNH6dzBXij+
Gesjn6zJYwSyiwqavOjyx4OxJ2qshRNIeO3P9VrpP/GhNnN9l+CpeXd0odyp3gXx
MIk03hGGQ9JVqw/7PLT6utpDyz0k6+NFl7vOmJbw+KiMGQOG9ytc0nvyUCzJqbLr
72+VnE3P6X1jF3KjiTBrMcvy0lZhq82Br4ZcnCW+C+Qr0wCdgzKPybXYu/aRjdI5
d5yVE0zm2NPuu4GggkSAgQVsbjdsf5h+Ch/oFd0pvCLct73yCiHgDxF+WrFZZFUm
tt2Crn1ll2f3tePt5fY/U4aJaP+QlAl5i0FhVn09Bg0WJPnYU4zNsKqdUJsNd/VZ
atIzgdQYM5KWp/ZKGnELmirqSQ55woWRmfpUe3O8ijC9EaEJrLpvZkbLiOpZEkoG
CWcMNblVk7oq5813oW7PeA7l7I7aVbnPO8ubunYS/MBJJrd7IYwstRf41kWm9KU7
nXUTGYEre5SB4bd9KCLYshUFLVrIhpL6xwfxU7ZYZTrUShaTC57fcykRmLWI2wv+
Z6eM6w4eU3lXGPJnfGAkThfDcbFNXQzdvr/nIrTuzuGqt9CMfo3T97Y2ElMobEAZ
InuwjCQR6lRLZeahLHoC6Sg9tJJa/f9L1VrNND5yFY+7IVZigWz7wZQKpTaADns2
smzv0KWKTuVwNX69LRL4RlqYVaPwJ8WMolrYcg1HxGdLcrLjmlrCWYWcgRaHDV4T
TtkS/JoD/5VwEKI29wL6HLHTb/lCy1b5ZKZ1VMAlVi6F6qKCV/vtC3N7FGFdjC1J
IuHG0wnHuPAcZdCyt5NRyAKv25jPInIl8mKWkfFmRakM3M93/TPxC9Cun2RDIb3C
3YlNBr89JP3apaw4wpkqgJehwADcs4eD1h7FGPXmpnZz+bAn0T+jDbRUgtLKLfRP
OE48sP/V4HSWDez7db7JilhZJetFnli//lnEgiTpBu0ilqC/kSb8FfrrVRa+3RMp
SHorg+Se0lfdAj00oER9waWXehkXeq/WPsJvRkDkvYlTPrl6vGHZFcTRImfi4CPB
Y0K/TJAHHSs1Kuy2hCmOzp3TreWbMNTKxgMEdKp6lg6eqxooPxGpKEQ2xPhx1wFg
NtM4dorFA2KN7WZ4+B6HYQDzgrMwg9wQWxrSZklFO7xmKDVWG+BVJLwc8t30t06Z
Es1c7jQBApwwjKbSdQ0qXjanDvZ+lcjnc3tcBgqXMtSJAIekA6ncrI4U7JvfwfiT
sbyseCGz3IqQtcvtUkx6IGIeLsiNSdfRGQnQCb+jPwFO1LBmVqUqdnXKWkX0oL3V
IY6Val2N2Z5bi9VJiebf7nBe+jVPrf7pbpEzIL15OTiOSFWolqbUi6iSxWObFJNI
TFCLJhiTyrv4+Fx4JLsdLPKNAtzWXbReIkD20kwBosroeBNQt90uVol+EAGyEXUn
+oyN8d5+rTKcxhh7+SAZFeMmDDGJpoBJIykW4CAV0tIXUJ6Ll8nrvXNN+5aOv7cx
GlOp8NWwTJnTmMpTX67SYW/LppWcBsBr4C8QmWLwpNwTULepPylDqjCNcsgFhUMM
a2D+Ow0tPncoxtCqGubqYmA6GQxXtD3x8eFXD2Qqwf5qSdIvrgZIYOmW/GyWjqxU
8kw/ETBTLQFj6GATFhVL9jvIAJnLHSto2fCbVUSJaT/MaHNAY6EkLrztn1Smni8v
fVylV8zEobsOQspk/K32pJQW8GPFtszr5TmvbZ8qHDZGI+RlBNv5ErYplLulaBR4
FfEA30a54CLeV51iZBBtoG6/VOngz7YvZTpm1gZyizZzYNoaUQZDBF9/jfGWNBef
1siIXMJvoCSXh9dWS3hIvEQ1yy154zKf0fgE+6l5lGeLTx0nB/BhfEruIJRQo+9W
qNdTumLS6ohgcstdpNibbRn5hRD8lv9FNg8U1TVzgJ/z7/aqOE1Ms3mXxZG6sVz8
pdQtB7eJTkhAVTdBSgMfeLOsV13fyGvq32cq1PV2LPy4roSTndo+jWnNGNgPjwN7
VynvjmKL/EASsSuAYDMM5gnbNtGaCUsljoGLRC2ditVoPt5Us5HnLIl40ThUeEkL
vj+74IPG244SKPXVazggCpG6a0ZuvpC9DHVrIK7ZI1jlCiaPW3TLEl1QxMT7Dzlg
yLGbu/vLaNJlvz30hMDPerf+ToWepid5QKtT742WBnIjY6raROC0fsU9Ez4pTIP9
/hPm8FuOxEpMFlVbrKkXVyKNMymXG5GHUnQQZRaLLUsOLad6MWW6A4bpOR7Z1FPG
fhfLi7piYwAXKZ8fb/tAQkixSCNip+h4zp0ZD/93Av70IIeApsGf4e9RBxFExeDD
xg5SPbt9i1paPCpyWsIXVazxBAWFGwlriSzbPcwLvfuXi8BCHcFwPFr7oNzvOlWW
aMxQ0mn2aQkfHpZ2Q1Wr+YIbrkm7vfYp50o4ylNVhQv83CSewC1CQ4kUzbNF94G+
RxP2WYMTJ77Nlo6vAwAKoZUD5a2Uk9dMdZ2KTYFPslXXgGi97w2GJGi0VeJZ6td6
+0oup4rnUjZP5QshZ9bpFa8WnY9JkgPfxYQgQxmsSiU7jlLIb4q2VwaqfbmkjrEw
x5I2gKUVw+9csQf46ZqBqEE0T0ZBKT/nuEwydSn5cTtEejDG9Z6ZVBQQL3JphYpm
6USt58DMNXi3a4jeXLmQWKi5fURQeAb4NpbTQupTuQBlGSRzewpVq+UC0CdLYGIk
5wDQddgoZB5BbfPZDVVdZNCcZSB9Ni01kp8sdRsDTlYqTcEa9X6+kZIUBQR3Be44
qROTzSYo4xbPk4B6/vnekEAFtVFHKmAdHm6eiXMCCle3Y8HHDgzTSk6fc5uWzuRH
zsM8evQI0n1oyaeNrrJV8X/i4TrNSBiQtrxnKjhT8pjGdXh2Yi8fzbcxK9c+5v+4
APC+eDqVFzVItVUKOJTV4yR7BfuZ5BpfLRerNnA3HEsLft3r3Zodk8+21MmJov1b
LWa1lx83/Q9Ih6j+LW3E0NFAPbitK3GdXUzLZ0vNOPr+lYOuCTS/rDXtW0Pp9p6B
I3IaddjhTIrS7lJ4Nbriu9IkmGowE8b4h5oZUU188cuRqzGp9xlCI6VufYFPZmo+
NMGVru+g9lAuLbNDywKduelQQpul/QGTtjYxuvXY4ZoTXBY7ccOGT6Kl3RVGL7ZN
kAkAHnpeXMIDas+4FxjWS2lgU30lKNDf332ZjCQZKwkh3R6YiSdmsrfU5wsxDMgH
6TApJQPS5di92k0VY5861JxbY3qZvrBzbRQJwvVr0IbnF/Z/WnO6wq4bXXGIosj9
LYxmgoBgZfn0ztRKYsH2NOGjqVT9QRZw0tAuw0wVFkcNBR0EL3hhDq0HcikcAyiF
3W88fmEj9A60P3PZ3mSXbJEMdnfqDGPz3kt6XOqrTeTM+xja4hvO4KpfuWf1jglv
o567q9/q7xQ0S1fz0SBnPCJJlvxijAvyCUKB6e7LfBzIY1bbOnSyqJx7Lte32a6g
eRbKUNaSn7IZYFCOpOsLFFhkMIsmatGRfUs4TCylXLlhh3cgcAvJ//I2oifeCB+Z
SLierekFGRZCsH4fslHQUqz5zdPvpSTW8Q7JLzeqG0t5dU8wMjBAvpfRtlCVnvk3
d1qiJla6Qg+FnBBw5D4Ym0FoLrXvsaoejh/qbkGi9lJTjTOue3wUr8Yj8sdmLZdA
aqSk5pIK1orCdE6rBqiTTcXpP7Fve5hKA2oWrJUNii7fp7jEsNGgGvK76UofzrNE
sEUKFEq9OZlhtrSXstTaVuZzjl/qmN/9i0PGz+u4/JG7yPnlxIAcbmBD4XsBigXI
48gczLQwH6U/Yoa+bNebpnA6xIeMCE5ZoTxCwaHMlGwlfUp2hMzqheZpeiYljS2n
RiKI+a7ExJmCWAS8ppD4+tj63mNT2/W1ehbbFw3m4vZ7DaH8i5BX/LmXD7M3+5g2
CrrJYYBnckrsl4hq5IQlOU/s3RKpXv+/hJ4nJ0i7L/Vzat+Aj+IQb4ibS7nbOPSM
qgFqKRNXciOVwqEZQLxH3KO9XnkzmLR91zvujzc1RbPEilmNFmwcjsaNOpCSR+6z
kuKUvBtL/yZUbzqbykE+wM6RxL6FcCRyibKUUseO3NsgZLpUnPGS7yNjJVEAYTrl
YX3gUFarVuT0PBvQ4nUHWGKFeur9GJbexh7yuJaW1WMdC333WM+034dm5o6noVfd
4U3oR/id4NjiDvZsYWCzHzr/1oMp/i12NL7Nk5pHqaKuUk+X+ZZZTA1ouzk01H1q
2uX9ApoWH4pYSWQfpoWjT8JiUt+eK4FYD2aq1hNp/N2utX7BBthA9KPG+YHxmB5x
4g46Ltjee3L/Yn/9pexTDtHkL0myv6tN4qCF9YOUCYFqJ/HywppHXVUFXrofXxJ0
vx6/wRRoS7zLTNiDzzBZzp0iACYCZA50uhQAnPeRO6i+wYlS5jJ4/eKRTZUfmXnm
iwLBIyi19jJNli6r8xHDUt6xT/9K0XXJCuliUORtPW1kjGRcxXdGEpyQnamGLLK1
hQnlujhlrGfcbsin0CSatTDp+Q/EUD2ZJDhA2XCXwGwNx0XSSYvszNUuBO/AYz3w
+JT3CbL9DvqoMBW/5J6jlXtyK+fzrq1d+pOkD8kczcEcNSXaj4Gox1cftj37kOgF
nIyI4YJexHDpzRdoGWODAMpnNR1sZd7+655xQYI5j2iamJLwE8MT2Mjvp2t/Rxxu
7Tsc8tCWMdN0dN/9TGhX8Uwbqa5Q3d9mKuGyG2AqrSfE89/Ov8gyGqKE52k7A3dA
usgW1kk5ogbQX01prY6g4BjbqV36Z4YhuSuJ4Qc9yWfEIDFxSTcsraoiklS2R46F
esWck9f6ZjlH5MEQB3lX/XKa8s+q/EMqnOu7GinSbnsxHUZAkVwbwqi8UE2skZ48
6p5ne2dYlHHQopvM42h41tQIt8aoHKWfieLLqsR0SE9elRl3rkmXz1skIfK0hOKk
4Lw/HrriPsiqMVjzUNPYOeK0KmBpm4TqIajp//5SNLMbnkEXYQntVygUMSJLj/6N
SySiZGdLjdgngffvEjhUAoz1Ttftk5vEtd/YU5qEMWd3QebyB1r59PJSnPhszqUl
oDtD18XxzIiJyELjORPxYdxqmbHmP4pz7ICJNQlMNpfGrOT//x9qHbIIGRa08Uvr
t0t5hu1eCTPI/QTtd7Hrxaixer6qiTIPBKNHz0Xyiu0yWqt3uxu2w4fZjj/MoQj5
LVEECT6kqjd03dzrJrMN6O693mhG19UnGtqsuYpXfKaGyzrecRoTq3R+hSgHhp4B
sF+7VvOmmo3nTz+ncrbJV4CWkg1JoVDHDo4CTWO6eFuMoOfdyyq0x2DZqLUKdo9B
1Oly0nzvcx7gFg0u5l1tdF59JcYL+c+Ahiz8HCmk2tFzVx54rTGNgS+QoJRwYWbv
SFZfHhP2klxNq1Hpck0nB2lhk7IQJ5bP56V3AlsYUcG7rnCyOu/UdG27bhkwlM9a
qaEhkSfARGMQxq/3b/NVJ+W9f8X2GLqtPsEvsMiM9E/qekfXOBcNV0eSqqBLRzAp
OX2vNl53QQDF4VPmEaTYQjgc4Jcg7POXC1RNuXQg/tfXMat0NWcQxVoJlrvq1ws7
1wYR0USZfw+KG89hLIIM9lUz/V35JgNvSOLR1P8B1py2KLF8FwuU0FdB7X9rJQX9
YJ8YcxgdsOS/PBz5WA015th7DOTDi/I5i5YHO6v1O87GHBCnRc6QNvtGOTYe27Ni
QetpkZKU3NNbH+EA19imCcoifB1HkJiE8/HBvB08d+kvZJfPc/1p/pR4AlQDU+aG
/usXCepior/cjuHRQB5vo91cNTzpNvGiP/kDQF6PwLe1TNUxC1dY5ffapOIfl6WF
+m6Chd9fok8cnXTXAGjVVqmDiC6zRQdEr3D59XeqDiZb2GZi+h68Lt4Z0KLSxvzS
XeJysU6JdpckIo815kGAyU7tnWZR3lHJvb5Z3tTYjxRw9Q06bcxO7+DC9VFHmOR1
UxKwsAinVmaWC7ASpssOJvs9fPHkTDM+UM+UU6vt6eW4ce9v1p9TNDweU9vxfDfi
Svrt5IOCVHJ0qG9h2ntNiGK+wlFCpbE1MNr6Cr4OeTDtLoNET211ZKC2cfQtsVKT
G/l77qRzIVTGNDN+vPJOO1hilMJNVsLuYbqAXzbPyA95M3/PTf4MS4a6E/Bz+2iX
TfPAFsjLLjwPfskvWjVrvAcWRq5LF4641uPBxaOHJ2/3EOxSdUW5NfVrckH6Fp/y
ikBEawuO6G8Te9zry51E74sNhT0eGEEal+Ufshum/W8sX+dEzDWzi+qXrUGfZAz6
1kU+WIBDHjkDRKC1U1iRg3UPyMr6korw+i8j8gi1KRUubne1unZnAagPSizoUpWF
JxmHhKZVDLkpbDW0fGFdhxwUTknjDsuxuWW3w/kn8tHNPaerlQEpLZ2vU20U4vUn
TQTqoZLjsobPHpx47OuW7+GJDF+XoQubvw6wVpLZ6SK3B0/HnayOsTjuh2gnJvKX
7e9eM3yvoCAoXWKJyoBMwbLEvyGncbobjOZlX0iXQ8LEkh1K0hGLEMtc/MtLzIyf
Cg1l7oyfW00kExqIsQz2qnEAC52OuSyy2zM90H7S4AN9fMsLRqYLsQx0xS+GYSct
xwD3d+XLQWl1Q8SAQvpVlsceSImX50bRNK0gYhilNPcK/aDhTlUS/KdKOhckEwAe
9mLhdEM80mOK8Z8FnCUnN0HB6v5d6RUdgxPWLpLgGVY+8QKS3A1MinAhHpNgyaW5
uGy6GuwfQYsV4U2E2/TW5FalmFfgGfJ0/V+TL9c29K1iZ8M9b36+RS5mZkLuQS1K
H6U/myNZPQr7dr4LwKdQ+U2ZRmqDGGgM0MH4Um11G8GBQsUp6fluQ8uublHqIx2W
U/HLj5djWy4MGe+iaAKyoYSxUdHRamSGYTVpD+3w7O5go63skSF61X6dkhYm3Rii
Lpks6NVmjQbVrrrthj89V4zOcQTZHh7AWt3XkZWDh2Tbw9h/BWAbaMl29y1HAmpZ
quUREaHWO1xChgii2dLuh6Ekm94YpuP8Jw7VyCWQxRuVrSHNK9t6OAO7mjiFdQGW
2AmJY7cZtSrZ93x05343zG11LQr0D/pMRiKeVhLYP4wbAdNQ0RGqXFZ8OauzBDhC
cXkuneA6cP/e2DbHitAx9+t3iBEIfFRjcd8Zr+c4+iYCTXhVoc/UUt5XkvikPHgS
e8otxiITNLZQ3lzrIF7Gz+8G+zVmx/5KYaM6kXcmyn9aiyqbgUVfCc/cJc4zdJlY
tt8brFoElaHl5SFMBZUt4RjW91qCH3EFBTze0xwIazvDHL7USGZVZWjnOa+vOWVd
0mGeyTWPa6RSjSAeBLR+NKxkpW7ZhHB6foKYQzJZ8drIJpIyTmK7s/CsLrHCdFx+
/7z1XVBgLvkfLRPc8P42Zzzud9jUuXghgaJyI6Wk1NwgnFMtNL+MHX6ps0eXStEs
cgYtdM8laWflYXBFkfFxpqV9Dmvw71TQAjilhruFlv5FFzhyZ7Cb13vtOlP+i/y8
+CsKdzB5oKbE0BzaeC/Zbdy2eWaFTnqymZ6bJPMq3AioNCTssKOeBV1afnUG3vwc
uM16OzYzpTGO5YWROdNv1ri49sUdOnhLEXjK5CbV4z6EP7r/Q1JFoClUQoC0RgrS
G97Jtir54DMd6H1svIpk6GTUgnbolB9YN3t8CiguD6zYN+g3g+S3Vx4z9V8IK4JB
Mb/UzU2y4U+Jpvbx06LCYqHIIEQwFeccRrNCa9QCuCTkDvhpi326TZxVkF5R4l9F
TY/g2OfzN3Ts0FepklOkZHBE2CUxr1efVNXSyqY4FWuzrKofILFq79cFEJwHwWri
oEgYrjUTyHINzBRaVqkWzQkRGYYxes/wp1V/0Www10giGX+9NkUPufWgWmIyoxWu
MYYVivDyq6vTwgyzILMydevPj6RsDKa84bVPJvPRU1uYDTzmB5vWXW24kuMsjNGd
U3ZZSxY/+gaqP5McSRy5R0shcmEjLhRWxqBz/qy3W+QiUHlTxe/3Avjw9+ZLw1J9
UgC4HVewLoD2rIrQFSdOla5g04m7pCJ/D4EMFMQqvO5iW0NLctLO0nezGZIGfcfW
DDFbtMTKCM2XH5fzgk5RrrjFfTkvsbHqaFEHvKyVm/s3fUpJFgdZfDBK+j9oqtsv
M2UTSaoOw9yGmBmTj9jzZh/6u8W61vylg2+k5mYJbNPlg/Usp8N5zrXDIRThPTMy
ERncJ3rEsGgqsoRw54cSgbBeu85BFvcJymV3j+wTkKCMre8+fJUihFMORwGoFWKM
bwjfLHuTaUJOt+EiBnaAjB+kKPwInWUweppWhZJ/5vblaKoKo5i0d2zufTKn1RsD
W3oOLDI7uMFfDEwslxTi39HZ1EzSuExKkQNY7+lJVFzTbly0/1xxPte6UWCgCF68
jJtEmYId8L8f2sHbziAsTx60jubsd3RTuIWsZLj5XDAX10k1QpiJKFU8eK6xED/1
Qu3GL7u/fYRUzZpr68DWQS+mpKAOPPPNlrV1Y34tfYpma6bI60D2zs2lPtWATbGW
nHh7tOmN3Rc0hQIS8psaKo4uP6oi/DFI0b8qkpp0tFwJ9jBYvvW/fODF/rH8zrMq
maPJdDEfkhDw6nL7oqhfCrWKqSMeXnZY16BgsdLKkiOLa+ch3TOOhsyDrZl8brOh
rbGIVo6zK6r7P6ZnSIQFKHF5AwVrbjQMQ9U314qG3/htMWhHiX949l0PKGnZ0JIv
eHZAHfu0NacrIUPu5dINxqjaXtAb4rX2sCP5X8yVhcWuB+ZwBfPTRLFSgfEatQNK
1Ag3Jk8BHuZv1IQbGOTX8DouLfUkb7meA20fdr4k3aHNTIu46Xk0FfGTNK0pGkjr
hB3IidRXBTwdLXsiZ57LnPs7t+U8XFn6V17fPnJt3AJx/htbueXCQH8yfwFR5OiJ
aecqSju93muNC3GRQJDynLQ3hRA1qBeVbE2/4U1sQRmn+pOD6VdBH8y/mOmEfHup
QD57/tNnGuoENY0qOgGa5Ozco0oD6sT5zCfCBlrJQY9UswopbbWA6q20HwS8oOiV
Ubi0VO/VpF17zp/VsZQ403dL4pISmnbEoIlqglBQYLd+RX5oz9bzRLn988I/qeWQ
Sgwx4w+4JI0OKNs54r2242+KnMqjROnn6LJRKiHyGXWnb+emcvEo74V6sFLrk/F7
VnA4o8YWXy58v/J5128HI5yRvQwmRUW+vis2qrVU506ZmixiaNU+yQ532tNQ5+9i
pJPsGPFEtDuSMseL/8QrL0+mq8ZBAsetSm+EN8nhEWvoFEntwARJEv2/4CGooXs7
A+WcJ718NSA2rEEuAjqN0wqymgvL950oC2AU52fx3tIfQSjGN9mqX58uG/B/JsiK
EKIEwDhLkttSIVo245FUUq8cP0LJ4jK3JUH8AeTQOPaH4SNT9OUA4wJGpaWNrzk6
IMU02qlaZUwUvgtJRnyQWAUD65D1gwWo9byiwRltqima7CE48ys/RzaWYHQhTmXj
4EO5KFhk4ZhEKHAk1p2BclqEthO90GC7/hfhnEovlYj83xoVIAcjPhf24w57qzeQ
RmtMBezwjv7doYr6k861IgJUkN4ibp3jxy5EszRncraBe163Z1tnUxt3RwSdXapU
ZwZOcIv8+z1YHT1M/Aq23sp5gXv0niQOg44uOS+PDvJPQGAzIid1MRG4u8zzH92B
bIqbtkft0iAoyvb37rSzsNdgpQ1F47LOZHtqnefpysWR4FDeUttlYcZjw1Jr1EP9
DvshH+FlbRACmAtNibkuu0g5XdIFxN0K37mEhhj62dt0+8wF7j4crs/ierIj4Fe8
e4dycDfohwW+z5EsR2j+Uchk3ZevRlmhcjphyFh2AAJjOvLJjbwvJf0t9gQF2FgW
EblFu9ZoPl+6m/l5/Py+OXkqFsofbKOdL/UBPyaN9qbmBlJiWPXKWjUdEYietS+N
K6EXGZDsEMzWO44IfNbdrhmaTgLVySzCylhxLgJC9Y8mZ8va7CQEdivZkWLAHRBD
xkRPCC9kv0Ic3z1Qu9O7EsjqyK+1Wh9UAih8D4CejPElHC0Jm88pZOqlGtiAcLIg
/khgDijP3i+8qKDPJtR/esxfDdLbMOJb2IxnH+qxUqIauzicXCxsZF1eJT0thpcl
gzyQz6ojvNi9k411BpHH1bJWqL3HmiPUlStilRGBXo3ofKL5Gf7aIj0Y89vJ66lX
zs8TAdCMAEXSFHQgTpfFOxA+7a5IbVJKi3Bxad0zJK9tY8EYWJxWubazWKEDEufv
glt7AfcDjPhCIP/tkU/8LQ/ocGCueM9QInrpZmyWFRXS5hkbqu8sLeSJMN3KGScq
31iLDRDls8tkBp7LK/Z1FkS3cdGzgc93ooIrDz8rVqGEmzfNlB6zvI3TQYgSmQTM
CDBV/Ma/otlnsJEKWExUuEG15x7rSl4LTOYJAAK0XNLqloOc05F2ruxce5qwYN1H
+5OyI1vOrgTenN15LN8Jq3HxMKAnF524IYNe2EOwDbaDCJpqC6roU6jIZlcLi7VM
SOsOEPQQlHjpizRmrAu4T2XjNFUYX6MPd7Pu4sgiFYJ/LliPVlDhoNoCrrNZ4VuT
s+oXv297gnzKi2jvs+PpXxBDkkRPAV3EPJbwmo8RV9Cwda1jo+poW34RyL3nOfUR
igs/6eEy4ptBM6FoYEqS+R7r7VPMvxuBQrZr7oO45xGvNFeJyl70nDgzu1QriAqq
upnaiCfhBW3hDfgvSdfmlywTC5UjqkDaQfCynLCjtdnB9JeG6JkzxCrSAUVNr+XJ
4NHVjQk4lg5yp1KloPdg3d66nykyyquJyoOxLUmevupohskIaduwDng9haMu4j17
K+djuBXV7BGaBitrEH/3Wfwym55sgovb9JH/NBAdrcLwv4xPlGQ8sLZlb6A3DB+P
JdIXPQ2OoCE/+ji6MKtERbRsGrO7UYCg+KsWqTkqpd97YM6Gf67lkK4/tPhTO497
rYAotRGP306nrzTU7jiIKHLKJQnFwIlQIYsbqLD3W0hCVXpzgLb/TXNGtl1tRaTM
oIeh3whKvbsBXZRQy7TmAzZJ91E3fto/sKR5vBgDjpRY/LyJzf+KSmzzxSC47wlI
VtevkAZCn07sr/h8CFGjgUN3vhFlsTRd/1JKgYEFVbFKlPsBaU4/qShph5ZOFcmp
usz9VQxQZjYpnq/W7P+1G+MbeRe5u1/n92xNgryvCuHuTWiB9E3B5pKzO+JEL566
ruIVQ+/bF3h+4qGM8ryexY49X5OR8/TRE0CUSU3nlncJGimuXmGPStJ1n+uZ07pu
mYhUiDrdCN1ocN9wrfjAs1I61XILktTi064K1pOlcroRn5zOflRzFv6gyXyFXMbU
8u4+5ZxWj1n524I8cw4lRArkY3KPWY83+rOWHdmN6S7q5SfbyzdTiPGJM583rDgS
PBRhYr6V7/H7cYwuMetEQeYO5aR4pLxqML7xfnMaJQa49OeSBYDH3ieTjqFIupUG
VHMs/LGNnsypiWm/JI4TOXK5xlTDDmXzbUgGp2tCXcAzpEdPSTOEaKRBMoFWE7GC
IKTutPaWY91OcVw2+MmyjChJd4UZnRl89o8jtY66KZn6vTEpoCaZK4/6zf0TPFT0
tESMX9mudrxNDgu+rQLedKZ5aBBNkrpnssUdd5Fjf/+hWbh/lZQvXB6IOPv2WIYX
PiKoVPtkcFzYhzZgM2JftJ8bB11Be//Vr7U2JFbfK2DN0lRDIXMEOH4N/rBnIPtC
DpKBB23W1Ga3+iPkmLpnkbLezJBTOHbPaStbDwh1FGumVoP2/ZJbnIW9a2ff/5SK
f1YmliI9/XZRrm/l3hD4zqwWP9CgINuF2o0CUJ39adwYFtSWG1TIHX9uWrMVB5v2
RHsHRmU8v0KTVtpsbAysRmzTDCixYHE8KSqpmnhP3ynUWbIwBxu2Gmtp3aN2hkti
wIoxKP9ecIhZ9vWuIpsmmmr9AxMiIN9PQjZsr5ahYFpO7Tam3vsQR16fGcskogYU
V3CZISkURK4uGrFLzfwInXE/xVwblGZYUYAsxx4xPqtQyNEpuWDJhx2AV6sPTmQH
XpNPxxDT8iYCJvigFYE8mzrJec9MVOF4MKLTkHx9W6SBOe3+FmUT28qZfntrr1eh
ko9Sthfvsal9OOHHMI2kkUnDXXxOJffiLW3njpWyavQgi0FZyX8a2g+B5gWcui52
ZyMlMvSeMSZVLh4bk41aADRbOAM7H7PhCwdSMDFkxKzTVUS75YDPmOYoPgV1TTnH
yRgZdVbSWzYuhUNdqUuP8JXTtuo2jnffKXCDCgh64Y800qAKrINKu5pVHw9jiMW1
gxgOH+khzzgebktGHfaMLof9kgeEVdlISgjzhYZUOIHHlPV9adZ4B1XqTTJm8gK3
YMpod2G/naMbHOiPxBBn1DkmowNKGNGADjsQDTBg6UtuJ1dNMDJtUWn1PXpwS81a
sqcjWYcfTfs7HAEZ4FAJ7EDgcd42pegTdKnBtA5G46lsQC/xjvLMaxz2qQInaxEf
TcBPJ+kXyF+IgrWmbtP4AWhcy9J5nTz9VAi2HJeZptW3v30UpwzAgI0lkdCN6/Gu
odwOcoL/CgZbUdYmwNf8C9sOkseKH39ieaWW6ryXvFb+QPGjgLPebJjCkhYv+PaM
hAHAQDuYkMNl3HqongaoSyuYNmfdTdqUYl293zoRZ9H1FjnH7Wi+glO4vZ/K9BzX
jFbhmZsnu8RVTV2NS9ESz0mGQoLzttf60NbJWci0UuiC1aMKJv/fv2NqJ83uomaB
kxNCHtYJf97b7BKzyj07oO8GClQVKPe3dI6dic6c+vI6p6jbK4Ocn4oOhMPyGSq7
rygJytozLr4WbIWhunZyVcCUioRgdg3sXfCgW+pNUqjdHbcLCd7yr1QAFJFAiWSr
0WYd7pfp8zkp8I2VgJW84h4BbLIACJd6kdNst+zL+hmaeyrLKaGY/tsGBchi27Ou
zsLr5vFxx49MMAqFrRlUxlaPQuHVqA4uVszbtNn+Or3SlybFSI18GobRCjefAFT9
f488ZUy4FOtIhrI0iNy38qe1ONq9F6Zpy6jwXieVu5RMc9iYV1E6839HehPzsqZW
1PeLJJgMV0/xP81BOQvtQV9Io8uzr1jrjGrEcMMiMZzY/SX9bjxGQYyuVrKk71uv
QCCFkyyTD3bIfKFg+zdWFzj/goPT6nMQeBmgiwOjWJzkqRVDmVNf6/b3wDkNDJ43
YZNzJpD5uy3Cmgm3z1Iy2JFk/1C2y5c/uCTbzmRb8CvCjULspP5DgNNZlTba0jd6
EscT0qu+A/MrwPIyHFBO9+20qNbWy0TCfYPhQ7s+9vviIT8nSWqGpht6fv6lih6j
wmtAi6KzWBOAsIudgdVZCzXVWWDtuLoLFh0a72Iiv5XHg7r+ViaVwFlpYI37ciHX
EF2AfW9cT6moAN+YepJU+7nnJB9cG8x0oS4NMAP9xl5dq0WtPEbEhvugXwwCz5lK
dahP72ZvHvx4aoso/JZDc3p2BOCOkb7fPuQ9+sisc4hVbJ78xpLUK8kBlnOUJ5A1
sfz0c8ArFDNZf+higr7h2x2ZJTMdRM5GCW9iRwpGln2EpLNtkjc6q9FwPfrWbt9y
ZmvbaaKgnpB1/54sUs+y5KJr61dBg0nUBGEAoHmPIY1fyN06RmKonlRbEVcTCHQ7
vaXqMoBsL1dFEtwDukThBkJEU5BErjNgKvMhjP4unla7vQqRjAhiNK6kL8DHOsyO
SFmE1iSOyb57Ol6LU3Sa2cbtImZdq84aXeW+jKT0vLIuw7vOqmv7685qNSW7U3QN
rKnHSK9rHh/Vq6c+37RVflyLCH1QSZJvhW80K93oYYgQUgEX6ziJUvLPIu4RUX1e
uHrZAwCmjeGLLHHOcHUO2FmdK08Qa8DDvaXtrsyrMeCjlKUr+n5x95kQkEjoHXUB
Bi5PBLOynE1TYOzK8PwKz8dl6D/1AG40ZuV1fhxTyRKdsqUmsBOrhcjuWcx52C/U
ixkhqcvPK+z7M2g5SDDkhs+OPH24jaPctlhstL5Oj/GsJ5tkjMp4u2rgcB0MggTd
uHZ4XTOWrrNvw3q05ftSviHAg0tP6IHCHOAWSVhuJAES7FJDuvt2ZUOa5b4q7W42
CpWCzAkE4pKulG1+DF2lIiK0BN6G8qqDrEUv6B617hjUcxeJCopmdydKYGJpT3OE
qktL9jWpfn1e5DLFu9Wse3aebBha5VJumCaHy7AfRElPC0QnuzUZxotc6tbbPreB
kdrJ1XsF6W7Xoi2yNlN3BiM6RcIaj1gDPZ5uXKAxfE+pFf54ixS2t6xgtouAKYUp
LfhSo2QVhK0YylARsFg6bVdQcRFNs8w7uPuvw7av+Z9sY12WS9EfiBuKumZYtcJt
ktr1eG+LYlEgrBfjvuea+/PVe9sRu6xFFJyt3HhChTnLpd9RuxYrcXwR1HiLQlco
MzpK9sA+N8SIWLctLUqT0eVJQ/Jif93Ync2pQK8Qu8YEzH7GnmvrS5lYeYPwdSUi
6ImNglQOowuGA9d7QExy+JpmQAZajSinEh+LnOBsRPJ/dSJNsQxhoSABgIlW/Snt
v+1geDqKW6lCkMe5/jvl1WKCyoZCSBcoeF7XxosfSeV93JT7ukk71cq8r/sQAqR4
Bit2/YX001dtRtrNcZzHsdEZakOB21hUuPw1SFIPI6Ge2V+p1BjOBE+OuGXB5+dW
qdAmTduN1C6d4ilKKAHt4JgB6U1UW5+S6kxfh2ZFsj79vkuT9x/CuzUmUzGKG+JG
+PzBFc/cy8yn5kS4e7u/geoDelvTULzotP16ZdhWX3ivPPcWnBlIJHka83+0Yn1Q
/lIzu1RX5LMjbB7i+HK74HHT8Xbkbnqu+7f39mRLpAJN/CL1fpP3Yc4wGIamLATi
nChShDzp2JaGbOp70l9+E/tlle2XRfsVu0vaghUbyr09uVKc34llo7HNNm9APQlR
+2OZkw/bcXEW9EMvvYF60QDwgVerJYRZpcAyr+2D0iqwGhhpNduS/2q4J3uRiZgo
jUACEUv41imbAegR13ZLLoTW3+CEg6MZlxD1mBiV/LhGab0EdGn2wQkAN9G4q8o5
eCL500tfDR050xytTgm9c9o0Qpz2lvuNroQNUjwLj6Su5r6+jMROT2HudFCXFvTm
ApvCiNoDei2sNoHtydElEF7yYJIptuDJsPJKJp0EA9fWwn9HFze7kSvJ4mcRJbqN
0fvxjtE9Gku+nJGFtOZAO18KoADvnMiSQexNdY4q1R91n0jAf2PGzR9NuEAmDaHM
7Zv4IPMOqypJK++fiauXybED5NC0v0bjuk8Jtjow8oy32k94oD8uqrLeIqUuH5GJ
TrK3uA3Y8H/IDHua2wx+JZNqLAdOjMuve/feBoCFoVm/TQypA63cVxGp5Y0njcym
vMXNwQjKWXbCb34ljxJFyLskdPFMs96pkJMoPhsY0oc0/6wpAkFgPTWPhvtNYHH8
RkPcaiKfGjuCxWR6PuBMnK0eyuk/scdL/q8+MHRjQZHDiuCjW7wAECiZZPTkI3Jq
x4MYW322t/hfTNhcemHNu7oHLoqlokqsOf+2+ekv0ViSfBuHDkPgs/hr6rb00+NO
9Ex6TCALcrieI6HCjwBk3ngl8+bC41JdWClrEz7yTCdZdI1K+jSDeoKipFCBZoj3
QguOfvq3e+opi7NsIxho4VBi85bGUxZeADoomlI+mAQyYtB75YQLU7G2p6mK69QQ
4zbt2mQbzogsh/sWpMMygsXVLJYhE9VUfY/9VRxLtxSwQtZ4l/e2ZmngV+T1a58q
8ILeqhDidfrLuV7F8LXfcTlHUIJfG1oDg3236vTOEtkcKA7JEvxlpZIh4s+XSicg
z+4D7BM5U0BfSAk3ZcmXWLlRzgVryM3tlbd3QuYsQ1KTnF9+rM6/D0WfojOMZki3
GnTwImSri8q0ZzKeVHWh5R5Tyfl0qoZpCaBBF0phKWAVKSVHi8JTKXyikJHCr9xO
1ka0iqiro8TQRN4heiFe9Co5FJHWTyC+Di0+eEmNMCiib8KijkBBjtfDsiNaSqCC
1xEpEFbw2zs3y/9XC27/KUNBiEt+H7CwP1Bwtqx6lAIvzXZ4qwwn4ZsRxpBbCWBI
qYL+AIYAyilgZov/cIYM44pIrGJWiJznuESnjaYcfzrrqny4W/Zw5ioGp1Zi1XfD
XwHKweV804WY6pi0I5YrFD/mrhmmV4X2x3B5TolSxr/fz1tf0la3y4+UkolohqYf
OaehS2hv6Q7rkNqMxOby8dmNzxDFh4a2vWGwLYxONNQLY4dYC1H13HXvx4m4XNyH
hJz73oLjPRkGG8Klsj9jONVPSRLzkDYMbWrtTY5CgNGyLxm1oS5WcXVasAc5/Goe
xWIPIQeilvZRA+T0HkAJx2ORyMH8OR/XhaNv7KdiG+EZEutJReUpoHvYAd22shyn
EPUhc1OzJRnvgGgIKJ8Q8OKhmhx6XeENVG5fdMSKbe3y0C8mFyQoTRk+5LROEesh
hFYomrgZ9Y+PBsftvfECb+Yn4AbS+njEnDWuiSonOQQu03ZZW0Maus/v3vtbRl+m
8kOWHXXdzGv+5ZB43MB2RjtR3hEImfh2ccxXQuc0YQVKMK16kxXIq/JTVMH0yL4y
kAJ/mW7ZDUgA1u+w1uWgpF65jkmbxx6+Fm8QC1wCe22nwvaMGWKR+pCESRvN3GF7
M+fYnyciYLsbzgmJxwEaxy0956XXRsbfNii9+XBwOVUEbpL+GdCWV9xKemkQcMCX
9DCAyivfw4Zs7UM8Ecp/mou+1pHsFUqBfTyQq6WV9j1ELq8NpXgCr2UqMmu9KLHp
iuAjTfs3GfXVNhcn402W0tey/7STdRLpSHfVJnZiHiezKm7h5YGqTSQ63J/r2TpP
1SwTiqgQwrFHCXaw3ClVbfFb+otsE/Au3J9oicEonXzDSRG+lPlPU2vN94Kn27Fa
nlARS59SMgEmAeYzJSO2BpiD0d+Ck542TSzxNAnWcy3mh9+EqifTTYTddLwchR4S
skS7WgcRCb628lHwZbRNHOHXhCBCtkJtLJEokTMwuIv1qDaKB3kYHqUgHvpnVEOX
K5tBniA3eiLXXYcQg9JX9zsA4qoYGu5sOdcqvlaGaooqvI2kbipH5vipqflePfYE
ywCESK6i0EF8cr4g5YSU+he4mPF0bxJ43xFTBHXqlRnH4cWRD7CyUwIZF+iL0nMb
LIEZOO0zRj+by9DUK02BV/XTV64mn6GQuMBq8EKZIohqwvvx1xA46xwtedoUBRvr
DAib5yYapkMawsZUEUJe5ABTweLLn2EP9YciVAcG9wKl7vBv/gGLckSwLRtYdNwa
pnJvAG/op+ErVpAb+L6mkGhTTRJW6LRzU7eL/6KQvcVZvgCACBsjuDMLsFhDA0uh
PDY9BPmDfddyhniv13iaPB1bzDwk6bgeqQj5UKrcJ8WLfYAng2IlgYz6+PpVkLm8
r04KuWBz9sAB50fkREAcwEP/UsIspqW0ljjCrPJ/pBPRDIxc7pXQmNBAxX9+6ZDV
kLH9Gytv77lGvboFRGD1N2S96bdkRH5ft9QveVo3epQZ8N0fIzOKbj7/QGKDpcRr
8MSXbPFEy+UxFXhznbKIgrb7sI+vI3LURNG42fIzvRvk49fdeAghbOxJoTRVlM46
G57bT3DYPfO6inFELpvEubYwmxiQ2qnebZ0L3hvuyxewBfgcf8GlUMPNlDhdmcYV
cIJnK1W5cKkdx3D8QJ0yPnHQd09Qc4ecWx1b2IJl8CH3XwllYOQ0+5SJHWXrje/X
P3k5+a5EIwuC6pUQLge7LV+qCNDkDdkRqB5qqpa1I/y17CtCJDyL54TgAwQQe6lQ
ohc2RYFT+uWARoL1GhInA7VFb4nytZGrl7ZdCNaBKq1BgfRL2EFZJ2Fu0N1GcbKt
rGdz/PnR6j9e3ufazifDcWRfv8PEQDzeHtRffeDzZe1CWnKWwfsEGITBkdr/8RR/
Q+wq6C21U1WG2jBqQ3xNBpVb4ljT3/GLwspTzUgPXJksUzkPR6ivT4THcmdf/dYr
2itO2vKQUACC1nl014XmhL4J4JXDragQX4dY3/Vtwl0w8ehqK+9IRrHTP7lZY5jL
6RRKAES7SJXJTgsarJGNKBDIDPNMVXosMnX1UxL2Uyzekb54aUf1Sf7oMnmP03xx
SIxKpzZYmAgx3YtbUcXonCY5zMxQ7naYtTT+aNB3ILOJcW/RmFNW+dC5V4lJVNe+
/A6VRh3rTHsJ+4nR2TkTUIm6fbIUVB8MFmNwnKd2Bi2hdYJUHh9YIPiLCx2kFmFR
qRPmNNk2DOcIQBK4LI8iFiKlcN4W84PuCn2JnURn/aXCat80t/15FbrxlpLU/GDK
DxkLI/vy6zFR6zoBVxdJOEeaZJWAYNuWsDmJgCgbEJuzPujnAvVXqV3161CGXwDH
y7mQNQCOklgNyJzW+TTqeDL26qVde7CtABzZDDFGIlQh2nmT4ZMNOMBlR4w6SiEe
Hoour29MmUyuU4wxQRYWxoMNVK+LdKHGYuJSpcKwMB4rOC2AGEB5MiWWD5g12OsP
mUkraPnzvP1LKWLImlgd2Vo8+5ClGWNLyjUncCFWxq8lWBITYObj6m174VW+oDa9
pl7zohXzXXK2Ejm/AnUSGXYtFI+xH9gSGYoY1t5k7HtfPl5hapDlwoAC2so2OAME
jcVXlsRlF/3n/nAxu2FfYaJmZ19MUMq/zLTLlwgXD5J/DaVp8SgpoEYS6CEoOY6r
ebXISQL7EnRfhkDxTuM8rWADtJxwWW7FISeYNfIOb/JcUIXrFAL7DNtLVaO8pszN
/CgPTJRaF+VZaiibQM1eKiTrpiZEgjSRuvK0Kmo5yAC3S039EB4cgyXAwBvLwX+s
WEOqmqo8nfyMwqIyAwxAwGWo3wRc04FzR3KQMHYYejUODNiyvNlJ3xkKAlCCfOkr
oSDRb/jyqmjnONjMrekj5qlO6VtLRdYnvdcW8M1ivyHvz/9OXZELfgta1ZNrp9Z+
m1Z47/fMqytZDAujDACmzayknDCSV0YafBt/5wGG8NVRyAyh0l7PR8b7nhgWFGlD
ZrJoCWRCj67Wcm1LHtSswUBfeBnyT/IPwRI2azjCCM132l/qkUmHBKcdGtwH2tRA
odQ0Nx4idX6zmoBcy3Rf98kzNywOC7/3xpq69I83j2VyhuOXci+5Rlbzu15nxmE7
kDuWXZFRjAXT9KlJ1zI5a34fG7LAlQ1yPoV1W6cIRBBQdxZUB6BXFAcANgj8cS4E
i1s7TZ4rzvZ7lblAVxo9mTsHG/EmMbJ/K9b3bgeIlqVXv/RaOJnUDYVWM8h58wbu
YC4rvGZOPQfNJIte9l/8vQv8ebwINzoS+NYV7eO74Mu0MPj/tCxj2zx3rfNoSnAa
hGGkg4Tm15xsMkrr7oGSOFzexqMslF0otXVatqyuvOKqJ/fkhDbYDnGoQeR/+5E6
Utma/xbSVUsadRJXKPVbHM+6Gm+BfPUzq3fvXIquhSY57h1KQdjQ8YieWuT+UNls
+Im/LkoT4YRDQLMGm/t8KAkI/QbDPMwA9dcw2MmFCi7uK+VhSo0jpROsxKVKlVUE
A8TVvdixUBQaZ1OHY7ZgzKvEmimdUZgm4bjTFm/oHEziLZ57ibmX5pPeRBJlvKYT
uYVX3aZoPBoLotpIkhVArXpNqRb9aANjP2xiBD3/H7Nq8ft5wG+O9Al8g6TvaLHY
c69+W+cplDSCOPrPgA2q3v0UT5DX6zi2KMJersLnKVTi7VzPuAutotj3//rytIMD
pxNet3q7TjxMVs3plkhu4kTuvO79O/wyODrX5qbsG24iFf44OcBAnDuGT7J1RjOV
JF8i9x8bfHsyYNCZoVfhvEnSrOdEm/++WrgviFcXVmLpQREJP+StNPZIv43vaVAc
LxkKpbfpA5FkX2b7PNFsOtlKzxb+9hWmsFc7kWUwI7t3nr9kcAkZMD+bWJZE6tHJ
4lmYShiXUpAC57ca3MmBqdngbbWWIO+EUY4xQlnj+xWUkSrPSpPfhI5jR/NoVZnC
TDrWKSeXN9ZRZi5D2yd5v7JdkUGhHGi9yeiVb8r9Aw6A9KPUiIs7y2x+AOX9p61x
3G7fc4Wg8b+dv2ANtl/a4Fj1uYNCDETS1kvi1SQ392olwGM/Pmw4KsV0hZ7rCXbC
lXE0nA9968ZIxMG91lY77UXtWSOgdH/gPsB+32sZwLkjLEA29RoeOaKVjteDc0gv
xwHmGxObmcXoiN9nMFw6VcPM2gCxAjj3TlJ5MuMhuoBaOUl4gtL4MgSVWGnzqIPF
UQoYZNwN5BSc8wDnKKR2jyWljGwr46ZKiQoZtqawgywV98uLo6zsdT5tc/y5yHLa
mR1gqJu6ngBcekLfsdMDfYq+GBI8QpSjt7/yu34FuTRArkxYBn3v8cPW5IE0YzJ9
pk93klUq37MmWNWeCotoRgJPiU4sXA5XYaxNVdWiK+TJXDqMFP61YCObWMwZRE2C
NVUEvGUZ40dsQBgNjb4N+Jrvxv/4k7PFYDfT4dWZsBLG4RTo4Dci+FRietXVoxGc
6nNFMLwrb5BVFwCb9g8yEJV65gokgHXnUZ+Iq7FIAXBn8h7QWKWQCGWWhcMrIpyu
xqYmkzmUzfcH1B+9TAaTbF06ms1hPkor3Dgu+dRF2zwN08jM4rtygz7BuJ0Pot0T
6vQZTdjdEWn8XgW/YWZmetQ/K5OFDtfU69hD9nrnzBtaeI57jyK3IT+vOuMLvqNG
pneslr54ZjpLvPU3uYr4C3lD8NKDdJ0ej2MKLBEmWT0jvbSs7MeUcHjjKZY6zw+g
PFMyKBvFq7YVXawbOiHXBwOx6TSJDxRAqwGXXzFoH3Npsg5v0RBff2ETU0tdXGn/
QdUjlEXc3aUcFvw0H3zizVbLiyRDSgxgyWuDyCGaCLIUiFCpDLjPfbuirZO8Cvp9
WVlxS6c7ch268hmCbGlib8DMgVmQ9/YIsJJLFFAx5mx7cVnK1UB+wanjVOpfH89S
j7oi4D28N826SoAIfxJn5+BKtry4LmxKrFxY+AFvYGBLi5pb7/7pfYPcFUuON5kj
iRtut8PpKOM33Zq5g6l+sYB2z2kMk6dHaEuK8V2IIHEuFktUPzJ2LaPt0VTN1uD9
6mnx2Vz0bXNicAHSbSlNDw7wqtLkgvjTtrwzhQH0Tyz4CRfxBsDwtzXPLfdIaW0M
zF1uNmuWeKtH8xEe1E2w8E5/cA876FawInfbdBWsQv8mLLavpT1Oa/adCw9/kens
g8C7GhgzHGl/sfsJnjyioSWhlrdvH5pItRv0uDjXDjglOZD5qyXIY3fi8MRHIcpf
di1wDfkxxRlsm/XOlABqc1AD4BpgJjXx/HCupY+B4b7KF/nPlg4HvfAvX8TrvT0m
fqlRWPz+3VEjYyUch21A3Xw2X1Spy5c/Y6BwphAq6ZYPx9bMA4OAOvt+rLYookmC
kLkaZ0NO2ACPeNPSPAoKYLv5VGwtowhjJ/Dh1tkofVY0opmDUS6zXiYFwTiqPR5D
M6c2EFXnkgl6SqsAsY2+11vzoIZ9/dc7MOHa/owCfPMEmc9qg9C/Ao/IAT4XNe5j
Pd9DbQSjnXPhROQypzl0J0bJVtPEsnr+EBSMV2Ox4nTudsPOPeHoM+OrGzX5kDZ2
buCXEkb3byU2G33VjtgYsCl1HzQJSJlJbiipnI8S60KWVGgge86Z+wsFxZ4wqeCU
rYMsjNlP83YVtSMAOHKnDfDeI/yF86PaF4xu0uYhfWfFeuCl5y7Z3W7r8gHiwj2y
r8ZIlkVET78TIAaCn8RNMK97R/mfOQN/O36wtKtM6q/JI1CNRu+bAwzinPyJd7wT
sJXbMFp0EUEpE7uBLHTQLnqPVhchRunvK1L/np9svILocgdUJy9jJBAXJq705cGC
jf9e0C8mdFnAu6JkQ+mkzkrRO7ccskY2F3Vq3QXhLlhKd3sxGBQaEC12sIp5vNLC
X6jn2AgOBdk5g04vmDm1ErdStkp3YIF6XFtO0eP//exav/c/Cr/A8F9GLTa9xlG3
5cpIqPMrGqNagseTiMz99vGUShkqi/bakgKYbRm6L+aJUCM9t+9giFo6QUixGUCc
JJysoOqRm44PrAYZwaXDmP5AxbeSYfxNYbM/bnlP9x8H5hLHXaklrZNCti9SW9Or
il8dhbJAPGxjvjYXf8DWBgjdBYnmuPjuLKN1F8poz1Xhho8GyvYMUgOO6JGkDquX
al8fjOfVkNazVW0u5IsdsntpbQbXTo6igLUb4vZ1vScipOq1epkqdRSPGGfOhhYz
tOam0oYt5QaBZQUfG3ggWhhhaGYwRqyAXrnTc1k5DKdwmGtmsUXeXtXFOophQJyj
TuAGq7/OJlLUQ9LndBHS0tnslboZmd5U5KZcI+aDSTnUAUHlKbW8yZ9ItaqThaQ3
qwF5WOuVPuYK7tJRrHFhYi8NFAfUlzxLBX0AH/auOJdO14JhfwdLA1lXzDN+NKrp
dwhyk87xOivrDxmG6hqBZx8jbN66bImzB9GdAOBcY6Ts8+7hua5j6kPTEFU0X9b7
M1szfBGbCNSu9+rLdSrCrqLKNwNdFXfHUwbzkC0wtjBhD5SxJAoWRkYvmCF1UoO+
TGD0hHdXIt511ON9w7XtjXHaQ8l4oKa7XvjnLUbvQKAE1cdF1xf0VRlccqydArR/
YTARRivcYyt3f8AWBEGcngIU2qZcBK4Eeeu0o0EfxmZv14NgIMiIS/9jOVX3NdBn
w52zq5yeOZWl5ds2JHXVPJAyH9qK50SMcdimGPJfzpca/PIyIN8EWgBYuzTThq1e
Eugczs2hKk+eaTMEXVkVmQXi2gT5W05Jut+wj4+XA46jKEwsLxLQcYL/6XbaUyWy
Iq1Koit8pOl/6F1sLbqRPZoLbSjb+wj2EPyF9TXOuhMJ5YarNsAol0KUHTpUccvP
3+jpXrHBxkB0ozFGLnG1pun931DC4TRIYEP8oCmTtFpOXhpPft0Sgx1NUc+WxJLn
6/txqmrgABKRaIcF18DrgArVz5TqjTUCtujgL13w+bRH+2BsGw4n+jdrR2AhIZYS
QnIshAkY3bhFPMfMO1DDiLf58fAynRUSoKFCruEY78Z499xZTZJk98RXLa+B2rX3
Bwx0iIsCUGpzXnCiyvWEB7SjHvEuM2UjX+OjjN5UKNjYspdtr2CL8aSUXoC815aD
+heLBd2I3LihIodwjXypCDVAqrSRPwTgBOD/aeOzzqHnqjqvoHzINFQRMqJHkb6n
ECMNKaBXGiTEcEdKfsaoR5upoxV+dFr+byVt9OJtdbqSTwKCxWgHk0EwJ89FkNz9
CN5Bj7UGI2BfYOyy+tawFHeH+W9wOJABTPg9svmxB0JbxufGG++ve1QTEkX9FaUf
U1Wa/HGEF/Tno98bcXL9E4w83iMlIMQ0rFqEI4ZGpCuRDCjj5BOlikklgZsf5lZU
JG3XiYkorJb88tii3fAsFMJ9fhYJrDbaw8t1wu97Yv52c7n/I2/z9m1qwaiKeyBi
09jtb+kyCr+ifz2bchJFiJ23+btYz4d9cx8RPmdtHytF3E0+FDu4WFMaMTdk3agT
egSClAvRI0xyVa3y3TKfKDk9mY+oMvFYSURtcfcmp+bJiAvrhrbRzS9m24kcS92S
Oq8KnS5UYD0g+avO2dSeZJ/YrSq/KSRkEiwmmoztXQfCFUNMSgkelti3V5kPTuPE
SEKGOeyQrJwTNjOkcqeLBiwmED7D0z+VLeVaH2N0oarq3cGyVOyJaFL/CEk6ugfK
3pXj4qKces1Yzng5f76UGwKXVjHqJRmS3FQ8LvdULT2/XeMtNYJTmgW17fxVsrgZ
fgffbAvO29LzWKWNKgrFRLVNmbZ+8NtxImlbnipzDk8n8i1IyM1dW2tZ/iDfzXuZ
DJu63sOHdjXkHwG8bckSQiD2racMM4YhoiKrdcnBQPSkBiA4jE59YB/H1KkgfVy/
YhZnZp4w6w1zZfQs4nS9+K0Mi3yRiW0CaITyWx1udoHV094rz0DgIU6v+dcIvcK7
mqaJljKqjW0T365dkvj8ECwLi/BGuILSsVYKivR7BfWHnni1hxfqnUktkKTIGyKP
NfQ/B5fYSqw/+kxQfzaLM6WMfnSsNoSdL1PA4A5SY0rn1lv9PHQFOEszgkn5hQw1
GODVVR0ju5KGSvaQ9UjQxx2a/iH859+BD4g2qeLTNnRe94olyuGvN8P30/sTwEJa
duvrh5X39So7dsbn00/60tDrKeVkJRVWBJkQ1MXFzW/erkwOdLctQ/0KBimU3Vns
F8PWRujEdNx6vCpaZOAObT4ikYyRJRheHco89rMBnqhNyK9YMvY6buYMNXIkdxL4
sihVHPWq+stc+xBQNvoIccaigpER2Rh11Lg+ItjeNxSLRa0NQURYziqVXwkjzNey
frSnIHkJ2koWhfggLIwuR9J+1sPp4ZXCLWSXGuO1jsEiDT61A+tc3QnBWdKWWXzE
1LkXCxHEgxHnmRD3eREGCo4gQH9qc3Dd94uDustf+4otDM+C//3PFheRxbIPqq8b
zc8ARWZQ6S0pLkg6yULtl60cJnvu/h2mpgRFBKjb1fCUtmpNMz0x3SdnABB1y3Ul
EaIOX5Pd1+XzNwqYVX/5pXEMM1SpZfAHlp6rg43w6CRUmYE1eS+ZQFXL1PzY5OVw
inUf615v9l93/6feReM0XHggyARI9dSWQY5yHT83TJJFIz1MC/DfI5PYHrvJni8z
wDeyFTRB9JV4VZ/6h+ULhvww1FhG0bwqi4h6d4oEJaAc5kHGIa+PJZhLnzq+8Ywm
rbXF72J2xpFsceZWNbjUbO92SqGWruzOOq4Th/iEfNEVA24Meujp7MbsJ2YiOtSd
yc9HCHSq0ghxONLu+mhATO3CsRD2dOaaXwUV/daDCdXJY65IV1gugkq5AcrifmE8
N96rRjI4lE1pICXNy23+xaaowgfugdPUw2X+8LbBr19hdvdXluWPoLA914t0MVfV
C2BRkbUiO0S2U2NfN5840V4+BQwu8k6og/JVjnwiOJtYZryHhACQhKW3FCmvYuT8
YcO/PL5eNPc9vP/WV8nl8MKFKJsQEhVvrKRUuYPaoJMoQqKSH7wJ9ijJA/R0sXbc
mRKtPdB2JOqGHQobuPNikI/ugBDVNjQt/D9b7Mk+q1wS9NohsIrE+ORjIm6MPKKs
K/fGGnHwfiBV1ERUWlmjIxHsPg32v4fPchHmWoMhrGyDTOcYvjUrce43yU2Lv4it
isGGVTd4pEaL9y9vTX4JzWrERk5qN5X8E1jIfYU9IL1NNf9P3Jl72sNwmrZ5KOUN
ab/nxuC0EOcjHItaqwREfdPmF2KdyDi4nzRjNUsNrGWS7JRLsPIAA5mO6PAKRLb0
PiQfcus9IZWDsKxS4k02NJNh7RCnp/jYcPjbnKjpv64+XiaDeMsarRiTdJI5HdNH
VCCOMLl8/Pi/jvrfvQjIdTe+Z5EqNnQaSzGzqAuV5KtBXZmWocB2Dp0d2dv3PvI8
5w+3AQSayKkt5KIvps7d9cYAsdY0qbuIj4SiSlQTcYMAKczGk59rpjaRdEkWI8np
vvHP4DruXQ0OJ9ITllRqboaymoNOXWMeUryt54VYUOwS012ATejhkCTLSuPKgPno
mwL8DL/5YN4wiTDwOJtKh6IV4kOuFugfkqIEORkdxF1lTxfBDHJ6O2afgedcRr52
iEUUIxRI0RqvFVs4af9IJMA6f+bK6dFKweBJICffecEVPKT++5xLojfffv6WoyYZ
8SgNuvA7J3zj2Csz4NassIPuEfbtBBiLTAMxTpLaPhiGl8zRurUdoYcF45B02llD
jBwXHtxd7n1JNTGNfoo+2n7XomXSHnb28dViw6xrLFZ/1KUhDXMo5u8qQrihp5/O
X5u7eVexDVp8990EU8GfC+DDI1I1dQJkLiLlvrB8VnEtdBbqkjvZDXeLlz9m3XeB
yisVMYoNGC/l77PGYVHe9fiW20HHmNAmHaKuFYkKpw6K2pIo9cBD/ij0OVPpA0pt
8f3JUlbQo7Je4BVC7pbmznkFWzZZf4vP7JWHh0L6e7OT+nx2HQd+5uyYRMQci6XC
OOavelP9FaYJh4nhBAa3uo98fGqEt6QvUPjbVDBgvJn77xYNFIppk0Vnvg6HgItR
HXjMo/F8vOlWWxcHLtLLV8gfHov6jJ7w9/8YxF6UdIoZvBfQWeGeEdGBwdGqUWPG
BG4HK90nihY0oVk586AHAWBFSvJb3+4URUFRg+P4UQjcdFQmt8rM78QPiiCdZnNI
j/G0xbEgC02A8N8jzCEb98q3oTHibPXnPj+ryS74kA3Uiv+EOA2n/ScfNXhk1Ejr
395KRhJP9BwJldlZmK0yF6J3WvUukt5TTj6swAs7M+vjK0EjkXQuwvfCImeNBLyF
OO/HYJgBrTKLrrJeaJyGPvnaRbynecIpZRFwLKGhnkNL3sJudhq6UxBjJBw8JR3M
78brBPQY+/wCFOPpXJsxLgoHR88zF/p70el0DYBlzhKWShXBsBH/XUD9OvkK2ywT
R/su+ZMeSiVDWIZpAAiYDXXkBzGi93KY6Wr6OOsPkHIMXEx8BVSuQmERnY44fXlF
Zctu+igXfORDt6X6WdwNy/Bf9QirPzQWg+OBo0nRXV5Vrc5sOEZ6W06E4OLPK8Co
BbpTUj1bLoIAzy4WuIWcOck5I9RGFWmf55dmFJCt/rE01W1f43+fMROhmhK/vmMG
zaQQ9v44u/c6iE6riChVVX/uXjiPqCJ+QP2uyjf5pZwqbwH425FUYl9XgviK1Ern
+XeDSOtRuRBgWqJ60LYaLAMRBsoO+FLaLlRD0gackwoXt94R2PDJzykVXxPErgQG
c5637/CXaTmmRNX19b/4q7WNG5knKPlFdUc4Po6NCTF/00R0r2KT0gvb4hw46lu8
JCBkWYs+jy2apijHsWugJGqwYEBPr/oLhIHYSouaWN56kJ9pekYcf9rBqBk9qxil
IJQlVhOqTMRiNoU8cTeiEmFmurZkP4fV50K3luGlAdUNVC8c3HfNp3aKlMm+UhMl
3kSWP+bMQBhG0tCRIaYZQhrTzbNrfVQLaud2IJI2XH2optX7bNIZSVhIxVo8k+rl
zTdK599bSk8sFKX6zbgZ4bLvTb2eTTL9NrZGgM0chJTeGNOtp33z6veNx7jb3e7h
hMH6whxapCs91pfq77l4i9LMLFUUtJhhplf2nFIe+XDoCjYV4CpPIXR9nGuAR+bO
0xOe9SEfFnhQ2q6wU52T0XiQz7XGAPfYUnIFSBgjkuTpvN9OLjmyAmVXQvx9B/q8
QbKuiX9sQfbh4NgtyQ2xLDxSVnDfIW3oAa9KGUQI8TM1d/VZVC7MoSfhXKFCDYnJ
y+jDM9Jry9guALLhgQkmni6i/11jNFr9pnymKbLINnRy5tg/Yk19/DbnB5SvTOID
6atdW4oN7rDc78QQk9rVzeCY6a0mnPQJ5z2Y+EQRlBoIepF/T4fJkeQrZNJJ5mSd
pu0rfs0k0O3ylKTab+L8izgdX84/4BkL5FI6XsglqlRJKdK/M5UnzR5t3/Pdk7Dp
eqeDTwMOFQCLqzCY/UdkjzhbS0GrzGMXeqtffaaQXLp1edxSn3Cpxu/WJr14/38D
0d0vaucHOCjJfGyorVE+PZnC3eQrm9Ba0RSaI4K2C1UDXc/9KgNML1M9nVqF9lud
q6r1DCiZjko5+ox9R5TBvEymVdRHBZKBK+GUNHfYgEPFvymL+fYe47JMgsR9adP2
Ua/KXzaMmsbAOGPiwq/lms/OA1wqGhugEk+O33xGJLVXtgmfoFHWU3NKv+22EbgN
0J6FuK2oVwbfPdGRUi76EV2cFp7T+6HazfBsM/tgwSqTEjFX5yrW/V3033h/SF8+
5w/k6rBTy9pqhXS8L8ctHGaFwZLQAf6ogNev5iyq+oMbYVk1cWcpTO/0WXI/A/KU
mJSMQ7lo6So7THgVV8gi7TSMcbh4Yi8dsEb1GpxWYpghrqtL5QrTGNzgr3gK1v4B
wOKG416kjakbgnVfbTGBGQQu5wuC5ytH2ilY94TLrJjpv2PcDrM3a+ZsF+mCeEMI
9cwHlfQkeuo3vZlIdh3DJBU/N6pRUQYzQ98trNssny4ff8aLcKl8JV34B8wxyjSm
OV9Ocxm8W9Td4cqZk2ReP0THU/hNtv9lr3llqbBUGa/usuJfhJfE0gVKpcZaTNMe
psVRsDm44xR3SwEAzT4Dm+tANP7UCyLnUEwD6SOeM1HxZDxa55DPUckzScAbJjGj
fZaOyYkY9WeCnA3Xn67jMQjYNwFZq3w5qTTF4pUVYEn4z2RMXFP7zGQ1OOm/P5Gx
rbiLWTIE298PXK7A5dkdgNpNeoggn8wgcZxll+MtiWRlSnsrEwkko4SJD5JyoOY8
kqLyzPo+N3GkK1g6aqWBKmx3rHBW0peOXpPNOaEn8ixgREOOlcDDf8eydgfCvs2e
zBQKiMJ9ntmRh2n7ny0GreIfVCe2qssoGV8ULKG6Ecge6qAmfiWwRY671/tFNHoC
pCLZbtWET3cjEngCGhlDhIuOTC+u6mX8O7WjIosKfsilgYgDkZn1w7OmlG4jfJvq
dbkitcgLJU/jUK7+6KG37ylW6CjSnznjNcfr+FkfYAofnoNF4iN4AYLCjq8pvIwY
r1wRJZm2QYCgua5GSIlTVNM/+DBx5M1mMjnkvTBRuKRPE4PgJdD/AM/9k4RnOvdC
C4/Nxg349OLVRCHYJ5SP3KoSEGQcdgRZPFLwVTlYOGQwhf/rj/zhX5IvqFsW+U5p
H1EV97+ylx/+Pzx1ltBBlR8L3ECfpEhfgqZfL3Pu9MSuTf3mA3xCKzFQKzUcIa71
kIKpoO3ukfOI9nSQrZFT48l6T82GMypo+I+AAxi0AqNwJFF7S/6QMB+RKzv0C9XT
OslnQTo1DCWeuxbryoV2F7oyNxXrNRoroBQsudLFRs3vOuHD7zK+gVbDWU32BGjL
C+jUqs3LHXBKKyYi3iPZI5w35vPBPmJVH172AOZW510yPDy/apJgMt828WMTer0w
U5Atmi1uMRuOf4kWnj5q/jyyDe5XZlb/8VYLqnUfx/plUCfmouE7lSMKwF/3Sigc
InZwhEN9EFa0CgEmrNGZJ53jWGdYNZmqtaqreDt2KSYNUySvEFbLOhDtvzzeLpRm
BogcG0jiAKgD5Rc/32mDRPJJU2n1cdQcQF/UL7dJV374adj2GquHwisdEhVkJ8Is
iCD5ZsqmjFjJzeqt76U0gDEHAZ7BBFz3deBEBVC/U9xCEVS5zx6LWE+1p6OEdN4M
DmD5m3zgfQhU5/BKg0uutHYcYIe27iGiAonuhod1/r0aUyJXAUvXrTixYlCsF5eL
ZToQ8r4N/wTeCwTVPxIgFfTx9uiRhhkUUAy5Pf4CW4katgJt1AHNjlm4BClKNY3x
O3xdNdR17CXLaIUqVqdhld1jxN3R+JLcKNr9L0h8+dLQqJtuv2aeHQ7ck9UclAr8
T+2TLFFwxAoITQmnsF3WuVUGfOBxp9bRBpY+MgzyfCd7mjvKvJ96pAfKWvimbwOM
jnRpC7iT5WAg3NrFcfH54s2coqqw729HYSY+vp9IEP76SUbMW070IXNq+ilksSbW
VZVdzBQ+06eIKxWuu94qVz9sCCZlBykND/lSCGZCIBU0JxTSh3VZWzj1swtJt82C
XLz/OG5zvT/c6VzaA3+bRiqcBCuXprbIUjGO0toKgNcbtIxgAGEiEfeQw5J9OyGo
94pH+x3heRfcdlgSg3zBw/vH0rf0kbjb261/N0ePmix9tWCmkF8Kj0oO5z+CQxck
LzIXIuNuF+njFbkIW45GOJ34lvkPEO7AedYuavt16ZgcKNNlomGhDU8lmO7pFPPK
IKoFL7VnmJyfsRj6Gz8bXPtqRizuPmYggDT0PS5+jl3sy7EYtj1+EBZtMKet8Pz1
8rbcNiFa1nTo3O4A+/y+qu4DKEUhvf0Cii3I0eVMuxNDszjfDSQ0ZRirf2GAGmvx
u1qwtUn8uxnthAqrD29wSo1G0Hs4zE0/dTaT1XASRvV7rJwTZOkdkF0Bdy+SlFra
iqX1A1oTw1v6orboPYntYvAMFShw2E7NXqYbJkBC+eI8oYFZ885/UdcbKM0cMLqZ
3uCXEBsDCzWAUUJpnJqGs4Qn0dNh+rPHVQ0B3wbfu5f18Q0oncMGsbghPNDBAmrB
4q1/FJ3FdZKfIm2t8ZthooMAmk26X2+uBzXSYRgqfxJcxzRXfud89/VPiPsJn3FX
mKsIrrAK20jCULswGgaZjRHziAsJg1XHao8rMCX8W8gAGdzk9I9G3AI9fuNktsTB
Vgx83ruCAFkTXtn6BPYVUnbUJNZHBWJpXehDEjfuKnHYJWnWaiuBP30Dh4aSchLC
QGGsAC3E1cB8LVJTJNONfg9jlUyoDMP8AeKhnR2wZ2WC0i7Gl2QGFevdB+1CTOFn
RDyMcnxHOgQQ/2w8kOq4KbFfZee3hKSPtVypUUJYYBlJ+P/H/XQUHUyhkPk4HFzR
dd50B8mWFePH69tDHur8rc+LZradvOinXQ7QduE1wZI25dsoopBrAKfvQ6QBlD68
yzJck6xSg/6ktDZSYEnfTrL4c9l0Bwlssw9CNzh2YUlJ2/8x/MOEifwxQyDqo3Ow
iE2DUqmtSqNQGtWAvc8z2njtvgFQaM57xRj7DJhegT+UQe5MOzMnq6MMYZ2FEX5h
E+Wm9sYHLy7c/NxQzyi3iFlKgy4OKTtYOd5IHuKvGXgQU13JFBRzhP/n/nsHdEcw
VzPDx1spkHcGZTf5+kfdvHmhahudGuYTuslxAh6gUQkL85/wJL3EWie2szZtTTaD
i6/RAnFrLfOHLGMRe28eDWeuD1Yz6ajizb5hWe/CPBIy3Ogs3Cc++SK5Rb1gd4Gl
kbGrEOtuwZcSCcKJI+jLiC6nEtLqpohBn/6HuGBlhSDU+5eBsVsECcJ2JD0SB+Kw
rdekk3yEKzHPxknr/TXOauQ8jmamONkbSvBit6chmZy+XuPHapDfnugb2/9lmscL
hnPQcR3FlFuj56QRp852j7YyIKoMmrmCwEWTAnMTlCfzFCBD/AenjKESts10gKin
LmaVoHXw9sSoSq9UOSZWuPUtlTDHTZyr69nOP71GUGj02E1UoZqsF9uNNDyIXdmS
Ldg0wSdOuujDqcwOkYHHvU/FlmYES01Mg4w+WszeVnLQENGxVZmUH/sE6Z/Dvf1g
QdRg1Rd/8Fbk94JntWGoOwokB5xGoFhCd7sDjC/NDV2+vrmWwlf3CB6cOZBHHM2w
H70zNr440TYaQ0c0s3tNHUOBlLUPczA/X5ZlX2L/WrP26cZJK5Nu8N/cwAbrsX8m
CEByYlacmLAUcsIpYLF0z3mq+wNKfdyCeUWmpAm6I+t6BU6GG1AK6AMRvRFhVS3z
BpRkTLQcjVG+oe2Tulgw4FbRo+vLy3Nn0ygphLhOkrJ4p/kLGBpCz9ssPAJyXZVG
4v1h7wtEZIM/uzyrY/QhfrKWHGq7NX/pGDFaNjYHUqzbFMvTi8VUkC5Lkv7XbVkm
UHk929Rz5tSaztT2wkjkPVRZWmrX4XWbDdBw5S+Eno966elkYpcb5MVcfRoDmtkD
gJTM+trFFvuzaQ0zRRU+2NKn+1oEjY4qZmEAM96MyCA3Iw5Opxjls6G35Nudwvl3
zUYTLX7zLbf9ZlwWnhqxylEfUyrJkYmIxMiPZhrC7vpKgX/huEG/6YFZJcuh6oGR
ZFqBNDAOda2tZXuszTv/XxBThb6xb/9FRN3AUWdKTDr3m0ufk0D7sBVCxDEntasV
gPz1KLZ9C7viVL5M7ZAPMMC0fCove3bmYcPTufaGo5DIRUjDD4w8eZj1a/dpMayb
7+bRp3Gtj/M9NTX00wgs+rBlQgq7DyJ7m/4ujVtEClEMjJ8wf2MzxCe9yXfIdg+G
JxN36Q5iMZMxtQaMtlA1VUDqbpb2KvqT1heg5xAAZn+F/M6ONsteMIaBsroku8eX
dz2opZs7A4Xp/UZDIumEjDsjkC9mmGxv0Qo/quXNA2yYujxVhE/+zdiD5xc15qJ9
EPBkBjd+DFzHT16zC6ngT4EbLynwMp7c4AgvnO3EYMTmuWoBtNXXRDCe5xVBp69D
YqUpWXbsywfPQEWlUyOeoQhAB9UdXMWOqDFAx1QIPX6KGKyM7HhMauPIXBz2iFIS
5Hlgz4R86TaZ5s254qOEceuloksBN4DfUWN3Hte7stMDffUahAeWhe2HXUxp8qpA
pHqy6L5TSFRUIBZ2HGGZmFrw0ETUrFL0a1v/527juZNVm4WgA9xr+Fz7G4L3T3o2
K9rQyk18TDjwhXww+jdjJDHcI/w1QsFiBvbk8y+ZBUbmGqFC78WLjXI3XEBIqHsm
f4vdOzU293gT0Ha2elcVUh9QgXgsxNoE+2Z/KDOoMOIXkgSYLvrQ5/+0RYKQzXnJ
yDF3tfuQKnvOLMWQfDlQ9/BnCyQG3ESCohIaLvDfuhdbiVpD8BDTP4tEIh56g3Zb
YLhatu17yB99h8NDIxVXF0M4MqjSeVRN/6+WEzs+RdNO38zHN4cNtuEtWjU3BaxV
HENpCXNfvPSqJJuHVAN08UX6d2QE6xdYl2R+ecVE8F7GPR2Q5BvCno9qU2XbpU/s
fAXyc2mevPX2B3/UkvfPPepyHj/go4jU45aMdvLhFtkiteQRMvH2tsXvo2/u3Vms
tx4E7yZssFoW/CrHdPXA0IXehn8mWUF+iW22jdr5KAnBzvKuleggabm/5omwGKFJ
R+BrtzaVttLNRonNxfrMV9oVGFu7XohzUOcmR1eKpvgw85warDsxUkvcGWggBar3
cRbYRrdeKl9etngdVkko1HOsdyGBfMygYzyR6aDU+Xbmxqn1iVIXuzLM2NEmwMoo
C/wsBjaA+rebsFfOUB/TWh1TvX45ZcHPzecHi3YvUUld/RmC1SlzFJVRzYejVEgz
ywcNo33dbJTkUA9XnoMdzNqN5loy8Pl62eN59RrZW+Q/Dbcr7e8rC1JZ5SLR8YGC
EUYN5m5iXObsRrd0WaYrqSNcVvQ7zUx89bMzQam9A8dLdNoHG8QDwFPlYreuPxOa
FpUqX5cGXZAxvqozD9bWNVGvqQqSp3YXlb9UvMs1XeRtyKUbOTHRmLoh9LGicXH+
EvIOwfSJN/o3nYZa4B2k1rzYHQuwGSJh+0NmeiZa8o7p9vKjsO5gc4vcanm+COvA
EPwCCaNFN77komm7az+ToY2dvqvQHC3sYFcyhvgJBqX94ZBGGitR2xiP9x9DFo8G
zhVRGbekFT1DPa09LS3h0esa7W2t8WR08FBI8qR6XTpwwDVIldu5qYxDJBxX1e60
59PMfKKDgxOq+RtTPOoZuenHEdW97J2FtVBMutY4G/1B+Iwr2bz22KUJd4rInr61
+A1JVKRo5k1NraxPsFPwh2OQ6S2/huvZQ0kChaoQaZGdZGG2VzUkxqoRLc7XL2ck
skGydayp0ifAcOtGA8GQH7pJHT30ASxL+wfVns9qya2VlUNzKLe5xoFYYm+vL/KN
7qLWnhPW7UNO94Pb5K3d52BZ3IElbfxhIwDxWviVT8qNP3EXWn3Yu8joPfR1ybH1
t60SLVjt3QtjQ+Sy8fNWhGeKwFd65XMFEmzEkXGkYosGQXQSPWRCsEovP0B8AVW0
TuTccl8AqZ2mexqfbieqoGCmK0uWyQ0lAwJBMwyrLchDmyIxc9eFdJkFjTd97/0w
MFAxQh52OFzlRJtIbVRCzrnqd6gALJMlzNuyaBh8gGKXyASszk0/t/wGi7YdvQpQ
6WQBlgX1np9U7tYK2DO4KecKVVHKEQ2xLq7GN4qXCeFYpZudpCIs7W+jNJi6UNfW
0okGxgmDHUJ09iT/VmvzVDLAFRjmxUvtLR5AtPPL6t54bpD1BZ6DAPfRKBKXrK02
gZ2JwGCRf8RiOhs4S1ymQX4O3COirfg0xP+xj5nkrd5yAg7xGL4/W3okWbiMGwLF
WUIGMofaVvLgDxen5yuzeubGopYMvi6rVZB2Dsdc8hTb3w0gRhyCgGpHtE/peE79
LGRIufgYVCEvTAPfP0aTsmc1aiyFAPnRx5ubvO9kpy5BuZlNaeY8y/fBkrtkUSkT
PtNIV9zpLP/fgy9cOxuWS1Im5oR4HeZ8Ntrbxn4v5wGL1EULZc496N1SjuZOuEOQ
cCmeFla4EZj4kZg+6orvj/4ZR4IHVxkO4m3zz3dl5f/38JqnCvXdzqmlcXYialHS
F8X/Jv1sXuG9z3AXe4Odr8Sr68R9c9ICoOCRV6+Jt9wmJC0s0/Z7DyIp2yScot3o
IYZI8iv0Ao1zyMmJWTkHGE5H0LqQsMPyqDMpnxf9tApTk/1KXSVuZVytiWkeWD0s
FJU7Cbh2GZY0GirypR8St/A0s+rpWWN9/IivwiMlAY9N0c1ax5TCg0g7HSR2nbPH
0gWt+D+e3tx3uscP/MxedBcVz56yAjU/sxTjWBn149xMC262eLBWJJVKQYvzfcPv
mdPh5FmggMP9TvQzx5K3TzTEfhbQCPHeCcYHN1ab0hyMvU5Q5/4kl89v2efHe9kr
GAwImOGWl1P+L+nKMvsno8uO53Dfv5NpLWfRl3SblzWo/bfumtTz3BPP43xVA6xz
0L8rP78rTOhPVufn2tBRb33C5Z9mchaJqH0oKDWdWwQYYzpUbGw5Dh/W0js6/Cey
L06YrGWuKUbNuWzNZS0sD8Kpdk2R+ENhnBQ5VzwJiK4/Ex/feEyYIEvf5Xl7hJ6l
rTneWp5nG2W4/Z4MmYV4hVglSrapkiaco+/SLagNk2Kjt4olpew5XKJ51tZqL4c1
UdF7hCFF7VNQCgbeIjz5ZEjXCQVEkdX1qmJOp1qNemrXRDPvHdWQxTdbHB22tAxE
UMjKdS2zY9yjpUGrsIV+JyGdVsW0Dq9rU9fPf/drVoMN6Cx9DXJ83vB8cINKBAEA
i5w5OzoMQZzWkobLPhXfaeqtU4bmrZLpEpFEBFTRftYfCtnnN21118ROA8qDY5Az
cUtq/s3HjmaIonQpFUAvLjUCk3344BKe7tkRKsr1ciU/c4G0f8BLbH9CobJbiJ6M
u5+yVk2fB0LFV62lTWQfx4ROGPgTwRL008F/aea7ChmhdpN0BJMt3JRFgjJnbi7M
fvfV6lVvGVpxxN8vy0iEfWWGr+W+YFayijVNGRixyiC4BExTjJ13XJ9twO7je3wZ
uZaltiKclAmFqDWwhP1vLK3soympqDZ/OBouw93QfLxUWtJHo6JW71NKejuLMll9
SEav7opxx3w85e8pOGMAbouD/brmIs3b8e6Wx4YuH1Kv/wgNT3o3gmUHqhQcnFu/
rSCqAgBEgmTB49lnZ+RKdpMtZZMm2qXnru4wtO2DaPnhnjIYZIK4LBeqb/7vdSGz
eCjQmFcE2AsDIBQt4/QLwBUmcBZ3rboosh3gwBwNaub0T7ZC2Qi6MmKOoig+gyhL
7b53psxvy44oIcm9NAxucOPbByDjwN04niqn2K8wXc/TAtgX3+GzzlUbDHA4HcQj
1o1HR3D3Nz3+KmZE5hLjMW+hA5UnI2tdjbUnWY1HySgy0NvCAIkEyZ4YdfJfRcV1
/m4i68S4Tthy0JxhuQlaA9U8ryaLvAofUahl+lyHt+fkUH+XAHeNmVP3obyqFU3z
lW9EXAl6L3SjHvAUyh1fbmsTNLQkkEJfjUxEA1ks9k0aPMY/hUZxxfE8/510+cmO
QyqPxEGnqjKTYqfVIXm6lMzlhkgu+aeZwrhkVrOI2hFu2pQ1rr+1hhAq8MCavnYv
RULXvTh+7g2rlZL+PNQbdtsy5j7nbM93yXt0qDYSrlDw98SEAqN6mUnwaqABZv7L
wsBJPhTZt6JvZ5INfwT+QS7VmT+TvpTSyrLoHMgcL0BMBBDFXA2/WmLrZy6zFuwR
KdgVtBtnKLzAHGoDsAQmazJLpaHaxGjtV18wF3f1XjEXixWVcmd4+sskDPbRx5Oa
t+6efS4QRtu4HlYAqBRLawFszE1o31eqLxOZJ5LRy42XjumanZzH7e3hI/q+ppw+
RA10C8Kc0Sg0+FlG6K+/kGeVc0h4tSikxVenSgoPyatO5D9yQ0XRfWit1gIAo9Gd
thJrahIyiR3HX/0Ro1MJj1ACA/H6aMXUPiAeH7XS11wJrfhuYH7fflE4ZoBwuNuB
ifExzFN688oDZmq4bgh5uPRld+NRj9OWqRXsFIPJB9l/v0HkkQWR0V2b5X4lluXq
IqUZPadO5pfiWQ8zuiOrPK5YWi5PzOzRTauVub0r+wA5rt/8+f0PYLauNlJFnNlV
il5Egj9gqTvCV/c2ziBZkoZljJf1g5scb8bo9maJgNrOrysk2WU60eI9OiO5Cvdc
v1ihy3PksSLPmhIdhyfykZYQU9QWXt/2Uc+WdnfUB9556G6iFM1BzkzKME0++DRJ
hpU3l635JNKAyuaaGx3i+N3K+6f2TnJxUrDcsEkQYtUUrqanyOXO8iI/x+zsNOI8
QYTZII4WeDnOhxNCV9gbGF603HzxcqNa0nyPyjU+xII7lfO5mdZIH3jlEyK5dfYw
ohtrAvHqb2SMiPnrPwSq+FSoLxvaIwNYBA4qmt8ksav9SltqMXRjHRzqRAbDKUKS
0GPE5R5VhhFqWXVM/kO/dgsihhhatxf+wQR9Gm6DAYEgl/BolhW/AAHYqBfrXm2i
zZIhRgUK/ks4EwJX8x/KBKGnaQC8qMwzv2ClYiPoi40D1UQyvrRFdvFuEoA1+iEZ
kXpIdjAqpbAQK0wOHmo2Sk8j00u45JI0D/DuLCtXgU9gy2bCNPxol/vpweDKsrVY
0Rce7pkm4gxlnM2qAXp/jNLq3HflaeJ2y2SdiIqBx8o+AOIo0XuUfpJVQ+FlgS07
R1LzM4YrHDQAS2zSEl9OaXgUbbM37RwHExb2Knhnp+0TIMmRIZ0UsIGc+dXcb7yA
fH/c/vK2m3iyHmlCeFvet1dnbdkbpkIOfiY7CwVNdArNFim2oHEuBJV/y3lr34RI
EYBnYMGuUen7/3zWG/3nUYwZOrKu1fnDlJZBsN1Iu/4f9JirVwgz1fEFl9NYsaKs
GHvShPt37oZWXHk+bi9X1cfN+NzfWsBhyx32OpqSTylI9M+Kqcts5haUEorDr5lv
zwGLQFFxsm9MiT3TOBVByhM7BY4lQeBGzRhzJMfkg503CVZ12NKdrO8wLcfiFTX3
cfh/qXD60jLl/iOA2jNmdG/RJLxD0Ik4LoYuajWExvoT8/KjDcIjhIKz0HAJjolB
XgPoZ7ldeEhJA3//+WHPXh9G04D1MjBl+151XkJLgdWwjZwVtaQNWoQeSDvaDLaZ
a4COltuPdlDMGOscwmDZMFBr2npJ/mdLTWPw6kknu4du8pjzZ96VNPiHvR3xg+Vx
jMkBXB7zwOuyDP4NEgBf5OiDTfpUQ1JkW8bnrGk3+yXcTaVVgwSJbRnOkCbCFR7b
LRazkMhNFJvbjHyOyrbCQPS439gK6gG+AVmbJs/EWJ6nN1GB3o7yKEZLkI1B1w9i
6yXIB6wQS2aigEKjWd3ChJoVNccTqaPuhzAm/nVZCmxuJFUudNdOO8zj2L4C9gPC
gLYOGosgpfuxFjJoSyqNdfU7FooBEVU7yOhHY44dM6ld1Q1yUKpCx1h2bwY8L7tD
k4k3Erhz13Lm16lpBzI0dXJjOuwSmiDsgl9Y6D6chfINWY3cLeTuZMo7BiDin7bq
pRztVpSjj/9E2YtTMhoxzqoqGGHtoDzVaXnPML+Te4zMG6SMu8tecE61kTIhRbV0
VqDJglPymr/RXHq3hQXSWY5iEZPBEJYxpYUPRT37mtU9c6bW9WSIHzgn9pdM2D/x
p+UYTH6tW/SxIYVAwRjV/6zrWKS8Rkd/mDrKnY5FGwitGnGXdnG5gjRJNpmEoGMS
IJkJ3eZG83QU5LVybWl5nrAB+Sjwjc95eiNnRqjQeJrGm06I2iazIoEWt+vB+kCD
qJiCdDc/3SEwWW2vQTN3bJ6bOoMOW+ak8Y/yR9Dnb3ok68rs28ueoq8GPzjCN03h
luOLMEBjZql9ALGkTspFo8ynD9jpqHRI9phaw8erqzs4JMhEU7LDZSKYJ7Qwnb77
YCgIIebp5aEGHR17TI3EC9xPXTREyZpDbIWPiL6Jvd028hepUtM/qzHyPt05vCbW
Hv/L4X2witvEx1Q7AVnZdpxs4fergnXYAGxSqdJnMfJf3vLM13SalVUal5RbKFTe
6R5sC6yIMKMJmNtlvkhj/kXaaaplwp1AHipYbQgKnghc19inHis8ZSFpqcatiVzR
Fq5B7r0xPHit43E1hamcCsN2zD20WtQ3qm/lISlqWXNq5pSnMpEUiBmqJMOQmHGL
CuCYKgfVLK9elsacNEIxAmX5yPfmeCRCz8jn8ksmujJqFWjMXRyi+Z1KxKIMdpyF
d2D1CWN3OuKHwiLzDalA6LPBbdZgICyjQgJ3ZKsLqiGbHw7zzY3jXZgZl6qnk4Xp
FOHfZIQFGQxawVi+5W6e7ljnpvt+dwNo2UpHw7xiaMzMYfhyjjvLpyHDptkUZkh2
H4KSg3RFM38sJvsEo8SY2iiZZqq9BnkujkB1O4SMT1B04zPybr0gmsfPNXIazw6u
rajNfL8R5Or3sXsRc1FYOONnoBC1kgomCEfNaMo0ns+UF+d9G4bEaiPeEewkIl5x
5Vj8njigp8xKXYaGbEwXI4JI+O5xi9ACAmwTYuLFib0HM00ayjgq1bwfYrFa/hQZ
QMEZEh+UHOT8sxuxDFxGmWBADXvVYjKHypEYBF/U+DwbeLBIQnly+0aNn3MVTD41
MSe+p7ErxA4pCzmkUan9CzysYKiVXnoJyWugrD0oJgPUv0Uh35RXrsI72zuksj9W
C0Jooe64rpVrkaQn6dj3lhVOnbYoccHpXGM2Qwd0J4FmacR4lQe/LsyMahZ8EMkX
8QoCv/ZUwMA8GquOc6ag/SFNugSII0sgiTSLGPJ75Zx8y3UgPz2iGyOWxB7xS3R3
Gbu/GnCoq/DGwO3OpiO/gZmObqz+Yu3gqKhSI4PjXn+WweATIuqzQm9Wa1jbIlnD
Tw0f2M5KHY2/A0P0Mcm+AhfyyEHyryf2h5G2tfQqYJeRJF+4fNSEAAJTx1O2gnbq
7HKBfVy/Lkotq7Xsh7odv4yUlHPaDpdb5+KeDqgICim6LYXsVlnfwqdPcMFuNWRs
tRQ3/s8uojAikBYARM1la9HdkjO+M4pmSrvyyQAkn+Buza3WaAVIR5/UYen0o8Ud
2VyF2rKUGnbiL897QhN1EWXG5FAHxq09jRNYPIEy/owUvd9mU0OmIkN3gNtQd+rW
8+tBWYmSi6w1i04rirqOAVNdEhNrSF/NS7XqouHXXhzz5fS1zx0UYqWhIitzWj89
wjeWBheoLjLAJas7XUuDkrT4U5eePP/4kARlXIYjy0zzpZKol9vj8NjmqBewmNxm
R5c3kh8xm1NtOdaozs5bCeHV1Ci2Pc952hKTZD4EdrK52/1qXT1vAOKeMsRyeNkj
88jOTlCmek5/LWQkrKulQlvm1ZbzFqaJYa0kh3R3gT6PIfhvkhDLIXsZvdOZKsTO
aZq6pCRYTidyA0K/+v+CzOMGP0I2LziVRUVcgttDwQ2K+BYTlkCn8LAUTG0wGYw8
3Z+p3aZhSjZPkTn69n1mm36fpvrCgzUqbVOoyD96uWCtlpIjW4HYqBJEjNwgkvKk
zZAFe6vXKoqG3EXnIDheT3TGcez5Ybiu2KFO8/eqmZrDHvcHjRjpWmcHD6vmhHzY
tItHD5yQ872nck3c2DBvosV7K4tK767XnLyN6zRx1z1NR0AjP9EWE0hrJeobj6Tt
1OjLPYU4si8l7Sq3ElVl5B3lJRt2xJJf9zCI9armWTIHuO2q9IXYq4zQ137N4JMu
slcYjzp3OpcG16ZGp2HQVfMmybvln2corHaI6O7XbktjzGJCMLL8xKXr0uIrcvW3
K7e40YtCPqI5NjZuo3vqyeWKFhgf+oArU8dSWjzTVDvDakvuznP4PMCaUmabwf20
/yQfGo3jl35HzV8rjtqkwcp3AMCopdWzfDt/X1NUQAcqJRHt1Vj+PVCjtfp3Y8Xs
j0E1sahefiFXqGAgbArsFkN7W6ShFiaBmCmy9GLzE6W3oVVHBcJeZSklut0qinOK
1WVk3EjSr88Tz4OiBDgDCRypEy2p1gXDJueD9keGnP0iJovHodwNhvw4zjpebsN/
wAx0tNIn/aRdFUXWuQ97pXurOjwcLUAlaIu9/F8HH8uKtNR07r7bZHwwSzKgxd0N
ewD2uS7oa/HMXmA1rd8Rrkb6CKjOZq1+6HeKLKM1uQrB+AVfb20Ji8J0VRqIEpxa
E/RGDLzNih0Kp9bu8yQbN5jgwfHG4mmvrdnzVxaC+FbfGF+9ACBujm1O7Mzkfsjn
uC6SY4yo8kRJSwBXgtT8GbZQYjGvTuvO9Ry0Mhuc1HWJ/ZJ6LD5AsgEhF8O23Wao
XSH60Hi1SC99aMtNwmk0ZdMmOrzSdN2w5J1fovBWlhUBqkadwbP8FUlphscI6EGu
LBJc/Us9NUZ6O9D3Jm7DSaDAAHuTlXZmLYhMenAaerd79ggVUMv03dnKO5uZLQ67
NJrWEUci08zqIEC09b7A5J04jKI5xKD/ePhc/tS76D1F+DnZYdCG3Xm6fJ/O4xa2
eBb2bewtrsRbm0NnHozjI64BGOEX+oxSeVOQYdLowVVlahEDK35y8gX0O5zXyGDw
D7N9f15ofpdgBfwWu8wVSvRlIaNXGJwl8EBOKVjCHWjV5d3hr9uBnOy/NVEvs+Jf
mJmx2/MCpQ8rY9310W518JjQ24u+nWOmebzkUhu3rLeneQVBy0ESHbwse+Wt6DyX
uUHuCjvNzX9qclmjUl5Ba1JHFqBBj7kOSyZiPXzNQnQNScYL9shLO9c5/Qq97WMq
E3PSgU/3DeaQE5uyWA83sKeDWIHI/qlNXfXq/RMJ8Cs+ffOuepgOSW5jU34p4X1X
IOH5x8E7L3Bddp+C9JkCVH+OYrkmw8JjGQDba8+2xI4NrNGP1k+BweddmvZCioeg
M5gZvMVshMwgfusFzZ1qa2Bt9PGRIAogbbO3atXY0FjrKS49Rt8HPbaf0b1z375a
D0sKPVmzeJ2yLJOaVfD3YyQgcxi/4a9h73Fg7gpUfejOFDn8xaIZYv+qaPCYXz09
x3MPdRWE46Xx+53QW+tAC6SBcPFPx9B+uCL6NXxY2P0SsWIPvGcEdsDVNgKKguHR
b2lpa6NDby1qnptz/iRBbzsVLv06SrAd4n4Hlwknva7PRbKsUzO20gr/BSJUYeyS
4BJEnCDztBc610+bPgqPUbwQl8fuVVIKA6bz56MCuojHYSdOAdEefvxIKgCUfq+s
30JrqxdTN7X0dm/O07kVpphTgyzC+A242cK0d4PB0OJL3T9HLC0Qe4yGrVM1fce3
PCbySC9wGvWaG+U+ieMqKvXW/pFbTE+goMRGXLO08Ol0qA6F5NYmBMzXwYnLziM/
N0OK4ifNIWqZBd183ASH6don4BIPSrqJ9NvU2WhKuIyTuj582hHGx2Gq9ij1GaEo
etZwcnze3afxZkjQh3OVdvMDhFQYgJ+jtThShf7pkPGlG8nLj9uPwabq+V24d9ai
m+5sf0VPeiuzNkyP/3TOTvuqvKWLQqB1Br65zq29nc3D+Tpy+uXtSp+F/TnLKh1n
AbESeDUjh6HnRL6COdkdJpmikd9CL2WJTobqHgU3qIGhCNzJutA6qxWiCKKGs2EK
nJigTttNcuMMV++oh+yEqRksucHJHU9fUUhtS6qGfEZ5z/G35auR9mzM95MZW6oh
6FW+dCahpS4K0zwEy2mb+8p4nY+W9F8KGbMvJXfe8JZJJRDSMOpI/pf/ns3hrO6w
bKzMrj5pJy/gwW6oCZNhGPDGw2rwuNKML4SHQONN447WyNsPRC168TpxV0zMaIR2
aA47IxTRuR6NCBPKl7XlqeVWsqCjKAKvACrakYdC4CdxJ6sB8U9joOrWugNAImev
AOhzWFNiXf03I3FX+W/uqKY8uw2G0cvKmvJ/+0AGyDDmb+d3+yIDrR6KGDw+iH2z
VqYHN6lCKggKRA80sn4+gpA9eKwcxCsh5LMd7jEW4VPS10jZ1ogssyu7Xa/rbdEw
PFqOMdkDAYp6uK1f1sYwMhOJCxTjVzYR1GSoo7WP6fsw+D036zmd0Kkg9KM2dTzX
uQBHKXx7buTlnSGix4PIYlmMPQF3JfP3qV/ga5/YqheM1unZyS/T7vedc8uGpoLM
lglpNTnmz9iIe8rQ0UYIcRNAKOjdM2AVZ1nrrDRunszce3l12wxZEfN8l373UP6p
x2CCRYB5WhRA5ing2RVGSjhM6VfEVGidMollp4fj+790BGNwbfsDaptE5emir12w
avDQ9VTsGSInjXF7vFk3RNqlRjw5N4yTqN/jJrcjB/glFh25tI3QCqcAKr8FpdaC
NzDhs0Q6p7v+aGWzLTeM5Kug1J63hp5Fm38+NQG6HvSjtUWVJlswVSNoldZdffN2
1aTrB5CZENRuQ6sOBGi0RxzsHzEj5N02rgg4dc2P4TW8GmZtpmUn0Sw1Czh9PhWL
32XuQ0Jaye7+J9nh+6EHYTTrgEnrgork0NNp0x0A5gRZJjp5BXAAUzic5Xji5oDU
51OS7q/q+pnwojy8Gm+HV8ZC+2zrWGuX8+M8SZteBHVXM+J3+aAswNutMHc1bhOK
/YFcOK8WwNu0dMpW47k2pzBkbLOO7jQ+6/CDvXgkNuX1DhQUqEo51ER+1v3F7l0K
UKtvLaMtdRTw1QURezfWNoKL3xMHnMfcd/KgeTAhBJKHspIMII04fdh8WegVtRNv
UQby3EEuITb8vPguHED5yYEVaVa1R7tbDh6YUvIwQEjyj2UDfh+/7C4Fkw+zpJQF
2HqrVEPrerczllSeJuCXsBk1J16a/QRWOp2GPIDiloICRVFbEdbDkxgynxDIfi9w
cCumQP7GTeVDEVG+XN6jj+lEMByJqyvTNL7hy3n/noFA07nmplT5aJM6bEyb5FPw
Wcywrot49msJy/EqmK/u7STEm+LRQ8dSscx6Sw/NsUXPPird/2l7NJ1aaRetvxVZ
IWJ19zIkewFOTpBmhQvFaDoidcswnzq5e0gl4MCKlN3HN7DyvZ9EpYFa/YVOSQ7Y
akm0GsxjA0Dzy5xP5WcfGZN4lAX3B8dIsxTgPJzL2yVj9I8qdhvfLODzC+06tZJL
IBuf6jMQh6pqulucf+Qi3iMR57ngOyO43946cwJmbxyao9GV5Dgufwo0oyfOF7S1
bjHzKZ7WorSUL7FeV7zrwIKREJ+bVvSEC1OXJCxzPaELWF5mOQMfK5mGlIbxkZHQ
GG2ppEfIDSpoZ5g08iThPLqRhxw/7hlW/1wBdUQt53q9+F/KiqkgNSSxaZLr9LlT
y460S4GLgM8EBN27Zlkcq3eUXPzPRNL56H71mUb9UBFx5kJ73XovzzKUaaR4a67A
NHSbC+6v6Wz1Dg8SYpVWM5trG4hUjJKcGKYK46dJwlxYS8XjkEu0YVyk0UTVFI7Z
LJzJH0wmtlhYAAdJiNk0iaoKAr2TAQpmScho9dwSS6VN2g0tdP3tqdbCsv5ZQkL9
OkTdZG2k4M/NpRdGEQmQlPDzAs9XS0SVJwKXH8tP0Q8LvQCp5ZRypxNS2nIeNKte
HCYizM6GAjVA+FlRf8EQKnYS4rM6RusQPqL+Ka5PJ15z09FNioh3Z/EZOTbe7I2I
MePMSgrGkiVZZt93orTpwCaDZV808hM66qZ4RsRUShNrkqMykZ8oKIa7WWi9dFPU
deoqCAOQzGQObr11tcnwtCwfwE2upfpz8CpulD64WRWKeKaSashjbWCAK+WR2diS
+p/dqh26yDtnzY0h4Jg28XEfRnfaNmmWwuFba8QZD9gCgvEsPMyuspnJvPaqHcwC
V+gV6/fOni5yM3EpIEKaIMv8rqzJo6YZwJM7cOg5StVxxnqk0aKmtdb5xH2G/TuD
yDRcQodwLwq3im7RA7LzQXWLYkopDwuWZkkKmVV6xZPfMJF2ID6X2i6prjylIcJV
IiTC0hQZDEGhMVywHgMbm2I7GPzop5Zea031xrN+sJQFvVZgY7TaTFdIwuumDHqw
QKEbA1qMmyi+iS90klVFe7zx1mZnf/c5/Z0RqyYKJz9Hyegd0OmKZBikEjbA68Kc
BeraR9KNLy0vyqt1J0G8iLxpOWLkGVj81z8xl9k9EOzgYpoRC6XbZMMM+vTuKGJK
HUWdER5zIKehqR57FLXpZXgWvNhVwqGvh5TtoDFwn+j30xTo7tLFTLe/4EJ/YUzd
nncFnPeetmRCGFYC7uoxULnWYBHgNMF3B5CNEzLS578jEYaaOcyLn980v2QnSJqw
ee0isSy7fTRynVNESthCy+Xq/hTFEeXzsX55dUmEBXFps1NIQG6aEWxrHV1saQnf
0zUBUUWZMK08osTjjIIhp5LPl+7ZEu5ZsiLHROgxkchnhXtJSfQv87DKh6GAYa0u
7BNfvqfPWeBrXJ0+HSwoxHhhtscqJjFhs102cWzhDgmNv8HA2bY7uqBWOrvaui8n
R0VFMVyEdaUDCguIXZmS4Zah5g/CTcr6CqGkMu5lD9NSyMLQOsc2N/FEkcQtxBuB
rQaGkltJBxL4B+IdTV4lfciJM0Mjv9gd2pV+3fp0cKS3dJ0gchEopwFKaAqWgNjn
KCsb3AsQSYtXm4Mm/4dmSFw64VfX14vae60EZupAAUx55aZxs2L6VDZukDC0X5Fh
cxMl6FyJvjB4yL8V+JqD7SIu4i+P0Q69Hl7Rpm+E9m5VPP5GdatFHsYjorUR8Qq1
zYLuI8kE/nIqyq7XIHrGGH6QzaypgsGOXLbCVcVkSaHwHVBkIgPieQRD0tgo4Uff
tcNCyKC8Qp4tcq5kS1mRFc4MGoEjKoi5Qkn6cY05yynvSVs4fyBzqTwPBJB7X33u
GsiYu7RhZJbU5ciiBoc0m2hTkeY+88o+s2KHEYnXaliVDUY2aVKlsd7wycN2qTd5
Etv8zgkvLuxvzT8hCAJyK19MMvq2Lt9yj7majSzBqahKvNcTRWyhnDTWiN52EBez
CJgwCBrQKB05gL64Se6omCgNQLdq3EOTexnKEyQv7az0bXGU+F3KkOjMCgH2SH+d
1ZVc5siCQ/OkKLaUwkDo3zglGfk6wwbEunaQQn9hxM3v1XddiI0C4oS+XiFG9BsM
HBbxXSpZWIjfpCiCNYAH4b37zV9KYJyZl7SvjOuanimhN/Jxc8gzM4KWhZXO1M0F
4Jk+FUITx5dPnmYMDHHp+bRm58sOx+Cc2x+GhYMqTPuXlOBlYBYfTvHZolrFVrQc
UDad78FyKSi5G0S3SyLHcu22T9MyKxbhW/c6Y6zI1L7ychqBVLDSSzyycQhztn3c
Wib9Uzf7a++/JandfqTF4lIDWOagbcHMY/5gdy9552BRONVHWciFTLPC9/k4baXy
KhsHBIntfzc+mk1BzYgkft+PS33Ucr2lMkhQL6KSORCvSAC+2HfLhQadpdq6rYLe
0hoxmsOZDsWkH1X2kGBFMAwEzJq/aQuWZfb2FQw7ogEpObOiFKOTiJ7jZnlPWobj
6mnJb5TIjGZC+mdeYo+ETC4bA9tVF0CffDbjR0OErshKLT8YMeZw96V9WfJZFYZW
rDz32jR/UhcOXv/oai6DWYOFlF9+mlF8OJLozdVrx5I1jnYdIGWLS7ZQbMW9bpkd
QHKp5Q8uQq8ygbVfdd4huqefrNkqiuYHRGHwUIlxbr7DQhSacRrg/yydh2KMqIb3
r87g4L88Aj/LHMEzyB5yFQAOEk1JAOgLx6CK2VLI9tJyYxCm3TOyWWYKPgI9a5GV
YTB/gF7PRCx0BcBsYLp+o5tMoMEBr5aUm54wUEow88qIFyci5klHMKBtLq7hJYsq
HiqlWKZV1reVl6RaLwiDBwSSEK/PwUX4vCvpOXeNWQ3Kvrc1juawOj1PXovgj6cn
/m5xWmjtIUvWsQOaQSnTEv7Rc/8iX4puk7bNZN0XwgGmdQhPbh8L+VHawiFBTU/C
R1zcC5DKuSX2Jbkxg+rjVZZG5PbOIOYSe4xdybN3M61/9VyAU+hGa+3/p5ci+m16
llxy1sQjZaX09DFR8ac2CLBNEcq85DyvPrNpK6/dte3KtBe32eHXOlwWuNYyaB07
eSqfImyGkMNb05Z2YX7GK4BRxxbKGsw6HRHnTbE8KdiVb0odFiLiZLQ/ZYJ4IBTA
u/KNvvYv2MPQGYWsbG1IU9r9uwsbtrB8X+HCA2uXQmFJPMw4LdBbuakGZLBgtzOr
h3YgYS4EOHLuSOTg0ETt+I9y3zKa/IswKf98WYJ8LJtfcFzIswjn2Cpha8I/d0g4
A6kTeKVv6sszPjSkWIdM2+nXOQ+ulPzlrCG0yyjwwUsGEY8zbokUTDvAceQshcmW
B+uz/vP+7R5aAcjgdWMXHDff9N7+HbPeQBY/lHWs5x9EdWv+/tONG/B0Yr/MhzpG
20SdYzapz2H6MZzm45VgcF/hVchrZ9d6iaCEon9ezkcwX6cPOvTZNaposqVUvK2U
v2PX+7oN4ppW8+3fGBzKYJYyHIfcXJwtMiuO+VxqWnidtig+L6ex4YCihxe5M4kM
wy4TmOlybk8IVZ6C50xSvu7xMKA3HKw08ev5gYC2MldcOT16EcWMwcYo+5iRP7R3
SChZWLemolSeVJiW73u13gLUZ0UmNtntHdZu0hpKPq3D3M6zPo9c0oWBewl44fTC
7PXu3jeJv7iqIGBpCWpc353jBxr/efGLt6LbNyXb6hmZumTiP8N8EQ/X8kR835nb
nuxGR9ewH2DWjx0YNGtdivxelkyrtWXeLxgExbcwkf0QkKzLq1jSn29qUIcTKpAC
bH+sqphxN40VSRpsl0H4IVNSzzD/EA+xiNu2L9Ft9Xo/lySgvRzgxN6eyfTPPQMj
M1l0aFQk6OKClDISF4ho6+9ojBLkLPYJqmDTkyi8z2O+EbTzeW8kP5jSOFI2XInL
6/6JpTj22pFhaLwHXBiasmOAPdGwHkWKCpRVDP9P7IR2Aqw53o2tQPdl/2DV8vmQ
sgDpPlvfz7K1OZfx1dAq2jge8ZYTO/JpbJgIBujKzjeGcu+SWjG7M+bXtYmG6F2Q
4id2+jC232oRmyr2zuEFLhhb0zOyOkLx1z176VwVHZJbcMfQnnebAM3IUxGHslJ2
vi1Pbn/VtvdOW4pH/OOKL02EVQputj5Nb9cSi5IQIGWpJfU+VH5UDK7ivpE84nb/
hhPOFzvH6cMyxa764ZUXq6/aGBa2jwHftleKPK4fDnJFbDxmjDw5METRrjmFsZHX
W83LMkZCx5rxtFEer7wm/IhEDFwyFgdpiXSyWMD9YEepJSixiA633+S64YtxLnBQ
qZy4Y1tU+Gike2BiKHPaEIV/sbfdWQFBurHYfnTrFOkkenDznc7I3CTgRkwyUWRi
sdbbYMxM6gwH549Eqvz7ZDgo07DRj+uqSKHl4ralF3e/Cibie7zpO8Pnu2rGWdWd
Z6JonxCZXrkW17i0NmQmyZ2lroVCxDAqN9f6fPYaa2iaLA/C0jhDQHRqHq0I0VoQ
U6sGJ4uEXPUpnUvWxScTFwizE2m4zQ/oY7TUrM3Ap6XaPn9AZ0ZbJoIzIf8ipS2n
X2m24vz51D4GPaweICNL0+edVyODKTqxLGYnV4kbhPUkhr4jXRQt5ZzHNITf3zVQ
a4FHmFLVwVyqmtEwhH4g7lQX4dl0c5OZApoeVff+GJrekr/P9kUmj2Tskp89ae2y
5EvzpMZKRzPR7WqPMDrDyFA+58XlNhmANnb+hjl9Zp/u6sA4xr4DTGOfpM4kSY0p
FeCi7VNN7r0myzfoarWfMLaayJHE8J/5nscbnPzYy8Dkwhy4odqkbDHB8mNle/rB
BIUQXCDIw01LlXjzaAG/nvris3pkYnwrE6svgjis5a3Do9vZ4gas6r8f95fTR1zp
OoyG7fhxAuC+jnKUCoa+nSs5qGoOk28RaHHrWNdESM6u8nFySkFWfUdq7ka/tIJN
7c0qP9iiDLyMPzqedpT+LnJz+5olwSecZd4iUUBIN41t9seHsJzxC2ZiTBC5yQlV
4nPN0E2ra5UuQ9hibWZdX868edPh6qqSaXnn2tkvZ5qEoya02QFCLJs0+mvUVb1M
ZO2jl8Mz789rhboEQlDn023ZnMbz+z1RbmETZGTTQ0Q65+5dzUyEbDECUJqnbKYK
vJilnWKWsSE+I+DMwk3P7CMIJNqApSZZEP+aXPDp+Rq0J3ub7Pn6X2A/aekycrpN
Wt3BgOahSzuaVkHDk198HIe3JZTNGP4cklOpEHPnJtRhWAryIaJXbSu62/EVzzGl
Hg/fpG6jCkLeqV3fkCfzxbl7C4hbiIFSnhO2swAugx08rUkOrcuZszbtCsibQTFV
41s5rJDOnah8Dl+Ka6rmyd6IYWfAwYzJ3ilPfCVDvYXxSMi7Di+i7gAsDRFqBSph
CNI1cqI4ZOZPMrDeNyfXR3GiEnkx6hQsOCtx/hbNKu315l7f8W7fDW9Pbof9JPHM
1DTJzW2aBlY3CFCdsT6gZZnleyaiXUoOu7YD5s+kMgHZfTvjqFZXgr2LxYKTDQl4
dqJQkmphWSakDkTgeO9jRg4AIsbpIgjUAkWZ27TATd1kbIiigl7VT+G4VcIxlIZ6
hGgP84/sHfFQ8eooK/7tWDPApZUbdHZlGBqT2Wi7/KthZCWp5fPVgHKHYKB3PLYI
VDDqUvdHhRfeiAEN92o6hv5gJlLebBA1qP0D+SNeBoYT456dFyTf1BDUub/IbJrO
lJWJ71PGiOahTAeLg8eXavWLcmzswfkTqv8kiDUL5V0ipriqOgmULUD743JQMFnU
cwcRY8Ny7csNGLHPBHcaewX96NEgCJ1mgCOVbhfL2RaGU9WENbIxAp3oEc1X+72I
4ePXn2nwcE83TsZUVe2hEc0pWb9rudcqfAVLRkFuSlmcaBeBskCzUrQA1/PDsoYE
rZxfPAdwcQ0PrlVFm0mg9+WwhXuVF3Z89Ucb9OPLVgFoHRJpZQG+KQ5hhcCKvc51
fNgczock+PDfAJCZuX70k/SMBlgX7FlKSbX+bmFQy9gIOPhDIv3QvB3gbIZ/nQHY
L87URhwx5mK++128ecYMb85t0TiHq2RBvJo+5doY14B0TpfpMzItIwBTrIC6Uznc
u4/woDxEFKYSLRAWSFC74ZM9ETrUsOZbG2Q0ofxILu8iO/ezrVL+4wT4lsmYhtC8
8LoPZeizko3NCZzhuvorBo4BbQGtFCiCdDnUGafV4QFhTHTH0Yr97aYrB/BjRWax
RcrUa4FVnjk6zcFViCZUCcsg6z2mw6sLzx05tumO9Ovdm8QoNDmOAcAF45HwJAFf
KCWk5pRz31K15KWFD5Z5lKdFP2R6JRoOSYHAnwWz1MW3cS/ylTwYkgdbgzG2NJPI
O3d3zcnnsW2ArDb/lfHsff5xoHev7snG4FNL1HXsJd6Babh1uFdHIZypg+RGTjOj
BpcVWOEEQaZ44PB6qruNOHUOdLF1xgzy/oBl4BD0ae6QTmYabmvfnGSVQaEeU5We
xEto1ciVNnmUeA69NGUU78sfMZnK6B0tqIZ4BHAAUUuy323/lov2jNb0c5meMhYU
jmF6Bt0nt8j60rZmFE5bUftSMpIPzhJTKrIoMlLblaV701htSYaCdd8yEIWLMRkl
roRK910G3oOq0yNHi52RFwG2FMpamMy8snyKOlJPHguTdbfAODXUunNdR5L8QchY
Ftx4/KiIQEHqeKv5/LFAeF7dm1LVaiUbTxYatsNPVbj6UpE4lf6Djo7oUdp+6AO9
AHNsGX5CkQIAt+japfC/9yE3/kJ39e0Apv0sD6xjyogQUIDqZTsGcLIK1ZYTibm6
p84pOq1PS2V6uXoLOxDnjVo0ourHwM7yNBZFe1Tm/GBgczEOdgUNnGaWq4bxzLjV
zqgYzY0+fYdrYzKi6gE6u+O3HSOcMAVvk3ZmgLpsILgi5yhBtBRqC3A8jt0R7Ity
hY8DYBnsjxeGQvzbEuvsMiU8zmdzNEOPZ90FJGd6VAfENQs5aWrK1pzRlFL61S2O
EyiWzZgZ2wXUa4XozjujkiajLDh6Fa+r5FkyN1RjB/PaHL4qXE5ghvGYpgINvbFd
7gOloUUHXmemRmWz8i91DKO5X6/84aKlpQqJH5fnpM3p0DDy/CSZMu+mmvrgQLl0
1/EDH4U+1B/6s0aNlO7WU3OvqpUU/a7Wh0QXNUWy51bUN0UpmE14JzmBZzNwxqyx
1wy9jOJXSCenHuyVpjIfz0pJSMWq/v99JWMF2y7P2dXdgACP9K/2BPH1SRLszRys
ss/J+tY/MRVn+JEUNx4xdZ8Du8cARRdCuLnwXzhFmDSsy52R6QbnFENZzQSOHHSS
gtWIGCFr3U2N6R7LJiBuvdP1YFIJCrTro0uWUmk8uuDbx9e6uaW3dF2+wcyCaOWS
t9dYKyn4FxQLvSlNpGcCkcSnL+pomQLNhdOlmja864g+XvOfWdp2g5Zcf3eK6Emg
t8JiSrB/REZAuZFiach0++BMOUQs1vxvfPkV2jD4s5+1ybVImx1ugZtkHPS1lj/r
LO6mbVJV8bTIIy8ApHxL3gBa2lse/j5cGgyjpw/t+dV5/PuGM1HdkMmUNrJMm+Nu
2i+yGqTrPYYFX9WRTq9GLK2afTpxSbfqZpU4Vugti/wQ3XhK9roS/LPQM1IRQCL2
A47jeAkaNKjTdvnCZ0LlxcLdtOrrAOkxwGC3WR+X9uDXxJRXwNYh4PuVUfYthdMr
WXAaByRAX982j8ozafkPIMZttVXIBegbwIpnzfxny4geq1lvqX3qU5wDBh1linKz
aRYM4EAELEToYWtLSpBzIcsZm7nFWnP+XOqacUWejQlqDxyKvLqhZO2hTe6j/KEB
dfj5eUQXMKm/7qsu29Irk6Oou/Zy+S/DpVmZohttw00jQccJ2kXngJBSdJUGdRiE
B76n0nx0VacFBFk8LT5kLveWlFyUxte8j+OJlwMr/Cz6NPa3ahGAW9Qk6FhZEtdb
dlPFvtamkHIqCU8q0XLcOMqZBnDC0y22qIc0j0foHhMmZgsKow9MBwqCZsCDkKaA
BxUJM9R5cOWYh+MkhpR36nhrOU0tLSg8p560GBbxVpAGacS8yqMz31db43xF5nVu
8VRPCwia7thFIRe80BvagEUWXuWZZuk3fwhrObySyJ6BCrxhQ29UQ96uz78/apJ3
bc58Fhj9lAxmpJFNiitGjkiIWYt0NNFWAY0C282lkzGe+LsC136/U7chbOwh4icf
Cy2hUK4+S5xv/TDdhLseIqv4WYLENBsVWXbV4dBx/VA7s8ilc8lTp51EKfsYJO3t
aRZbEc0M7NHTNcA8vTaTMsSSkc3M0SFPMqbg2CuSxNrJMkd+ZFLH2ia+aKXUA8Vt
LkP5jpvVH94sTP774f1MDR3xayuRIoK8v6OcoYKDAn8UbAEA/slAuxR2su+bPRIf
ZAjJkMW7qcubBzHQI+U0g5sX+zj/iD/JWDxL/p/o5U0KMKU70gz8lJRi87DKdJPw
OYz0DzJZKRtDHMaQPh1dxrmbOghcpyuUD35JufTsaNbogQnPHpVrRCHhaMsK/nv+
Hxut9XGGd4V+19QXs5IIoGY7RgAQKr1bMaEHpYKTLSGOeBwDoJS+lDwOWbqpywVl
pUne4fhYdyfcHv2ftN5sd7rngo7vqrMKz9/CituH2Mx+ENTX74pj3NuyLgda4cvW
KZQDsMrQPZ4QriOoqbFydGubmAMoJ51irnmuJflSmVqKHwPqd/EYvx3OlecFTRPw
M3hAPVJ2dbjNl6HdTeb/FCs5oZz62Zc+BCCllzlGlG4XqSueZeTUaKRc1DfFEDWc
2fFTTyNCbGM+MeC/LNrlhI/Z4MibkxssJT6cwo71rGexU885osOaYLIe/FuImJCi
BFsJ+VEntYWyufwS0NT5lkMwoQmGCE+pJT0jclGokADnPu1apSpE5Akk2mePwaBY
IwgIsbB5G7XiGDojuCxUk7brNdiagsXrfxjA0OZRpEKmFQPFgyZ8RRsZ56pnBW1D
56l9n7ttx6+r+HMrP8ADDSQH9lRjk1LzgqQgXgaNd1G1cGuMXxpW724cYFvCrW15
oHgkIEHmAp/RxJqPjNAINU4INsSXjH4At0IQDrmZ8ubhWAZJIgp8F/abZohAwbu+
dkO4isDyRw3Nsi1irrZVQaRiuVuZWiJON4SP9klCQ48pRTU35raLtnaC1odEfQ1F
q0IwsaZELlJvxreL24/PafvgN+TAQU9dq+ZqNsJ9db5zTczK51Rmh5PyTdsVSo07
Imm9OfYBhl2eNongaVxjW+wSlXjAp3yXEloQRv//VpLjY31fPe+O4+AHBFzjICoF
pLj+2gmRMuX1MBEgSTJJiTwuedTpdBEOtpWOtIZ7FeYi4iocgMsO5NCF9EG36UTC
cgRm8PniU8Tlsi9NkZKj8E1MFKYegqF0kmCsE5W1amwqOySUN7Yh54aVTv7kGKlS
7ndi/VnWt7GplC0Ls/yVbDxJAdtJq4RmL/gSvS3IZ6V7TKy8gTkFpmHS/Wil66BY
KVgYh16vO1Bzkx9O4R5XH9ju+t9UA1LZ52m5xT1PgEJeJEJKnTOnmu+W2qcEesBa
aL8/hrXh8d+R1XPktsGAL0rYUQpwQK+UrhqoYLdRSucb7GIjjEqMIku8dAPOenOm
cmg+ji/dibFv+JIoASVKIxb2EhKkXSPbBljmny8pRN5qWrxgcNympwo9WCpMMxhV
dVnrEM/QT2D05cpTUlUmSkAVdM3K9YrSQLPIkjf8Tbchk0VBUG9NqLiNtXl+5eRF
dlJemkNhSsWkQgAR0wWwVUrFIthCivQOfjVxwYL3p6P1JD/eW+dPQaCy5klDBNbn
GBonKNFbdgkWYlV5gO+gLT4p9KybnpapVtPYTE5UiN9xVc9NTzDj50R6Kl+Re/R5
SZMAXTsODSPucjVxVoNmLEdgd5noS0eVDXcsyXkOhovI84D0lygjowXGXNtqfWba
owQKRnAkLCHH/RSLZaOqy7wd0on1ZMX/BYKAK7G3ZsUVXqpvVC/R8KTlrd4ngdO2
Wf+Nw3QpZiFaeKPflqWt22OVViOjK7DlzgTE00wmzuyhbRM0lkhexAZjXZ1Gu4os
LRuq5T3MzlmaKp2bH4UrqXH6MLrD4TmHkUYPqB/z5PBa+nh4mXz/CtCBr1z3JTnd
cyEdm5On3vYiJZiW7Fa/qKEyU2/DnimEVf+XjTO0+dPi3Huy5p8FFU/ZNdtUnMh/
2JuZ2RomI6ar6GiNy2vYik1V2rsi2aeKVAqSa/MdpUCf/T1kYzmhS4k5jPM99oO/
3nSkt/ehvOSIAbbCECiAvPG7stXNoHfDyBMfwUKWf5S0Dzez4EqQV7B66m3vOrrQ
OTcS7tgd8wlDoxkg1YtPGkftNG3nKNR7i9w5mkt+74s47QXMtSHQ/1QXK8m/xhJS
MpUbgZU3B9p+H3kgphYPSc9zz+roSKbIaiF2gDkD/UeGJrLsvUAML06OJyi3rHxc
VU1T6HfTqKupkFMjOeULxMAD9X0JEh90UfdEVzvdHlLNwO4UyjIZEXHXLaPyZzoU
FvicHKTjtrakc96AwaS/+IFpXNAYjRw4P3y8UautDlj4U85ud8T3D8r2tMm0xgmb
NiKE31Xasq8l1SBp4Kdq0tb6pjXYVtFN/XoQt88LZvoxzO2AcCo4AF1jvnYp+JcD
1R+qtej7accbEoykcMoXewZCiL8Rc7ph9OcLnDogHvWBJmnztFAGa08zKQ7mwppj
hfKiQGoXFPJh7nFOJVY0gItwI9FtLzx24R2aAd7eTsTjs3wRinC0LVv92jG+WmFt
3WwNkTXRxsStfaxeCVvdP/5dSKI+I8Fgx2KoznTjHIiSsjYFSe4mZtieEXLLZdOa
2+TA6o/5+6n6qxBk7f3E/tm0JjLxHrLFMtJpnOgmIp0Vjt+9G5jJ7qErpB0DZXSN
CYoeu9G4pmBRjkt42sXxOlEGMU91DO7CgXu9uj80VMYORtmLMnqUldd9QMmj3heT
BjZA5Iuc6tFyO60MvNybLr84OkHxNpDaEE1MNZgRz+g4k2GX77C2YCLbrYCBPSjj
EYJSz7rbwgiuxcgzEtH9wIr15CmNaQfm9mtanXFvRbJqZkMC3i4188/Kpl/voJS3
jiqVFbg7+AGxe6r3ayIX9i+XQIRMewk1zcSQm18hQK+E6eR8PBMEfgIDNSV+4vrq
HpGff1JOCwQEcgD0ixPEHmGORlXU0AioQmfjUCn4gAM3f1Xln52u8rvDVI2tooe+
Cg9kt2mCG/V3EoZ8Hb4kwBZ8FRxf8UNMBjWIwFvxQCw7hhBHG22SsW2bYHPqkXcY
jyVMAinigzACOCJSCSjNzrgrkQ2PHFPnVUPjSJjzdp2Wys86r98SqtUHgZz4MItm
Zr1xFuPTjWcGHKKWN5OVJmcDsJsO2Dn/zylU2wHDjOgjRZ6+c2c9WchxkkpZTTfu
6J0FZJ4f6JhDdFXmiQ+HI2cTQcgOpgTdwIS3wQPkfPwIsipJjjCOfxQL2TUIethQ
yj+UHwC3asrgouqzW9yztnpI4QG3yIn+hDcJQxS4niLMwIBW2W8EV9nKuh6UMt7s
T3QNke1p9mwhF3IY+eumgb02zqOtwKyzhIuak3z23c6cFPcVAiQGH5Z4KUD0bNvx
+Ogy6SFTBC7V50ZICfbndv+es18gGpYpulbXNv9Rrt+CG7cqkHgLBzsp+7G87El2
ya5ui+Avj0b3UFzT7VKSiarIPa9Ha8i1CgMhfos3BHRoX/djDEnvR67Krfg6cvYV
6L6k0CTS4Li8KDbSz/cRZhOxdJTXWR08LX2ZXbPHtrH1BXY8XI6wmcMI51efiRIv
SMspMjYOuIEEWgJLyxq7PPDKH+53Egr4W+qm2WIEEff4uxmMYuXii2Sf1Du7Pdce
umSQ0goYxX+LYa1u7FOKVimJkLoEpzFXoYhjSsylppbhqcEeXfmQoh4v3DBFToap
OFnrEzjMt/uPdXDzNV6pBAdaM92RW690kiXTiyRwQFxcoETsjAYjcq8cA2TmtaEp
Y3ci/HlI1hVEGchOzETzsphI1H5AGSxDByue9yVBnVCmTtmtXBdZODmBB3AbC/AE
mZsDv9ei3rCyehwHWQq0GIJknghvlE16P6pPd4HQvmbIVuXujmgfmQsvFxyjknpH
OifnelHLYBFJI7qLAu+dHZ+4wBKyqoaJOA7v/077kZtLsuGIB/vAjq+fWOJdnATg
MdAoFw/FrradjYBFMRHwSa/wYyjfU984nyUteC/TguChU4UkK3Asejr9PAn77ZH/
niQ6aR74uF9t4zYg1EvMsHF+luMHs3poaux5maHMfAbXNLiiM3pmzigfaofCGmur
I6ie1lVWrVTJZvUdVk/cvZ49q7Cm9nP7I9OLk/3FBtdMtYN0UjRqq4OKpqoIjh5R
XEe5B5F3jBhmD1VSkJ0tC2ekeY+NRb7+PBlP4EqThsi6TJ8lbC6GFZ0NPEsEdt3M
HRw41XP59g2g0oiK/jJfsaYghbuXiUa6Q84+ifGe33dFhtVdeYxFdBXxAX+hl6ts
8ESxKGpnxpquWWmzVy2ZnGCIcmKQ8TiH3Ey36oLntf68VAalwpBw9DI19EqF+fqv
i1nUAiEt6qJOW//+T36/Dy3Er/6gaQv3pe4j61IdaKu9yjUm/2WaSS1s/Tdn0V4y
0nZW4dmSUSthS3zcH+05Ncc9ALcO1M5bkan3mJj69z4wOUWaHO6UQqOYH3unk3B0
2v5TaM7ijzA+uHQlmU08Ixk8/nH30Owc8MG0tXSJNvozJ+75dV2/HdjHvKwKc5l7
Cpt2sdklpcosrr7Gjf57SynBSP8mipJGiack/5bTGptWisSaI5i4BgeyJ6aw7yfZ
WzyOU5GnZIiHmi+G/qG4r6lplvioA6iKzR+oxDOpcim2zkdETM+JpGfYz0fdhBwY
Q8zWW3oiiezBcCMYKt9q7RujWj7ktSApnF6YHxtrCgVa+n98G+M7x5j5vAs/CLXt
U/B1gFuWZBEc4gCBHriQ2AwIoVpjgYfAKr5fHb2Hl7fYuNpcaqr21dIOsy2c4x7x
hwGTBnmlcXGGL20dJQVCqDDxfmQJTgcx2hsMQp6jVpPL8kL7RfRpkScsy8rdUlQx
4wi1FM6PwuCbX6whMxbqbL11ttrIIsYA/7/NOu2/zJ5+OhicjDabPVlOm3ZhhLO0
zh75/sQmfycMnXvisSNZZ+bRL0hzFILOXjRM4uh5u2yWjU9J5lF/vBuwl9tNKOEE
g80EaXkSJg8CPUVBY3vO2j+P/uNOLtSHUpgfy44jMo3v956FRemuKpnD6x0GVZXs
e+c4QFUHfxb3sCcf6xDEKzhMeK9gpxesi/9//ocz03G/ipQCbdHonKmQZOsqDNZw
OebyJPVE6qcq9XErESASyzK8kIo6dCxRg8QzIMlGmoZ6cC6mQ5RhC6YVWifTtI28
2p3+v4N+UOF5v77xdzzhBSe5H1jXBYbYcQqbsXuZDAkxCu9pt/LbELkntMH+9vmN
DTL6wPMrXCFv0jnRiAPMljGuCnZ6E2p4vDM1+7zhRQ9JteRceZAnidSLWSO3a0Of
r8Kio1G23AAR57B8eVub++QA5sfLqZy4woFohSqzCN4tf/zZu1lxT3X+inmtjb8T
w/iXh4LLVsfGiwPYVufw+6w2PrT5Gebcj1WebqSONgUDFMyKAjaETD0K3agQHeIe
wAcrL+3ztZ9bZKW8k7wIOTuhAOkaKEGqtEXVAIJ52p9MtmCb/kIXnifh7xEyJpPE
JzF4ADMIt4c4AgfQlpYZV3tlpAVpAWuxzSjgY+GZPXyTgKmZfzAv3rR6/EWnnlA6
YP2Ql10zkBm2/KrR53V6c2BlzBqyYM1hjbPyUjaENrr/uIE+4O61cCpsveTJ7W3N
mZXpJxlj0D32pdTNjZ+EfPfgGYK1JtJ1TYXa3h6qp4YJ00xM1aPVyktK6mb+37Ti
/IA+KzJ+KBs1r+GsN8QdPaRflxIkhxB7cogVy5pSvnJVq6KzF6dtWesAsCp+av6f
FgYL0xcjrdzVk9yz8oF9McPpQTvf79S478+4/2DCzN166+inLXQNn2ttrR9jnhnL
OPM4uv3bRFF8KdltBkG4thIGQZUEXA4bdAwCNMM2V2K4IIkNCbnRzaTwlqAqhE0a
ThYo3yTgPMtw8oAQh/g7vXYLXFALxCLEuoMyLKyM+Id9ysWXJOUAuqkLKQ1pbG6v
IZduVyi/4AkfboU7NbSKPREMgGqFLlFKw8ALLgFUsxJLOIhP2+6+kNwBnotflxcf
GovH0D4Uk4axGD3BMlCpQoGd5h2j84xdyzuficec1VeIStMAa4LAuVuHxRKe3m/a
dHLj9XFL4A/NmFe2usZE47uexQeaoFJNK12EXo8DbIJWJzxZmSFWoqT4Q+EvWZDr
Qf9TNbWu+QoaTNHXlFamo4PVUtGMVizZtN5Rt0ohyIr551by7hLGMctz3fj6rScR
HbcugsOrh06nHbsL3VIqy9eoGwqiYXiqyjyqV2chjvJFV8y8cdCoH6KntW2719Pl
4RxlURa+G4uotn2FkRcn1hbfkMLyakHzocBDPDu9Jw5y90POoWnv5f2G9WHaOs2x
OR6wBhtErbqP6JPosz42KZMdnLCwGhkSRoZtUfXl2R8yRJ5CjZsYV5k59453btjn
7VrcIiI7IvKyov6f0gfIsn4Y+n3iUVMLbF+z1B4dgCRpzBHsLS2eUdMYkUUc1y12
YqqUmB+KN++lYgZzmw1XCp9yFp/rBIdT5Sih/K9dsyIDagtvjLBNZ6/cVlqiUb5p
0SV+Xr1ZTa6FVU1AdcH3IaU2ETopbXZ5Wc9mWoQ3sXxOsbzzNheoDImjcXjBI3O5
iwPGBP5PqDFPxnKu6Ru4Igb/eSr4jmCXAMdxK8E7fVpbQ0TKa9alm1pEfQrnMGjc
NfXhYM/yWxXuBnSotiIFPSrulDHJ6QcbtGNShFVCKSezcarYzq9GnJWb9bA+LhAq
bfIsArGFukL/68OySsVFTDwWSie0eKI+CoLA29eorRPONCO7adVAk7rWQiVf9LNH
l8eOe+7VMqvtWZ7RJBNUnDxL/g7pY6TwQagMJBcG3R+/MJvs0Hloj9RoBEx7nb2D
Uh9MlHdE4cwUfJMOsQdTIt0uSM+sYqSE+RM9t4RmgnJUiw8t0+V+PctwoD132IKd
NpNSlHrXsRlQd8v+dpyWnvyt1wmcpOXCnNN8r9PvJA5sco3nOLmKumZ5EKpmtice
KWgBIUoOr+DX2x6ab/B4kRxu3t3VjZXjqs6ONtAllW7GyLURtBS0bfS9bdCLouUr
bAPaSm4aIZQ64wjhGUjCIazJiovps6GDSOUMt4kxUEow7SZZkV6MGkRBos5kar61
B49KkG0JGmUqQo03YC8z1JWZ1HibHUk8mLST2ucANzLaaOPoxQcpeAsk7CTSLw+9
xGqQzGeD06hJS6uB7e8AH2z2zSllDnKYYOMMp4aYGOB+e+ucLYDG3NAIhEKP8OOd
4uMCMMbPs0hg5ebkNnvjyoADm8A0tx5jQ9Xkf6fYNOn3s8qoiG335BbdC/Pemk3j
LW6G6qwRYDW6YAWWZhw+BHpjJj1b+qilgkMQ1ZG+XmzBkerClg4R7akTJEXTtY6T
MN0/L0c0KXaW+XoUaS0mIL2wn69w7A2/0DJx7pw0DxgkMtSYStItAoeaKpsq0KHe
4p/l1ZvpNdrPNax9TEIIraS3FxEy9GVIUWyDfMHqPSLFxvl/vLC40ijevMOk0lpB
cfej07UUpdyfPCh5NdxVhk4UezUhyltFa61u0CPRUDOYTmry8QnlSHcPy7cIY/g3
3/Th9r51JnIVZTrqn1sAdZnvQXvVqlUjnEw8C/OcvPcQyJx1FMnd4s9Dz98jefxX
0/2dDjS8pLGFaJCYPNd62rO97SIGiBtJ7CMvxbbuFfboV9jYbdYRhpi0c6sEr/sD
NmNHuEcA/wAZzpkZoBFw0iqoDub2H89qeLzoliaOpFl4hFpIaDiHLVSXv5UqG7e5
Qis59q0iLF8dBxuBkf+JmXayfsgJFAiFJtLNbm6NpO/ZYXMrQWadDC6uPlvfj4At
YIzvkf3ItLivRx9wZlKG5QYwyLuRBxZ+PuNiIerb2VK877Ki6h/y/GcLruDcaLMY
MsRJwXAnMIKe0jObADD8EofukSTj/8Q4Tabq/0Toe34GRG5OQv4HGZoHyljfHt7Y
O7Q3uPDSpFPAjsWjtWgY59bt54QTn45pJS+yrUQPhjGem55mJBpV7+ygf2XRRfBW
uVYuCc3ZTz03DK6bHnI+knjo30La+dN7NINEEP5YmWL4+eQZ70FqLJW3xuHUhoBa
/8MQ9KB7uaKqCYVQj4Y5HZqxUoYOsnSBsKizogwNfjP//8Ge2FHRqnQwHFONo0/b
z/kWS6kCrX0lX0ZRyRp30Z2T5n3srLGKyreSBvmxCtexksfrXoQQkIDM+jrgFMh6
lV8d//X7YQVPNHUNzqdNC4V0a/YRj0WkiaO9gHt6hh8k3Wv9n6iHbN4nDSSbe0vK
WObgiIN2dY2mJdDKr8slb7aLP3IQRJKXBdg2MdHvutI5/qm+bf1nWcKDovBR1mBn
D6SDVWxLnMg3qDImuKee8O4+uoK8J/V8QBG422v40xBEcN54AdOUUlwmsJYNNBQm
SOMB3TCepBNcrW1XGRhgF+ya2P1KO0tBvKk8xk9gt4ASOxVQoUZPtXkwqeZLzJfZ
odEtqXczgrccLxIKFLw9Cn0u02jly5G7eRVfJQnjat6yTjbyacjNQVM8YYnBFkCr
BAwwXkrGr5QoOrQlyI3m1scxYjpxJjAq6gbp+xKKNjJbkNXYgBxH6P+GKm0lTDl0
LzDGDKun1tyO9Odh/zXmSKyAdw72M8fTCyIIN2zUAJRMdOT8erRKVLw41dOi73VS
l7laigCz0/3k51qklR+XBci4T/+z3UVziuzDH3fDX4lu7lSgl+kRzvW7+Ng4dnZW
jOGOUEKqzAlJD8sFewXBZ5u7KXzFJOrKoTku2wU3qKEZPOJTKcy0x41m5DlqYPnN
ebyeDDmkeXytSgt79j748HFvTsK4LmIKXtrrpsq17aOjdjjupOJ28dc4CORuDhhH
LA56fWk8rNBhXqSVsRBd3xkLLbH8S1h5WJPKckKDTMQB5CZ9Jo3MmAP7OdGfu5uX
LOxXKp49zHQo9WKGXGkbvXlQ+8DglBxzMIXnmIfmj7uKO7tUihNW5GzYpu1Ynnu6
hTdnT1x54DO9b8bFcgtyHcKzX2feCW1CK3FB0WQ/XhfIpu6seyTneYPey4w0YZJ4
J0S8FeSmmVXEvrISy0V0dr48ilDGeBDN4YwCbE/lfIzwzOaFzpMAcWHwYMkHjZ0K
tZe6ItbF1px0SuJQwQYsz6Otu8saEv66oBob4oIjfa0BEKyrEoQY230BmHxrrqL9
2LnM8SZ+bWNGFrCzmoV4gZQPwxgnuStJ2z5kIeTbum86OuUgLid0xADo6Dwz7FQO
i0l6Qwrg3BrRLolKwDeHA+86xCJTm9hf5USWO2fwQ9Fo1WEzhthxvoCEvPwKRIwI
Bo2C6ys2ZKQFL5ByteD9ustYCg0fUzP8jUhUcx0LZ1bXkjp51TtAuR4ezeq3VHny
7wW11c8EKWDBrDyWH/K3HfAgVqEVZE3yihu5+7yi/z7CdtruHIW71Iii81oJR4PD
glw8+uVJxaIxWUHgFVK8kEUh99bpweDo4ZUKwQLx/xnYT9JBGJRnqubthZnu84LD
KUL4ET9xJxaZyqCim5IW9wPh1lkU3ztDK7GjBSNoKxFtguVtqeucZLwhqVUi1KPX
Lp7oP6kpSCxrAHGUVE4eSYcjWZhrD2N9csxiDmNWkGWk/mylzWaYWpiF7edArHfx
/X3uJWRfqx6rAPwXmXQD6U/+zQkl51PtwF/x25cq8mSl8/MRF8fmIoVn3wkKCnIV
Cr3HlKJLYfnwks3rUhNqqNV+qHjoItyl85IyW682M0iQbxzNGSear5ua0YtxPR2/
cmjRRCkGnyE6mjreoCqTSq3p33hUQjJuGNoFdKzw/IHGqjO+dcnEap3tm/c6xPMQ
2ZnrtYIjwGXAhijf6mdzDigAoqMGoi2xogNgOAc5/09GRLpz7S16c/il48FnazuV
JKYrxjuoP9dXeUyiAvHpG4pmj3rSz6YWMdxHyWSATjvUaUFu5/ayM98KfhLxSUTT
6IYU1lj3y8+Gkp9DECVEss9X5X7Qj3hH1O0zEAkCKEM5QrEyBY+XVKZgUyGN0fa7
pEnkH87JhcG8z2bbwDUdshsJGIyx8YAd5LyIZ1n0l/eBrBWomex5KP3TNLTmM5DU
ZQgp0hM1kp7Mq/3rUAwC+JbTzwGs+axVvx1eHsHx4HYyAz8Je/AM8htUkNoPcIGi
xqRWGQRz3n9+yInc90p4fucnOXey9h1ayT7FXyWwZkpRngeftT+Ld4d/OqUHNUGR
WKN3ONyLpdEnZ3qcSjT2WCK/EmR0kcrp3Ex9F64oH0tGge0BdIBNnk5TjOcGNzSC
uclccf8ZEqDY6mtuKaih2/s7Fgim5jiMqNglKGF7t5ygXL2CFsfk0uQhLJTcsZLr
0tNX0+u9CQhn8DN4lW6yS9JLBbY76w1/Un4EJKTqpZ1slQRlwe7w/WeRWNK5FIM/
unQXfP+g/DG91HBtcCE0dgeTX9tg1cra12ZYAGG75gXvfQZo3Q8O9z7EmXUOQEfL
ZCP4AhMd+vLsSUWbnrr/EVZyQw9OomrDSVb+NhnxKnNoKui/JaM4Iq8QXAOIspFo
s8WuNjSU96DheZdCbZr7PfGiQN76Tj0LvWWIxNSpBlXxKw31R9jjpiJnRVZeOoa5
xiWgXj7pOffeBlwvLHAOp/k7AtQyt5YQViLbG9k/Kb+0fM+7qA0CabZaexTQRJY5
/z0oUOYfR97qqEP58wco2rJ/qwTGfFyLpVV1QhL0ZnC+W3v0c6uGp8C3vM4BgsaZ
kuYm9hnC4KJdR3TTvmOvkXYGie43ECPO/1jzMaxv91IejheG7WyTiAMNYbN57woW
6jxMfgYPB7nqmTIRFOExGfn+8260MKlQGD33baeT1BuoZg6wSLu/SEmyhMY+q8Wt
0s0CzkYryCRtnEqwve5OOu5OImqvbKKdYKaoHMOmGm0AvwEhtjYICOLyWayJhSAq
AFadrtnkhULGxVJ5j4vhIYJeeruh67TX+/8pHhkQsTVJGpEEsLe48d9w3iY4Op9H
qZpeV9YmUKAQQF28ND0hZKYD2msHOexGZjl8dsBn1msjRwhILQ7CQb/ZtgaEuU5D
05QrGmQyQUH1EChSiUjEpPyNuYkm89jKAHnsQv6Ba+Ub+fPF7CfR5jzKpJaYkay1
xU+LNK6BytxWWXdqIJjMgh9c4LWCZtnUs3ndUkqD8wdMQ/PMHBzNjMZUwsSzLt/e
azXztwjx13SoKZgZz4cjDxFyt5SoD9v4LeiwI1u9S5nck9mv4fd1Hd6NuUJ5iXUM
BuhGuEPTNilEvcNp+RX/oAlIdthcvwsScjLTUDSWmeTxjH42HjjX7bRjabaARTPf
tJ5/P3il5K+ramScZEP4qPJwCrTRDT58QvQ6jqKAWxWfzk/aoShCjA8iu5EQaukV
/DAoH1aH0URHwRoQ0MN6DiKxrz+kPoHy8YR+MHS6+8snqu/vsxIVSCIPM7egI5cF
nXu8Tu+faNz1XV4Yf6VDz2m6GoixKhSLD4FvVwLvSVryop5UnChojVLnVx/aN1Z8
rAZyjOU9iNbU7oED2TEEwwh88dyQVT9XfNFZ/1hohe7uKI5vYtNUAf0cJTrPDrYE
1ubZhtipvXOaYVyuM63KUX5B9rqFHvYgfGv3fH3JmjIL5bK/pYfgURfFLvvk0cW3
cqriVU0nsDAG05KhU6Fa7M35K6RqieZTaXOGn4nkNFWCRluR7ggyDMz4Fd/JLLZM
oMejQnN6ipe8xl/rSrQtKrzJ+2xVECgFnVyGFBcOMi+MDruotKCQDhsRbCYpQgxP
1SxPNlAvjjfaOPJz+nJxro2DOMM1nD/b3jCkox6XmnXySmBa3A4gcsgJ4kDVP9Pm
WWm/qt4OOGmrRhDas4jCaFFeamgRJZZCUD/jpfcVB0zeVZYbNVRfJaBlmM3cs07K
ZdFec9w+QzOh+s0+3lxBTzByKfQK0EpR9jwkBFKTeCIknzhSXn8H3J4rQt0X0qPC
aHe4+83m8hQHCZA4Q7RNFB53l23DbMmUJpbRCi9NpnmLD+O3syKcqd107gnRo02k
cGD2t6jH3FEF+ydTB+3OCtk0SPZz9zxFKpzn87pVd1MObYPr0Zy6fO5bAbZJpvFl
ss+BaTda+UXGUfh7UBgDC2FdcHbG3HvWAYYXmCUloLp+YtUuag4RPCqZHeOZMElQ
Y6f1QnhfFuuiOLhnFq1AByAtxZe/CMgLRKm++vCikNOv2V6/W17MdaLWbyJGP1T3
gEQ4hKnfSSO/Pg9sZfkqbnys/O45Sinx5rkIGDDWT8ViPbVDk2YKDKO5XOZZQZSm
WH4VNXRKWL6F5w0uavaEiGYmHJ95LpssRuOCG4Gwdu4WOl6UGqDU1f/8RZbeb6VU
at7kcq5/vdANq2SdbVqzyZzdxIvdBd/lYDzx8xNChbj8x6PGY+VLjllb5xfb1B0n
i281PBop7PcgsejL7N3fGCn8LHpp6TYNdVCTeWYVHeWajWZqD/weref2Gd0Lki0d
sShCgG6HlEq0+s4NShbx6/+vsyyH3HfjKMgA6WreZyYyngi7JM0BQepoUPNHfZUg
xRTsW8NQ52YONrmtRspD6HPzfZIanAEBKv6eiO8VOuQIN1OMIBULPm+nBSlshLiz
nBy6ujqc+nYX7qacfSyLV3Emo5KqMwBvAj830hyIgrxuFZOqCmnNK0oNSmESL6oZ
1vE5q2bZbjXJK7ZM+RR6rR4NiruWGfWg6x6ED+lC6lx0H42I2bzKQFpSx+lrPqCz
MFuStujsk92WnuCZgmX4r3U/9J4R7UatO+6oFPU95F5D1hqgsGXk31PG++ZiIyZ+
bGCYkyl5VHFSBrr3dHsnxlwC+zZj6RVwUsHmorT4NLMrUOzkWS0gFcFLR2J6Xl/E
WsbhXllHW3B//dWVj2pDiivxrv7lGTIuf8TSBXh1Y6CcUNt+wPRY2VxocMninatg
GyAEQEOjT4Jj3HcTmydxE5acDLdsRzj7j3a/EaucGxhadRwg7A350UGg+AbyGqq/
kPEZaL09uulCqEvm0X+yIGAFO4kRijx7q+nz56jwMmavjt6tfsEx+MrnrcjOnx5w
070n02+QAlgZkWo6ycvW05Huzai04Ad89J5MF5iKTEtcW7CFtkX9l6eBr3ZfzuYo
gU0BNDh+ACJNKH1JX60wfxOtOIt6/ow4OJmQaxpnmnCnqhgxdB+E6GwcM0qfWxIz
V7MP56VPNMnb2hjDZPYlxiLxRERAp3qazjQAiDeJf6aTQ2tiz1JsPu+4G6bJtxZC
de9lbdKx5VqOyNuQNOZM5SjnrAt+9d7OgFwulSm7dbRmJv6XnQ+EmZ3OGiJOxb4X
6r6C4+A4Oun8LjZqTg+I1NUUdNtkrA9EtmDe2J2FD/S0Ne1n+wQU/qIu/IYBoNqO
5pUVf3tV/aPP3g37v21lpQ4mC5x0Vm0EPkShlpVQhdG6SDGox6LHWeo3NdADts3Q
AX0CRZrnJBqod7M4aaGKeyJZar2ijbJLQWcw+4f4Ccctsbs6vgMG5CD7noZ7Eh+q
xQeMV+/KcMaAgqFFEpGQ9dwcdWBoySEpQmFAn0z1YPjxs9LaIJeQfWhZM1azW2dM
RghAE+htKuZbmRkjgLOpWojhz8l2pVowZKlVPW9o6QpnrmGgnRA0WEwxm5dy0h3h
jXcnzzTdqlUqYYfAZhGP3ES/WQxOarlU//BObl7Ekso/af570MVZCbhRynlgJLb7
odG+R0WDz5TpI2vwKA7Np44hPzJN2JPtLnZ48mxaYxB/7GSuPPPWxC1ADk4rUhfJ
8sJOfV2zlvWg12Vymel/Qwqki9+W7LRVMzUlXlNAzjMKWGuWqEbUy/dpww+lBrrd
MfKzUyv8MYqomwIURe5dZ6YJ1ZzYQXPajif8oX6WZOcLFL3YDNyhj2cjuK7TiAB8
Ix+z8fcZDHRUG13bYDOr9OS9ASOiaWXDRiOVm4GyIDodzM8zHmga3R7GHOnXrMLP
LB5i7sYbLzIfeUWo8oEqxpPBRlatyb/2OPiL0ILBua+prrFePPcjt+bDC4/xTv65
SZDZE2fHDbLffXxMFRSoYhV2tlm+cU9R57oi7GmVDE0cJ/24g+0E8ouhvaiqdwaS
icJ2lsiW5n7WxhoB1lN1YLypEF4ctieYkgH3MuX/sQ4CmnTE0Ub7dYVLFMi/muw3
oqzDFTAhhzGf1wl6fmo5nd1hgt41Ciees01IeCdEtA5CRpgo250P0Qrk4P5Mm9Ov
fQCng7zhAG6neYuv7qwH/xoMegWa7kiwRBiOCaNU3oUOdUIQMPuICSojdGTcgN3g
YTHxE9Dd9P0KsKj3gaLKBpaI01d4Nk9vHG/IcXARCRYMla44wDfd+rg0rjEvl1tq
9Yjr/O2bblpiKNqGx0HrCLxgYU9HC9pyg1WsmnA4z70gvh+v5N01mBjDfy/+Rhac
roypZL/BrmaJbkoluWhXuKNpB+6JAryLCnzdgdYnTuYAJMtXs3+JzwQ1rx0sHp0o
O1cdGE/sCCeBP2fydtnFKoOc9OezSqmV1EhBiUHobu7IP4DnzhCePVTFCq4Vkwfs
VJ6eMNq9YXKgJwKX6kwEtVl5b97LmDD2VNwAuw6j49wgsXtBraCO6K9K6X8E7wEf
uSwBVY+e56wyf3syso6nYM70NW2307+D66CfgWzBzk7jssPUbYzoWH/zspkLJrzH
Li29YMlhyH7bRI3IU3g3P2GFWdGwWgl51gTBmOVB9uH2WKBWF69hNTWA5vMt5+fB
obrkeYpuh4GkeiiXryncuIs/fnwGsELIZ9BScMPhlmIdVDuP68C/EquU08w7mYRK
bNsF7zSLsQ+Q/GpTUXQ7nvxtWuDCmCTgNugSLzeGnOe7E/dWG3sUNQZeIo7OAaS/
JiYkGWoOD7pRHXeLgOnPcFEOfuC1jBGLZ7do6mK8EqHPLoGje80jPHXXyK26R9rr
ppoS3iiDMn4H5sSsCWedEYSBn2+xzFQiNQBjd9Swkto/aKi1VkDQVkWi2uZfuzd0
F4lgzfwVrUYI1FeGphNlruizjgyCUP3iBgCKlsdN5D4LB0HcBRyI1Ie5ypNkl2zc
0worFRGpKNCTRTxZ4oY8ufKYB1KY+jYxE1xRuiCxTviizGIRjQ3ap+CHraIwYhHD
0v3KBn54XTpoy+7sSs63BigAEiZx0S+rd5/ge0ljkcOfTUuClzX3MSYyzVk1SJT3
hburgU3ZFmUP5jzVbhtfvy7QvHje4mGLtM326zAh3NYhbM5VrF6bm1EE2wv5nvvt
Eb6WnTC0WZ3/cV/bXKogyO7fUQFpKr4q/cF6bryST+ICpz5L7ifyf3nvTMQ6sK+4
3jus9E9MuEfIahgGtc0NEpBY9L+Kgx0T4EfqAvGJeYXZCefrae1roSX5j6b+0HUh
hL4MCxCZsRdGefPXhNoRWfuc9beJXRmhslI0XUfDSsNNz7UKYLmMAt5vyzZa245a
AITf0D6WQMmZjlVy3Ab6v8da1ysTRZIkkcjf+8k8GhaP7kqWTac7tJdEMJ2Z69IU
B8fLdHPYqlxsMq1TRqy0Y3fp7smbOxURkwAyVORTnO+iMwDp8hMB7P56jIUMl4Qy
6Ts2e97KI5O1amZiUOoQEyxDPDE2hU5ik7n0vBDH8fedxH+z25BCdA77tSJ0eILN
lt9jJ8Z7UAkoTO6rdtAAuCvNIQGOLnOn7NanFWwSogSG8QJsasEQiuRy8MSkY3TY
j+ElPbuBylgV7nq4r6alcWYt1Pts4YXG2MNW3KwSy+o/66dAimSI05+SKfqWrAUM
ovzlmmesXYWpI1DrdZUIJfZVgoLp94P/ATgHdAk5uawWQOzVW0VjwIsr7ZVSBLqt
YN2ea7JZYAfEqRBgduNoYZT29P6kzAxZp/lE+Cg7YeJL+Yitx+J6U6PkRygGlyMH
/Ry2UpVJUYb3YCC1urDRxiEs7vjGPytHw2DTPfnShslQSQ1ZOL4MB648EjZ/MkYv
h433glg2dJ3TAYWIQGeZN8E83nMu0WIByywncMP/sdiEEsQe46Mz8YvEfGjFZyOh
dwZsr8+uy790SJJAuGTt4etpDUHQ/d1ym/F+rYIujlohrYL5txmnB0E0t3GyNNnu
EZ1NpXAF8Rm0CDdTqpxKQ8rJueuR1gWanyVzxX/wpyOF7EHmBHBfMilgdA7vsLj+
1/TzuIDYXTH+h/1cpc0rVF0agG+vm2iFpEvPyWgGu4dbkGPCJiLURZhKY6hsIIzD
CKYLUbA7SnFA7U0sYMr5Mp9fskF9mzuVA+12smEo2vvRXuHZVqvptgAt1wtBdel8
rwIPSVTsXI7+e7FnWvyFNTjgsxV75ETyjFckIpKgqzzi1DwafSsOwmJK/9SBVTn7
4Y09e1bE88kYZCbJU5tnTsjEwCEiXPJTI58yYE7XYpaYgycj9CQ8Smu0FB5YcAyj
SoQ+stTAxRX+F99LI1f2RDU3HqheCXEijyWWrcLhs93tLa9u0KkNgGC3pX/kGYZu
CpT+gQz9f2HzTCSu9IIjYIcZowbJmbvs944LJEBD0T8IZKaX8/VLHUlI4i1+6QGV
MTChrHXO3QwHsuiarfPyXvzqkYT/4xDbAGeG+p+pWG+r0Cw8uXYfdGevpH5ZXGpc
H7q1fYyZ7N2kQ+m9ObN0b8ast7mJ2B+nunAqtgs0DhkMVrL3pLLPiTXcz6s8wNMZ
1zD7Vw7+Z+4XDl9JiY8GO/MO+O0orLmUumH6LVwz4AkgG5pOb7hXvLm2nFRrrTj8
CKUHETpk9nzNurkLo73OxOdN+GMZF/W1tEe5c4DszPHbak3Rm7ZF7mo8yHW1mxx4
NVsR8RBtpp/xPaG46YZvMwUHI0mDak6/hR4bB0M/OvPllQ9sOQpYGt+WEZ8h/KSw
2qLuYsPv8ZBKN6kx1hwCid+AQ4nJf4aFkb/68WKqu9ZgpDiNvcfBYWwaMrjyKBvu
6slGOws2nwCPMHL5l7Bbxn8m3IaLpSl068236BOay1J/yZHUJ8vpgMP0UUg3dQ74
SvOZSA0PAHr8eUmfiHAToaFWOPRowJNCkVZYT9T68QZZMt4o1zsVp+ENT89+eOS/
DrXptEo/Cy6OV81VMwRHPRkMFU8OWF7pSEUyASiQC+aHeHDKrNMB7DXPZFdos/r4
BkwyDtz8KY7GEXwBVNfL6IGl/B3tPAYWBKrudUKZ/MWZf05/PtHpxdguNfBHoFDS
i9x7DclLlu/bfAdsUIzbxN+U+eUta8TYgm9vw6Ba2w6k8XrBSKeKICUwPne4V/Ru
4bBMzGm4+t7agHh99O1Tg/3njYFb/c3SsQNc07n6yB/t3Kje3zsRujOSIeDF7x+L
5jDhnNMlMb8mBdaVF3gJR5LnOHXG7htsYsUdBVul20G3SskFCyGL21p7azq6vxdg
hch7gEJwjTA91DIQZvwGt7ed/zScgAzlmiRk2FNj0kEUMJyDUxrfY16TdlFa8lyx
+e31jH5SgKj7hzpZXCVMCss38XTNb6DEfTMTRyfx1sAgWw0SHDYJrS4vC0v44tz7
OGsemrDjRoJ4XKhdN/yX41r5BKjmgXxfUsqrdlYbYmLFi+uMFk4JkGmKfcas/yMS
h01kDY4EGiGOwdU+f4iecwkmn9PfL+RmGCIdbeJg0iuLYazk3h2QwlAqv1/R/EvP
rH3JCfvItmwIZzvLB4SUfiZKvcItwrGnr5CB3qXsVTV3v85SkRYT6u0RucEBgu9E
AGld92QuMqWVZ93+zzzWKWvEMu5uSo9ZMLB/Wu4oBYZt9XYl8Wa4QDKzGT+nj5zQ
4P398Q71yoLH4lxs51d6i70qomqL6Z18KcOXBTk51xi0teMfEqYXgt1bCZ4gZCi5
/xIOAgFKzgm7KBDKxut+PaxwCveNy3d3Ydl6W7iIi5eSrXkrDDYfhqoimz5dl39B
cGI9DEeoFXDMtNgOBY6bouOizsQcm0WY6kENUXgVxlxM0O21020lIn70vK2WSIWi
5jqTm14ZTLNa2C/9srUrqENxtEKqHWRcwsYwYTqjiPPrdq+AZowz92eFON/khGER
8EYlWWLTmw1ROpH85XeRW+8vWA+lkODDyvKE+ML7h7nGXrsWKAEMn9HbkBQfo9bW
9y7kLAWfdTDqJ5hKIO4a69nvkk96s/iauI+eD/Dg5MtMyd/vzXVZ7TVD9vVuHKKI
eOfUDDAzXi58KJ2ARwThm3tf2e3Ook3si+eqWJTEwgDjKF2OCfTKL9JV8XnZkCAV
2LqhKe0N9oicv7WOKI2x0GyjlNjUSKElCVkMQJqmtcpW6c9cl09/UHUyX/vfMJRY
CFxMaFvpLzXpSbdtkSHEurag20av5DH7mBkkwAVkbfGpQKV77Br7BSJNHnh/mh/1
HvxzU9gtLEcFi/J5o/KwftmV/Qbh98Ea2JDBSWH8ZnhJvUd93002fUTfos8rI3JQ
UivVAcHZW9GHXoqTSrPzqX/po7HHCO4DGpUMWlJQy5j9ihxemq5q2GMjcyHmvscd
CJ8mlq623YL7svISy9HYCVLLO3lBD8ls+EUeEWG5Im6juJAf8pxwmT0kY7HpqTAb
jgWLjeiJfb9+KCc5d4BYAUuwppQE+4W5pbocy2YCi18xsg61qz0io1G3tMHE1nph
HmjiNLZ7Qfdcqta96iLGn/s+O4M1LqI8YixLHPZ7h1+mPNKWxkCz/yKZL935u4UW
gEh2g1EqUfPxZMTuJb14+15dnshIfnUPZczOiGvdZLYSn00eR6+HeEAqFzNlLbyA
mWgilIIzAha91P7RpnoMuoZ5ziW/tHefyad0ShZfOQX6o8ySPh+49Puy70Z4Akc+
+paY+MsXC8TFoquCIKl070KoIOIPbjeLzZLiv8oA/Ylg65oLJiaDamdeZivshhSW
3EG3GO6DVKVO4j7KAjKfs7sAzPQfqlYlwQvRp8EMs4oeTpobLlmnbuP73irC+RHq
u17nq+g6PkTNSROIVxNmLig+qMxsoBOzHO7SOuY2VVFKYMg2K7xylL83WKsFrzcZ
bDV4McY3fZYdAkPtHJiGGSifZS1J9hnjIvD5q0kilfv8WMzrwqIhd185jEepBDP8
OhefBYkNnM5VVbk/a/sfBi2oEoeqMvkORDcbI3UllClc5KXbdNu9zr8ErCz/BdUF
DkmjF05le6zW6PSY/O5sXYs7YukxOW25k0OyI2EKehotbYGto2ALYkwbTGZo9C/s
YSpMrhUKFbE3e1/co8/wDiGNLcssdcL3OFLhuQi9UVBAJlZL2tcXip4hUOuBMShh
P2qEQmGf9eqwblEt8pZl80spTeGYIEs62tnbRFwlmx9474XCV2kcFH+vOnPJYzUa
3PG8ISQMFr/Hsv4BkTHyGQORXRTLstjP3vLryXBZ2hYFwfnAPWP/oCl8ETRfO3E6
cM2Ka4kkT/q8LrFv1MPvGKbyZM86O+cxoDTM/iyg+uRZ2RzTrRzda4K6xJwy7IgP
xP2ozSMESbm56Bkx/ESnjtl2uH4lTSMTI0vastlmOLbhcO6YPvJlHjw9QyCGtiQT
96y+JTBH199e0zrLGlizbc9Z/fWDP59c7gkXujxpTX2ej7F1G3TNTIcRW0B2u0rV
R1XbV57q5l6zlEzfuGaxIfpY/sP8XZ3gFzbkpzD+QUV7aZBjEMzXplR3m60pRv2J
B75Z/My8+8VjFYSMKe/w+Stof2tpAdkodCow3GRkl1CsCrMqmIX8wwEGQbPxcWvK
oWuMvKrVtoWvAxR9ODyiRstYK0/JUgWesQeHIyrOO8Sadt67D3+CEfHW/MXzLa7T
bCcD/fIv4XyIyzveawS5iw9MDQctTelEG59QIwSVyaHesnN2AK41AFwCwGMzAY7A
Dg71m5GjCjC4VOhmEkqeKjZ0mkPHnmdHqe7BHyB91PFwZp5j8IAyNXB5Rm9rg8U6
W4658AzJxSXQlnRE45mw8qnbuoLZD5idLzwDK5aggFI7O9/ctH2WAYiDyqzQPnpI
kIqV/lCPQtbtu1uObvCsvKB5eIPSnbZtgyhqof0auvQCVDrY2dxQN9LfaT/SMjLs
BoRg98ghnOcUEy17BCXuLBtYsq6o6gTBGEvxAfnZj2w4EVKNTbk3ls77Ct6lNXu5
c+WWsCd9Xiar9ILJhsj36YUe+fNSOyRM/Loa23pNe3hOt81EQj6oKFSU9tVvn7Xd
TYp+LGt2oEZ2wuA5pZX+KvuUqvGvMwtB9sUMKL6FXwf0pHOSYp9ZrtIKFSZcnhck
1F2yli0vAc3m61DZyT3ev85JWJuVWWqdrcL4J0tKwZxTTQ32a/4iG0xjcbqR+fAQ
KvBeLaRUqQA9ciHSbTIfXdN/Z+zggiFQ0WsqIVtgbyuo6CM9iheMVWRwRot30LfN
KxFq1Md9t4ih6xbiWCC2GZjcJ3pe/hEUWJjKBRK+p3ZDrUvOaR7RGxffV3ObPDfj
ts9A2FMaVx+s/biqy8wGezixCTDzT0MJkd5DVtzX02DLfCJ8H9xkcdL4K0b/39Mi
lSGwMzN0yiC5+HHHdzh9y+lgIrGCPjRwPBoo9BT6CsyUWG3EUr9/ooZQT39HSlYK
Ix6iA23x5eKgok34zsiKb3rXJpf0Ti5NyM4VQ0CMWgpdIEog4LJ+FRl9TJwOfvxq
2qZyxvtnyC+G5keJeFnZHMTA1ouXr+2zF82iRahkevqls4OMQNep8dV/Yd34Rkzu
JA+0ve04tDdP5SrtSrjco3i6jEW9u1zqdrpcf34iOtR5NQcDY0KR00067w//NTKd
8yHwUM22thVbmP8SiT9PETUlVxNV6hfV3DPgvYxhfT9zNfw97Pf0CqAqZ2lnmPcA
aGirPrQhjbdJDmrho/+IOkeBXiq5hsdlWiDZXYSIQ1ITTMwsMQyrRxIBJ+PLq7GC
OzIeXadPw7HrqMpQbZN8ctfXQkCtJOjOXDlNqtdJVEJmltoJYbRQU5UO6ykljI2P
GxE7o/5GYKXOpwT4jsJyEMy/CfUxGb5FLAPnvTFQQHKCRL3adoykvcp7VPDpyuOk
+QU0FOCR+tla9rHRh2o3F9ONbhPkDSwGfkzuWgh/HBt4pJtvJEf4+EuAW55yxG4R
+sj45OA/zGZv9MucuWwMHeZizj/ZmP0H/FXQOpoQHSISjI2Lwwbn/CM6nkm6DhOt
dKpY1D0hmvR1x0SvfXOQWA/29/i2YQDyES9GXNdlark/wlAgBg60ciUa+p8JtnsG
P2WptDYlt6SwAZNroTzrLM5OT/GDRg4RoCfmPOD4cxSozPIkCDIBOPwNKmxk4t5Q
M2iu+fx2GH+tqhLqEXnO/uZL5XlpH1RhiT0vD/gxhcSq9P3ZImJ9+bPnbWuJxiGi
qqXa/t4cTKp2RPIcmxH2bgoAMq5UPfUn2i/roccTkOR/z2jK2LqIqr1vry+/gMLO
UT4QneWYDN9CoVmljEbrw1aQhpqEE/M/vVus1BZNn9QIbx1+3imeQDPRPSapGRA5
oVqjL8GluN3arMDTbqD3YJQw+XrrA5yHqEnqEhrDh3MH6rutKqLEl8gzcaPG14ZU
tKWX+pcVM3Uia6rmue6+vviEZbY4u4y6zabNMTuULkHL4Z+hGR8SwhngHi9Qy6If
bdN69aJiyYULILJKG0E384ExMYytH5nipRUJ5UM/R/sz9j8tEGbgJLpzWgCfXH5b
/li1WfO/f1nXtp7FHcGpmN2PtqNs0imzyPKGaIZXJIxUcJA53+a4EIRT102ZJHtu
HBE2ArUkK4lREZHPXl2so69bwufJw1lvP25sPf4mEvDhgY1Cob6ux+zzud2hUNBd
pLdm3bL7fTOw3oQurUk8iZ61pYGS76JG1sTPmQEP3DwagCFsbzdUUFsqX3fAzzzw
AMt1pQxEw2jFEiO5hw9kwjhTyVmzqvamUg0xc3OV9g1hCdMYuL3t5zMxJ4jf0wm3
6EvnP993xYWhngSqB4rQHTMcDh3YjPZLSLWSy0cJFMy7qoRn37kd44VYo5mDmKLf
XZdTaEXBdAvNglKzlnk/LkCCr/YMD4qbLTL37v5xZKymF680boAZuQjjJZHPAlqO
qGIwA4ukbSo0j7RCuXtQ+SfYFsHttNhB8MHzuqa3dhU/pWK9XrCczI74bbNYfB3K
cB/VoGRzNxAFx7x3O6cA53Pd4vhhVMSnuGhPjGQv7b7kO8sek+1R2jFWuI1VW4Kf
YcKq0g/wLgQc88tl69OmmQ2d9YZdtvh9Cv8klkQiSEX7pOeRyrscoOWFWDqDtNlR
E3joeaL77raeyJmRH+eIixs+hbt9tr8DjsPD6tTYZ95iMOJQuFdEi7hgrVAlMdeH
ko0JKij6q1YH+Kret/0Gvm4XNsfwpZy1rHrTjzIuTIGotsx+/+3bZ//KoNRrzYet
6uTH9wAbHEuBlUvm/M8Y893aau2r9moI8nCKn5nEYjO/K73Vby4gxU5vI3KOGgyK
JeWjr7CXSSJxa+Jii9Tbjl5B1Aifr2vdOPrO5EFwFBqsYTFWudLMdQ7GToK/iFef
RAqG3oYT4dsx2uZiaJd9WONf9BDSPDAyfByrbRpetGNR24jpri47o5Kla7renD9O
NEZeGATM//p4zeKygiBzqdh+l1ob9Apb6BVuevHF+qwLyLQDIgczw/JX3C3zvpe+
c0sm2mQnC5ZI3FgRODSTKZ34iZmBXtBL/Rx+fiX3EwsWwgdW4UksKD69cTX87mQB
WstNzbyBFx7+fNqIBUw+w/uZA3jDE2ACZCoFibI2pwSqOoHO8j5rBhQ6Ib24Z+kQ
/tYbHRtyTtIWuS8PiH6JRR5xNCVBiXUGVLD9vrpyxMflCI1dovSLWtIh0vkgYWm1
MoleDJFnvV/cXNdKPoApJsaAzC1QYaaOmwpRyOgKLkOED2Qt6m8l9mPJerEYXTU2
+hsTaBBlgniGIY+T7F2IgoQVXLCtZF4DYzU8llgrqQqtfBwZT+u+CS44LpMvf3YH
o8Y039L3ZxknGmVryJ4SuAVTz5LyazVM6R8S4oqfNZMuCE3nP3wVNdMOL8FncRsH
sCBdjrAy8SE59bZZEmCxqI2d7jU0SXSbBtZGnd5agfLXiTFrW4ToRMKuYJ0V6kgZ
jAi3JmE3Cv2mqa0FuCL7NeNISoLYI3tRfcfyhAmuzt9CXt3/YdpFbllUN+K2Wsvz
U5fiIqJX1A1jNNjRG8/AaH6sBLLjVgnJ83z8xJiBJ3LFD/sETK9tw0t0QA7c2wiV
18v8iEuXGBUlrzqEdPD0ORAffVz47bA1U/z/Rd6aG+hsIeP9w98c1m7r6JpCG1Jq
MgWmp5bpCVaxFBE2xg6TYXHTGjbz0GCApVXZIG6r/eJJIs/ZIJhYFC40sIeht59V
yMuSysKYzbgKSxtxPzBT0IwVeCOCDiPn1cA7EWNTeTBnlkJ2vO5q7ydS75ptFPNQ
Mlj4XHnSCQjGWM9DWU9Rd66AifkrzyYw4HQghgufTwNri1vd97wTO1oUSChYhuaA
f8yJtToiZ/RT7kPXDcVhYO4nOXoZVQU10c2SJXJatkD4OpecuCc/Yby2ZzZJBG2y
yfF1lPQ/wVqRDjMN5mJ1ib1xB7YpiMKSWtATGI+QIhQm3cHp+2KKtZsUXfor0bCJ
XX/XTA4wCv4WwO4ujg6vkmnf5BUTxXYUdUpPSU11K2v2sRL2ulBigdX+8E+FAtpQ
6EJ5ZBWJeRhuR3FJ1yLgn0TxHYlBpvTT+ZLxCJeZDG8vEgjIoQ7jfOKPoeT4tvkN
f3GypjS232l6yfPXWx9xfQAky6TptGP61D0IUDDdypsy1erQ865n/NYdlvGBmY1C
pqep1dDPhkbH6zhc2Zjvo/uWaM7oP+IM2AymH5DWtr3WHv0qSncve2nn3GplYeKx
PeUOm3Q0T0McU7Y8mqLgFOfYSg2xiaFOUYTW2w+6Z8mflkR3zRBL8tkh9mXFrfef
/jeQLeE2A+Sj3eb0SzYtjSDfsiusW/aIrhvGSGS+dIRz0OkcuLrK1EvCpjvV0BmM
3ENnnH/eIDXIYbEev5W2f3zAeNqC0OzUme1Tj52kynBtrFT4kAC54LMU4VeNk+WV
+JdVOLpNrgSmTvXO4JwBrxiXfQ6OGPyMX0Ln4a+MsHv/WDR+YJcb62HbAUBjSSpE
XMXdprJBFAh8S9f5+cXd4ruJRymyFl9YK0g9Wcbz2WqH3SVGVHNqwTE95Yf7I//y
QPua2IFBudNdoLikszaC9WcyS3emfQo3sXV4sapZyDO6GeQl1oAKM64XF8Hm+7ud
zJa+YXmm9k+xunEy2PDmr3F8uE1wiPS1Wp4Km5muCQrUgP7lzjKnif5/z2VwF3Ww
IQjuCxOY+c6nmcpCY/uUlcbwu0eXhIyYvTc5qXxAJ0caC2ymQtOgT/Z1vnst8U04
gF+i1ignFvMD7pP53UOiiqYSQu3emDFYb18ZSAalNYhIHEnGRc79E6rJf2e+/9rI
Lztu6aw0UrzgtLUxyB8LQ4vdxQaSTEAv4dUR1ddPmnZA1rJ/8yqoDq0H3GH2kEy9
iHFO99RMgm33s4zYLUI+eAAeqrkGQvzts/2gpSsoytpptkSSXix57ZPMV6JSNXI/
hMIkFxgCNUBeYR3I87xHFWJmIaHBXnezdbGviwvKsZQEoYOky3aMGe1vpy3+o0R1
9jneACO1Q1E6jG8MRwbkwIz1kxMKDxkloOsD/cjowUrxWmrLVx8Vi5ige8wcFTdp
SYPVUbpg/MVB6kLjZR29NnjkEM/G43zTaaZASjI9J6sLzWcAz4FO6Fk+5GJd+V7Y
1EPsrOLHTOO0MaOzPWwLF/sw4D4oPoCMxusBLyN/ysLCbWBBAeU/qdTkh0KptXRz
3lY9yQ/icTO4+T1mYtJRTzUcJwUKk+KTAwT/heFITAEw12L2OFAg88oFwiOsBxvE
75AWiPxAZcd4o20pnqlAOswMlnsRZdGuigA4IED7QS5qGq56A7fq5my3l0UAUMGq
b6kBvvjYLW2i1SnaS0aegfiRhzTTNPDyRJ7fTsSBPyDdV2a4oEz4jD2/moCu9G6K
ojRqB28v0mUcvuXMawu6EHqBPyj8d6daJUWxvDG9IZ1c0WKIen4TetEq7C78vK5g
w5+W2wApRaLL+lx/U5HwL9EDA89hfj20DpHez+l47VAx/+TXLbwDmYDw7M0tNSrZ
YSi2g4l3XS4EXwLI2BGTZh/OcGAckMin7OO1IgnOa0C1g1f+19vV+JHkhvOEL+GT
DBAyCNfjzvjU8/7d9o72zgEnCyLaPD7ZN+O2k0preIrbBRBaGlauySTdSG7VwSKK
o9ytmFEaQmy0YNiTXjEA/z+cNwMEvcOOMhidUbxI+b/4UF8eAT1ZWXhNy1Vk7jcz
pXWs+yLJgZvOyLEnEBCED6k6XUAvA9oqSZu/YaurECVG0+24tBJB3P8Ql9my8hJ5
jpC3+l1w4frX2/Wy+HpNbDKoWVh3kTtncro06KODX05UwKa0k8whJhCPMh+j2r5r
CxqMaxAT3hbZbZkBnsHQJemNbBYuUa9NGhKXqdSIY0JLlkHtc3e77ZxYR0pukqqg
23RFEEAlgebBnkknAyqmnHBL/a4xLS/tsYncub5Pp/ZLxn1QjERsnoYgYp0WGfK5
Pfg35akB6jCGGQPwgrpstcYrm6cQFrQgtg7M1zTHX9tRNS53pHdy1fwJZv6/UDTb
C4eYp72ADlIvhUbVnqTnNMQi7wb94su+sdIefeL7R+2gWSNS8yk7H3JNXe9SUSN8
b9A/36xij3Hu2gTwAiVucHyvQeS2ZocCqPMWyo+UR1scaETPzng1zIoDWK3qXz4B
gbTFIGAr23kAMN1ZpZC3dvOegawAGfnoH0yCJg7ipduC4EDzn7Q1q+lH/y+mwDU6
VqtQzpnGfIg9JsHsph/yRdmr4i7MOWN29HWNRPpZlp18msBww6gzTwn0teuP66p5
EM4dAwv93J3I6K/JYVMJH/IpOoOhrgXLA6bGB2nEbUsgEj8jAv3vdSAU8rXZZ8qT
rRS+oKGFWjNB5GLMB3VWTMGuIICaPbPZwdNT9mseA0iZmyek1dMJweeXybuFiFkx
lF2LH8WjyhDIy/kEh+/NBC7RHZ+ys+j3Woz7jqGP91oI5i/mo1iaKdT3s5aYB/gl
x+d/Q+fNcsRo0PwtgPPQ60rgK5s1EkDjUWcxA0E84WRDlcErku4Vp5TJe4b/QihT
TovkzZ/KpHG6LRnfh+xnJd0vuiBldPQ0WP1qd6TgT6AzVpiwHm/rvYgqZI10kIuj
V1wMR7BB9hAgiJpruF+bOK+fBz1UwlnFdxltF8JTqnTPhXgNrYZfEh8WHomxf5Jz
2IQXwbYyMoZ0yLZCQf5tPwgiJRLU1mDXUZZNlGKb6gciqT/gLUmK2oxqBMOE4jAt
4YtAG3054vtl/X51Vb7oSNl+CG2uZhZBWCKSd2NwJcbuWt5Z1FEGild08hYScxy6
S3L5Jfk0eHdZX5WYxP34qhxSHgl/GeqxcHO0DfBiiYyexx96y1EKf2OlY9+mVtA/
r4ugrF+vSlCEI9lcidYzTOVONYUdThgO9P1w+M9M/tRsEXu0/kug4W+wR2MrIi2T
lWi+FMjQEpiTRf3OMNYEqX+7mjeBoBqVvsBFA0pWIrAY/Rkg8R9OQB5o6X+pmnK2
E6Mh7W/nw3M/7RJhGkfjAaAqj/LXt4yIbPzkz2QWSs99fLhLPVgwDQoJG1IrLgvi
8HdDgoF1T4SO+c7CgCdUrZNoaethsricGfYEmGpQjnPqxExYRL+teDykEou9bXi2
9cK76h4pAx+G4yoKEMfFXIlWyqbr5quNQZzy2Ne05bLiS2LvMs2f9XEtttWve1y4
aSy6KqsayERekZlA7ij3p+bUCfQcwR4vSOaM69y1jEN6wARfMr3oIEFTghm3CE0x
OIXdzZRDzDRNQ3NjfXOVzxuP25t4pmKwoszc9bylTWgRttE/BoGD5S2iwTkSO/eK
CkeIWutV4UPHFQeIiMLoGd9QUH5ObhKa7EAHepJmpMrvJkslpwgCwpD0qompBuS0
3JOkjlBqXejDv8sOTQ+JuXX/AWpmajd78F/4XjdY4cjSK38zc+w6hrXiHd8Jezjk
MA6CdOd2J+A3CNeLaRu+tbyaIe9JjNmnkRrnAaQAqD1QFo4QbGk9YugFuJ2VvmYV
fHQU5thEArBf0Sf869NOeLOxjNUMNjYmJ5jBPGMONtkU6wQKTzHNQSXi+qyP+eq4
OVYNbslgrpNX6XfEuHuNQ8D9LuKdfj59Y+/AfOcqjIFSVmnju/Sgv2Qz8sr7QZ2E
SMqlwLuZR82xINlV0xm/wGw7eQxdAtsoNssPdihG7jgTS+dmLSKrsZqjUlNKoaJV
mfpFmNH79ow5skYShVLiodcM/6WXPrGSB9GWKuo1PTs14gRQu2OqYzrscHPmzodS
PCiOTYwx3ddD65ZQlGq623Ifv8wabwmORO31QNA37ImefcNP0Jvv0fsdkMZ0/xNj
4YFmU9C/AP7ClMycx6cRNX21teg9IXxf5LDxUUydsXYInW9v1sMH9mJdxkl1bPy7
HtMrLu6KwisgTCUZkGIJVBp1VrBdNJN7oWGCfbu721yKkxkEvq1uYmXGmxHPGRq4
I1dItz5ppVz+XYCze5ydzG+ry9ss2Ud77NLWmnVSampBPDE3p+P6lUG508SLQmmz
8v7FqOnwGclpzQtElNl65EQJYZ7DCYQefQaVWg/XcqhPZMMqqfT3yVyLSU2N+jRI
64wVdkMGTvpi/p7Q5SRA+AAq6hpgXBbuKK777byJvj9nqaj+qElZn4EhcymF2OHy
8vyhf3+butAQsn/4RoaMCfdH1qKzY19jtqa4ne4B/2htNI46vwJeLk3YxTcPDNpT
tGBdCYw1DJR0D751nB5t+pYVTYxR2e8temOC1Efn6CdFzfy2pnAgYQ8xfEIdxjns
l5lV8VuRLQgXV+eiEXim26j7BkOYlwRfRjOA/flnzNKRD99Hh85RCCDKX7dSH+SX
AXhizW1J2LO2Gt18qDd13R1MDW16jCbhCbyVQO1LppYCkYCS7jqnFOrW4hAG1aU+
zElkz6nMT826d6ChHMghsCFCrVQowGzv3OGKJ5Qhj2p7XFdmyNTQgMeFXTddNTck
gk4FMMGXnH98QhUTms9X8owhiJVBUAhUYpx2gSvS1hbTqZ2OrZGqOQpSWw6G1+SU
hhEziJmE0OlLILCNawn6FZb7rMnjlBKcHHz3RtwwBmgcpvpgOfGuEL655hp4f5XK
2kfhFYtcRG2ZHGHEWACVPOLxyciRVwDtfAp84bgrOukOKzkG6rPLhxXgL6zf/cDV
1gf9xv9mQYEsnDVt44LMzi2PnqvI6rZy9SD8K2vgI82Hz8fzRn9yNRxb45yD/H2S
Oyv2OhullpJxEbf8mf1AJ8M4/1hPNqpA2hZXK9R03l5sdJ8e9MnKKQMKlMgZo5sz
gn/JsT9EVLreeyFca4g80KUIVWDsVdhfnsaIOPIdLQfhjLs2DZNngxb0xNB3ZiYi
Elp+Sz/QHaFaQpaRyo4lDV2sHO6K1IqS6lfg5eeTmVWEiMuONGHywzU40LWY1gb3
cEq6cnCKT8YpszKiQLzlRpxlthEjptZ8e4LAjB4qGRl4eH/KGoYEUmiHEs2R+jts
88sIhr/T4Clir0VCatc6a2HSwp4daAJaDhAPV8AYdoH8Qkj5g8zttMC7TjwJpSLs
ezXFGb7B8ZWhiTZyBl38v1/lbbhor7TpHGyxWGMSeKNh4gWGfjQwq15bUwB9l85G
XUOd5bEOg+CKxB/YA17PRUI5BrPm40s/AwlkfSxNrDcqlhmolLIrknXr1OgxGepR
idvPaAPMvFlUmj+Zzdbum99qenUHJSP09qvJ1/t6RnTVxybkiWIbQ72RgJjBQ2Bs
a7oXpromZC/0IHmH5h4rrw++gveb6EDZBt0Gq3xpTMdSLUoPDeda3XvCvksKiMtU
ljmfK0cH1S2tVPXROaK1ok1HTD1idbStZ/4Z7H++7ZqhV6NuM3wwLhzevoqyA9L8
RhFM0SlHEKL7kRndWE78CJjnpSrHwckfLlUTf3dvvO8bbYD8c2qkrBDt15KkuCAl
h4E7I9wHqF7Ut+V18uHMoyOhhpLNvaLT5XlysX4VGuCzOxJDe0lu/JtDK6nTL1yB
I/cHTit/U1riFYbPvRHYC9qDTWaKhYMuI2IPgl+oS6YkK6cMNVAqeD55rwGcI676
wgtv2+oQw04W5VR2UiQddC+qKDjSaCqbJvbngxHmNnCdT3FQDqI+ObTcW2iQ7Vzj
vTF2/Dk8IRiTodwIpNz7Y/WQODNfiZ1qKQfcReILQMUTY150WBF8L4TZODDYbOOo
SN5Eduj24UWWRQvxWQoMceSMM6/0caZXTwBwlMN+YbtGocipzCjoqedtcrE97g8i
G+XtyOXLI2Qwy5oyc6sAWcIU/cXKmfL46WcNRYJy39KN5TKGLwq5MIybGHveJRHq
pkGmX8BlUWyoD5Ox7eJMiiht2Fqxl6ry3q5ABQ3JgSSURk7FYR3qPu9c5HZe+ehS
bG25RGVJZNAGCkni4CMTYHgzOVV3VwSWqmzLj2fOtWgjKVG0+q8hwdMesHP3ho2Q
xj22mGjKiMU8s+UYr8RoTKMxad+orrYjuN9ig2av3KTp+sK9oH2nWEBTW0inBXZP
Ai9iQ2qVz8fSwgQyvxzmOEg5zXRf4EvZnKz+hNYAwUMAWcdh0uUg5Wy5rNuqLLXL
v61jcbuyJIAYHNFxV5ZC9gHCQ0ledglW83ZHdnZWH/9Fmj7V6oRscy42AGFBnalB
9aE2ooFHyoiMlrWdc2IKLSnqOP8jbBWU61dUQfXgFPJ7vHn5dRgEIboKGQCNc+3l
6zkZtIucWFPzleQwpk2uuj5uTB95Clvy9/ioQkE/jfBm9ZuI2ki3O9Mec2DMYO5w
o7rGW9/gLToxQgJZa0/0ug8Id0iIuQnwCXV2n50XoK75NDt6Yu3CNSIWcLqtSqZP
86vrCTtEl7RXpbTmkK0qSWjEnTDZUKLpxAwFEanOkmLlS8xk/jSYIiSAqBq8xhqb
OtPO6jNhhRwAXrKZWVOLnRkg2HXAtAak/ZQejXblP62r87eh0EV7Aaf8O/xkeX6d
RwiP4F921bqkta4Kjoc7I0BJK5vIQ6Cw9LAzVNCQ6svMXmvLhWdBfLwfz9oMGo6c
8kCF7nxC01+Jh0KZH2+e1Tk9OHOTwdVnM92AgtVXE4cRRHc2jG3t4w5LV07feJ/V
fORzspHVHqDQELdZc+Jpu679NY7MkwstpGsfm0eXTAPBKi1kQpwtxGzAtTjgFq55
vj27NMAJe0HsAPmJRrx9rLPn6VLOmE9ViyWxwxzLnSD2eoAMJJO3juLq/MZW1wNw
9pkzTDogZESOD3vgKYnoVAc4+bnaPEqaTO/PNxdVFSLvQGf7tVLkBp94QsIcW52l
vV+kGWdPeUBangDLq3dVq21rG8tbRvt+8rI6ouaRSh2rnlhRF9AS6bEmgQFoN/vI
yBJu0YHLhqj0YDVY+DYXtwtJIkF6CFg5FOE3I1DT3uHN05mkx6LwRKYAHWVqG6rS
RkuAqrIeXkuYVpJbjFWnmETZyD1hmt5vAaxYkHXAHJ7EV3o3AWbAMEqGDvh8EQvp
QAocfmSz4dZDHyGd3WfloruorUEA9LKxuFEhwkymbVL67oo3giQKTMkc6g+7GATf
Wa/9+ziENtECtLyAqjOuy5oUA8TnMz19nviY0SAcM98hWwG/2EmCrLzl3l+g+TqL
zGx+zhn8SIZv87ptPy9Czy3z9oHYIAKY2NcWYQ403+nbDqUQu4M/XswPpW1suD/8
kAq6AwUlLuY1bEtelFbYbbAs/yqlmcSnmWIMsBc2R9OSWL5Kbn+4i/rX1m7dpW1g
gKQ7VjJlXhlUIJgRp20sCuYjakL3ofh0IMqpZU59Ov6WkmOZcse2/8EKGIuzFKLk
QRv1/qygdQ98WtEcTASWd4O8x6b1LHVYX9SuPwMAg2+eli5W1EdFU2hblndQEteZ
J0xKOlIngRsMjOeE/Axa088IiW0yRWjQVySZFs3KUTuENmtvMtRdd81HfbXFHUhE
gmWC9bHq5QgBhOlzjEs/jHm8hagkZRmblSdR9wNa7Raw2LBVlOHhBhvj9Sa9VnWF
i7XfFLCeSYukgX96B2RurYr86xwC6yy9s0uWojV2afVksJYk98di2wcy6RUZKDPb
vW38NPWLnNpdIp/ol46MxxNK1GvcZulMP3H0wZrRPyOOtjs86fjo4+uHkazxJaDn
KJzAgAtDNK3QX7bsNf2u+PQqFd9j4zC1CoSxArhfEXQqv9SPedZjdEMnYq1Utb7v
+LpzF5b2/smKgST4B9M+t2TssOCQH/I+mBpfMB0jX3ORIQluUxswc9xyzrIwQGo7
xWysQTA4ntmTgVfYUmw7Ph8F3QJbKriFgCT52iWqUj3FPJut/GhLqyFwVmDC5VNr
m56XaMAM1VebZEIPYpJYOXcuYYFt+UrQJYdvn0e9BHiYYFfUiNdjmR/v3fphEEDM
mHH+/YiDg4K8JvzZk4EC8/EPoNjq0lpTDQfua17Z3aSnIWlsqz/MjAQWo9kxSQzq
b5taz6JMwBdqfBvLjqcVySLArxco0hVU8Y54LP6JUYStLVAdImoG7zHr7FxWcj7N
Sy5zZ4OTL7pVdixMRGqHgVxQxrY6cELzPJN8bgm7QQaXCP4gsdnzfqlYzoiC7cUP
Flx6LDbFqIx5UhHkio+z/ppqhY8MWQPOM3IWt26ey75v4P0rn7xRwUE8Oxo0KLzw
mOKwlbSn7Ta4xRkmec8MwFFTybNXGht/Nqy7armv8dBm/jaxjTxjhzfa8i9nqXhS
okJC4k2csi7hC2H09iJgkk2kEQob+M1PAuHGLMZDkE7yiOYt1Czg6jlnDW3YguCf
3XZb7unibChSHbLxhlijBgJa55BIgkunaJHV/cUkU8n3YUHYIZC2B6HCaHnPlfhD
szZUclOk2ZYdZkewmQrnHVPt4J8nSphanZ/UiGkS5hFlvDz9k4JbMHa3Z+GXf2JN
1sEUUoNvDdRKVsvg3hV22z1OT+dcIoWTNVN9mNmCV8PyyMR+8kLTKXbSez/io33F
SnpM8AMP4xSM7D7TU6D7Z8yz91qL0shx8T/Jlfn9oTbaJbS0HCdTug6aTNxJ/guS
edf72DECegcq38Rgn42cVnb+5mY7UB2UTvbxKkx9wP2ceRrW4NtAbWHK7a+RgYf8
yLEnl5sFI5sFfSJ0YA4Zo/6y93F6KkgI/cmMY5dKlwlUB2gYk7WlL2+EkdLwJkBQ
oL5jCF/CnW7UhhMLh9Wh9P8Rj3RVsqGrNB4zeu4YnISGFOy58IyzHQJc6/KH6kT7
Kduvwng+tL3DQGtsp874n1/DRPlM2wG1qc6rS+pG4qm+eK8iCUhj27VZGhk4oCcV
QS7126iJ1j+VseFnkAijQi+nyarUK2/gNsdUIlvuJrsxOcgs3c/UBs966BrzIzRZ
KZhyffRS/HMkIKa4DKrfsHMIxg0BSbFWwEXgTHofDPzIThGSGf5verI/HXGxHT0w
jvMbLcOX+/fZFXFNmPqD+eUj6grdEIhcG/rhpYF3AfmMW2lIh4t5a8zLAtndtgay
7Umj8o84UEVFluSAkAcDvsIREPbO+oZjJhhP+yumvwNIOUciHMXgwSPv5EwDjiHv
li/6DXIQVLx4gUjRztVOtoiqqZyBLQMtdmvFM6ByVyPlJlW+pd6Xh3sZUmzx/j2F
hD1Sl6U+hOuiomQYNjnaapLrHWtqa7N0oa4w/+Ry8EzV1L0YxPmfEMwHhrzmP/n4
5Urqq4rdWYjWm0lu5d4QmOIeA39aV6yoXMZIXp+2uOqd46XA7bb1zD+Z4QPidqL7
+BdU0r6+QhbXgZqUHgoaS+PyAnynOJ/VCbaAxpwU2cHJtjLxgvYud5h4ZqPiOVtv
5OSElpWA++uobG50wXFgO9qZSwFdT87ELhUW2krmw+b5CbA5kgG6GHmyH/mPTwjI
xjSVQWtAnwU2CKmUfRChPztAahJK8BnNTHOlKomnqXTh62xpIPAMTIlHyc+Qq+G9
6U1kr6HgjNyB1ylrjhbjhVBzAmJYVYnfuA3ByURQMWHcnnsTUWfJaT1hZ30QfSsB
N/PjgRPuDTP33vrqzKw28Hl7PiW6yio1xcZfzyCHDFJxJd6lts635SJmgT3VQRD2
pkR3JaOumtHvzDfVTS3YeGZ5bV4cmcm1DDcQ66p4NXLax//xkT+/cBegy7pgDADT
ba/i093bvSzIqKEMQDyvuT55J1+xt9Ejn8p95+45XCGg1bejglLNsD08QU2J2Cjv
3rOa/ZLoVQAtofboA2RhGAy9+2zJytXieNwSAZBfkswiABKiBgqsSb/fmbgNhaSF
DO6BS1Rsilbrm1KiMEYx0HN8autHHQV9Q23DorgUoZPyFukcjWahdsknohfiHFoa
3Rxe66z5uXaYmM5eWfOuW8qsNk+nJ5hqjb9YYnQUHZyvgqxbjsZtD7ZiKLB1NAGU
vKBP99C2gKyw03pQRZFxTSW4I6B+Ew9o6EuWoTj1drIKexquPu2nrrCbn8dRG9/y
YpchzorifCVSN/0tTHevPcJI5hvoEcr3VOdT+whm1h+nyvjPUlCwSuqobeQo0KVy
a2KNYd8elnCv0SAWjAGgU7hFgEYWfIFOpo7f6KJoJNqowGRRWyvlpxz1JIzD8Qnm
QLd+sDPdCtq/woJVDkZYTNmq2qAWAnpZuxQ3Une3vIaa+a+2t4rEm+ZjMcSnEa60
0e+e6Bidy+ozJJE1ql1tCQNvS63mds9kLVYU5BvI7nzgrQ7rvWChS0hrw9qnAjua
umG+V/kMYyXCWQlmgFxuY/+7h9udjwbNQV2JO+nWevGPXmqLteDxVERfpvdGA+nk
FnV4Qr9Hq0bn8cPHU+4sN15o9jI3Sugf3xbBWsEus/ElaFu58z4B4MJQdEC9V0xG
bpoRGQpXjzZflC0ZblwUN84Tni32GN4X5pIlOoLpvdRsrHtWdp/qeIcGDFhmLgbg
+FPZEn+FC6dzW8Ga0bP0K61F6uoux91U8ei1k+Af+syQnSed4wfBHQ79iw1Dms/o
vyZJK4RebokjTXYUsBqmXf/CC+doDZ8UM6Bsv1vl7YNyTz7yozRPzXL1FT0WBIHu
O8k2QYqzkHBnqGMSsP1aDX6AaSwSAevT49MX/iunxFa5ij3ta1MPGADYuXfouegY
tOJpejrF4ts/jj2In2zMCkQzVlGDm77qL4PRfUFypmC2w9iSnHUoYp+osi1Sd4F0
QQZit3ollBEuLdGBvSlUzfGK+H8yqRBq4SZEepTsktqkkZxUGqF62n+r8m+kNnKJ
9joxzjEZyDtk94GERONqiiFDiSrVVOsqHLN4dtpbvozmCNX0Mtz8kAibG5AqN5HW
DIj2ZAuJ+3oB7M5KZd23AXFznSe2RSDS7d8jrRXD9Ug+VEvTo22N29qZnkfPmUVM
kr3bLYoZeKUQjLVc3di1g2uANosn3PotDFekkMsdtUVHJnbFdcz/2X9Y7Z7ELhDU
XvpCf+myWFoinlc+4aU/hY2fzlf8n1HtwvyiNOqRiEpkXJHVgUKCl9eM1veX3qHw
0u1xS+6hZ/hdwcpzlF9ZS7IBTeKkYlZfDmAkaq//fEAw8e/ePXz4qQLDcR/rrdUh
v/zFTQ4CpCA05js5y9CtiOQNI+o7pH5WGrwlozivU2Ig12trM9j1FLphUCcs58sW
KG2tgz760ErDHukVTLLhIJS+Eujs7+Ahkx2bo5hz7KYzgVKFSYg2H+XTCc/J5w+F
U1lHFl+u/pI8y3CM1yoUrqBlTWvs1Z8Gcah7oqQGfnIGELiywP73CiSEFVUmpjwC
h75OfFyXXlUKCKXo2MB7ygLHPIJaIUnppe9p2Jkpk/3STxiowJtwxv+z6eRU3/CH
nRcYNZGK0F6exZy0TqkEyizYm9H/UdLSJ3gvDGU9Dr9F7lqv1hV6Ocl/07TWGUAD
87eIn3esJfFMu/gS35HtRY70xYdlRC6D261BAXVrN6M8l5AugLyYqVzP2Qsu0A3F
N6pzsY8zNWXWK33vCy1dNoJ8RoKyqsTubGy5EJh3HubuQ0/MxrYLegVJXtfiIm+h
5V7G9TXamQC2417eL2xCdnd0p8adNEECDwz4idxIeQ8EwSR7f3zLUEtdNolJgvBw
PM2rpALYBqMQloN/VShBap/xPxLkKdfvxrGA8MCYfm5uEWLJ//7/QZ7iT3t5Kd+/
J0nVOLpaE8yZBmEIYBM4twNJ+EILtnnZDupVj7mVtWBHl/lvepTX61ozB3F3GmLM
TzVljCv+YZYqrbnKBjBvFTGWSbZdvTrH/nS6GjOmbH4u1hmYLqhrCEhbLiYB8ont
dGBVehakk5LSfpxeg3sOrcg90+8IV+IffAnOBvFexah/mDLUUzBk6/5XR1ZXEndZ
eoe4W4dhwdHFn4HQmqqvXE0rIYZ6LOBHQnAOnq8nLGNFL4bKdX75orIqyp5jkQ0l
/Tzz0DuOld4IdK8ZIn0DLFfdsGtHIXmkra2dYh9qOXZnZWkRQVyaEeBuxyTkA/aw
/Msjc7hMAidOlCGoX3odQ/8dz2ZzTv1VHczaHshBk/+SmCCmpHUAiXIYCj7+2InU
WTAgSvyQaIy7SeLcIWrXD9wV1e9oUIScAuJg0G10oX7mlHQhhEDkSxHunGpcFlYv
67DcmIAcYKV4ViAdAi7jiZu+wMMEZAd379xGrHCqJEx7D6KWYV9+3BjM3qAB01jR
TygvFeGKeDF7uFHX1D9NXoHQZ6iqeSEBasmvLVHECUx8MDNDbk8B8XsmVXbdOp3Q
er19LvAOg7JCXnlOxWkA/PILDclmApYubC41ziyIpfGJMzhddsbDAGezjd4KaAhZ
oXxWQxc4sHm2tmGiY3cCzDVCb6Zxd9CbVJUOQB9noKlK3iFog7KfUlqLI9aFlHGc
00Bkue/9t2CLOrDXwrFEQf/48I8Z4k39Vyde8ssVHcwh2aFfLq1oz3B0SxMxIgnN
wTIBG6nQu2wNF2YEYy6MiUbrgbniIXAD2a/b9b+Bm2ugI6orf9NfERP8L9F8ivta
Kba7ialiICSs+uiO4Y95ei0pY5SXb5OFAkRxFTeW3K4eu23hdZDCuDe9H1Ce3av7
T4/HcJTWAGZKBNID4XGiZ0H6H3SQoJbbekNw/4u2gjQEcz5VkK3sWhYALYOTIK6k
T7xC9ayB6yAJMdPS8FdX0HiSvJ5fkSgAX8A+P8KXmaE9vzlZ+/RT1NYM+ZHXS9ZX
HJyC2JS+ZTfjO3qauQ6wHwETHfzHGVoV+KhL8Ke0hHRrWTikKoKgCAWi9E1xCUfU
Xie58ij5YTUT6RMesKnMSQ09ypTQG+oGPIWv3a2Ub/y9KayGBdR2f3AnuyqoqE5t
wJNJjsFWujkzBjknKuAc5Z/DpjM7uTd98cuJ0EGmfDt5g2BAbjHAqlmjCEOMfTVo
WLGL5O4giUWQJmk328/Y9UEwR0/+kaWWEU/Nccz+xc9O46rsJFhv/UAf0TZS7+0X
ErFsF/MbMjrte+ek58FdFpeUKnuJXkO/VdngRC4aOqHHr4ztVVhsWhEZ+LvilJpm
BM71td+Y7V/E+c5TAYlqpW6e4+enwSRhwnxLCCPv2f3iPxEVS7rwtOALg1okkJ6I
9r6rGJy+bInnY9CPReWbxHh+8w7Nv5l4xPE0zB8/G1H5Iv2mvy00CS4yP5ZUNNP7
jqAFC9kdlXB/Ld3hn4IgClNiZLDlX8bRq7GWnzLPfecnO2+Upw4n0er7Jcj1sdzm
K0kj9RQVPglZVIfCmD1+vEuI5JAQ3JeP8VxEIbMs3+Z060eeJayStM1WdoYbW0ba
P7bv+NbttJVAB0PS4lQxXHhfQ8aPSZuWTQmoHDTtyE6aShVd2M/jVLWsuZbZscht
bVrneN+nXWDH6BbHbiAV6XXCXGTYmsOAy+jkgV1tyAaLtpOtF6mY0XdltNDiSQsc
KWQz14f7IuLO4rp0BDb554YYcaEgjHmst8PjLwgTH8SGb92S6XjPka3z89twtESu
/Yg7HHJOCoKGD/m/mO+dzdkzutr4yA2bQo74dvAz3Sc7haw78n5Q742j8uSbkT00
z3PAAvZahsE4AT2jmEt0FkoXzc94jlRJLrYaFW92sqIehvhvudnur/seewufPILq
LzIy+nSq3IYmuHP//EbKmJSAWx606zx2twDcQcFBGxG5gNXV7hiTj/TjbYXVNSVF
wkGvy/SwcQOkwwm+DFc78JUQbHBo61HAT5s1lNxydAspKKLxAVAqXzBVDuOXCrvw
V1iRQPwSdR407V1Edf0F+5imHVtS7CcZAVw6AsXg9neQDfrorfFqTGk+Bi6awT6Y
WhHOcsPP8C40q6X95n9fI+F67rl5+d0wSleotkybh+Ut3TONHUEbOkzzKmlUjCUg
zCea8NkIHVdTksl2rHhg+2LLfbe+z5lazZI2UAd2aaoe8b6dZXhh73ZbFRVW5pXw
idig40kT0k0Ug2VfMy40O1kWJ5wNXJH7v9LIGTD25BtuP9UkSgu2uWuWaQWRz8kU
tPkPpWBdCOM8Sqcg4Xh0EjAPcM8CyGdKYozBx7espoiT2E4qhIa2OI0HoSvk5bff
7sQbqb5xkWDGQ5WYC/Z/1ieHRp/591m/q1w3ElOIdRA25L9FeuYml2T8bqQgKc/k
YZAXdqVMYLUzKLijLJ6wmlIcTpaEsNlNxvxUEV0JG5WZGRqKLLC9VFJVi5TVf20Y
EI372LYQf7UksMM7sUDkryxc/azwPMfZHmTQyXWbb3zoMorQSNO9WAtSp4hvyGej
6Qh723voFZ3Lasp67V+ycSURtFIJ2UuZf0GymT/QGqaDeOhoQQuOMI2/NrkaMNLQ
hZiJ0mFjlZFaqW4S0mV8Xyp8XzXpE96by+R5Dmw1qkTN6q5PsJQWo1234W0ARr8P
3P3d1fSrV5YUgpM+a9tG3uTE/3xVrfXIThFoX1y202t2j62KazQfpovse+2d0WFb
P3bhQFwcdD1eaJW2/J6wSafNcdnWro358INtWL+zRz9+5ygwsp58aPGqEg+LY2ko
DWjsHrwHI/rVoJNRD/7Af2iZPW/FMTjshz3XnnJTLcgd7zlM+7f0LP4psc0Y9jr8
EjdfqlSS9SoFdgW1FRWfVK3LVg/Vs2l9H+mkLmpxr5WcfOrfVYJ0pZDar4J6qZdQ
gZLrhYM0Yl0R0dHQprjHfnJsd1IF19P7rbyJlE4YdNEvPs1yPB34xKhYMnotcRvL
RKItSk6yvC2VVJI3I/Iz5oYv7vU2/HRvvTmD9fzPIjpTX9GeCCOZ0TD8UKlZRk6P
HOtpWiAMrr8z3V+m/VAn+emYJzZ1/H5rGDA50v7oPDVq+77+2sbXPS4iRbhSLS7S
M3W2zqAO07rG4zMwrRYBx5NUYkMvBuAyggFts9QqElI2r4GdDYtwNKnP8gIoeL+d
U0fGiT1oMgcGd31h/GwKrymZXWtrNJgI7fXoKXfa2uWOl4GUhwYf54ok9bFF/z3r
zyt7aNLBtQjTo6q5rHbdrA4A5/TIlfq/KP0bqGvmNjJv2yLHKAqIJBhIN6y9Beax
Qdmdt7JQsdCe3SyE7AMxZO9WUXe6+MjPQLxqZt3aNdHtxMk4zyGRPpqWYTvTCAsR
NegtCq4EqRiBSInX1ckt5P87++BGXDU5l0CwjncMKUU/KRnVVD0ACv66TC5pT6Tc
2gdhP6NjxznfuqycOMl9Ey+ZA8WlubvDRwMPTK/2E6h8tDNqj+1uS2aX8iIODoXF
dHsd6o9hqctvVQUTWMOL1q5lcrlXhipBhrZzH9AAEGQdzXqkJ+BFNfWv0/RfPg6s
8gwwQSJBBJCO6J2zRN4TukGCvpRToFnHuwZHBJKfwS4Gh5uiVKqB4v40xD8h66FL
PfV7GCF8Uynyn1MHOyRw4faSkbiogaIRG1O6isDX4ug7qb4/213Vh20XtWDg24U1
aHL555ZFWwcI9a7b0fCAzSkC+BzRGoVwYoq/wHTlVE+Nwa5iBRfEVYKiGBeX1ycY
NKOYT8QfhYa6YKgZcTIKKOBPk3UhrJvQRxKCgmP1D121NuciVWexSyOsLNMBCp3+
Tj/eRkl9UbxrWEtxFjqEeJXZSMKvewragb5QRYCrOLY2LNONGZxfB8TOuDLEkPzR
Qdgk5nwcahqgLWEo2J+2JVxt0ZfFM10KIMsQ2ZFLoe1uWfy6J8/ZT9Ky6Vmkc9nt
FvOgX/Zoh1tmpZ8pLNSfA09d/Q6qSQqXFgRtbl8nyAleAx2nXK0+k5BOlUX4AlCC
iuFhgqEgfBAVRcDeF964/qX/UuDm+XBr/5PpOmpyBVYGfHBpJVHV2ycijFS9F1Tc
Uz4RRo9PrVDNk0lq2exsB7YTyoCRgfhfjenkdAQJ4uyJRsaCiG7Wl+zq8hS2JvJP
ERUpXArw5SEu1mt9vuvZnq68oHTl+7FHproTXUGBu7RognsL40+BtPUY3crcYI38
w5QzoLXcOvq6118Isv7qsSIC1H3VKIUA8EtYxkaW24PzBzY5G4/cgSKWPga2oFtv
yhsG/KD1GgpFSZEr31NZz1a1ZWv+uE/l0yAxa9S7F1t9hD5mWK8vTMPhgdmljQku
8tO377ekFyDLZfyR6uMS11TklqQJElBO4EC1gQhrM+exaoFn/9bFEeyCFRUEfJQe
l6rbTYpQJ+Z1eBBxPgK58xEOe9zDPUC8Iza6PLnIEZL+hF4zQKjq7R6PlqSS5NNr
NMBHBDHzyn4zORgMX+DKGIPW+faovgsm/5gthL+LtLjoR8wVWeYuVJrHEgMyXBkK
rkeswl3gDhNPxz5+Unz9pIKXClx3AENovwgRPepoqILcrhHK8rNTZtQtlOSQ7f94
ZmmyoiT07V9dCiTbNzp1dxMrwceUgDayWSDBCwMRZemTXI95ABFdqSKiBY1Oj2Xw
eld2Q8ZUjJqMahwTRKIo2iyf4IaywT2ORaFlLqESXHcNE+vT6xQlZwpaMe8Tmmp4
LpZ3huRJv2twHqB2kpko9JiXySlWCGOsEYkz9DrY/hGfhD8lEUaB9gHNWrHMKbnL
FUeQfArk5vsSFqEpYbkTCNf8RTZbx0X+JUMxbshZXERlJ6ZsmKVdggxKpXauttgk
pWsWawCNMhtx2JW99/tW5pngAIFxqFwSKdGnJmLWaYPAqLAT1W6OlI/7lFS79BMd
SpNZ0ksSvC2429JtyaniAf4uTNJCq2ACxPAqIJm4lHRoRVCuBCUO5i8VvcZXYIi2
phWSz3oAQ7wxTRHBS4N28ozaDxUeVTHfXmt6JuyVrQa9v0MCdwPa2Yg7r2jpHEQf
E8BzlDCkYLAHdBertp8jm5jkCGcl0zRpc+cPSuC0uVSSLKgxCgswQm8UAxE6Zv0x
ygvFa8ncBNGIFWss2x8ubOL0apzySZJj+T9hA4pkGPOiRDTYzxJ44cAJuPu85+dJ
nZwBRez/4QhoOLO9c4uZFld/dkPlvehNJvgxNdTOgBOftKqqE8Uq3QmhUoTJp/bY
c/KjZhlUhAfkYc+s6IerO5kxZFjgtjMhflc4r9lzj6c/WAY7yckj9BaXiQ5zyecg
zn7cXeJIUQ92VqZPKbunQYs/UHr+tz7ShFQrl6n/88mcj0pV7lmU2pHDJVb5Z79T
pKhazmjHlVxOlBl+nOuXKA/czV86CejlvQdpClBXo1xLUIQDz4/sV79UM7UTzRDE
E65XrMq4PR4/7I9cC0NqCB5wS2/RTz2nG9L2KPkU21nJPutgcMDhaxXjw0rJjxuM
xTyOhtH83pkj3dnubTAbXEn5N1BcUTVPfx5WeQ/iUbckS6FjuuGHclvTmA6sRyo1
GxF/O7jnMDvYaCbL7JHZNZ8BPvhdmH6+3/XMsD/LjIwwG0F+QSui10MP1HabsfQr
y6hHfhlE72IU+hZ4jjGqOkDFFrPfu90D7b4csQRsUIo33jS/o1hxcK4mBBQTW8bL
yil0TkZgARFBbcr2uQRJuoPYNZ4NzK1FExvGq+CRjcyInrAeb5nz8O7hvkDUlhdv
jq78zrJShzPniVTN0G86o5BqMS6DCH1/jP9xP0yRYf7nEaURjXX6454bTmvWJvaD
LyOfkGnw881Ukayn2h1BpRiPLp5MDp+pJ6avwR+ypSj1j6IoAuwpNOLGlogRUvom
SAA1uhhQjxHAHafSPIC1iBtmpSa9xLuE/BVzGcZExoN7X53KJlMd+oojbJg38VVh
ibquU4+GLTWQmmPbnZrPy9UYgHX1neKWa93SEYkNRRXRARvuwlPzT3wjwdtSTMFj
IKmZmsVd6JWw1ox11Yf5mpwxKLRYxHBKxU4YB+G9LYBprF19gr+T/BiPK4lGVQZg
86TUcbEz6Xvr8pwoK83UAQXXpNjL9SyB125jZvCAbVhDGfcn9Ot/J/obavRqs/5Z
ms/y7Vk4x2NfAnwxKNkqrhq3mMsCqCYNR8XPk6qAjlPuCwOy0mryfyokWaN7tvqz
7trelQtbRYp8CDWwalh04Mk0n5DlI4gW5mplOeW/m8IfNcMxcZQAMWrJ48kkdg45
bLpBQQmjeKfoaWTkgf0GB3A1f3ERbLyZqNK7I9H/jkz2I1AZDMaSnMz7pMaiq1rx
5OkWMTZflMUE8cINAfDIJVxrDm/tfy769gBzpFcZp6sF/oZKbaQPsK9MIYZXBFNg
QTClcOCjZ8fTuBNIW0/4QNfz4LdjoU/2DAKS5UsMJWjDDidyWotXr7d2sAA8UHJV
PUNfgc+dsShDdFX/3Wdf+4oJYAnl95gDfh7zLaohriOEaKJoV+o0v/5dNk3x60Sn
BnXrOPywsWfypk+lL/8bAdKcLFX/qHkyv/1yxdbFcymtXwjf7dI1BFydwZ1I3lBH
g0fGs7hlERZND9XXEoBfC1YJoFam03O1TljfTToOzphiIqWGppZaps+4TFMsEaOc
4HQB6burko/X7PzBQpllt31B0CDAlIf/ESzH5FE9xXGf38z6jqydKeQYmrKnMYNn
x7hqi+epWWZl9KU4n9w8sDz6tD7D9vtX+wUGm3Jtbl0ZjyndzaYhomYbC8xwfNzz
PIoyCkuuIQecreR+R9Yr1VyDZXq4l13B4XA1H7UgRK52EIILJV4o9BPF1O0rhoBH
hMH0HyeUXRvXOlkmCupCjgm1w2SE+XkwJkRZ5HNAO3UkU0qyCz3ZrInC889i+icv
KynSZAxKF7NkTNTUWrJs7+JrHbzm2SnSF6lxZYbVH0jVWQex/b4Hk/h2axMl6I1F
74Z6l1iLkX0tGUAFPZhm2HNPY03zk8OH58K1v0Jk7YEiYvjbuYRncP0AkVXszPui
PMLkrlEKpjLBLkLUjVtzg09ChWMZ/SSGbLoFo9tWbyjVYte3flicGkEDQvrIYCK3
Rl/kE82o0smevcovOqvXF/5maL6INj/OzAYdR3qKWHPjUnSAOOgrPHLxuIE5j2Ze
jzbSApuw0eVjYe/GZ22ZicVskEfkVIPxGSpetBwyogGZ/FwsWefHQ7JI60FaniFg
5mo1ilx0wKOR631zRqptMMF9CrpemqxCuSascUxDhWk7giO3UDE6Ju61TXGcsOLw
2q5D68l4gglsDC+i/WSxN/dK7WIN32ZU3ZL/y9yTsbAH1H48Fdf8RUuNq7XqKd0K
YLp0f0e9zXzkz2aR81ThUVWua2WhKv9xCrfRvrJe1j7o73qHZawrOfD7kBLFzmGg
dQTEJJ2t9h7oxdRuX/UPkHRm0XHBR4JCBM/cTA7vn3phYIUSub0bpdpTjzvHPIA9
iDxbC3fRiIUsjlA7NuhQEf+zBlOasdD97tSzlxa9IiakozBPg9B+WbuvoNG5Dk/b
u4SfpXS0h/jy1FSgDED5VSUVRnTZrxPqx5T0ZfhSoZd7wn3IheO7GW9ZhDBYNzqT
5PqJJWu4AMrKMAqcNRT894suaO6+29FlnvnN1eqUr3JTgifGIZRxaPOuZ2a/hFYT
LZIVEyLcJsZ9WX4DYrO/WYme/X/JxDJLPwDLDo25udR5c1IFY+dY8a6S4+vWUDlN
YaeGGF9Ywo5pgWewALNySFapNDyz1IzYKDoEXvluURUwHgHB8tJGfLkj292o40lo
2V8AkK+DZmIFNAZvMi6hU4wVIOFvY/6ugRARiLT4kyhFUuAqVvIWP/aIXLxJJkO1
L2hV2W0Yc1nywKquXeHewA/jNpWQss3O4F71dkgMM/gepRt4oHbne1d4qjwqwInK
FxHrONBYjtdJ9JzFahSXEuV/7wUizluI5vyL6sUjsu2Jpgg/8TZ+quZoCWm/F6h9
uFyi0hCcMH508ut5xxbewq1Up8ZWj427gt8F6FcAUfOfZfTFdzG77TG+cBjR0j8l
6RyluQGValOrWIrXK23iLnovj0tQph/lKGbXNl2nZMcS3djdW4k1HL8Kn1KYEpdw
OvBDG48D11QOG8dNwCOEGcuSsQ+rSGizEnJJvmWE2IB+AaUAHmfW9saf1k9SJdTh
QoX6Zdx36yJqkNsfIkmljYGFHKh6TDEbwaqPtfmLjVTbj1M7nZ+2T3DVPLkJ4C72
00qNkoDUxDj01nuVuxXmkns1o2ZDEl3c89Nha/5Q1uKY5xaMSKjPkR/aYbV3VPAT
7zAlWxAaJMUaedhMrqAKk3SmodgE+BPW2fW3h6QtEBU+beEugoUAJ3ttHFm5wkmX
lwz1mWQDDHEuTueSH+wJwnKI9amBP1ruAd9NDhzm137MShqtXORiuRIGSve3btvH
tzANbm/qLkKzGlv3KjQlxTFqcKIMY+Az2QGr0lD7nk1rqgPTO81gefau8CMN6G2O
rJuZfeYkAuOxTIMzcnH8bJ0X+bEOLZLWjMGPUQuiJepU/Y8QyKzUmhQC822Fmd94
VJB8KIS1httVf47MJ5qzN/ge66bAOPTnOIaXiN8ZYO1BaUpeBL4lU7f121sVKpOP
FMRVA5VwjPcvcIDRxgy+bQsFCXUxT0m/JzlIqG6z24D5DaBTtqhuP1QDJ77gGAN2
a5apFtnN2LFYXw3pMZUAr11CN9AuTuGg3nJ85IUfQRAtBtyzJMSfw38kr77WN2V6
ZhkKVt0wscTE9a1RsFZEMRCPgKcgfLoBzsHdeoLb2lTpLFoZoeNmcF/vHusjxy1b
fe0IMNVNUzgtBpLCP06ElnWwNJNTO/gyp3/Pax3vzisTtCahSsqUmi+dLtFduDZ8
WbMPijLW+7QCIMGMrt8wTMM4mKxKoDtrx8yXth3t0TxxAYf0YRxhohucatNj2uCp
DEP3g2UNyODJ7zGih4hZOPSuXgwW7Or7a2M3Yg73U2Umeku+mnKNgQhLrILZ/NjK
eWmRyEbHlyiYvxCyc9VLWDa6qyohwKjzBgeUQsLg3WugHFRvOlDG2XuwWjbhskkR
emm41vnor+H7aNi6R6jAEmRe8P0wIy7FZvqVWrRx81pauYXtE4obbzFVCgsNEmc6
/LzGpmn1DjxMtmfyui4aOgnTt8wdvH04iDVpyVevl5xTPxSN3u8I5ocJ6ZJlWexg
mJW7ftooT4iYTW2Mho2MHcsHyrnnssDwOnMRizCCpIXbUsRXSFf0mRAev+ptMKXX
LPbpqq64NMUTpwTc6PWGLgbHu+LZdPOdFesw8J+wkrINKicaE/pfL9SAtXvUCAHr
zOZjTqVyqIo38jxaAdCsPIu9LjpMJlybK6fC5cq8nAqo1y9M9CvTmo931ydkp+O2
DMdDiaWmAcoRRVrQR9dcjY+5ZRvnErAqgF2b98bIF1eUuMd60qvSwo65d1yzZL7z
F0pN7g6PhXf8X4hpPgJ5ZtZOZsYGXIgEB9dAfp0WTtmUDGZlCxM15px2dqBDNPKB
7ccEysEhJ8bxb82LKKjn5KiLmLT8mMZT5mAZxbBdDCgP2BTAIC14K8gvrda3uOUM
YMY+QB2vFBL+EaFQu4apMVGkfGq13GMIcrpSbAGzmv53C6hR4WdrCD7euInefMcM
q8fNSPhArbSo0DBW8BZa1uInJ3SPzmFZzEd6cHPfUsepP7wdRGXKIBLm0wrao2WV
i3YUBAPPiH0W71WJiP6Napkhm5B2VYBL9fHRclU2yWGKdGCjnkZ4XzXyM+IonynR
THWAOybZAy+YBd2w3srbY5pyaYrVD6JBbS5KGXtZ4zzAxYFMxkw2HnLpH9m/8xuU
cVEFDW4IgR+lKKYIu2pcZuqc2jitRFzv/G2Wt5C/etRUCw36mo/xx4DQqieXcOZd
cs/UmSLSY43o0hk81Z7znL0+EufhbB/ZVDSXrI0GtePVdgw6QxZ2/ZJZQApDbD/5
XFm7DXFTqJJF8SNYEj8Zj6y9fty2wGz3hQ8yAMby3GLQbIz6UOkx2rq/iu6mQmP2
U/q3i72ES6t9PjGhXa8hbQqjpLorrqjqg7mH2XQulKOnttVJU1tMQomMkVHHfyYY
GlALYKPKuS6Pl78EJk11PBT8bwf+uU+7e/FRX4rl15WYERMkqmyvNvk8GLP2sspr
VFYvIMCy0YPPN+ixstHDl9yZZcKrliWP2N1XvbF/2kBHJB/4vVM5mOG3CTpPxoRF
k+5LKVcXofeqE0OojeLlFGkqiTXjRDKYgOf83pCElbjZGvJTFOPtV1TKhF69tZK7
Ogj3xA/y/aYRO9D+nflou6Hju+qt5z2dmS9VhMDKESqHdYiJb9fTQUoEVIQJG28/
bUySUW4djdgrRIxZAZvAWSG0znXSRi3/ipeaFE+WvEFVhwwvJa0r95dxCo8Hw9HE
JcsWu8IUCziE9ew20WyiVsJOgUaaC4WtN+pWgBzDr7hK/dSqaBQGmqLrZirzpIDS
p6bprKVxAVOHr0JHqSf9la+ke8HAn/vZrGqMnc0pSRYAKBEg3tpO6Wh2RUxuE4Do
a1mK2JnwsWMp7rSd86qfh/0nshq+OtXBDLyGQEAsy2OdDd08vEwzD/TL3uEiH1XN
H5umfVuJXRURywqXYMUJzpcp0tLa7j6rUepzJHcOdh2A23GJ5UObUGPRM2gYic3a
vWhvO3L5q/PykRO+rEmLjUCZ5SZntIu9+xPpZhQ8Wpyy97RNqnST2GalniLxc+n7
Ftz+Qe34zfxJMfp3JP6eKaMZjr7V2nevl4iHjTDti0IkbEoIOXbHWokgvsbTctVE
n7h8TNyY+O+7IZumHAkeFCWFayns+ZHMgQE4tVapkoV+orKh+rAbbPIbGOUb5N5N
sOBbdW97gHB7GtO4mMHSNeAhZ0svJJL/yT+ha9qq7bkhW3ZeSXFkk/wokaGLdYfp
KoZTu0xihw0qSDmAlq7cwJUCq7QMZiEllRuMRIrYC7nJpMBZTV3wDxhWpFtZhCVl
zpd6V6n83J+TSRuJKoRVndqAO9LGY1OK5OycVoXGIDWgp8C+/y2cPG7Va5Hs+n5R
EWqeVTNwlUccn+dp4eJZyvnr+qd8/ZULUldcPUMqz7nDvgOczy6kKXPM2XhF6Q2a
8/jByUIH+9OV91rplyR97ANQsLI5oTlBFLmHqQhqxph87mIDSG+GQYrFMn71y51l
JBPtpJargX6FPk8oCadp40BYW6ud11GmGu1ETVn05bpjtWtrFOGw3N446ZpjNwMJ
5OSdhE2pFAeVAdOjlSkss23XfPlh4xtdGi/lNRVcB2YYZugN1EnviUTIVVIc6TQI
lX7lntCi9yI8EkFjeQCKNS33clsCOg3tIZZNvyrB4yL/r8VeWVekubhtJlpgyiMk
ldJ+f9kWroVEPVa8HF5k8GUSZXK0dw8V1AuYqmzBvAPK/rJ7QlPG1D7kENB5rb4n
H0xYN+WLjMKjoSV03vGSJmIT05WZa8+5nA7PGQ5lj4BKHikivm4f+KfC9RD6otsm
TektriOV89+MVeLzEc9V6TzlM3EIaQZobJWlTplLBPOHJuz6lKj5yfSQDAjej9+M
40y7dp1OU6/pRFu+TakcKnitKyLtBbCB3o1CAbgSIZ9eKgcatBo3ap79kbP+2/ON
bPWn8xTShyxprfuZ0Z4CBei59OG4yIc8IyjTkBGeKBtJS/+uunqKtqehfKHLownS
OUxc0AuigltMSwatjxDYh154R3Hfivoc9DXqomqoYKWyheJEVGJ2LLRTtiBAxZB2
aPsFtOA/eQOzt8EodAR3sYMpC0x/toyPS0Fp8h5tYlTzl6rq6AfbA8L06G/D6TMD
/P7YKJh9nLQ3y9tx/WoGpNojAdgH6wobEcwTDq1voBCC318Xn7QDlsR3cO9vY1jQ
hCI95FY++zhqN/PjMG6FOAB+jpnE+X3XObAin0T8cthH831O9wyRRBCeihtiA2dS
Un0ab2rIesD4C/+FGoNSAijATTBTMoV3t4NacFx26qis6A3PFA/rhAweR5QJn+/W
4Dgxs8FYOWoJWZNugxTy0FDdhrGlbfJu6t0/alG6dyNJAkzcKDmX5jgDjBInnFJT
rIUBYAn/dpaRYDKqhv3Wi1py63Nm0jPONMNMBcYWgX2aPyqVvpZjyaQfizSL3YCI
MlkTvQL2YG+rzogRY313GJjsVaitSqvsl6hGK+FQKDVO4iDfJvBwyzcsed2fuA7V
C6R8RJ9AD/GK1JhIDbJ/qh01mqZVV3XqKNphEjEN4uw3X3IZl+rcwzIzrPRxLW+h
3BRs89tO1QfM36zoFBw313CJqHcusKw1TOm+x7ubxDCIs3ucTJiCuc43TSRbhspm
S/bT0wgTIdLJpQlGzl1+T4IWImQaTkmVcCe/+t71eeoaSneC8an5+KrhTvAM29Bz
SRrrIxLeQ29lcDd0pu4i+TnbmFKWI31Lfu67CjTu84eM4ywq5bgZySe7bI87lPpF
07xC9bwap0/tN6FoNHxy1SuwEhE3fj1ochq0UGcypLnX/WYi7idEjdf7UZ+EaAR+
KZpGHBohkfgTcgSxaR9wJ+Q/Cy7V5A142xrstMmuAgr28fihE7jAgpKMlThp+xg7
k7E6OfeBh0iPdvO4SInAlsnfBKnaj1sUrasXEaW01+4USlFEynAArDGdJ2x4QAIQ
0cklhbmVB+xvgsIZo2Np5LGxfEzVr6Swt6WMSLoHQ7RQcnp83U+y5RblrI+ZR4cC
3MTekwnC5m0UDT6xcnLXawtsIrq2XOgh0gAApeJXvlcl91UbvfCArmIsoulIWaWh
WWmJIVJhJokQk21jQMbI1shCxPRNHmYk+nUU0RPZ1T1OXpvWJeD2u8NWcwbiXHB6
rZB/H5YMTvW8bhOLnzrWAUT0pKi9NrDSg/46x3AUMKA7iOTZNVIQF2UCWl2+zWQU
0IOStOcaXuglwEOWFq235SiHldzQ2pLDMRou6aLHdIp6Z/q25R1OGGVx+Xv0fBVh
0SirIKdeZyxn8W9lEBS2msmHZBBBUzBogzUYVwVmVscOLAkGnr3D5tHxg53mFjO2
0+FbuSU7HFXRrk6+KgN4wGBMr/rhKxp7nxes2Py5E44uRz8mtsZ2qsuKLNdcA5kO
/eOT7MqCWloLmh9l/8BYNUokfb6Vlna8Ell8CatlFwJuhnwY7vbDQT7ehZsKgBL6
pmMk4tq4PmlKiJK+Q2eNnnSNEkBEz+26C0tN1W+zZOMVXqeMPISvdoZIVu9xkyc4
t37ufYMsF74npH2dPB2dKM0aACpF23CLRrS0BpK4nPOC7Ouuff/CResH8XqJhEiD
KUdJ/AiolhzTz1EM7V3ZQ2YHAL4JYPuIYo1xSmpPUhjYwvowR/kvkV8KBbqACETp
rZ4U6Zpe9ecpzqwggInn7KrHTC9+fqjZaXkZGfiWOKNj++Gb2p4YuS1bqlHkhPXa
GnfZiPBESlwS22fGR327pIdT51Ta6lQsg8lnjVFqsDWPFr0zaLT0cDfIGUKciSKW
/ctDS8EWvm+UJJCSjBiyJWf9DAO2fK1nCgjk0n2ddVOk8EWa2t+T4c6mDZAttPze
E7oM2TYrCi/1K2fUKBO8UjORwu2gtXZ9jwoYeAr3oaoWl3BRynaig8EqRrPHJPik
JFEVfHCvABd1/HExHbox/0X11Xe8HwPNxsGGXUP5HZVLmkhpEJaj0vperkW8sXih
hIvP40BoBvW8nY57+Bct5a+zj0uw6Kb4oocozWSURYgNJTZXp4sdUpVdHBCnCkIg
k26jnykKVF/F0sBbuJtU8uW0fxEo1F0pKxeoItuW0/fk8vqiesQrLEG8rmeZ8dOe
8Twofyh+nkJ+vdIetfI7g8NeTvjjRY1a6HPIiXCGoMcF3vNPVCv3asKZWFjfP4we
u1dnaB+2ro9p3nnNoZk42At18gcWEXOf9/XX+Fdd8BbxhtUNv7rWM9oRE/hjWO4c
gbAikNK+fpcR3v3r0ay8eq5g527BdbMux8Jy8KbB/cGASbPvsZ7tS65kQwvmEOTp
RooP4amrVOyAb3vK0LbB4wnG2EFFi8FTzz677zr+K+vACcukdG1patAtydNa82KN
+WeO0mvaz4VusXwzXFy+tZ7JvDzntoDSDtIaeQDQZPgHKi75rpEN8wWnaNXBkHzp
HuN4K389SpQ8lNqV4mv3sg3eLWodHNovHJfyg2ggfXKPN1A9mxS37C39dnZb+GXI
EojnAS/THaWfqWUFmThqgLjRYPcmeqhZy5GBHN/Uh596mXXrBmS/Bsc65p1ZEuO9
CAl9pbOrIVQiMqtaDvq3m6GK6KZaF1N2/RJnBqevc1jZs2n+y/fiRx2xxRnrXe9t
/vWvg70DqrLvKxQgVfqswA7Qpd4cmOJP/4SrNgWjHOM7Dmy4Hjl0VdilCZ4sSVN3
TEw+A2vOQt4RakqreUfF2gzpE0TbIT38k7Lbx9OSRHPrMNv9SzP8U1p11wFGLmXV
Kiog6s0wcjbrp4FAu+JrL6x0efIf6/D+cA+rD4K+cMk1d+DnP+iUG6KhAfazu5Wc
ZDAmvtf5tLV5Wb5ZRaf927LImhghYV/srA/7W6Hyw+rSE6BRibp5aMcAGtFzlc7D
DoLCiEEJ1U79F48tGtfB9G46KtiaH6tVTTwmLV1s3SlBA6Q059bHRYxBYb/Cy7Ln
THhfAsqs7FdPsaXO4SPogQYwSxVnOIakVO6xKRLywqSKeTnTcHHT7k0iz5/4QByB
hQfjGeOmZxeZZZpxXNKPJC2TKLt8V4UTm+VsuxY1ycxrDU3MQ0uGwbnKKUwkwNPL
SI5adHPpyT9vOBra9HEwfxHW3Q+O+3kLoE27O9AaMl8L5uCyfXgDMpPik5muCXp+
MOL6DTewqHKN8NV8gz5ymvYScBa0xdQaL6vQDlGD1/6oJlblFI7WGASWRqOIGd2L
3Iy9L5d+pO281K6cWZcUGQvLHnW87b0MPMXwUmyTmGbTGnw+eW2DD2D5XduwtD/L
ju6kZRWtrrDUfeJCy4FaDgGPYO5DHYYwjUBgtwYFVwXd6ruIgblcvmGlT7xtJsLH
XEg+59qBoEuxQiNqNU8QKFfm3+rFWN9XpDyFSmpFs97NyMCVF9cuOQ1Ju+lsDQZE
G/CE6tQg0vt6F1nvHjUrOd7a3MTdtjCDR4VY/Ia9NqoDhpHbCV086STJEYR+3yV3
7ye8no4VUCfW/s4awVJfs57mzhCCoxrwIVtXHKyEH8iBG3qZqLp6KNV9oAUjGE4a
5sdgb2U4djxDrcIo8XKMq9W69KLBK7dhZMXS7tgdD4/Q96f8vj0LtooVd8nxhHXx
chvwoFqk6gPpNhi8eMK9iIUlXqwl+v6cyjWcAdOHj2cepDNop/3F0d1tKkDic/Uc
t95ROJW7ScybMQ5PNcsjIJCWVoRef4GY9nt9L/KYAdAMsTqGAp2yKA9/Tn3itFNQ
qvmX4/uZESGc6mlPKxWfD1r7ckwfK+Rj657MLsGWwVpsGvFJ0c4URCLxk2fG4hpM
V6ZMDizD098wLEEyg4v293eRdKjKK7NL4it3fl6YjuoLUFqbBmfAZNJxeFoA+9+P
4GXTjHjo37gzuy0/S2lOQzA72D4zaQXiHrfcpzoFEvNSJfpBTiwizx612r23/Hbx
TkUCKQ2AKkxe4yv/wCOa94olF4QuIhCp8NkOoOUXxLPAU8w6d8cpZzE08xVjLfYI
rs5h+Mz1WCr8q5rM/gUBoa+VReZkS/Erh0j9pdaQw82i2FtHA6SW5xsl9Ajx4ExQ
iZeVLLqycn0uVb/4fUyXYMQJXAGfN+7TweClNG30UuFQhvUGHKeciiNyZSp/tDRt
jd15tylLlh1p7MVWz4i4ILsX5MEHfXuyTc3YuMDf5sJFS36HBx/ggi9F3gwxWmK+
mHsUGqZ3NY3Sb1z7Dw0+J4Pwtm2OCgD65Uh6QVy8S4a39wpqIQzq7qo2BuM1+eqp
NU5VMDA/BPnIwlAxqKmPxtUUTORcP83FwwAi76IWo+K6CmAdrLpXcUPo7w8eUEe6
Tprrhsjd2xPN23EL6saqQ4oqmZmDmOGD7cLeAanebSw6EA08fW+X3ADDXiph8C1q
ghNE1MoqxYRNyZJzVbVy99A/8agv6pfEGtlzwLT8HMNMU5JtBaA9U6qIvFQUIil+
89ur6i41A0XZhcQSZkAVEHxmaxDMDiz0pdSrHcAmnoZIQao7ZwC5Fh4hHDVY4ZOL
cRuXb3zUkAzghbYROoeksZ4hJnoj3GJUOK4BPuLt8Akmzh+pazuHwUAseQU1pZfs
udfAHtLzMQ6ULQJ4hygRKoCsOYGpGAgvI3MqPpnw4CJgl11siSrj5dEamwGAQ+JZ
ftSx/7eabZQvOYZuI+62kJjDFjPFTHBW4MCKXWcnY+HyRKi/3QL68oUQccQR3jMZ
MA0FojfA4O5/RxK42elt/cIhfSCsD7y/akYd1SSMLyPkIpWD5CXLe2IRKeAvETT3
l/ruPLJFZk40Y+3SO71fm296MSuvm8wOasG4MOo4RFXz0iacKws5daDjgv5dB0LN
G/TsyVDRRDZKiLsUoRjLTHDpM3PqeWsWev4pu1qJe+gPbf0gU8/JLknjT8mTVelF
WRpWKqNkNjXnI4PZ+3IcUgv9ggvicZHEtJm7ek5SPCPHqCCdztkY0oW8SGIJZvCB
Zfngyvw7b6qHCW/E/1QKifeqNasom9e7wQdvZzakzikFKsiL9SmkqFNsysjIM6nW
LnyYxDzYw11jI4IdcgPSgbYNiuhaeWv0jOECWMRxSifjx7NDWRST8J/hNnE/fRle
qNzcmgfOY1DLQxpuoSLdafh8+uoshxZ634GOUWnqMQ7wqYuGdxAm6Wh0qYWRdZfn
dxGC++W7IbEWbfwLhcsBMEh1+0Li0KIUMUTIXNONb6R8WVm5ZeAR81J7eWgYyNV/
D4pXVK6PC1Ya64scV1eB5YIzTdgJV3zg820HGtJxivvqtN8gd5BMzrEelQ12zPsi
VFfO3TwgSe0FMWTvg1RtH7wc3jnv9ykwKWxnMIQ8pDPW3lWaQh8tuol1+EmGhpO7
PRm53tEnLb+BKNP+WNv+EKWMrTFKiM2XQSn4B75cjyEuqfmSa1ZHa4Bg8ZlX/x4K
QBC9hxDaRFQrVMZdHgxL9hEz2xI+HY5Zu9OsvDAvmdUrCeJGMQvZXDYQnFFXdfOR
EjmdPJDJsFbRoq9EapeNwd9S+PobauTBs5mTGIn6dzrZy21iHviiHghsrOTbnlzK
iEKWG1IZ3daQOMbyCU3y3MDRPgVcJMEX9NIsHDenHVGba2VKQqr3in1343U0xmMY
tnEJUUPBe4V+/XGsxREHiUdujJTUB3aWS1ipQooTa+lgZ/a+ZC3tZVzu8jgaITMf
VHtF1XVVg+Q0CDHxPh4mIvBSS9f67Ye3oS0gricmuDyZAml0bE35dy7X6IFVhgF7
BMxpLrXfLjVckPiI53hJ7mqcuEtlD0wmNYzlIUA4vgFy4ynkPGkupYXNQWT2rXue
bjv/q6egqCeGN0nJ3tDh/sZUsg04xShTNZ6KBsRs1b/wyAr0ecDe1u/8PEj7iZya
WZIrUvi1Abn8XkIHwsivD/A0ll0JMCIj4RXVsxfUu6HLroLZmmUBksRHsyHF2rc9
mPyCg4x3iDVzgSzw1r98BaRUa5862VWjascPADl3VlX16kJXjAEKnlyd2tldEP2Z
TndsAiHLuatuGOSc+wj+srsZL7LhEvMP28wcYlWy7et11+ipc8Gp60zP/8YHBFzd
RluuWBQbDvitTWWH+0T+WcXt4CD0kO0NOLkzZ2S85BtaewgnRtWb/bmiQq5thnHE
IgX2MigtruK5MjeR3hxD9C/ZjxlGUhZRrkYhUGH3Ywu/czCJ81jr9sUIKlVpINtg
4m7ftLYyqT3I3hHxp4LkdPeUHdZNA4TH6KhpjGjKxNWw9bzI83BrCSjC36osviik
lojcZKkX6KjET5xEVCeJTLVzDVffqsxVaujtOpxyv4zYPrrk8HO89h+rMBNakIIT
YBx39CT67Hg6qOs6exGs1nA+jxbfAKjbirkdddAHraoQW8cSaumvEA/IGh7FuyR1
iEC29TLIyUi1FiHIFmOoEohns5MSbyrbqYIHjos7xIIZYTvgi3ECdJ06LGbf3dlF
symGzDPSyYWgDSdwInsnrB8YEDqO4Bpm7McUPTI1jTYsgVHpz+4agpEjFJAJt6s6
nXFWt3MOnRTZFqnJw+aDgtPJJg6KZm/kvb9YwwSIS3i/mlQdaXnQlsw4hEbKmdWp
qZYTNb1wzmL1IQj0nxc5phOPGzESSjjOIzqY40NOVKc+7Xb88X4Hf/pqIjgaGbzW
EuuTRstUX56f1Xnh4mlPP9usWouVdDqe1QYkFFKhHSssqCJO4ejwdRqtR5wbVKlr
+xHaUcfKcCCFxAIihdua2B7SprIORugA4zIYIzbqqE+D1c0sO0fJL1pzRbYpkqzm
ijqxxuyfU0yiHRDM65xhJZ+dMdOeYXFDvVve2P0SIZu687xmvV8DCo5oS5j7+8wJ
0walGHwzAf88PID1K2z+u9i3AMYxPBANfGS6ObbdrY9Pbj84CVjHBiDiLlrfWQ6s
Pfp+l914Mx5ge8o0BIiztuWB1d37MR5X+iORi3NI5/q1i6vH+RgDi5Kpm+gDJhzf
AHCLY19RLitdKsP2wV1qGV6KvIsvS1fNLtD1/RjW4x9oNL97BZ6A/90I+6dM52ZU
ta/JktsuCjH3mUr8tkNWSgDGhNygYjqGhCwLIxsclPigDdG/dsg5t1DfYikzHUlr
nd25x4BCA25huURgTpBIom2omy4fFSmWhg4W/RQVwtO2QVMSTeU0Nbabrp0XCKyE
Ezl4Q4MMwunblAPstWM3Mi1XeMAtK8Hq9uixdQ0hZqI4Eqlu8vu1WEUrwB94QEjD
kX7rEG5+lw4hUdEcDNv7KwytrnDqbSuBJgEjJxCCrsPQP0kiYaySGN/3DxLKtKSa
xennb1z+SMoHHBZBYuzp2lcUvjvJuCFOFhHrQe6yQ48evdKNOznGRFLXW5e4a/DW
O7EDVTChwedNEDjnsj7nJtRwwkJuv2icH9UmC1pTCmwiiFDisEVMrK7N4NBJ2Gyl
Oua2ut2161GbplpfYVV0tLQJwTVlkxXeKHMYekgADp37LYuDSp5EcQjTMgqXASKv
ri0qormDwZ3NvjrEn5w9mnXBRE5C6UdlVfatdsR3o8Uc9Cgd1drvKMCceKmbkMcc
ljvA2RprjgskZNHBOn1lK0RBblYRVD9zPZcbK1+JXtm/u7O7CsgqMD0BmfKR1SM8
x0PQv2ojZHAVY0VnF58vHMa42qJ0/GyH69TXsXGQGnY68wWkDGkxVjsu2Jsgojox
mo9ignb9cL5AQpsvvr7XFlAIe8U+Ua70tn4NpBXAiR//3QpFLsbStn03d9TzOm+w
tJULQ9Ci8hNxQKw8iftlbNSUv4aSISkdWkneqA36F8ZabUifEcPq4aeiVSyOCtW9
ewN7+Mzdixsjh3M6N9xNm7NOGmSgXLCMEZX6DGxRuz9X4eGIeVIoBq2J6J3s0L9J
Mfx6CfDpbe7Fp0h0hGrFhaCJcKN+d6W5Yc7INKzOvrAqvjvw3t5nMCBu1gPPyQNr
k84WWvUe7lYRbaMSBW0nwd3dFK0KSBCtyxiQSBtw8GBYkZpoa2PaT9Prk2X+0z2E
jrmWefTprLO7C4OfYYNyM5eiP4t8rSbQCmfBTwY+JD7Q4o0aP/nqyt8/w1R/ZN9v
tgaPZyBkrZPpzM6VO+qi97BfCAVnKzj2wXg4Ei/F2BxC7WRfCylrSh/xKbytNkPE
lRIy2kVp7sdH9oXGvxIIhd+hGh2p7fbDceTXriI3hb4dXsVjRPd6fCcKDommgTx2
VYMZgEnx3nEvHZbeErgBE5ubaJZSTJZErp1nKotLUZjI0t4Tl/RXiPYLhLXCHr44
DOiSKD0gp2Hq1w1Gb2KTWBOtVoV7SJmwVdGKXvPqeh4vPpZ2JXZQS5zVUH5x8kK8
+jE9Rt6jvZRcqWs/R5VYAFMpSv7nwBeHU6GUYckW/JUhm+pXhFEURFb9sYiuX4Z+
fQoZkzcWqk+5p+88rWuG3spq0ydHNR2kSxipfBraOhoZKkHQO8lONZ19ipGtp5ez
V+M7oOVMGi1J7fbanhMVzS0bl3U3HtwqfjuBfPO7yvfxOiXVtjL6GYAwR9BjT60P
wDsp26/3NWWYvT5Y1sqeyHrk6JdUH6FqJvjJ300qvLWuFhH4Is4arOrj3mpOYDhG
Q/nnTA9kPWDIzTUcFsVWVpTKLn7ETB4p0gmpP7SUuyZQ+TYRhccdv1hGKiCMdauC
XaxeHkjmxb4SKY1/b/UY7m1suMml0ea3tvCMrneEW0DimToSGbyP7OTb3g62cHD0
gmAOwlbWHV8SQXadFmvYGVVZZeGPS6xjXuf28sNei3QngCM1i2nsIzlRW3x5B11S
KBaNcMljQOrkc2D04X2vHPLlyX/ghq7AgOWTpr8Tbwzkd9b2nHyurhhOv70/v7Nv
i9GUTf9ZfGPWzOdNBYM1cnuUr/u7qK4Fir/cnP5ElicYh/8Em0ifDNJB42zAbBh9
gxnJirsO8r/JatowalWExzs3MxjwYdKA29+y0CQUSbzTW1p89qCrmoNLB94AbyF6
YR1LNSD4S/dIiW0wU4CUrQLTm8+R1xiomNMtAcWks0K5IgH+snD/MyrDH/HvrAaS
Psl5xwuNaQNYwyqGMX7A4vHV8zu4921W8wXtOtAvvHeoBh+q2RUW4kchiDycSuN3
7sAXrw2YFqVe6jPpkPzp++JnJntFGUq7rldwY/aZKVcWWk+wxn3yZRQ7H+yp5Z0o
58NqeW5BTRalmEx/qxMpS1qOCme7mxPNM2sqWU+a/jzmwmknp474ii3gqwwfJD/y
Oe6s3nmUnLZmjkF02FA6za4bOEZijQ2uVJMuQdrPga0Zjc1cjx0ErwJD4C7meOxw
Vzs1ODEWIyn/qn/XkBkGGqKmMFvchCso/4VL+zOPmJoIhySfd9IJOtuivv5qw+dO
cV+i3oySpyTM8iv5JvwaoClF+wNmGXBNw+5xYXseixYU2dcqo7h3TizFUvs7xsLd
DxaY1h7fNtjL2BfVe1sI95lbgwqsSUr52G676piMiiiDmbKda86Pbe4twC9Xe8i9
xKZZ3MPhCSnWWI0WcM9D/FVvjSiuWH9VZ/4zCh2+EUEqj/GayrO8jvdA/Cg/0V9k
lZgHPPbFpTc+PaxZQOdpwUFDickboz9NktVPyaIL/oXOMLqNZXOnbsNVzagohVi0
FEdd+YsNN+6HGWF0CEzgxO3k4akIavHf5CJCs9yhyZg75rAiZPgeJc+5N6/+vLy4
ulQvV+Y5ttC2wHOapuwGS92ww3VuslCnIFdpEL0dzL9Ld374tulza+n0BBswyo2t
0XqrfG4760MMnsC4rRyshStOp0NzBfSRiaSyjTWQwKvSCA7te8E2U98ZyFBaLo2M
0MU3hw8e8hB168uL2qgJ5GTNHQl94JVuGTi0ANc3rxn7YiAgna2wjPX7j5hnwDRU
JyVOFtzjHW4khvFqtArY7arKOb/S+i9STf10t2c8fNeJm6YkGo1RFi7WTjve6iHo
FD/rp3P7F4Tr13AaNNDT1tqQVjqJDwktV0Y6Wa2U2HaMsgo6szt3xH2wuCcZYI0B
iHqcBeg/55UqVnevOcJnbKIl5Od2xQf3jkzFEbPD9enKuij3sLyGco2WLSzjTZn8
Or53yff8G15yeSt0U2LZwOT3A4KGiGHTPCJXxdBhDTjc+HGDyK1DV0xOU8NciqDU
2f2wXEb/Q0+O28xGFyYaPBbTefeAHm+QZT/vrAXoERGTSSlLzrSXjlO7m3cVyOZ5
hezRBmgj9SwZNfo8tdv/LdqteJr61q/y5m0GLRfxdNVNx0aauHde6qtRm9CBD1Ze
BmlBvTGBdzM3mD6BOOYPdN6p1dS+h73lZs1EmJ2GJ9gKvfeRLv1tz2DvcdOiETlL
tm1tn5y2ndtxv4YsuZ9DHOpjqHdsLvAKKFcGPXB8hBBWoAOGR+Ek+SXa8flk30U2
+GTF1JPzPJIP3AXlrMMe1zmmfpej6wh6qNXkWtc3+UeXSEduqQoZb35oxxLbASfH
7ljV6fR4XWVRZWF8d0JUXhaz5H9L3u72ML/51aPW6J2luOIDbIFm6Oo6WaBurLIf
LP0UwBOFeEx6M7ToR0wWx+sEmXgNNCY6pUfe1dPv1BvIOrzLLTAqq7atL1rXh3RK
fB77nuf5ctEHQhAtrGTk7qSX+bcTWMg6Cf2TIrD+CqZNL/SIVENpYgX+CtNHhJ2S
ihzMSZj9HMEkuLZaxK5UZNk8XInYVDJwFF8fWwKSu1UiSyrjuHzOXQwHsifAabkw
xKPqDu3gz2ePDVmDDJ44SQS6cslB239B7M7r3adtMZuvZHXRoGSxTL4iTr8OQz5q
MO2WTlhOK0y5xsV99pdDWdPV+hG0dcgnAgOQYFYg6D+9IZWRNpN87fBsDumxPlz7
U4kIRFIllkZmUYeI2y6x4vx3VQ5SPp9rQDziLyx0yadEHQk0L3PfuB84jVoQ/66z
dBy8vZ3a9t0kj3d8xkZcfKUv7h1IZm6337fE20MWKpElOQOjxNmHPxIUwsXKhawi
VElr/HvYSrMTDTAF960dGWwtFSfTBq3OVKKYq8xG23MK4+xFheDHNyKatU9afK0H
5tO9HWR+BFyNT/GXyS+aGH9HHRWngxQiNxWEc32i6S30lpNwOz11F+V8muo3vCQ+
uME5KtmtdEfCC5mrx10mB9m5shWoo5Z7Iv2TUbV3jFiZMMFaG8j9y2bV1UwmaMEY
LyS+pfGVMvwwWccdv61s5Onls96DH+9U0zjklzkWImACSYTgEc7yprVQE9fOvyvR
LmDRBxsVH+DLNTqBSR0jxGrlRWdafdUNxep1ozicrLb7FEa9bLnQjHL4RnHSpQX5
hWPtmAXCtd3L1VtiVm12N1XH7q042EGUJ7I6ow0WP4UtKQHE8SOjgYRgCsz3sPfV
CoQkRjeXUK5Y2tFrb8zQJT0QuAbW3DTWRBD1EI/AO94QPVoug/zKNIIS2fKluRY3
zj7aWtyJm3tbAaD2o+EzvIoA3/gpab4fwZcg6acA56i9XlRSyFaxI3jxPpyliwOv
7tjlEmha5HJz2f4fHGjGbgomKjYEJanM/kM6JqrrlzRVWaZ4Cq65v42D2Y0zqF1U
lOWLtaQGwfi8papyOYA1UU+9zmGygM2HCG9307bdca4Aj5LBwl8OCzS9YMoDv1HF
4pRrk13rxVEPn5ch2iCE+NjE/pcChFTvtcV4dw6j/kQMfXy4bNmdX3K9mt3A7RB5
/9stkfVgiDmVaXABExaleyuaMrVqahNisZJNiWvaJjovZg17otaWrNmgA8GmA5WW
dl82mchzvyhHELiJKZ3FujvoVgl/k9+oDOpgF8kKxJQSrMbm97TMHvXAU+fmdV+T
2DHRNu1RHTG2+4af16afQp8zSZ14veervvKUH+6r+5T2eoPm62xSMxh7zWPD9fTZ
nQAj/ZFEPejTtiY04uN32bxHgt3Gt7o0dPhJBJIuS4EsASXZrrA2h6x4eCsV9Uea
utKFDkTVsuHHKP56T3LoUduCv9J+EpFsYGcGpA0S1eBE7jSI5xYmKxKVFEoiod1C
xZirq/6ZruXg0Uk3CqmK7/n4ff3IP5K4dewUEDusK9QkQx0yc7PAmJtxXfwwlBD0
T195g02x421X10LX3FVwwwVX/jPW5UDmwqAIqQKAqo0eVkfDZNOZPhduH+cHIPbx
SC905Pgt3AiJ4hACnIeQkSyxUBmoh/OcZ5eUpCYyvUqOwbDefFshEmcca78gaLvF
zEJguuCrSszgRW4GSL3GNXjxmCVt7MHxn0skG0lLm10SV3mHgZrn+p1PUn2yOFXC
Vq7ZsqQTU3DO1pzEJFOlh+H1N/h/fsujzDo+c2NJC+EQ4yY0hvhfHIVZXBEWeqU7
tudF5/7VdWAjZuZhqA6HGN4RtNKZOoctLVIoYbMGLU1qQqF/aY3nsvytU3oPUDwd
5ZR7vqGwN1KROZROQTWPf04RjsWgd8k5XPH3nd1eWymxSBM3ljoBxbRkNa+d5T/z
LqD9HZoHj9TZkxsOie2AoJvvVaOmr52ArJW0UVgEkuEq7eO9O2Tue8/3nsjAjzIk
KFMiQjwYoqc2IZhCRUhGxjuANwaY/iW3VAXefZYMRKlMENB2ISzqpmwnexMCKQ7p
kPa434F4+UW5gZpOs8/dFIrbL0tljCHqR833YHSLhPn3iT1vcPyTj1nTyFsn1WV+
viNfssP86bTe58dZnZP3+lPvz7RbES68VvKDL4vlhAv8JnHNfPdPPxjcZswG4DWa
AuD8SExTNxePcafm4LjDZ7cFtc4rRVHP1EghPRCu4+JR9Ikphu8lN+13pCzU75sD
sXLdBVI6PYNpYTPmCH7/UpULhIF9/hPs0iafSJIyYd0jrY9zvmqmt0xuqgNpYLKs
YepajSckfPPSUmfQJakybx29GR9SzDdOsUyKr9JppQ+pLlkhWivfVDGbAh5KK6kE
zbeWpVxqIzJIOj50semUd/X3+iDeVWS0WDyXIWmoozpi6PfzrIStbbZryRWse/if
9K5SNYw0fz8U22AB20CCNsKyfE+uyYvnx8wudch7vN0zGixG27D9VxjQ7H5JrT6z
RPgOCNXWdQ2MKL8ZSQVGh7VHuSgERM62h2r15KSxmAn45zZMH9kcMdaEouaOCJgV
Wrzoox6tx02hYmMUztGOzdM5e3HbXzgQ+fJZOuMV8NWK9s/oj6EYiUfzeEgRiVaZ
TJHiclJUeuYPWTweBbJe/bzLk5SGOzD0OdPR6dCE61VGJgdSB7RDs7+vhbw+YyjC
O7B8BgHUL1koshRPAEpIUbwG6NhfFSCkis0O6HbYGOxj4w7Q+PY5RS/+wD1U5c0v
QH2m2+FaBbaoReZZNIMKukMflEep2zu1kQYHHPFgXfAaC3jJkxSV/+dbLRINqeSY
vLDJcI/HUlTo1tXLk9YvZz9k+ONWWil1VoETqKJgEFyGVvBGAlMlmhAkKVaC9azr
qBmslPDj0lm4iJULYD+g/gxWAqkGf0W0c9QDuGs/6Xy11WXL4xdOePNVPVclmCzD
socG7TqKcemPAfPP+QbJl8FJGzTOI30MycUiB3pMAOdFPLM+afyaOMjPg+JTvlmY
rYQpVS7WYaIgSiyLlCOVVwMvMraE/g0QdfGwbgE7jBCS43rB3cufvJwSro9QTdy0
PVp56p84R4Xw3giNcubqbaU8vD7FnUJ1tQ8P2u5hNDQOsaNGF9le3yxtdyC3EteG
w5jXRa/hA6keiDDjYYBqZRd05SSAQpNti99SfqOokwt4VqqUYVO9jCKzteZFvMSK
SHwlAiPz7uEGZrCP29y6MnZUWXxJjSu0WgqlH/TNshchdF2OPwHJK2XyMjSihgAY
InAuaOPEE17UHUoP8aqTmCwepFWeUaPdGu+euvSsXUFl/+6aE9sUjafEA1kmcLtY
zX+sT6xSA5Ar9syveuq7E/+RG+h8BahaoSD/+4YzZw0JajKLewzMfsw0FPHPjaNA
+LPqAEOWttkAeUbq6cpsgsYf4BoFWb3ULHm5YJ5OaUcnV2B5cxO3KjJ1DImy0JVe
BSPMSsxEDaw1qMHLqdoBTuJH6FTEWjv3L10hsdKqyB530MLVggMd9VOuSIJe7n+I
a/+M04Yex6jY9hupFb7roQxPT10nB0PaE9T458ghH8RjkxMZRHznEEVVr9tfK0kP
8+EFcZVMUdBcSNQyucoJuyKzg/UgXhwyxP0TBcrtcDcd1TgQxMRB/llug7z+rSLT
dP33eUD3ZpPMRqeP44i64u48C1mgoiq4Kh6ZX9JP0RmqrzDIyBezW4CVXRWT0cCV
9MQHc6nud5DwU6bipIXq6wbyfagqTB8iQWimsUJ2UL9z55kawrrQmqAV6uEdHq7e
8XqQpm0hNlCjDdPVj/nZ4XRdXiN8epnpJXm1YCHrMOnPyY+p8CzWYWQ9/O9/QbxV
0Jzn8tFm49rcgEyXGi9GKU8Z9+LFfDjtPHd6vtA74OVUsMKHGqgD6ZCqJnQjZFOF
mQHN0iE+Sh4Y0oYcB0NAlx3PQwpT5vWbVeu4JguvRH7AF7V+sQcf4gvKGRJ8H7JD
0HCv2Mj3TYES4zmcGQ7YfaMdlC92yXeIVwtnIsDgLvGbSGoYoxVJL9XaoEFJZZKC
aAqKXYpU6YXSGPgGs7NMg4yFnNtDsqJpMAR5e+KFClFBkKVH740+ZNHy71Oe/MPv
79LSWi9d/dniq7bkrPiTDOTfXQBzfHqn2cCgufY3+zv6YgW4PS9d+PSDJDyGyo02
zirQEmhU+CxlZepO13iQyBFkZQQ3TMK1C2eXMDXzmXKTqTBqnwb2dxQy0jZ16kUb
V04JAJ5ogDA6rjwi6666XxT/urhFyFUSAZtoRdjGWha1k/fwFXGrmYw93ifKm/WY
B5gl4oV559XPnB1FTAIUvvkCAgnZHmb1GRsDGL9Japxhij8EwkrFYg3+eCKhCFz6
L/x8pCyldC7cBsQvnWqE3zwlBiwuYaMDwC4P6wxtAJJ7b0tEUYgqCyhHBF3zwnKC
qxMSGgsRMJ1ABat2TWD4gtSVEuPYnXtffL0pG19rglU62WPT8ZyDAcqYDRH6wDBS
HZKvSaWUvxZXWVTAPognuwvlE3GAkSwoAY/0RlExyGTaTyIbKVCg5RIR7b6s5kQi
nazw3lbXU/hZ773A6a2ra+9q/+Vo6giMVkDtlXvnTtwEzncJ6mXd7x46EOBqQpi2
fIRPjZkWPh3qWIqMh3r9A9/xtKVWxSSSR/Z1XRIchNeSR7FUtK8L3qnIQDBel1ve
FWITPOte0vjFK8S7FHAu0d47ZFbxoQFYyOvEoFuxTFC1FVjjLrfWpESTwTE8xgi0
5zJIpbxCDv7A8XijxoB26yWyWoAeQVfGnpXwi5Q+S8//A7oPMBpyh+9JTz02EZyU
yBVCmDyJwE9cg8nusMlFxP3gyqkTMBnZokCbJp92+eC9ELKbuz23JUcPnLcMBNZq
3NemwFHIvrHU0jShBkd6hvGcW3+hOm/zN30fJ+i9ZmgrdrnW8U8Wa2vapURkyXkT
fFjZzR+uHLG33qS5H8h8gZf/nl0Gx1Y0hTA8FmTM08buvkwxiqlLGvXB/O0eJKTf
xh7A1eqqr6b7AMZJs3tljII8u2xCGCDzDDVxvccr7RFz3lfK+p+OIaE4NPyBit8v
TT0EdkZZVTfpK9Pcpuzznz8b21slkgtcsErxzkqn462JVG4mnzc+JbKkH7OcTHyn
K58XqU60S7J7F9BKJl+igJdi4gzEixnFIUGDjLPPSDNgyht+LxIU1Sk+MEadIBSq
bKIKaBqL1yITT0FkSxoNdSnJpjdSJoDaJ5EAVc5Gts4bNs+Q4/5cTRUKo0A9P7KD
kDm1NZAe7XtT9ML/6/p/f3mWwyxBG1esl7vW0e01RYiDWrdiZunMRzt7vq0dQiJP
4GA7fBOmi4x7s36AF7MH8JrJnt9DS6cYWJKQe+ojOBEhsEM3I6xkd6JztaRij3tD
BXp/aVEQOwl4R+y6YfP8Yq6H+EX0tZRS4T9Y3Y6XBx+MiGf71/lyL1q2cAZlqHm+
tv7K2V24HDQ1hwRhwnU0lhEJEcfNojuYxTU6FCwxBwv+4yEajVfGhS2NYIsdeciP
fjsvzdxlJaW+JBTKoztpR6YRepmidW2+aSdN7hZ9Fe9L0Xnl/7Yv5zMthinfDLiv
Vk22bcKCIQ30R7mAQTcOycM+GeR+qdmIaG/HrZuoEOD8jH+CjjF5s/Ygu/FjvSw6
HgA49U94MvumOD/jTTqDiIT0xPo1JWh1KURzWh11zt9u3c2p6efKLe7E5R/9N5Ar
kvKetlD7Lu1HlnlV1yGFWzU4LzEUOaaD/8sWby9floGZqQ442E1Z3ScFONKONB/i
Jj0s6UjMfHUjOy3k/nzDajR7Pw+qtTaJ/RD8jr9dKFMN6frUGcTzTjfEscl5Q1/R
LVmE8ITetWUgGruGXsghOgGA0HCUOdRtdHZxa2WETGjX5CgqElldcLA68sZ5GahY
XJaPPmZgLCmTGky59L2TrSSxGaSTW3ablQryGSZDOZhdXvFfYAlKBfyE4/8s6O4i
2V5ZhMKqONS9T8pbbAW3w/wdIIrAbxIioFcjQn/4FoGLJQ8i8i0bpJGz38L0y31w
6lb2yeY9nYFHbzwfamXgybdUS7UmLA+WJXY9gxqBQ0VvcZ53e9y4jzQ9MpWEa83Z
dCEWqTE1uLro+RhCuCDNk+/c/hM6BG/mQxXQfiTDWetoMzR9djLZlfd9cPglKsTw
pZhnKtI38KwA26GUc8qOmvWrT3xzYrT32VS99T9gUmNbFgbf83zd/ey+0mrtrAci
xJVj8H1V4jgdCZYMoMss0fqgpKq5QKwTfh6oqxC3+sgO2lz1NHEJO69DAAYKPbqO
qu3ndLISDCIJJaL9z+1fni5w9OfBy/D7ZhlVkTJcVDboBn9B7ndhdasclm70xNCu
OCrQaHgnmwZIdM0IpsziQrOY8S1O02Qtysv2OcwcyScwmyvV2Z8SRw9ZXzYY0k2K
DTJk8JCQd2XjNjKfdwfpdnkxy4z5RBvIB5iHpXmm03DCTSART1d0k9gvT5l3YGP0
UmeS1vD3KjxjgdEQzrABUCB3WBt9xuZQHDn9b4jlnMvv969obEMBGKTEhukjfsac
GfSVgN7jLxpuIfOZnwZevJEnmGrASnwK3Pq2X+GMLMmnJ+KmK6bLjutYPD8b9gCv
gtmo2Rh27Qz9fd5laLihJeNO1+RF+LD/sytgN+dSnScImkwV3aZ3Xi3Y3CGCxdS0
3v06zdVzEuxTJgUrU2T6vmdSvanU2IKARJTlDXdJSuToCH4G2d/PuMEpmvBAjXoD
2yWHb52w8JHwytHqfimzvWUP0QyvDwvR2zLVzMrRPOmJXHnpeqXlJ7Sn8+6nenlx
6NamwSgFeWmXwNRvxoR8IcLL2iK1ViLoNYE9U1jGlGNPY4cFtkzdIgxLYITXiuws
2tsHRspfzpEhnSqAn9HYADVdR2wVlsBF8d90iGBpGjSGaFhIgAh45YeUj7DlBvww
YPa2iwPCUZEklEwFTWmnTik+1kK240YxZFkouH+jpupgSOwLWfl+QJVMs4J/hBaJ
l/l8dtBJOc/39LU1+kaysayjHiP7wlRqyAjbMQNIUULco7Xj0iIvRER3Mo8HRYNY
awTu9q7QFuy8GXFZtVEWArCEg4lp79KwjwkG/NGIPgRviP7e4PL/sxmb9zlofmfG
HBEYupJjKVEc12mtE/zEi0hnJzvM0l4k7jJnhCGV7kpbxsuUrAyXSwcwEr4Jugus
JgJ3wgP2Xdf1DTkinTx+sj1aLbReaX68EZkz8DHtnIWAE4i+YNFOhnqRfuz0gPK4
EfoUXI3EzbC8Zy3e/WixN32/cC4vd4Lj2+fWUR+9E3Z85SpcppSmhPXalmAvnlD9
r+a61HMQYyICg7310pjvo2du/EYiXZR3eHcTgbuj6QOfFzZAkocaDX4TByYKeP9X
K9Vgs0xEM3YOU0+pIlcQalKOBiXp1iHf7t1EaUZgLomJSJiKKa1cpaEH/IFOvu+L
8Im840vfQlsII+mxIXWCF1CyoEXpW+wMjDEHW56+W6gd56AhaCSL7oBuRLj9aqKD
YxBP4m7n9raw3zCoHnqDzBH4cMPgHsx0f5KUVumm3/yTMSNKbs0BVrdNijWsc5El
rGX7oiboWzap1QWTFEps89mj7eAkYJl8QKK1SkI1x5LqhEShbDwWrA+dJmonNLTo
vKnUQ62AAtRBsCmN5SYMxEw3gss8ad4tMf39laDk7slqiKu8m+axTXlsLRHQ0V7m
AhfNstCogNdjTnjZ5myTE1YKk9bnaaI9AqnY+dMD1NufY7EwHiJckf5hpNJd6NQe
uJMLHYYikGIrhwwFhNQfujvjv+oOdv8usNWYuKaNx9nqH2+1DCvbmNrssZpsNK9g
+LqOA9HtygNhneBvaD6asifbmD73362kgzITUbGbYOzhUB4WpoWFpT/smTw3PdLU
5dUR4P93jOMOiP1Zd3LWBMz3zopoRUv3jbz3su62YYGc9nozxjFk27O2E2IDM/ee
Yt4IqypZjTd5HkaKyiczoLQJWwkd8rG0kEXgVQ+ePq5W+G934WRUYuj6oczIGZPE
UPhOBCkO+e0qtM/jMD45YKVwU4clniLBudIi0VA5/5F3O8RBD/O+LXknq9zVS7MI
pjoSDcI54BBrNIY6X0M6DeRiH4RxyUsHwV5wnzArZbEvtYAPlO8Fkl7T8GrMo9Y4
GPt1TywRvnpAXgcl/OijhvcaG3HsVNv2B/1POKt9YKqBZ131FSc8T7/YyLJJkdYm
ycAVakVI/6VjZ8/8GdThzgj5p7JTlHLBcYi8/4wK+iFIUGWeUPy5G05aP2ZR6lnm
DINCWx/ODMeq/yH81elW9GdumjUCl2ZdwC2JP0K92n9m3WHSvymGqTpCLnCiQ/f2
VZHqqBFwtpsFEfPV/VBYEHmYFH0f+g+c1I4saQPyJgWychzAi4oWpuFYhfEbjc95
+cbbeVpvsZKM3XpfcLlO5Exrbm4P+lkCDNObFD6rpgnE84u65cAsIYMJRpjerksV
f8sOE5rOJ5zJxvdCWRPHUT+gEiBdPj6I6zEQbGvznlt2Eq02HgLm/N2qEURjbbuO
N7HXnIenctKzg9eemc17P4MiDdSFborYk3t7iNQ8r5G8spezHCizf+xwmEreBMWu
9cGE/w7yraFKsUnRosdnYQtpbnrA6UlcRMTZ3LUUKvB+MH5webSyVYfu98TaCnbb
Uj51Ei6t3ZY1ikwDyQ7srGjnmvMZfj+FFGtaKeXtrCmnhWVP6ObPZI1hYfQWm75B
f5Kba+ac1Lmq1966OP6jbEYLEHV5QKGpP6UNkCvuYb3U5yUeo+/tMj3u+mG5mWpB
IUDnHWm2uhM3Yh0TO+WP7vjPwi14Rmx0tOEGuOqGz6zeFx/scsZDfvklxnJy0c45
9Qzf2sNCW57O3JgAdNCqrEn+Epnw3DtSSMmcaQtFeA0SByS+o/z6DPmE6jNhWNLo
6lg3pDqgBzk52iY21l8CjW2/WB9Qbcgwh6vbO7jvaNtwF06bnKPiJhsL7eT3wDew
coNZ+T82ZdkwyeGcp4WriOp7XVOoXrIMjIhwsW6jyMbk2vTjffUiQctAWWMlfXe5
RF76nx6aTpCRr3dFkCjDjWSEEjmsyzOVD3VL+evPLWH1VKVQw7FYDkV+01WfTFAB
KWAKdKJWl6Y+jeaHr1YM8nZF7US0w4xNZF2B8cgrJpL77SEo0ixniSLn6o3rJPC2
BYDYERqaYZ6bq2LskV/HqLZ564rY3cA3WPSXHcwkr16wb/wcOsz4q1Rpn8HWMVZ3
yIqV/6i+10IhOznsK9wGDrYGSucGXQCH5sppC6/JKJbWC7kNfKH4rSfzCdCMm8nM
QmATIqLbpNaJtmFk8l7NEzL5eIhv486/zEhKewDJDk++C2DFy5SRtDu9aeDkBxCB
FXIZNRyzGhQou4DkOzBaDEkWwsaE+QcbU1UCZ0bQwdmD125HnQax3WO5c7u2xbpA
q3HxOic3U/pK0+NoCLYg3fRcnqWdruxf4plLnuxoKxtWbgbOyKN1BtEuWQdcYOJO
NIdV+34BMvhQrlYmFHwbS/3DwP6nUnuhQZ+dq9vjVpC0sn55aYUrsjtkE730FMyD
dRJ2lcmDbwasP8KwjRJfrxqe2X8/rTKSaJlbUChZtHJhpu+wqBFrPZk0CVD+vWTx
ISmgnyC2gto5WslZjYVzUYGCzI2GuIpvy20pB20bCsTBxMRI67yvPEwDlJeLCq1O
ipVVMOVJcKRP7KHGvSYOSs3b5h50rWRVQpxWlNzp4ki4lhuTosUzh6ZAKHlkx7pZ
c8ETzBYnEBkQz4gicbiNnTzrJ/kus4sFtXpcZXqROTiZ0p68WmlVNmI4FO8ivy4v
ZpKhHx7ZHRcFbUR9q8ejifZOH5w0pQBkijpvpmWBgND+19bEDSUzZtGU/NYWchLQ
WZpjObWE3VBq0ziVUYLKNNfuJ0ZQUNrhMge6/Ec4upttEEw19oghms4AtWzq0TGt
o34KvFXlrnxdo1YvOZhPxnQp+n0sLPWh0tUSgcv7PNJmVxcOh2RbT6RLMzzdJ1Qb
79Mesl8H55ZiDv5SutgMbNH+2SyCNJgcH8XvXWXX9y3CAVKTZ8GKybmfmv1k/lf5
Jf35cgcB/PAO2tr6RZyWCETN8/XTpKRRDcEfA/8Mjx5SCqQ+xSLLqH0qEMz9iS+v
B90JIFg0cWQJSWgTzHpLrXZ6FZKHnVu7dmpyF+UZoKYnq6rB537iQtb/LsUOdY8G
7h+j469YYRFe6KSa9H+WNFUvfvaQV2jrk0/KcqZUhYu6utqUsC1YcMjXUqUiBM3X
q8SpUd2dVenSGgVq8K/AqNIoEWu1w1Y2TZMiMHAhqFFHdMVd9C7mD6eC/fAUIRwM
lp3BmBw2P0X960LkfPs4rOdFW1XP8T2a/kbXOXX5matlN+0bwU97o7ziTLBqYCMb
Wm8k1MAQ1cEL7MJclRo3DjEfBMCJKnpbqBgUVZcFHpdPjnShy3NsS5HYUX+KVD3B
kh4Sc2Pg94/4WnqglARpluFzFdS/EUJN7gSHFq7LfngW/MfBIzHThUJrkdTmdqbO
Wx9N9jx4t5emMHeW79hLBwVyVtkdWeKWbd8eZ+ckv2ndF+qIlsJaCKUCJfARkYNU
uuhL8ICf3RehV9McUmIhNH3ky31z9oeHeo1mcnmVe8k4kR2inhaI3fh9p3wtcCza
fOdENE8b5NKxUIEuLvwRJiebmgflqF+dAT4huMzqRPvgAVegjcTQSDzLhjS4AgeB
vm2xxaysKI/E411YIKhvQATGnns6Uewc5WbXoD8I5IHQfOSZN1s7aFS5hXjkNZdv
gLfzPcABRKmGXOeL8FhLUocTSYKnjGDlc1otTgRKEuMzNl6XKWLiQG5O6n9Sf2hk
NolZ7L155XP5G5s+tuBMxiZDzOIBi/zHt4XaytJ8PgJG9UxMsI3Ng3M8gN3c0+GY
xPsNfxkue4+Zi9Me9RLhqITUsyKGcRvTEAIzmo6pXSiblxP7SjmhNDuxsVvtwUwc
7niVboNP0ZurruUcNKzcK0RWQASpJzYJyRZLlT4X4b9aTT9FxEcFbSCBX05T1rDr
x/MCOqzbDmG7STGbwnqa5dKLI6EWQ6c2xGQQQKOioa6FH20yeCE6GmaZ7XxM+aTl
8rmRlhMIrX2HU+L9SwpLwXE0qDBGTmziRjbVVNp7kyXlS1xfWvAAvJpBsmLd3nES
4/IguDg1/F1JWFXWaHteyNHQBtqIprGS/8H/77winKkcsDc+AfU9fgVetKngeaEx
b4uLIrIVcAm49yJ2t+o7WU48DxKoJAUiP1BkJ3OUSC5sTY4W6F6nzdUvT7pY1HwJ
abvaM+o3M+16Ll+pdvWrzN6DE3MFw+l3eeQZToi1JLEa8cI9KgL+WfeVPMVrtlos
FGV08b/Zkvg3TfXxKond7VXYyAF8Ey4xTlPxlIP2XdB7+0lrJkECm72ConZR7fTa
tURA5TjEcDMk1e1EmLcPYwjHQL+gvxA6nkAHf1DFOnJMfEqry/Jj5JksbL9hN4/x
p+sFejKTlsuJ1jUuC82qhV91RhXymCpc9yxd/Ovec9ahwRlt2EruDpB0mBNH+PRM
eooOJEDs8u227CRim2Ox0Q3KbKNuWH9LJ3OmFWs+/QQp8KsNkKmTxk0OAxcwNrN4
mHHatjBU/RgUCIe7ZML0kJIBsDJvuyQN1Q6vs9Gk9WMotmy5QyWCBWnYwpwJeNZo
cRkcgYhzZbAV3JBrRMd2SFBo5exM1OdmWTDJIiA/xdkuHgS4KyrruQzxxP2piPA0
xv2xRDFeYBEGiAsw8cgPN7aq8hNxnY7FJaXXzdMuzvnOd/4ldDO67NPW58L4LaDA
RikwUDdP5L/LPpvzcF760m9+wolUKVOXY79IIbXju8CGBzHNBgiz0eqwsj+Ps5HA
A7tsJHMJlnSU6paLGB7SCN8yUidBfF9iBKD1RDwO2HqmWxcqGHhTRtGdsTSqK70t
8yxDv9nYYKPjM8W2A50FhnZhzdSzMCN/5t/87REc0lSHgB2PhZK0rhb/Ak6jHywe
/rAb8t4U5zzRAXYSOKQNQmPixArbWtL8I4iIx8zqo0zEVjdrnpF1l+sbnMPJ5mI4
w2I72KpfB3eYGgckbQR93yBNNoxllRkcX5Mlcu7pMGt8f5fuaXS82eUYTP+dxb7H
MaDjuG3oGDytkrVbOx6eF2Pk5IgBGoYFlbkbVwiP8jedi9sZQHCrVG2Gt7fRh5nT
8cvDWTOzIoO7bKVQ96Pm1+rFYshUnS+DGZ4UnLj6P+AZW5zh1BuaBf65zGrc3Kyf
xPXy5hl0vsukxIHUMT8rDTg3nmQ4TCXukOgWLpM4DifWPB0/b3RFBOJ2BmXJ95mz
aQu2dmzpCFSGwIt6xLRMm03E1Mdt0NR8nG9bn9X2yp150YP06kuzVE1LQdA0n0+x
Jh/zI5n8/9QVU6jiXY9Z0ulLbFQmFyKY7yXa25oC9jexMWblXhAb/RMRCxwy+PFF
L+kkQPejUQfeEkHrqWz4EtANrarcNaA3wSUezVpEZ4Q2SJaW8BkKQxV4QTQnbLtI
bRZ3jD0ujyNNrNBbZhsHbVROKxvTVxgclbxFjeWkATAiLakygwh6jhvFyEWVdsuV
O6HIGF7RqOPrVKsqsP0nnm3XsUSqPRL1ygPxQUS6azIU7oUTbIj8v+7GCNXHhRjs
qyOWgg2JUO55tXASRRsXa38kQuXGCxEssIrumQ3I2xA4H7Vvkq5/4Xw+/SODT6Un
h3tnu3QTpHR3rO3nFBmMO6tzT9R0aKZuNO+M0r2avuVA5yM1dTnweQKaEC0Q8HCM
G2qIz0Rog9GPcoUkTlGoigdHx9JjKVR5xxulM9Vz19QCBLKCVzHPXYVx4wfUBnmA
vkbyZ8u9DXVd3CGZ0GHK19SYY5U+aQhwJCvsxNkqMOtiriEL4NfIF6xpzKye15U6
ThHKl99Pzd+sChA1aIwunIvml73GQYwiukLaAOJYbOcfwBkKdJDxpxlhvXA21QX8
ddYA4ZFsvAz3Zd1TdsDaioEHc6o3NoRp57bs76Pqklvb6XfSvDb5M3wzRIbr+inP
J4Bndd2IB5ZB3e10iuQtokvVUT5ln5IezkvISRsNvb/xeT45W8ASWUAkkIQPkb7C
hC7xtk2eVYjGt6tViINfD7sLG0GR2mT5bixQeyZEksMYbiNMx/cpUlaGOB27HE06
sGI/F4xxL75XWRaWrHz6666ibR+TwHKqqohYkpV49XPuRSw3JxF35ElqFy27y9x0
gjK5crxgDtiST+yZ8oLncS8L9bVKQ5ybuhtZYV1+aTO6ab89WI1lTLT72714QR1w
yXw79EFFX+pSNmHRJ+eqcjEp12uinyEZJ+a+wL74Og/qTyCwEeExYlS4J8aTIDP5
niu+QquLivOcf2zis6XSM3LW4rTE9ubS+tHGLUT5QTvfQ4aVyJuciV1DpbzyDt3h
wFKPy4vIIcav2EbnTGo0brmTgq+PAvtfIsy7NZEjdDXqDrazx90/pxxYzUPBci78
u/IuBSOT9qrVbo1xBB/DoSd8obqMAMw+qY7fG8DLd5tk5I9D3XWtBoZLSdWMy6NF
Ne31OPyxm1HTllN2WAKbfoGrk543H0kXnSWPhUYrR5oh6P10prxxg4KWSyHabosf
A3rnbcFJF+Hpjodfm0/EXSWmiPzoZEFhzds1D3CVnlw4H6cBOx9vjZnnCfcsb5g8
exlG59orXCuEvdhxoAQVEvRxWeBbqOpGYGh3Socm2oiJwdbCSmDMLCPCrSO91j+d
VQT7Gf1uwoZxOb7wcEFj3RocsPy+zW5HSZTDw3eIFw+MsjDApg7iLrDRMtAP56Gm
BPyDYT9TsXRt2zCGxwXpdEMbU+IHV2Iq3c2bsAhNHqlvZ4nyYmDDBfMgL967VbuB
2Bwa1irBiEIBj0TGhUiB/ZJiJc0+WNZTE//ORD1NYGuEyqfVqM3Y9lvap2qVEuAp
Um54wJeJoxdW9lfM11hUv+M4bfLOb/jMmtO6wzIkgXe3Xl1SdtUxwZCPPVrv8UpE
BseFpjbAjSHn0ywk8F2zirGOJwwSQwoieXjV1r5VcSQkj84qeOaLgWNZo0AX2DgS
Wwm2O+eUfgeDqhhqBOeZTX9OKgoyBj4PbJ/4AJPNCydFzrqRuQQ4GfLV75v/NSHC
AQ1QPJ1rGDq+s9ORUghHlR8mKxWipNhgDSYWwF5GWUhQox8yYx4GE2yphHBC0q81
vFqisaIga8+Id5ktWZ4mvgCaBVFxjl6Qo/R/v8ReSIXdjHGVVsZb0nTdzpqGIdGB
ZvMLCPXYTWDYXl0OpZIkxUWFdkEo7NKRjI1yA8VQmtUVDL4TQpi88iW2vNUCzR8M
FBC/24+4HYxrPhmmt/0+KA8yNM9PdVsmQZt941HvnByoyhy8punOCiocVvhPlby6
vJlU1Rm5JJbLXLscwJmdYwwsAjkEPj0vYfv5po3hB6Hn9kABHtMIB7w6MAB+BUd3
Xfz5tve+XYCf4y/bAIvu4p6cwxw3AvJ7fAkGT+2HHlwf9FjMwAk338RXO3ET4pv8
UJ5sGcj3JRtX5kAQ9GDdwN6GJM7y/66val/G5teHr6ovIl9cI5BBTxUEwATvuVyP
ocZDs9aYamtqFvYG2IiB4xIDjZ4AUVDN4g+tzgdkwxZQ3rK515MR0MfZF9tEGOSB
UpRwQ/LQ8J3R+tf8T5ZIt6JG5/bYNhNymTG91jtvB9OEtlfSbED+XsIzDe5qgkzM
ibaoSkqTH9DNKsBHFdwrYcvFn57SEORUO4oZcScrtXlwqDR3gvRjnyQXfkBlcv/E
TwKm/ll+mQQlr7YVw5fVbsVSpcvJNtKESWdOvCsyKWYB0qz8280ZaHj01R3a234u
p2YBOKE/OFY2TFRAKddDHGkoTjSLCaslqNKZ9clsn62IdWmxXw0KA+E5OgdkxtvR
SRRVEvH5WcYGML3nsgIQHmRbhMaCQ3vRiAG2kXGnZOKVIc8VDOqTTL5iVDHl3OVF
RUG1cQsP4Y9z0COYOJidxt7q6b58iSxRwbLNWtUMEdLLJ7Q6LHZZFY/jK9G39yLH
HwVGgNhlZg1yxrtd4kQt8oKG6PEvEjl4lflqcReCUz9U9sSHVz8bkqwTMKyfMkXE
YV14Tpt8nmcMrsGLlV5hxhdCd5sD7P2p+e33CieAIeZ4q+0BV1pT3h1LcOIIYPsa
N5GuhXxAXzEKuMG4Xnhn+E1XpUzYUhmJf6unVSxXqoBBqqiY7fmExolhwJUVsECB
ka3w42ual+hgkcZEYvaDFSyttr13X/8/AHkjlze2LqLdbm5UkGfI9yKl/B/8tkGc
cB7NGBQame3/cT9xE66ZgZhU6F+qYf2m6fFWLo76n3lSQ5zVg7QirFzDYzFeI8Gh
VTNbOitsd/1FLcpyqUvdD5c0cGvurAfTUDl0yoZattN88yKYT2jQ3tFup23Z6Jsf
eH+mF5dWFeVvJ2/i7Q3gw9WZhO3NW3xZCQNyNOpGCh6tOlOFAUbiBcfZdumWJ/Ya
AB615rpsvw96f9627ajoRI3u8DstCLaultMuC4qOk5Of3ZRJeChHeRP/qOjxKLAv
sSig4jLi1H65RNDlHw0iSC26cNPkIa/FtDnISAoIP5sQSe51LJ90ZmqxM1IL2p0b
kw6UudyGVsK/6py6TJzyrBHjMO7UL87ylyA2XJ8xbkINjZb4we4l2qlhGoJ1OxzS
XKWu5/8vyCR57b0Uug91X/MnZQkrDgG5fNNhkSmzWAEEMRuQUsuWPUnbyzirLJvi
PwhwHJUgPtghBOQ/k/OfPBC8rnmY2vg8BPanEKjmBcHsFGQWpbLZVD7F68TBU01V
LNugfgtAP4UcyN1sJ4YfSGU7FyYU7Hi63ZASV5atWdTl01ldM0/mH7jJNarWdVys
kN9WsjO6YSQm6U7ueK6gZY7lWFSKhbLxNy0jlCNAAeZQnMaEZkP7BsKJtAnRPryI
OeuPet7DMtuOiRVGnnmbvzw+MxDMCytx4abRpvBPBeT4fivHdCSyn23v7SzBPzmH
jJ3R+fT7v/YD2S/Dnn1PflKd2iG6MGXMcisC20ddh4m25bDYa90n5XgBQstZ1/Q2
foKJFvdDUc8p3stBFX5YJLlCSWlUhQfRa6BHbyQIBhXZIltEcrEE4x6N3783Nunr
OOGl5t84/mEbG2THp8cyL81HfzSCVvntOjhQboWuIGAHNsW5D5Fs5Cj/XiHlvLy0
+7hsYgjUF7JyRfIGZVkFAJFNcRqxzUDDJev4IF8aM6VZ1QXp3kXuWMwEuDMivQp2
a6j3sVhziohAYVWylRKDOlbEW0xGWstWPPa1fpniFYPgJLm2eSNMgPBWwRdhtqGN
qRK0h8aq4kiM7m+gv/+wN+nP6Y1NsGlQLvNo1qI16psBLmAlZsKbC1Kqa2QPCqVY
tQ2ra+ID1Cv2RaomUUIDawPhY585toan08sY2W6hozFmMlaguKEnGfKAs0HZfAhB
ruV3bvqZ33n+nmFjfDLtD0ezNfYmCMF1uEW7X74OTUDJGAMpOV2M0CC0V6+efUlp
Lx4/MmRLbB6RQkYsuzzoHQM5phUEx1aeP2mM9g5wjHhIGFZPgHjQA7xaySLPoQk4
xo5OLXCvw8o1oPb9KSo0iX0Kb1bw3dT5LUsN69Jo2TVJizmlBMa0VVALgacvlVR8
lDSn+7uCUmlAkPTYEHSaaeFwAcSkqN4J6Kn1nYcC+AOhWLM+XSmln9KWy5CRdnlW
hM5jxZog2u3zqFt/Dv9/QBsrEwdGBTPM14OoMTx5fLMJFJQ9Uq8Leh3U3R77/zYq
EfuRxPQx13g73B1RJwISZkloGxgaPoqOSIfqC3+MIfTVMgWHiIxiqV8FswzrdY2V
ZWzlXNPi3r92S+oU4sexHo8T/KNdxk4OJEHc4jwWrLjgyd54RskEKvnURlfFnt4c
Th/FuXrzqqo0G0X2ZWJ169itJzeuswvNVoqeUlf7Dyd6qhIOCQmj46c1/62mKZm3
BDquLWTfAF88EtAyMJO2mQFXbP5pf4D9brc1hlA4t3O5RK3YQK3Lf7iIxdJgD83w
gPQf6K7knD7urAtXvl3igCcVyhJsRVe49bLqkyw6OEpMSAE/eafiXS33hAujAeGR
JgxQSm3Lg20SFtUfd/DnEN1blHCA+5/xPQGEv9W+gHcFTDvB86IYIhF4SDrHwUGt
5I6ACsxUgZm2rDHnjZx9ZqKB7IHR3q5zEFTIePZG2Fid0xZlPFc0diAQ05iJ3iQX
lCW+aez1Y/w+I23ffDExm6c4Ofi2ku8lNXydKeqnBsm5m8OxK1UviCDfQvHY4nBU
T/voPC7aARf41wDXA4ANAyR1BGCFNduRSAksbJz2TibGSPw6LFbCWDOQ4YFnklJ8
AM+xaOQmHvJQ9V4/efCeJmdWjcMHxSCO6YE1PrrePjl3Huv0pryMtdhd5NtVJall
W2mG53AmUEMCJ1d4h9l6V3ubNACG0C1M3Jz6UMwR4+VHwCbYdCli6GEAZm/bCdN3
C13TCnaGfS8pI8prf8tg14CH5xPTzPgSZ7Mq62Hby4EyiNYf5oPC6nlr/VTM3Xic
KEnsxz2o7ArKqiH/nvQc4DRc7JOJEJ++H8vdw9OpqU+XeyfLDCQXD5KhyMW675Be
Pmr2qUNq5hh783TNrjlfRW7ys4hju1gsDJK2JEN6UpSJBUkt9wO6eNtz0dDsrJfd
Vk305bTD9YSBS4bwzurAcQIh672cJBZefVBQumwtESXYV5LGIoF1ga57Ng6/rIpa
p9gmxXKN3MmR+xYqLeNrdspYLL2IFDzRHMDVMiByvOW8U/eZZylWvgGkuuezf5ks
HC3rwA5LUmKkriY5KEpcWAqEmfNI1hfG4+dxiUNDOtE+5QHcdJ4Rpdq3mY21qMud
fcbW5RraUFXvZRbj0We23WhMb1qmfVkJR7PYLoz7XbQK14aOpCuiOBlKM11IDqYF
T8NfiZHd3PcE8i2P1GzvCRJADUuY7OpZot+h9SmrmqY306WDcAij7aqoKd/pT/bg
waErJKLVt3k9XrIg4Z8Bf4MD0UShp1Uh30udWlh8YMT24XwnfpBiC3lugnHJ3Ggo
vbZFpu+sq9iv1x31LoRlQ+mi51KwqqW4jQ1AL0hc9bKE8h5NiAu/r3/fwxoNIKJc
Uw8OIqAtNTnSFOl5CVSo9xNoxC5Hdt4+Cxcbrk+h1P+1h36mN8hg3FD7WmCzIOrR
8g4qiMMI2z24sLMVuRWKM2Wp2WdQc3mEDPeHn5+OfTR8p0pHfWtbaeTUST2e4qdu
ZDckuUYsqwa9gWABIWYnuUZ77rE2Y0AnuGXUfpftzTPBG483jYtzDVzX6FshmRkd
/5PpVaje5Y6fDe/3TvEZKLjuSZzcJo4BpMOqxU1fuul/k8TLDwcOC8frYae1ikje
JrfZclbKSobQYdY/Is1x74Exd+KlgHS+mk7cINxKGjlLm5uUeYDFWHq6EZz4eGj4
oG3Mgv06vIfC3fWcas7/lkPBAkGkMACcfo+NgYYzwRBwjtYaT3yDb9d74/ReopDi
iya+ri1FklpiUPGNozXpZxSzMJuK/Y0JQypt6YBKFE8iUjcDtb2+c5COWkJuNn0z
73fsBSrUtpy49ylvY/UP2xczvwLBKpam/lwHGkM1jMxfZXaNsduuHD9XFvPXsW30
PQWNV8PeK9zmjhBWmanSbruvBewq3pvzg8PnUrRiGHWrLRh5dvLHDNS6anecLbx+
4xcZxi6bkXduXLoA8CTf3PRtTnlqdafRUZAFBbCdEtKIroeA/jwnwQxvmEOdKnrQ
WEYEP0kX3B0152Hh5BmwfUbXBChdn5RLB4/V/SJKgNZ9TbSOGuV3KssI2dRnp2mF
/HA5LiIRNu6w9CrpZdLcwh22b5suwERNuVuCt3a1HgLYltt5rKpggcQLxtoADuKW
6ydFnG7ZGnpy60uEfG5D1wQamNgMkuUTZRm+Ymts8QEVzle4QMlK12zU4GUIm99r
rykYAUiZzwdwL+fpghJZP0fOPt4zdpA1NMKog36kEkXsgkZuRlo44Y0jTvhqQSPK
TioKLjPPQ2wpuDu6Da7+/aVcrZ2ZX3XeEDuJu4iXL78F+sXdqVDGDI2Llu6b8NQU
IDU090s8sWhTuzz7UBge4HE+2s36+wUbjN1CDV7O4oA7eEQu1zYFfVhfy2r8sOgg
kr+1XIx0tuqwpV22i5zwih3SqoU4HEjUilYoZWXMvoOZlp94yJddTW6nJeZ/N1Y1
+68KeHzvHmRkD+lZb3opKiOcjFtJk8o98KoMMLo8vqflYmp1VsPnpN6GwiDo8JSe
Mbj8zD6PX1XrD592DIllqxzMBgJHjQDsGddBEUGnkEINSvMRw1DGzw76kIFMrbkH
QYTxufxlXtTd17vw2ywNHj+n7B8cu/JoClsxabTRTZBwRJ2T6OLA6p1D+py8wOXj
60uokDC9KeuLUhaRkha6BZFi+uMraIHSEcM/K/pE+eJB4d28+dmRnCBng2bTE7GQ
PK+4GY6QJKFCUGcv50mnU1ieAa//Cptkjb72mo+Zee1DAd1WEwZRnrnheNbzC1z7
4SqGd0y4Z17rrIw7C5Oc0Srd4uVa6A6DThdj8qkVZv5As01SLPTFVGrSKrUOYZSm
OAGep3l36qmWOEc8dnwqeRnPqqptqXsTewknt49+HWiN3zYETAQhwI4SFPmfgmqG
RkgpYOc8v9u+NpqrLraoxaJ8lzKyt5ESqzAq/Kg9F2aaU6nPltEDLfg0lqRkVjcz
IWOF5FwUxwNvMTB1mWRVZzrMZvZdzhEA2Y+Xy21f5FPZKctTkFWwFPowBwYB+uvI
ymu4gvIQoHDNflDjzeABb0qTDIpaaQXVFTk0HBYgcyYaVaEFE0ecHnfjFVtpm0Vz
RTPLN1bv6N7P0Pu6Gd88ksT+dujQoFjGyCpQs8fdG4yq4TpXeLDaxiOHvA8Am+34
LqU9ElUlo8HkBQbx7wICtb/wP3dGUeRwpZOJTOjkxBPRx0fyXPfkBgYa13b91+IX
cJtcD+xOfDXD9VxZ0MJ+MeiKVGt/g3WVMrUDuhhpntGqkhhX3Jo6X8F9Z3ZYGrkI
eGtTpSXecp2zCwNUk4jQCK/Ga3nju5E5rB/KbuRaI8JI0HyTAOITGudbwRUKqg7K
q8dNyA6Xa/5d1owT7+IDita6HzOvLM35qQxrhLgQhSjz2yFHEiorgVpXMzzrak04
wB0QqgS0k1zz1moAYRcqZatl/3IC4epqXweejWuWW1ZWbix2y9QVGh2asAfwCg2u
W8nDCnm3UgSdDGvgQAzK5jS2qOhQlvzD1UOG41VOAe4/LiCV78JyVE7At9V7TZUP
5+MDbbadlV6/FEpR9sRyoTuv2llBfJkwGAnRSzf/U1DF2sEN4YFnMAOgai1EunT5
C61Wxkvhy3pOBib7KztVD2A491rKhgmcIoHU5d+mw0Sz9jF32cDeeOue4frYfwhy
eX5ZAV+wdJruVN66UnJDHGg43lh3BZowOMnidt6T1R8dsclYe0aWD4M7tcq4V3lu
zU2rmV3AxrHnmRygBNY0sgXz07k+hhqtM3YV+WUYrPJT/zSx7p5y6Z2GVbUGdCID
o9Nln+WmiWpfPNEy3b4QM6DjwIg7j82IP8d19qO8J70FuMIWV3JJPXnUv5Vj+m3j
OJwy/ACOgYNYkAIbcbtZEyWBpnAIOrwJn1pRILTuC4DInrfWh1a6EyZwHpZzJa1K
LWQuqpHDhlU59fpt0xPYjDECjUSlo5g071ttyhAaYd1yfa4l3q17tNQ4/dlYn/ZM
TqxKfYCDM4JoIfUaQvYLXINK5zivCnjKVbfkWo+sgt7B20G8tIx0oGjX/r/2s842
+1r1XUUACoRuoGn+OQL1DfIY6zmHQYg/Z7GId7FZCUUBrJXtpuOYm6WCbNtS1GbW
raw+N0HFMI/DM70L85KtO2ZOe+ERprxyOsbSARkdcYxWiv0840eAoIROIMT1+qIU
12lL4pfDGDjD88iLV2VgtF9u8IBNf+GzfGKSVk/72FSlA8pL22o3P4IKSh0hN/zK
KymnuGrbaFpm0992HtjISX64aVyBs5A1rsjd2ZLIXobI3EqsfEyPAbe/Jb0lYn6x
ccq0FFLH/iGXVGCAnMz7gw9Djp9VYcJZH6n4APgWUzyEAPMmgsg6FDVLAkindggr
RHjy9zRNgDAJR9JwmIIwIOvO6i2BIBwCY7z5npP+0+cnI4AmeT/oWwjN91UOpaln
HOuAvh9yfG/+ErNPcJyZnQdnxo6HsV65Db/fwn3h1TulOLacglS91KM+P2Pbg6I/
ch4kTl3jfE7qUSdbIrsiaqw+3Gnvs3Xd8ohDhV6bKhAS6HYy9eVoylZKwKlzBq2S
dNQoiwZWHTONQTdWUMHEYiDsLXTJcWGGIMmcqMqg5OS7PpHRot7/5A++oQx69tzl
THhRBloUoqqKFWxfMVS432ZJbuLmX8Uz1HBwhzOUY9Y+qKJVIkWLydjwiGoOR2uG
v28HBRcihFga8zUGyQcA2O3DehJEm3P9pjsfod8rnbVLzPTCrImVKc9JFg25HI4I
8TDk4QHjVuU+CZZoxeR11wD/AFE3xoBaA1yUfhoI4ew6I2p43d4ZuvQXvPMX8uqY
LOx8rVqCQD4I7oRFMPi25FTdU9TJ1rH0Da414SF+Js5eXvUqo9vQvAFgIpiukJfm
1hniMYwmUT9mMLflMGbueTZfKw2TDuP1jM3Ahl6YkYtQfVePZU101aIVJB+obUen
mThhs1i+ekNl+/B9q88K9N7QiMCSpkPQTVsn2odz9OM+iGanxubUne1lrMP7uVuP
4Sh2uzMYXa+yM98PeIM/jeEqXJkpzlOtIxXXDnURHoRaoxqjN3HZXJSisKQa3hh9
MMVtcnt/ucSsJ4RNGIIPxVM4ZJnIdmQWAHV9LqFSo/PldOUsGacW54begGiv/UFX
2S3rOhQU/Z0i3Dlj2hN2n3EtRePvGpQCOuc/geNtXu9EZaPaBqZuH/StrF1vIPwO
TEDoFHstxBZKhm5kISdzRaB3yUhuO/2DF6yi0pqljLw4CxgbuuA3AE8oFd2wUWkf
bGqmmzmzX70caNtNhmxb/OiY5eCeaFUpjGnyVHMFioRy/4zPLJrBtVmZcN6uxX3B
BIrejxErDAIQTmu7D5K4u1sJ+wCyHRQ4m+PHB8hBPAc1+IFFfn77JMkRLCu0lbOW
I1+Yc4f5Bl4iwhgeotJTw8ONYT5eZyIpppDKOEpNzdAxH5bnOZqzu0QK/wWaQRRV
8DLtxKgZP/J+4VzQ7AfaRyifFPd7FSHAmxRD9SY6N91NV6XkG29brpUc7BXdIfDb
Jyxs7by58Mwq2WX83IU0wFej3xsac8xFt8wa/WQwtQcveXN763ulyGeoer7o5Xu7
awySMZtH9yWe+5xE0LGPuvDk5TtgNtM3j6INp0w5uO05J4Bwxape303iYB/VnxZq
qodurTkiFE9cIwuwuWYy/Q0XtCHMw/PcWlvJ3Z22+EHYy0+wIbDnueGQX9aIokWB
p+jsDwvlTyUku1THBGDw3J5RQaillW5wEsSi4yncvi6j+Hq+CfFnFmnXdfXWJJ1N
zfbAvQjmKmEu9q50GhKgXdBrFHV41qzCRk5rxCRpy8FVv9Nanda5/oJYeEWq0O1U
ByD1zaqbrAUp3Z4fwcyJzwT+tMyBrKRf/mOybRTWNGTNp04vOIxCOhcbA9zFK6Qz
byH8fV97UVrwytSIezZimHlZgbTEe6B39dSffyNEUEWGtDV3IcUJd48CQ3Us2LgH
Uz1xa919BBf3FVfWlIs0gHpEbySD96X6n+CH6fOmcbBHYi9k8QwszTtzxj7DXD26
gwKt/mi2/UxEqx/dpkAWA/cjGBSrHNCaRu69lLP7kCI2wXhSDXCGQJYNnfVOQ/ua
zSh+RvOnCu0wn2jk7bQy0OmH088zDQtfBH7tk170MRPRmktsXRyaf/Ny4xEnz7kC
LkPDZFdFIwUMpEijpa6Leo77JTiLuy1yIjwj8qJS1VUeT99SolbrUnc2YeNhDfGV
on/80CNSQqo7tM4xMmFdTe78ANQLOfrqI4prC5fIfI+yhpqD+HWAGQ8z+bviiXuJ
Pb1ZGG0mhaWJXQ6e6wdPaR1e9NG8AU/2EOSPFnJ6zmRidMHys8eGmasWvw6FS/g0
yKOfYEPIo7ck1fyo7emSEpwcyd69OOsRph52Sj0vr/tgQkNTazpCgLEiFNBG1v4B
WbAY7H5Qyoohl5pUd1ir2iLOBnl7uYtKC+zYUuUqvPv53l0x0C2SQmcDploRQnet
qZu9jcrNRaxwlphLuqr5zl7/ofj3TNFWH+q2LBJxXDryZqo8SZFLTyez7eKX7ozA
G+ZRdgWvxbiOd3UGp4yjK/y0NW80oDn+xEkNGJfKL/p+TaXFNIuPnI2CoNcOBn0S
LojGMmkwvXmGINk1bdS6WVfbHAW97cjIQSxc9sSxYxdyvTN+Tze61DfqM5RxUHT5
pJ/Nwm8lzbK5MSAFiSFAru2Gg4IlXFbmdIDKS6atpCH+Za4Cq8AqLZnl2LsoP29l
OAVoLSZr3VBWpXRx+6wJiR3Krtzr6eP6zDg6epdURu2Y9FwIkG9JeJ9tRovYmuhb
OD2BDP2oI5ubk9HDvvUFhU2m7Zj0oqHWxZS2yJOQCJmeE2YA3neBelMLcQqG8XAk
D6oQOZA81GTlsfjOu4I3EyTmJYoIZ0LJqBWlHh3+hopZX/4Yyd361Z8JJKJJ/gYE
YzkXWCxmLIYj4atf41kJDbvD5MuG/jnoTJ2gKJlSRXdyVjYPAcYmm3QHEHZBj4ch
BKvSR6xuQpRLe1b2DciLNpSz6WyfJEtLeiBHE7GPdm7hehTUapJg8Uke4Y7Xd5pi
SXnix16hgz2DNnansAuRyJpTyQx+EOE5Nm9TQys2Oc74dCrSsVi4iH9HL7mxNk84
lArB05lzyQSJmbZpcaRayNM+hG/VCitYG8O2TYTFUoPeTF8DBe0YKRuC5auxmfzD
kV1FFerPSQhsz6EMzv315Bor0fz982IqvjuVs9mDQVarusgkHujH9MyNtwmk/ylb
ukSipZOSphxnkNHllr1Z0MJYDh8PC2LGye2mXnarjlqWYnQ9zDqEz82sv7OPSVqu
GT8hp+qCHo0R7EqYbVDWG+16GzBmsyiadJpqLtksulYAWizHuSek1u1/7HsSOTqz
YpRnT9kUjaapWxzuW60yh4PCm2/jxpGbMRf0jS9va7kU8HrSLYwKCNpQZ+ZPcsFr
SzMNYeMPAQfedLnsVQ1l9So3cd+WRU8eg96su1ZrHgILF5jx2ZKrgeiAV+fTQSfl
Rda5NQL8mreZJNxrvi3h3X0xFR3y5tpQiOurSyaspyN/FvaGFdGk76nJKvMe8LVu
MnovaBUT4Z1fhqX4y8w2pNwCTRcoAh6JgBhWDt9mnQ9JEM+uoFNiGT7HwmYF9KB5
pCCM9uQpH8+IK4Sl2ezyqPK1VXIc2jI8ZKrx9wdQrDXU33Hb0zNszgGZNSrMR9YU
EqUDUB/i4RYKage2zYlkMUMOLmKnMfDFkB+IQeh0w9c7k+Mi7TC2Qx2jiT9GRfrT
+o4oqEYM1QHFeTdW+muxR+e0nCpp9gTtHhfNbumqdmA4Y6pekGk7kH9s8T/FPI4R
Z5JViY+7un9LZG8ouEwQJ2CwZp6r6T6BhbDgG+PLIWwCdjnzTWbo76oJ3kEcmlES
AG23pcFVRbnSP1lrC2+iJ0L/j9S4E1r2j2nhHCOKTE2i4qFuw50P944Kg/gCGMeZ
06eXaH2cPXIk/VU7KXp4TOE1106OgfUdKZ8w/LjWxK6YSB8l39lkzjizswghEOLl
5NYUjrTTwJvGUix++pAQ84ZrsFPvJ5cOb6AA/tqiZgUyJukdCsvV/1pmjmi6PLKq
pX4weNJqEtIVYf5ofKJR/mf6XqZ99Gk9mlScHzIBmUY0GovZU4Ayku5BN6P+20Rw
x76ERF/dTF88wObVUSfQ8H+YuUuBbS9neBryfI2WpqoWv6cuLQcjgafQ8aTxcYVx
hXSYq8+X/KCURB4yZcSQ/4LX/muiJ/oPRC5P25xVGxk3ba49O+/AK1vQbeD6BKQe
ST1SNibT09LHjmrF8AF+Pd/X1UYrsWURMj00rCoiZLkAgIzRK/dnCT0fW2zdxNeX
inePtwTGsod4L5Ya8uiNaowCTgwy8MK+0Jv1UU4fvPpIXU/uTil+EG/ijdyAQev2
29S7/uHJC3ZDjuBiXHJKhdSrcZPPmJrGTHX/A5Cv1wCaI8K7hq5OjaJNfHAOQOPs
YjUjtbjfx3Y8Ks/RPuknXsUVVeTdSvmtERFyfMPaz2HFuBjcBINtmlfdYFa1NKpx
gB9l85iuLndywj+T6wrf12oe44+iAwVOwh+rY1u/7Gti0horK1fANSgQ/Un0KVeP
7vs9i81LbmI5HHiBMxk3tEhTe3Gn4X9/wnf/JCPBixkRR7YJ3G3tk28nsuEum88a
lUGw0vuPXMUC2RjaDLrFMDw0OvIhPx/cWFH6Hg2jm65+pwce/kpeylkvCBJePN1C
MS8QoIic15PCiKSoOMmUpfceT2rGzQ9b0ZWE3J07FMnbY75bwSLwJ1mmhh3YYQrw
jyNkPRBomLbP9V52S5hzdo8E5ddU/ywPXnX7cBChHz5rO6vKnvhYgEzyeh8PVlQA
5dBzg/0CZf8gFnRvOP3MNAudHMeKtdK5iR+WK/MX1V2YV/AkuN5mwlWxN3sRIYVd
rA6ivsCvyvqw18FLMiPWfrPePVJuagaj+Fljojjh/IUsZsoYYMC4T3kjUAbBkSuC
ei8BgZS6PW4WKdTHoxOhNjj3FhdUHaAedqVw8DU7ppB1ieOKEvWdvAujcgo1tROv
CF5IjoiB4IMdOb7T8waaKUwprbbF8zSs0/ZJ0mKt19cXBqijct6ZvaQEUnH9Uf+v
5HzJOMtDjg3dZcaZ8+pnRIStLw2ql5VFpuHGo2Q4/Z482vfCcgptiHOEv/i5+qie
0hq/UgzFkP7KI8KBbhMviAptP3ELzF3mHmzs789w8dqYB6xhsJl3A6Yl+cew1l7c
LZ+l0dNGzSpbwgFrkVO6phmKUo4e7FAGoXIsRNNRu2EUBl6TaE91MWKPRlOqsUwJ
bI8tJ1/p5Gaz6pwjadBCNKe5eVJqgAproA6yp7N+aXm5/l9OXhTKxzsof3rqqqyf
yGs29WWaeMoHoeB7iEJqCBLIibulu5JP/3jh2J98PGgks7hhvf7T1yOlqlLkEt8a
bkU/8ZKvfthmV2lExwHB3qCQNhJmAOyhVa1EDmiE61CvgsMiWDufFumTAk7D4YF0
n/gRCb8A7+1WMrHiATMyt0Sl5YaYhBqmzr22OYsvLAlB0yRnKeisARJrwjOkl9uT
s6IdOHJ95BSDU9xOnOLu1fuG9TCFMfAYqoHYITWs1XUyPINOgisHYzVaWLLuyGZE
EILJqxNhl/+hboWXxJbe4Yd0VQmlJBsfwu9kiGFhRLquyeEGjD38awvP5fFlWn/p
PDZkQzcOP/xC6O5cgy6r5ZxBavTvzDiSB20vW0Agf/0PFJEmhtr7OKONhpfWR2E1
SzjNZ8GebxOzk26EQvq8vdyIdUClMHZAwrlZ1RM/35vPASwTqc3ciblECNq9EKfB
Wdw2KQU94sUDWwiZm5rxQEsSk05ntoQ2cz6IHkoN7jF8B/QQQkyKvUxkHmmGPeT9
+PFwVkeMSLwEKaSMVoz6gTUCx7JQxn3Iyd4ztf011zJzoHF5NBSnbkCaC7S8TR3x
KQ0qUzCuS1e17iEQrLZ7eGszGpE6WgsURldrY9xUGmqL8EXU7WUzF6L3je6rDrp2
PJ4nD+gtDHC3SyM5u5nD0cgBIzZwbIcZiB1Ene3I9FFFusdW8LWlXJa9JEcHNQvE
WsA6fTMAH/eLIXBAwRtBU9gKHWzQzvi5R0wFwmTFGrsC8Ki8C9L/HPTaeKIZqpSt
UgW5H5+dAn3fm5gvyP+n5ag7Dt1O0yv6qO84Pl4HVEQ5loBGHDQChxTEn2AB10u2
NjhnOI5IX1qVKQKrfay7fHB5Hb574ZPcrvsABuyx2mCwYHHq9mYrURT7dljF1yhl
GJuGCgIp0IQmU4xpJT937qXIG99kqJZphQ/51G6pxTLgwMNYtfZ/NNhzAVwnVLzl
`pragma protect end_protected
