// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:48 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Nbyg082J7QuAz+/isyScxk0eFtkc0RsTCitaJpgzxAdgSjDJ7Kpo4+TB0fNvYd1Z
mw8dKGF1/Xcicb1Qu+JVOtwUER4buWwBRiUOiMdd/z/rzyWnjYYcmK9kkRhteihD
58STiLUhP1G6D0jaSZojMbEDDXNQeR0CV6RxX2L0EJA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 131808)
+1itOKHRqf30UUNz0UM61ZuSIkorlsp6gkaY96jVOyEwPknsC+ZkOgFjDChEZmlR
LFTk0YeOTfiFyXp1FGhEgzDeyhMIUWL2XXkrl3ofYSvvOEAl5UCXtNaI0tx8fAP0
gbn7vAC4WQ+uM+O4+B8W8hVFFvqah3OzekzhtyEc41CKpce7MxBkh4jFI5Mx4Oyy
sAhv3VupI8Slgz6fbE9YojE2t5RICqQH+xHVSlPlVbPRmFpwfkQVYGzsRAQX3Qxw
JXlOnxddJR+qG4dSUwBzjb3ka0wfuTnoCFZXo8p8U7lOiaZzMCqGZNkyvvAffMmK
tk307uM43feTk21+3qLMVRK9Jl/a0NtLllWGf3CbODhtFoTtN9cEw1cjiY1/37W2
wEAlY+Rejx8zB867Cx9e1U2nHn7mLyZvBRUDjSJepRA0O4J2TAl200xEw/sScnxt
TXXV3EEAzAPUOhQd+hp6AHPOZeI8Mxd+zApu+mnsXcvHuAtEwkObRL7xj+Xex7H1
nSO4mR5v0e75THX8aLzhA8iWssUtnSGzEvG7nEMrc3OgapU1YX+R427YubFPA8Kr
kLQMLW40sO7azRnmuUH8GQpOxgKsz3rrs47XvNJ+8MO+dgacsHqkni5ZNpcmywqS
d2xRI/EQruRpxC0vqcbij5loxt/5nb7XDsnwsvXtM74vRRm44Hl+Zo5AAaHgxyhH
Vc9o/q6JIZ5o52Xap6tvvLAF2jMlyIxhWUntBV1XCqq6h5HlNcjjZda2sVin+inO
KQOlrMQOcBrqeJ0yDLFRD/AyyiTXk2QR7gM/8ncSQllbGMQukRtVkXHvHTi95jL1
VdV/QZKin6MyTeKpMZIQd5X1f97xpGOCVAK+L8fO+CyYqOWSaYnfjb69UZHVcUL9
NIUcqWbC87A3XF6qg6Vv0ZjdT58m29J6MV7HZiDPz6MC6VpoVm4a0nLcGb5s3gFH
wwA35UywA2jG5ziJY43if54F1c9AzuBSyMzUxbu3MfM+vlGGnw9DnaFo/fV0xgKt
6LgBat4MRcA/i+qs/C+hgADE2WX06kFUq+F+S6fLy0iQJYyUXAc5KE5WS1Gpg9mZ
5/NdFY83zxNl2PQP9zfLI/ZcRF0aiifPKMtK2eMwXf39NiclE93GLZfrf95zypA/
GfjFrYV41O62/IJCvmkT6IBGXhHIZWq7C3O6J1WfHN1tfuvFZip67d3oGGwjauBn
eAm23GIzVSZRy8p0nqZCFBzSrSlX36Fzi7exerA6stuYn63PMUib6o6LiNZDO6yx
EW5hSfv3cx/t7RRrpyishZotYqsLTx1LAeim+JnI1SEuFkrwgtseIbqGy0ZY0nCk
mY6OlbJcXEd5MH+/y12RoYw7zc15FfNzw7E01AI0HAYwDsGegMT/XwGvy3j6ny8x
3C//h21XyNjVQsEiZgMQcyjY/lTd3vc0s6hRHVP44hDjKK+N5GjSr92/5f4KF4cp
h6+6/vCpoZgXJHILNm2ziFBGMrsqR15liyc5FU+lPBFwRbLFDVMYzZXln0YC3jhi
2y+1OzsUtySmavb6L0OA0z+xb5tgpRhVdiF50o0L1fR4PinS7iVvM0ubcLHRnTeQ
QUDM7bh0BMVoXJwJ8yw0KtujfbD5tm2IrevUlArxknGLvEyjVAGnrpQb5qaPF13/
4bcmmI9AJOcNn1Da2rB+yE5C+NbhUApUjIyCOLMdrAd6KskDPwFNRD6TPGPADPQJ
C77Y5eoLLgJGhlMzQVfebZ/p+le4XADK+cZ/5nYU7n9cbXygTVX0yuEXvqpbKyWd
8PrsVpLewbWjt362gFWVHruEZ97BUZGktwyt6qXyha7fInVmEUl0oa5F46WfYZIr
axkWX/AlrbKPbqqMGQbD8LAA8FuMX6Vv4pfqwASWBAbcV6SZIQkSKgPm32xt7RR4
8NRR9yMK5oE/NaJhCO451xTPhoJ29KOGfKfOxbjCa6jfoI4QC2ZLlcUzi3ooK+Dh
yhhUxft/+fhdsGgqjAPtTgp/NrnAwKNXKTlW7QZdkPI66iPiKr1sL3LV/UgwcKZR
35wpzeiF2NSkuHBxwjn/EkBshfEfY6T26dxbxqxHN0G8LM0z+XcbVdbJZc2vtPRN
G2Sxe34p0xwwfZG8cpSeyPTvyn1xJO+9cYp6SIcJOinyOYGiqmCwsJp3vX2SzWrs
ceYrYBnY/cOMyYcr7gcYtdJhBJflqlK/OUrkrP7schXPS26XIBz6F9AgihdAarwV
nGb/iplum0SjV4DFei/qf7pijPogKMiC6B/B1tfOiKhJDxuRyjYUTIspsmu0jq+s
sYKhWq7JBMnRM/zB8GvlpuRtetEuvqJD0KkLLYN7Fr4iRRiInKq84f/6/qURKGhK
dlfDrBHzJ+O7vaqSwJrmkVRbDwFRw3nsNnEZ0HGnOLqI12+8ryLirViW9xGe1fRF
X6InErBNHH3xR7OsUTYI5e2LUxeqNEj9zx0VFcyus2jEyE3MYdCUK7H1ByCbrxUG
LxU4wFl8h2+WPSrh/tVSpQVfkHiyyZxVVB3dBDsX1SoTl4PxpLElMJz/3McT5QL7
qneGo8F+PyEitxDeycKme+YEV34vKQFM0fbG9hwP+Cjg5oSiSJN5lZyYFWuNUR79
zW5fFLTbHxaY9SxkYzdfRXbVX3cb7/8aRa+YDBwZduYyjlMH/f9Igsb7Wkyr+dGM
6CjWVVj8T5zXqN9o3RSbg1wtEx33G88/GFmxb+0LwIC0btmZdZRlZh+pbIZk4Vh4
0yrGwfkqtzOc8vJUYSIqrm/5VsC9sdyaiYznV/gX4gHmxTc7VyAN466VbwP1FWJt
FuyS4eCTsgc6fFdhh3d9k45wkPaTDaaUJpBwbMtyk2BRj+DDGA0bKnm9MvKauG4I
fhZqry7zbMiQ52TlfaLVKbV0M2hzjLPSazis/PqieEHPTYsnZ8OumoZrkbHIg49T
6p6t0vy3Cc8WjNH1CuVNuVuuwMzNTkEwqK+bdaQah92xNmemjdrtwFX7fTOo4jHm
v3TqHgqo42F73BND1hEkYxw9HgJJJUIZyFR9K8GjWuyUB6B6qaZJpeZd2Edfoix0
KCcz4bLB6Qo2OWrll8ak+P8La8kfHh2D+VOay5hUpZTELpzWHudX6oaUBwUaWBMM
wjTt2E7/dQExsZtJLJ5gky81Jrwy5lXjoB9KSvPK/qE9jEB0oWf2fa/k/Xw48q6h
YXgDYsdANAfz6o+imjzkmS6v1Ez3SHaS/tIrSTM/jIHascbvoyyWBl2Tkk9Pm8NU
CRwm43bH/9D3zraL8vvPg7zqhgc96rjPxecwnP7ICzSxT+3X7f85tCvckNzzK9Sm
1ilyrq++a1sdCf/0JjXmsfJrFhkAD7f5vO2wcwWtKNzDOR5PrMSdYnZmIXME8kTI
lgDyG+YwZzPlZ23OanDZaoOHCyIHqzg95CO725VYcD+Qop91vBGezmYe00lhBNwH
RO4NPyyZFlIUFJy4HISCBOrg1zPJZSdHa4CB4oPlHx573cBg+SVsI1Lca9Wsa5Mv
mln3fLYl0OGGmDfoOviKf5WrgtAKdNc37B2JnS8DB9YK0d6y7lj1+2zDV1g6Q03A
qYRMzjxcZiXRG9ZhMUm3wMGw7m04hfZSDB8i+fHofQKLQgpAxVBYK//9Y2ayT3Wo
sh7FLuqF5bvVmpINGSBiT9TxEM9WmS5p5GsogeKSZr/val8FVgiCyNhxa7a+7BDs
tG2Dk6Cwt6exZ2D1FACDWLa7XcD/Y3nN6Cv4Te3Gbpk5KbT0rEY32VCHziIfkbFl
+utuqrZZ8SQbyY+Y5S4Qh/xQyWIYWcRWZUXQGUXOL8K07OOk68ZbdtGhj5eoQGEB
2GMF22k2V7gw7E6st9qcv75yLiBsJWtVq9pB1GFm3SBl96V27AtDiVjUZE10NtMB
ScagDcTQtJAQgX/L1JBmY9kvESQh3+pUrYB27ZsBbZJu3Tvvi7NQagKz0KDsLThR
vcI7tbxpIFlzs4p0PtbNdI5qHKogX224TMggqkKkQ7DhqVW6UOd7JmmMhDrRkHGh
rzjl40cFZTZrbR+Dulj7d27bHmKg8zvYIp5ZOgDY965lwpuSFjV/59q5CmV2kTYL
JDE87/FxOAq/WFDI6nMMNMHO09Y3NtpsUAejlpJfFzUQnBetSk8Uvsy8uKPDcE5E
czwA+M/3SygiQyaAXOSm/+dv3eBXojV0/TZdjJ312aKVD7AjeQEqkZaKDzmQepGA
soWzfXET1ckRBKLkCv8dnSl/RyV/2Bvm2rGIzTq3Hur8Gf0/Sdg8v4HzhOgQfJo3
VsGHYcmXKxEf12M3lXnQkzrhuClxa5XLEYMU/I1yo3OPG3u51DxrXasvbXyxUjfO
RzUh1/3lD7dJhzkhKR1gSt+ySWmb9pRQiG+9CJuQeQ5sctT83g6ECQLM3qWViFIU
GeWCC57vDNZfol0MaOs74PF7O0OvxxmjH4TrjvwuECYsQ3Qz4vuVtlrqU4wgf7GA
Ay87fIWhi7oXslBWEMMiGGiGCbzzZ/xZrabju2v2owLWMMUJUaOh7yc+7WpC6EIc
wAbWKj+QWwOkhaRZWKaFtlxvFneJoJHJoc15t9QOe17Gm9CWf98wNeKu5xqFEpe9
YmcCoEa3zchUZbKYmS002/MzWDKlrSchNN4wvQvVnVv80w/J5C1VJJaMGh9UEioh
V3yrCDs5K/TMFNPNUHnfShajPkwg2lTwo4frrHTfOEJFYdptWBey5QT6wWhYXnb2
uTW1sSwwOcGddFfpB0fo4CX+swKQ9y/aVtcLVoMfS7NMnVdDim/G+0O4037huMtX
2f66felycUuMozi4Y5NaIwcH/5TK39rjfKdMiTnjszL7MyXGAhkyVzblz3/N35Om
HsmTu+PhMIZN3R9AcdPehdQi69HcUvrJu7+D3jiqP/ok0dIh/gJYIG9aiMkGKXib
EG6ucdzZq898dvcs87H6SDGwkDtqIT1qE7kgbLfQK/ghIugR5VCXnPEH65Ugng+7
HGkoSj5ieBYfta8PXVACG/EsXF/m8h40w7m+wi8qhOI2he0wsdXFvPg0H/KGF95c
KkTJsZJXlbSoURp8wkujQ+7+wv/tdVvjKcigzkouW5Af3OfewcLtz8Q2plV9/D+/
JNA6i1hmsToWhfr1x48d5JPGHdWXw0N45pzUsrc3B/SbSQE71rLn3x+R0F4Gh3fX
oSgidhA256bNQvSlJE1l0U/TixFy8hHvZUpjrR1BjE0SAS0jvYiN29+dgNS69R4E
iW+dThrFD/LAdaJtV8P7rXVfT4lfz1W3lMpnC0pjTdD/bM6FMlswUKBxwyc6XJ4Y
YzjG4/miRVvlDVnNnBz9YVtP0Vk+t4P2LdrpRV25BINaO8/Q9CEHGQtxdDysBOWO
m5qpZf7fWa4GwfI0HsZoJ0yegSf97XgKppD1xjf7xVbv78810nKGeFBhgC07JBM+
lPgnoXP+TAnMFSOh2g+6YM1OfAFx/5oUVqIEpAsCoYPA4xiBUDqBSZGLyISQ7PUy
0pNh+1YA3JjMTvUMvlgccz4mlPT7uRNax2hw/FH3s3icU8LLLeuiuhOg47MS2KRL
mWL8dzQT7KH6lT6yJBW2SyMk1z+P37NyTVcKc0ZC3c3Z98gUZWcrDWn/fRmL7wZS
vsa2AP6yzAr/lZBUFH0Pl3HrltQOiZv0EiaEpd4nVgEnaV5akxZOtCEhIgmeYz5w
OcQAsn/1FeTbN4cefhXrMv3De5dHkKu28wRMtSKlE0MLV3rT9ZQD5MZBe5aqgVeD
dtaloBOTLK/YfuriXGlrmuw/7CiaOEahRMwYFP8TCOxrsVT3m/8z+IDYEo0Jpyho
cjtIsdhpKZ+ykcfB8BCO7ZU1zwiIvph6FM4hVIje5si/is2a/xxDXCHjUfp6Wa+W
a0vwoZKovyllB/uG6I8n592qrhrXx5inmPyDxt7abp2tFc8IrLXEj5xiloaFbMu/
htSLiQaaxOS+9V/kASJWuXLM2Afexn4N6JpSqJ5isPi6r4HWrKGLHQtyKdQyQqCy
SCBUAolP2emkWpQbkesGU6XwxuYJ/sISGszhMpD/Fw33LeuqQ/Ei19bAi01HPYBh
Mg+YuuqsxV7D64qMWWUsDlmvXXb407tJNFApYmVhdePuyup7Iz5pbcQCltgjbuMa
DlEiQaLlK2ipR9xZUt4cYJLGLDo4a+Wgm4gezW5Lqeoe8ErgWKnBgG3yah11vXnb
INfr7QG/pgJ84I/lqUoycH3nzDTtMQraX1ha3+KQQQ7PLmWztBHZaSE+VA04zG5C
5D9TyHCKkm9AXhlgh9Cty+0e950BvrHy5yqHzMztfIoCTA0aH09xNi03uL6EdWh3
aEakSjEDY0JtGXPgXYLGeNKRnOtwUZUTLwxPrRVNqR4ZOy/BITHknTMSVnr59vpb
5IuIldJi0uaxBi3+D1NUAYKmPHIFjSNeXQI+vQ9tEFmQISQtiHx8RZSOTZx8WqO7
rsLQeM6vI+4fsArH8rSy8gaMszq2gUMj/psvH3QjMet1BpS6Zn66eAf1cWngv+mD
tuCjVHtdTgpbyzplTOeaJ8fpesR3mJMUzUKO8yPyWRX5ZAAudDYxj7qxUp7yK3yE
9k11hDx5qV3dYSUENekIe7IXYCHHTUybjY8F+xHq3VPUIuRzbY/xf2v+OmB/N8la
zYKeg+r3yjk2Rx0ZOKccF+SrO4hibqYSND6IwxZFZYClVAFuy/azcUJhDzg4DS70
Jv7DFGcoEdc/dhNrQDvHl7D7oHjUl5z5OMEpMAId8IIy83WEz6GoBaUvMkyb+hN+
Z7Xh9JCOpH9mYTf6mg7lhC37PqcfQ+jX0hU2F4bsCWn8OEFkgNADe45oqc/dyxtk
ujGkW93VXoDhEof57KjhomxG3SKUydlXaahAuTIhGGj4oyQW39Ms6UUJtdNC6y6J
EV/Q3aYXpkAmzkoaXj0mM4IoV6ZpU3O/uaqfxDTe8UsQ3vuu7E3vQQvCFZ/wtBXm
SNx83o/K6SSVhXoyggFBQZfXyGrxpV9Epq+LV/p7+eZYQKSr0bRbst3CDKPnvn70
id520tqQremekF9Nl1LEQMjsbJmk2g9yqg7zhliABZc7DmmsDQMIr2kdfxembtZQ
VGqQr3jU1JoI7ab5nn3NmFkLLmM0nLkSXrZYAAwIbjo4FGVAE4eVZo4cyqYh9Aw5
7XabDlLNGBRE2gOcFZ+krkIaFjirqwGMRPwuA5pKWCLL1V+Lp/Iq6HmjIt0wBE8y
G1XjVFO1T5Jw0t9VyzZGlOsJEVsCQc3x0HHzQVqW4lbU7+nuwxKhvTBG366mvHft
ggAUFyh4Mka5ccKOhBh63hJVv7zhuzQQMeSTqIepkAeUm3+b7uIuGpchxPNUM7Oh
3ChAXVC/lxCk+BUa8CWHVKmp4KmFTeT5mAO8DHr8x55zXn1cDwJXGhgQ2LEmdZM2
31O5gOyTWpFibElkf7yWx9CgsjqgamBidHFIFRRq4Lpqz/TxS97fdnaqkmkfdKiu
tVtcuJ209PuWpydQ5WJ/pMRTGDLU9shyw9osnDq9DLeN0dtCcpMGWtUYo3PpOHd7
PoAOjxMDDTMn13hPUjmBu0K9fgiOWzYhcmbJmP0yvXx3McGlbtKOoc5oiCwjD3g+
Gu3WQHVqNUVFBVtrNvQw58YVZwkVFFPW0mVDeP0dwMwORWjul2O3/4Aa5y1FhxLj
5XHDugDqTuycFRH47BDo3fsOJFgGJ2u6LLa0iHJAgdGPja47cOD9igWelOgnumVf
i2vXXoDBNFxUZhw5EECYNVkB8LWDZHlgdmOl90dow4pxO6IucpQ5VVvkCCl6e4Mm
E7omhPY8O0pZApR1aW3fn4b7BwCyM4z1xUjF9PtgHVgAlsCwz5HN81017S8s4lv+
RlmgaxN0LCRrHi1jD2LRoAiAdIEkgkiqpxYTHI8m/zTfMVxhLhd0fBhDbDV/Wbxq
y9CK093H1y58aeaSYMuXHwLloz8Y585a5ZhobpPrsYsGL4dk7CHhaktpxsGl7eEs
6Y6hZYziQ7c70D7pSAZxDR4TOzHIaHhA3DpiZP9pg4Swsx5NGYjjUb8vnS7Yh8o1
zmEFG9MLE1yWpg+lVwRgx61YUo62tINVIIrYRfkuPNaQ48tLN18M3pVvtDNWD0iQ
36Rd2tNlVKoa3UkzvqyBP+ztB+qNwWiTVUUqm/MyjdS3etft057vaRTcwiB6OAgp
3jsUd9kF1+fDpvhM9V9eCjCm10EZzkShP/g7xCtBkT96Bg7vQUbAHgRYxBTL8sF+
4AH+OkWvKTKuMcD6CcK1ScYAeXbLDBGZ68ZBCCHGF8MDAT4SguE9xMaYtJe8g3gV
6jzRtndmy4i8pYYXFLP8NFOY8hGjulwgsXf+h6rV8u1gM9vuOHWbogdfGbEIa+tR
ncjZTKpQ/wlcjePpkI3c3El4G15l6KHVeg19I7H7xBjt6SPsO6tx0LFGSw+WCKJv
32db1Pvn+9jL5Gh1PdaLKQMEJ6T/epk+SzUi2/SAsqUDwNs7hssN0XZyIflr4KBj
PDf32xkcKcsFj33f2ZYVQeKT6DOKVtXo51CAQKoZwgYcQnvipITuNMZkYCFXQhqS
c20l7fZbNIuyMmsdxorbHu05QZTWz+bqwYxmexNdQwe7LKqrfElASoGgtf50pwZB
Vh9kiopStaH800UESmaKPal8epDUkwV93PNHVz9XIsZpM/hm+/uZmvOj902plDH9
rhrImyZ3ZEhnQliripUHtTstRKhFii4LAaE+75w1q86M2EN+mVyvgJkJG4y0ik7l
7h/XohRID+H5iBsmSY8AqKW+7sK4MS3pYudlZq0pFPYqU8ci8NB0eIBZQJyy1oOh
GnkoENsMyIhNk91fnmTkULxOQM9LOayoRi05HZuW/1nyJYrqvD7gMiXvq66TMa8p
tUT5wcKPn4KgdwEeb39wqbGD3Sb+RY2otDPEkv1dvRdfzYykTGuC2RdszvtGglDt
3XKLZJ/37yvAdXbtKz0+nFZ5H+pv4DhYANwOhyyRrpJsZCEQdplmDlTQ58DXe+Vk
wN3x2057DW3PpGlnGc2oSJXOhho3lWtxEObMMQcaJOA12/5WD9LcT9gFraEXZXyf
k9NCqPt/yTIHE04ZCIpBxdrq1c0FqBlQlBNH93SZGcMqKN6dfYcyMyIG1vqtVMl3
JO6+yx2uIdRjAjRTVdGhdJVARkLGFPvQ+foXTMlzTBF8e57vCtHTBYlY3xdEhQsi
UOPHo4yWeqlGVw3xnmKPCpEe638jZXwAPg8YS5vtJfgKm7bpTQyczZkAVVwCkXlc
9/qj75R6zXx6hkweK3DIkPrEmLgVE8me5UoDXstbMFauKUo6Cecmnk/pVW+dstNL
lbC6NeA8PyVzg7FQg9FMxGsG2ai4eeynWAkHH3MPJEo74q0L0RywaN9Xne/thN+w
p7OBt/owLFr34a4bpRdiYTZ4wI6r5gI7cBZMfdvJej7us2E42hIm3Kojodjtw8Js
jwrHEW32ug/1jXzps4uZr5SqAwuHue6Vwp+w23J+04AuAxajx6gyy0+MaFgDG4xv
4bLqXwgx6i/FWW5nZNak5U/pU+FQqFzaB03TyjpIY5SkWa1WA9S4hTemAn9LMl7o
exO32yxpepS5+ISGu2UATJxtm+nnqtAldmWykmyQbbkC/jl+lM81xBBxOZhS9eEy
H2kOk99pjZXpG7fj/ibNjDlLgqxRPGU2E/gwrvEXCp5GlTE4J6/uxwAkau0HQPov
ljy+429GxBP3grpkKfXmEh/0rGrLkhXxHA0yfPz4KfZbZMx/3g0lCkyHaL/n69II
kg5aSpKVo+dS+9NDLk03U68V84deY7QSNAWEH3DSbR6L1mayO0I88C/B5DyNZnkH
sP8Jvkh8PXbueRizpRnEYWpJwxCWu+PmqLMq94duPINr9rf0TlbVFiVGXN/FBu8C
reXgf2ae4oI14m5Okm21frP+INCfDrRur3Sr9j8mR4zLuNtqgylSCAxz/BJRKAC3
O7VB7mSC1RJs120x/UW7vZHXb74nTrtySSRrDOsezdovHUvvDz4nkfD1WKjohqn1
C5VAagAz5KLgL/O5RhwTahj/OGd56XGaaCXeHFQd/EE+z1NVdFEBfWGV6qyVoSh+
zN5cTX3ZOUPvaNXroBRj8xzQpB6ny06mjxqqmpJIcUjs2JMHU/n0DP3A09XsK13f
Qw6pWmMk5jhO3NhZ7CNqg9xljPBfvkPZ5M1WrfLmupohrJ+v41dQDq32TG/CqZxk
zVxNl/RCR8VAjL4A8ssugx20K793gq4EZmy0BXV1P9AEdo4Fdd/GjjKHZeYDeL2L
CIW6kSHIdXlg/AJjgi7gv3AglWl6abZa/XtVT2taXLhE3yuMaB3hmeCPnTop0o1t
xpxIF6/2/UbaHn/YzVUifo+kONNM41R71jla4iXIt24eHJZ8MAX9tCg90VONF3YA
QJZEp6PO5n74A0wvU3xQLCJvviaseOi5bTIeEIdOfkc+TaA7CWmDprHrhfcibPxk
L3IuxWIc3J1LEc3Z1Z+Ruse2+uqJL03rlAhfCxmwtrveAMPB4Mp456q2GnxCrBt1
pwPHLb5RKQYGfwKV0Uz2hIEDDn0MhV0NyLAGg7WgBFjqJXNtpyJanuXmXlEDCgxB
PJpTHSLI+AjCdewPlLInEkN3UA98xgepZ+cp6OigB5i4LmjIzxVyJHlWAd1rIbSr
Jy0zyeMeCcz8YyrL9OEhtzDsJkgWxAWTHq5HqzG2Fn/YoQTDRwKEoToPX8kRkn72
nrU8cyt3Cy0GBnLqj1wmF+J7m08EfIFY2NUzTULnk6h6m0HZPhoPCt0rPA91M3Vz
NTg3ayr4M7/5vTjj+ub5b08whfPWPorc8C7ozfxwIb0DHLZBt+9B5RciC68oZZIW
YhvoDChpuvfXWkGymkR2hRxZECap+FPf5EQz5+VNQPJIsPGcu+g4orvsGK3Pnjzw
iJYv4PwLcNW10S1Tkbo2VTYaz5opNfAuGyAkocGLsyB0FZlOmz8h29DlUD6/msm5
feWYlxhkoZRRNfZomprJaROhn63nc9FitfNLdsIQ8vWb4/wYvDg5S5XIUlw9RZBM
oQIqWVekvT5AoyKSXGAK+kV0lcpBHNGK/mCLkkPXzlxdf5a2xjeZXnPAKxaPna6k
7LDNlS/PwSdT+4F/hutSfOPhMCHHCOW5UR+dsbgy+0C0LSGEmcz2FlTAol64AVIZ
3jpNIBAKt06B+ks0BE5GqbgncPU7giqGX0YyWVPrhCuCqpBE2fmZBB0yOslQIJO5
FQzNDsE2dNQ9DtLF8OLW/o/IEDUg5ZIDhjT7J5AsDKASA3/Y5nCz2s7phB35UDc3
h85UO5rQd8TCfLLjALbUh/Uay2MZbnVOop+8MCnTAVa5TE/H8Y2Oza5kqBKOmLIy
x0j5oddTi1U0xL0tkjdsGQhfvuuBKIpMCEGuT6IYAdko3uf27kFcSf80Z8HfJLaC
yygts9FgV6WlQB5PWinQL9yRVNXBdXR/mR5VRr7cPXCptLGsgUOEpgYJvCz3khrz
xOv7fFCOhVLe/SJ7jqEpf/oCxVvaYWUaue6oy9yhXqoe+yz6vqpKmp7YkIx/Q89B
NAAX+D3QCAEHTK7i3Jzxo8y3yjOyXAR1JYivlhlgfiLpdQ/8jsvLduoo47NOmWiJ
duNNdK2WAJRrENxbPxjsPitR+jk+VS6ZhUjeTZHi1152hL1lHXafR9K3cKIYapdt
/+oRQbYhazx+oecn9xIG4JsVcl75oqKSyPygsfyLvxwi6kiqW7LYDQIc4h0WPYuj
LeT7mjG3l6KPQ+YtaoA2GXXbROqKzn69dtPPuL9Op/HxR2QYxCKCQNexXPAJnZdF
d0/TWpdo5URSDpG7DDzczMttLr+qf3PSHYDrcWBz5P1Xe7TmGGXiV4a7Vd2NqilW
4wgFPSuLtKI0DBoRX5GKUI2zPg3JeGsKp9AmlxsAhVRmmBwTeh7Jf2lusDk5Fkd+
A6p8pE4fWC28NocRXwZK6nJ3dExhFJWOgf56rRA94K94m9/IgcyhGrb6FJ2B8YN+
2E07kSJ7+KPE+nHKpXGGbImWp38LsqaIcsf3LsIjX+eez68U2UzCUlwHf/uJiSA3
Wb9JGZYZ3Pc8gNFbMpVarD+hDkj65PTtupsgSA5Exi7utlCnaIo1km4i/EsO5+hb
pMUQYc/de+N4hFPRyLFFkQ1Vk3M5J/v/qdIetta310BUB2yjt1durKkVQhqJE5yh
Otewp4+GuIz/HJ8vYUKQ61IoBbUNSnn81qSnOvQ9y/EHV16RPz6i3/bRkHihWS9R
BUVE2TV2uzuwSi/4XfZLNqFzmBZunBZNrllAidmcWLsCy8LMM5wqayEWU0XmMBD3
QcEyfVw2Kp5bu5XJQjgA2fYSq7ERlmcNW2YwFP3CImsjeobhsj+Tyhwaww3CsjX5
DoZPSW7cSIilytNDHbldHfMA0cvyxKWbkYXW/GgQj6pW+LxZ/SKL8wTkRgNoZIpa
VUrk9O+0q2deHB/TO9VZ8ELXm9aVnGFrLFRjrnth2EoPiTIJQY8GsygTlMwXON+b
KU8s+318CH/p/kHghn9p2un0VTBmaMc14ithauFfN6TmibIM5fLAYaeFP0EmKl5a
o2aMlYVQb1Dr6AkSDpPSpMj3rs7syo+vXZFy0qgGNYmT+5oA3gIMW4rPcpGqeGht
oq5NwnPvw8u6EeO/vhzkkkf20bNkmJG3Ak01AEvg/o8nFYfE9NHLfORc80HsISWF
oBYIILR8LLCBQSgGaJBqMVfbfFDAO/C4/oDeyvS1tEeV7EW9hh2P7uCAwjEVAJ0C
lJRQaKZb/3bT73l4riolJWsTOdB98/zyvTqh9OvdBLAO/RtL7Q83e36cr8FwOC/S
wzfxNQTI5yz0wBQOg1adFJNU3pIM8TJVkK5OXPSSPZbzzkcD9IXGwlcZdcqViVuO
6I9rqRMTn7IU9Wb9q0MwczRnKYUxO2mE/gwWK3iwmVJn54l5hcVj9lvJbo1QPOqN
3Pyi6P4pD0KlPQXGCzI02DaAyfgLjWX4q1BdJbeflRPSD/LHessEBV/MJ3G3tRFb
lcuTHfsGAY5MDMMaf2NIw3dZvuxOdrOSU1eCOIlFg9kyQS2wttoe+r0Pr/HywUaB
CygusNzLYfCjnIaKDS64ZxAzINVa3AUsWcPp81ZwIQJi0p+WNermaVAzeiIIVsPs
J3+pN+lldfFox/5N9Ka0litcejowhnwhReSiCE8eMEIyN14Nb6x2RT5mxL4OVAEK
Csx1F7i5ncVWtxj0DNEwcr4W2rS3pr0hOUTB+AoUlea82lotVAk4QV0bAl0rHzJA
LqUxORAE093zSkaVTYckFKm1T0wnffpPcWWCy0BrbDoAPn0e8IntuQqUE3yzLbaS
JjR4Bs+kMyCpoJM/aNDvfKgEKknylyfgreURsULQFN/Q9jXF7wrtxe5G+M2GUlbU
AfeoJvPep/HhE8MpJVbqVbKkOOmOA0yT+fn/ZowsepicsTlRVADvEmcGpQQAdRx0
gUjpugNTqxTZifXWIciRm3pHNLSx6tKhdscOcjGusNb31OV0ItfvjAF8OO3Etxpv
48XsmR8uymn6NT8PyigQiWWiLY+lZZgohMEE+ySWiYJ0VGwDfSLc5iucSVkq6Lpe
iWgFUMFS0uBSl1WWU8+EPRbB8i9f5pWbZFQH4HIcvt/3+2VAVeDye8aLSH0HTSS3
wrHUb9gGHjMl2cS1UaHl5Ev1u9mIxDO6zFaDM4lx5Z4rM7EliUkm5g34/0otoTkM
2CaAvzT5TF8yp+PoKtoEjNEqXmQWeTewEoTlhcoCHWUf2htXMdn6cL1NrsRjAevy
YJAlhfSZ8g5fHVQMPNgbOqeH1ul3P6+xDSjUShujIZSVc+8KEkcFAMzQSH1sVsLs
cPWGUsCA2k/o2xvJp8VQ2yrNGXkAzXDtlhtms6oTaQyDaZVmLq+wTsuDFMWhn5n1
f4nHtErFf/RXPy59LRWxsA0II+F2tyDUT7qvJ+bcssTyqY3rYWOyAIBRbNjmJsX5
0C+lw6N99VQjjuWVrOMwyiuRgcpBNfzqsUTgGkCP+rirUeujW5V1Xv+Ib28No6tY
N2B2rGLavmd5QGjOsdn+1wBnG48M8c8qhyHJEJvFF1B4nR7IB5ox1WE6dlmni2to
09wPAoP8Dzo2DkVP11LYHwQGNq73YkMzAaQn1HatUHpYOaSaA3txylfT8umbCyir
Dith9ISC5ZLOomzDUdzHI/u5qMREDSqvXZuB1/+hCUaeWq94qtieviJJPskGvZtR
a/F3mh9330MCy1Z6b2+4UVnEQeek6UvWRp7Op7hm+13ZM2CdhzFAAV54TNb3lRkp
ISaRRYPTR9Yn+3rkFnhgbySUUQY8F5xKFauxtEogloCT2FcsHicmEjZxEgmxessL
q2Nl8h8EhRXwZNiQEivey0m36xqCdYRKfpEu7jDPWr1jv2CQku0YEe+mJg9zgNGj
xvPBY7bf4vvlYmNMyi5+2W8ncfLcctWoAWOZe2b5DvEAKHArIQvnQef8YVSW8vHU
wvibCXv95mEQK20wkSLKbG+o06fRN2ySZXoTLGU7t+mhjgt2sxnax5LP07aaHG2N
6tpYI9Szmv6phfJac7fUESWS0c+S/+eKjMndq29M7XeIB0xXlq6yYnrPy05b63bb
KfqVFX0eq2z087az8Sm/IzHSqqwpry0VauJ64xnVaaglPk751RqwDCd96AGvRG/o
R+8YTjesY9X4pw/oDBmo59XL8Rfd4Z0gHYG+J8OVUtTmUH/O1nJzimLgcJTqWerV
WL+dbFk+GyA7E5QbMHOvi9vKS0QGfuW83Lt4k57l9XiGtxV0ckJbwxHeWv7pr0Sy
bw8+9H3q/WXvwtGr+Cv1PfIS3kVcpK7ix2a0SENH4lJVQLGkcMaHjP/400e59b2j
Unyp+Lf4FptwJhaIleLCCIpRbjGPPDjDRS0DW+NzB+FtfTTPj4/LCqoWry3fZdCD
T8CJ5UWV9gthbrg1wAtzTPIYWw1sEypAzpX0aMm7/dBuvVa8XJ92mTwFJL2u4QM0
UzaOHsZDKtXCWaeJRjCcuQET4AgO2mwaFln0xhvGeDK75b5CFSRL+JCNH+jiuSDA
AVBgkdE9QzxZ4rWBBY094g8BLKgAKypcDsp6KB3vSw/6rY78vSkw+DejWp8h/Tnq
BV0lMstqjPCXFCN3n6T77qvW+i3syg7DdDhz1GRmqszvPDl7b9mxRAefbw/Uup2C
YK4sTqKghna3igSDYSN5F2v3GuNQIn4C2crtpuH2SaOsaoxjgBpuvITNeauscvl4
CQGdPrvSxO9HOYtHPlYNcAxvAHieAVlB5fTDqFJ1yY0qaQj6zopXJdYc7vy9zmLm
3H+tvEWtW0oCRF3AKQ6hO3DJp1FBVbW8gmhsbx+U/aYaNShPrPcXnvXeWNaDqbJ+
0COb1kpSHK7dIkpKzLRmjPZRxPLvkRkS4SXZ19gC+YbPQDSrhUAXxtPCiSYwtVOv
cHV0Feyhmn6oZX4ysWj/OzLeE4jkzK5lbrWmyex/Rq8ZROoul9L71cDvjiqXWCsG
VuhkXK6UlaLoLgN/Sntp3wsfyt5pEIBuVoOvUzTtdJLsu6DM89W44bbsNr6kM5fs
5FxmRsfVVTzTR5QuuPyhkJs79jpEGxVaE2ZyZ3/BXpq7vTR0TKhAmx5Hc5Ijg7co
jnTjMnn5r7I4sTTP9rTw3kKzuhssnmU9edIbvkyDD/XAOQPf/Z7sKvZ1GT14U+Sd
p9SdkokOfa+K7ZSnt3hi6wMSZ54lwRoKzvXBxyEgtvhXqUMW/dXQBmWe+jnj0zcU
tevUy7OFk8r5iHXNlDXhNTg2rNmIy/Wp0nUc4pvWZaXEbPPzEWsBEx1C4R/0KcxP
dOmaAkbBhxgXh2xkYidNnAikqxs8NibXYBluTIa9diaCebV82CKwfczFFZi22cio
vUw08cEE1aiST/Ka7jzLAkDusjbLl3VoPgenUVlzOC85g8aIv92R/oToT4cfMjht
WDttbYmS+DA6IxGDQi8h07FAT4kOmHGClcQbBO1I9hTzY/7cf6li9euu6hZZZlNb
TASZmsn08V+kFSqZltjfrPVLCcdNi7gbh/w58JeHbw5t4ukVU6s66ODh5WLN8Dx7
j1MV2g4OwUtKGxjO/qRPxQq2U0geo+x/APup9L1aLg63P+/E2NsBhmwaN8lSj8Jn
8r72Mf3JmYQSo+9GugtkxYgemTKMBxPLna+dsYHqUBzr6USUPr8UXSIsnF35v6xY
F6Pwrg+59uX//iMZHWU1yxBKrFs7KDJtj35iuoEKFLDAzZTfDfs7h065jbgqYYTj
EK0DoOnNbuMJvzkfQOc9SN1kGwrUYWfI0inywEX10JN+dIsnrt/mFrPBJvOM2Ne2
caN7KVHspNCYgGPVM2LdR30rAihfw2sT/d0G/ME7hDXJBGE7qjCftBEjze/wbQwt
RcXPvD/oAuLp3GHZRl+QyK4vAWUWZCkxBZHEfRMbgYCYUMQiLWOrBCsivnbKpsK8
OgMug7dAPkaC/6ylW9hdmebA4CvfG3kVK4CegPpmIu2MYLAdC+fLzxfxBRXqALTo
hp954LM1dzHB/2+EbdToeY8BeRcqB7864/1VE5B6/loAj+LyrCIe4BqLd83R1vkj
pK/DVJ50JeKQzNkIm1jE+NFqz8yK5sBC7Mv9/p4uV6L6aiAyeVZQ2OJ1sePWNJvP
hnW9U/yeGzMmyW8Yk+lO0ab/KjQXF8gSD59Fw8hrL+SFgbshmwTJzJm8k0wyLu5P
elv0fZXKEZW2P0m/aN8wtcRw6S935b51WaLb4QicRnTt922wE3psKDlefifUCHLx
w1IH8a9UXUaQd5I1X7b3pfVDrGgFMVEJaWiSqeGeRTwVvRNMk5sari9Xg/7VsvFD
iEfn+u0jCCamPuEauiTlUl5txLUyuNRwI36zzjNNvjunnr/N0x1ULSoeh1FeGlBN
BVWnScWm6igWKWxACt86kE1CmCVIfsbgTFfk2zex6NZlMWDabKlZbrVu1LAJGrKX
EaF4PniYXcpw/xAI3XLAJHAeT4bdq5WaY44YOVegl58TxmzbvXSdBNS8oexE9Bmf
bamyxT897wr+cBZyWfqnrYpZUyooUyer3YBkLVJZcVsbmWpoiec4PjyiX1MXOMHa
x82RZ5UftiLPYvFiPynwwhNZhAZvxF+zNRc4FP5c++ZuXXY3k1WC7Tbb+UGb9ErD
Mpkdi0wo2VN5vLel+vb9MjKZv1Jj4EjVrBiGTaLGcf6BG8yYKffPnG/1xLi694y0
htRspd61mAKZRAkCfx+qxuGCQW+4e0S1XziRlb+rfGgvGQCth5h4GZ7n9VNWNJeP
QXP6/fhJi053GMAsock87CuAZ5vCnh4rartAyMvWxUteIxNdO/QJNuLVawXVMeii
pQa7KhL686F8z3z6b01yT7F6N+ohowJPeD+j0qgCaxUW2CosIs0d15TihbLqRE90
CvF3f2d6qHwerQYOanQ3TCgr/lTqHbRYN+/8YGyrRT+ngEuwQbRCDUsRuQ42RtrR
gWHCBkzNxOVMvsjlTV1CZkhVjapaQ7dm1c/OBTfAZkdY8EkXajAX0vEZFHbI4MMx
B1eRDwbumMU8uHLBbyaoR001MI8sbYYj7KSBFauu3Pk2dr1u3qmNvr15WqwqOAO4
IpWtvMipWiSsUPXLO6jvQN6lgMqyxy6dmOOFmKUo0KJywdKpBL7PgmQG5F6n7edX
M0BocU1RBZRZt+XoHGKpZcL6ym4L2ffcGZSOGC+/X1EYrYpuZteFd91AjHNul2o/
01KWU+UojHNMXlYSM54TOnl79ObfZEGxJ7vv72d5O3FAFMe/8LN4RGjBAFMV/qc2
3RWSc4AmJZPfNtsnlm9KYGnxFFP9T03YGTWL0DnGS/+69fEZ8+YGdAq+5zOW/Gh9
rv28gXbXs+sVjsYyEpZDPswPBXhtWYSKXFKWDu4rcIj2XFDu8iXXOtFE8hp7UnUu
BZk1EVBhJQf8hPZ/kYUHyB5WiuVyKaQBKc5VQbDRT9TZ6zmNrU9t4t1NoV2FcL6X
Peed00Ff8SsrD3eOzAtKq4LuX9pIx7L6wgQWtINAiLLC5oe7+hbHpgGelV7IxqCv
qvVJoggx/OKukM8nlj4rF4tUyHj8KDaZ2Pig+RALz28SnOGspwXbtcU08dbVIo/z
g176BcO0wU16iVsc4sLNCs3c+9mpjcu35eVaa0qktyVnHPlMbRnHJGz2F5kEJZPq
fn+9ypECKn2m36wuCs8kUyqX5/dsYUVS1Ce6PJ99wbMzDV6n8NcurDyghqlgibwK
to0XZrWNB93sVTFXMK+HzdJ4xwjEa1n9E2tsx5a/AluYtBYoFuaCyveNqUO8Kzz4
v/Gw/FW9fEWxQ9JmgcOIUwMO56LQuqCI/t7RirhC11VlZpu/13aUQhWFnKUXLi0p
0Ha5fkiSZdnr0KLHe/vwp6pi5Rkogd9WSzGG+QvTJLXh/0EbLB11RrnkTWqBUBll
aduKLuGLCplL7fWx4FRLMjQmwlnt3+/C99Nazy6NFfqiY7xAiuTazZ609yh9yRGi
5MTpbyhFvofPyVrrma8nsXrNIJLOM+Ku9DRiRECkRY6w4zngwOrzwbJyU/JLaV2R
xIS7LRGLJN4oHqeTtW8JLQ5GsZtprbyG4uZTWGq2DouI1x085vhp+1EgfOyZ6C+f
fcIvnCiNSaWc30fNcIVFJKWC9HJP1MuJn0toOxV4Nnd/ezQoy3OXD5GncQ+myOW6
Erdi6cpJN/CyahhPxnzaXfSswTnx5hM3gWLkiYKAoE1irxh6n339424KcW2LkcBs
GBw32IgdhgshZ8/g4LvIBif2vreNfOdbjlqv2F8l/xqNEtviHyvDQG0jPSKAZMJ0
JhsZASk3RFhI53eltu70/aZ4JVnYFDwkYWazmOA2+dJeyG5+LC/zA7JT5OwQpRMS
hpRzKw2HFksKTqXogrvR5VLOMiKCeEP6mHus/4/ANeoGf9OvyicS35LlFt4+exDE
9EGSU9SzcDZ6vl9nWwdqIgvBTzHAUL8l3cCmoaHWToI+pCh1deHTdbH5ugwtemgq
J6Hg8kDUNack/l5x8nS3hxWBP5fYtdorN4eZg5bu0n0yGBGn3VxLG/wi1I3CSjeb
f1ue/zdkJPeL8y6aC9gtLfq9hH1wMx5IlcW9UJxRbGXUPXTpmUWBQoOo5q86ddpk
smoWhMDPap7w/D4wEDnWjf07+ETGXm28+GMBAVFYTe9k3b5pNtpg9k4XmfeVUsOC
hWA/6cahe75HbKyRrF879z8OI/cq3PdvLgt24LmZri8EOuAo3cRdIf+cJ+f+0e8o
DYvaLAEPkwvH8wEPe8eQ0I1PgWSddrGTR/oE1OJ3ZoBsT/S0J6lGht/ixYn/ypgW
ax20NNPmnV63r9xXNBsdVbzc0ZbTC22EExu6L/rHjprSYqGvN27/reL/u2A8rLGp
EsoVxHBJOSlJewcXyQjfQKcuNmdULCAKsYvuuxHgC7ZCAmjrEUy0bALZVx4RlmR5
aXsFzb/kfFnLnTYGFAHKZkMHolypcUVCIWA+1c/KLfAiXLvWbzsTk1/43LAZ+YFl
by4nThouB9JgWgJvQFqdcPMDcnljgKWcr7iUuv1h1pCwEssTS5FJ4vzbzw/owwd/
p2eh0mQFgqpDR1BsdYdCcqZh0sZdYZ5Au5mwDCrmZM5W9y8PLXhbiguumeLaFCY/
RNGsiw9MwVu4yE9zHJ6jlbHA6VxNpJwEJtGFQa4mnctdjL9zoJxzEcN2unELvPQB
Q6pG2qsxm/LBmGurYL4owZjX2ADPVWzyntplz/wCDRQ+fibi9GImmPI05QjnsB1r
+V2mrz+sStNcbAzCKeJxzm7SwGMfGO1sys/46kwQbcMw9R35YBHfBVrMR17Fdrgk
Ytt84IyJLE2s1wHNXU2T6+fjnPOJ/XHJrkm5EYRHXhM6u4VKrbcgAtTzjuMAbk9q
pxXCb8fKQ9IbRBgMa01P7dcmV8stMfkXT9BODlF/19FsYgfsemAxSn3aTewU5K8r
PKHmprOurFxarqix4CmxyHxjHeenzsAm/Kv/b4CeQU6t9RNtaRnZ9rWL0OdcKmp2
s8CTDsg6TBcFDZCnoqV00Lld4M4Hxy5hDAwwntMAlXycQPvhLSpvDq87eHeY66DM
fpj7mKoGMdlLlzGjr1l/y/q1uEQC3U+1nyOX5zCggqGRzyip9Y6/sUp6/xPIzF90
sx6UBbDd/6Onh/3YFhLph8h1RsWhUGGD+ZD59HZ3MUFBZg80uX76a870a5urGgGt
jyZAZxOvbNMxqsMVTqnCHT4gVjd2/rKt04U84lOdyVdvMk7fB3m8MNlkhtXcIeIe
V1t/ZoH72aofM9jBezi/fhC4dIOwVzPEijOLdyyONb6VxFz0MkRJvsJ4Yo610hl1
eCa3Q1FQ0xyDFPD68pSYI6kUAEmGquvaO4uPcBbW41K3E4kRsFzWsYwd6lWhdNi+
fk3/RH0mueFeIxoSDc0F3k82Ro6zXm7Az1uh5y1E+x4NBeAaJ0rA+q+7N02RFuVD
F6zS4KdaCvRHkoXxLuE3R3P0x7djBHa4hOWQNJMvMDijsCfE9CakiR/A6j3Cu/rF
72ytRPFdjh6jCxb7vJwSR+bA9Ck4AqBY4+eqMCVPKbvDNV/VcCClKR9IhNAjgIkf
5mWVCfXrsKryjwXphbISwebOOOh1ysBrbfA8SCfESS4scLzVwbxr1u18fHiS1AZk
N2g8ot8J/aMW6RRfNvH3tFeBkpIxZwGO4Sj0+kk6x4TKbniPP5n58OrEEklPbMLx
ycQ0hRTPDdBhKlNWtpLlmznMc5dh0NCgRmYTcGJ8Dwoa0Pq8OmYzjOPcilI7uQV9
jamb9scx/Tmjg66y5wjvePp9n/2aqVROyYPjNnSrP3lJDFlAiXItWuJPxxEYwydJ
zoZGm9x+JjR4uqt+oJ2+ZKlH2BzdzDSi/pEr0ROjcQlzWsjnDN+mh57d3dIozsZc
uxcYw9Km+lm0tKoP3ojQFEeAvDROCgEiG/eOQC9wtv2mIfC3kkbznhdrpYfznWB7
lCYqG+AXCsjWYecLj+3apeLBwuyvl8jBwnl3/3byugeJqDwOndC+dvPVi4KewcKM
Nm1t88t1MvnuDqeUx7oLUUygZ+34U1X+T1A7r7ja9Vczldy9j1LQP43og7l2p1wp
+RDA87gFcVwmX1BLrTYNBsY3/HCtggUUnITPgSgHFyPEcXiqrgf/PQhM+oVTrUB4
GmT+/sljfUsA4NowKBn6xMlj9JXjw2qZ2CNT/YyRcvzWFi/o18U8iYjDGl3nNEkv
OcOWNTwrpjV+mZbSkIZg8rpIqdKW3qMNlZPd1OlI5qD/sYhs+4N/hIoSNAgstn+j
91eG81WjmzUUaiwd51s2fcfOJ1iQqL/FHTU68pC9iQgi+Fi4oY617rBEcaeyg4y3
Ivs0cYb/hgb9Pyw2aLMF3RXsw7mmb4U1t1pU2PbhrNPqX0a2g0nSE9qqc0BW9MK8
9UsRxgDxXN6BrR/s11R5wUzqqDIQGddPb1okBc7OAeg7taSx5BXX3mzobmwqRlt9
UsGcA6Wi1DAzJ/W0DAToNmMEjQtqtyLn4l+NJkGfjNIDSF+CvLZ0zbzNodxYoDmj
vvS5PSr0ovfd9rqMrnwPMi4x4KxHl73brqhFStVTJ9rKJE3sSeoc0KHSu1LNde9C
CBT1cQgeq/S2Z+ICuJd+PrQGUHKpiIlZTsjNGGqGkpu/vcYjfOm4r1/P1vUMqgOz
+M9GjCu6nX5Xlv4nvjVpYwj6cCqtoKM1UJOVu7vIb5DJFxappWaqrl++qoD6tzm+
+xd/Z9UIeIu8lBNQOK6IglHvqp79lE9sJ+CtqNXafa5fmqZnmi2oEk8td60YCn3g
fOT28yB0AIF5XtcjpDon3T1qbxsr1F/Q6QrKkIt9w+Qjyff3p8AK6Asdy9igYJiY
8H3682fCX41W0iTjtWKoze417ktqs0JahlwNe2jGrRY0HqCmifu/qOVpLorz7fSr
ozUDWycq0bO57owl4HIkdVF6DAauARmFlwb72kpvMHqntNIIN72vGH2se8AQ+I/N
6mxQTDc+PnWhfEDXC805J4eBcuaSrd25zU80oc+/Fgt0PItuOoClzoFUBObDG5Cx
H2yTvQT58sct0ld2QOUduO2Kjo98haPlcWsJadGvVpWXmHFHFZ3abGQ6iIQ11hyN
q+N+gP9IgVzT/GHw91YE+2+LDwgJrnZil866F6R8VJzu31w1FDgIKJjZ4KhQHXNN
jpEZTwbSW1RFwNdsiNHTpQvOibmuPHwYWj4vYlOiJlontgSULRVJ9Rsg2BcWOiQW
V5sbthZdiRtq0BIVonnTPoYBqj6pwOUAGZi3BPSjzU07RuJ5YeKLGX+zpEWdSLsR
clyA8belm7fhiYN48vz9LQ47oVS3UJe8JBiLLkyiu7ogEzsHOzzjF/LuQInDdxUL
IUT34SXaadKYNoZZcFXlBDJUKbYzBzG27I61rLK/WzlNdCRQgKwnMKBcy3iIP8bF
dCKKit6dOHah8n8uWduXHWXCWvUAdMQp4pWD8b5RJDQYZWcBroajN0j2OwdMJBHH
+TcXX8hTTCSc6Yiut2HM6YKfPvGB4xGTt/Mv+3wF9ccQvhDaU1t9zayTR4cZF7ot
eoNZ73d9FFSuy0F/vzrFoO8ojBmlLcrVl0nz6Qzevv0qPGb06YfiUBbvyImTe5Ow
5idi1Zixn93ecPd5OBtegWXO//WC9wSvOx2smfYKh4byTR36rzYgugoc8QSSYnLo
NIc5AUHn6vArM9SkypoDl0TenFKdXhkEk+/lMRgcEv4/jKbFx6KvFvkj3L2Ufhqg
IF0X6skdwcIeUNbxdQ8JlbGkdWJq2kCXpGgdkK/Wx1As46ug1HC2BFxPpgH+GN+a
Q2HSwHKSw8XXK3og0qmP+70FJVVIEd5T+vRFTH612W6NVKPqPkIp7pARrEm5RUrD
x5EU4reTOHgvvBtxKQTapq/ySi9Ce3h9L4VJYHtBgHYmdreZS49PLRlehvmI9kYH
9bqRZOvL1BR4JxX98dUuzoQ4P5szfter5MwquojaqfVHT+vgGnLovOmmGFKHkDxG
s0bGYgP58QYNfgGwr5Oil3vCmAgc5cO2MCTomLl+cKE20f8GoVlom/0JnK4Ny3Po
ejRgpWfD6/10ECfkrYE+zOC45H2xvOOPLS25bjj/iefFkst48TvTZDuVrhZmuZjb
5PwkdcobdyFYuD0azhFhKDSI5DsKYhycuROuV8X73LBVZxOu6Y4c15kfNr2dOuoS
025L7ys2TmjDLjN5N73Pn8WcTPJcC9MJPLiXmSkRVimhSAKQg7ekdYfztD0z+oO3
nILGiKHOYrMmBILdopFXZS9+S9hxX7+NJ/Ntgo55mm3KPvoKXu/QbTo7kX2x4jej
kZ5Phy+7AIkdWlBbjXQrqkvoUfV+uIPCb/WZY+nauDlYAGa0wd8l4iLWJnHZ8JHc
MKAM55OZIDEO9uUNhMnUVn3ZOqW9hyZZqwl3KjXuZW968+MTvaALEGcTTGRuApZQ
O40yLaH7wj/AT/OEu7taNJMKmKCirn/OIGAm7P+ZqDn5lTQvAMrUnw3352B21hED
TgXLm2TIpwmmodk2VD1YCUHlIQ/7Pav+rKcPeotugVXhcihVKLwdXqXw3s2OfVv6
6w4r2ecKifsXKWPzgvqTHZ3s5zybjPZo4gYQkK9jLkv0m29DF0cqVm1pXcmTzzpW
fNg/bk/AN37XZoc6zaSYP9IouupL9Atj20VjMj3iugmszhdMnT9BYZXhvJcQ5LEt
ObBgkgRDXZH80y3TleIn1lspNS0ez0VBJ2FZ8Z9jiUZ5lLYtYjzNGyKLrHPFbbNU
dYi0Nul0Wxk9TS+dIf+N4fCuS0Z07yNdWJ64vIrhf/yhIG3R4iqKsLNs46CpaGzA
BBetvrlab0/i2flyBmuseDa2YpP7r7uEqvAqOR5B/29P5qfe6LNvrV8uxzyEFyOs
EZLEkbAVWiSEWDYkoHJvlJGKbnk9qiRXbknxZP/or7pooaSvSMsh6IWVrqjP07aD
eVDAAaIyIL3m91+M3Ft4buWsw+wN1fIb3hSAQH2aFOjKXgWjrD00hVCIWd29fttu
FA3oHCO5J9iTC53fhvxGsKq5RCJDpH69eRDHCNSGsTwfFgjNznn0YfZfWCtNRlUe
zNccFDJ0tiFBh5egRDyu5LFoRyIoSyuLs/Gs/R/vYK/2piPtqvtp7hlvBlYRDFYv
K/kdtFUAz1/insFOxH/xr4YOGgE2SOvuPXVZO/i49cNF92nMq5zhgRBy98q+AVd+
lwlDRDWPuIrlbNYtwKpRnCTrNwdnt6+RIPMGOKvbEjZH6hpxdIr9llJqHkGoQZf2
n+Ktz0hL4Ge2Pv7APji1YRJ4Wyi3xFJpadaGpyVodS/7lt4wYbAmWDFK8HJFSq0y
Xs2KwEOm3ZgAPHJZVGEHxqlHbhQbSdK0dM5BrAi+VsBw1MCZQJYRQlR8W3RmeTiS
2BHZsHP8DSVqhIke9HOhgCAgWRT45jiNt2A9aM7uNlXWCJ7023l7EABVuPPSA7Tb
9LXCmFL8izmL69ktkENvUxIQf8Q27jaQ28xJmsZc71ekxqw/qRLV5CxsTu7IcDXV
XVyZLcXKO+QmIie67XWeG7zop5f4iuAnpXNHwjos5xhKP8lyc4WvA0XgdgbAbSzd
CzhMK+JFg1q6GKycD/GM8QZVH0PcPC0fafKeIN6yVKyniqrEUbpOAqgb+tVlpcuT
+7dc+HCHykJMYZorXkoVpssgz3Y2ojPAPMObubg2YOrso8opGkWH43zwVGeqwx/T
+Dltci+xgDfpFCD0lyr0AhizkBIcHgZiloRHfUQHcfH3r66ifcf57+izbaLBV9Oo
SpnQMvJoqLzNiDzhc0kCN/wezrSpBx0/VfldV/IOo42pJ+AwZElvm4Ay0wgohXre
nkHDIpKQOQ86J0unacgd8eHvq4EELeAFYLPbWmDeJkt9HU3uQnRMr1Wfl1Atdxe9
+pQKadasx1G+ieSqliQFI4G7ETZd1XFLPrLYCCRDmz7eyF1YKNof21VgA8FJvQR0
IZMsn6yAXFallN3/iAddqhFesQA9qRqd8sMgYN/TsvOnKsYNrvmB4Xf65raybU2X
Ln0GAApA3AEbanmEwRV67tKY8bXkljlrb2W/aFkvQAJQffHtsnQnM+N4zR9OCKVH
J5JSiJUyULyKTSRGI7xTmSCieitufbSktOyTTlpSt0kVipDaoU/o30u0NZgrOBHw
Z5TbXV2jlrMCBAlj93TpzaDzQGLsjVnJt0u68in2qX2SNoBejcqrvAN7oTiTcKW2
mmzQ3xKJomfj11j4IOrDfSpTny+0vOn0Aq0SpjSzQPIkT7uXtwMsHdBpaLs3rb5z
v0JmoH/7IWmp5k+pxxK5XN+7rSVhhJp3f+PP0ZvnoKxbJE2v7Ouqb5OgEiD9dp94
lg3tvH6q8yCDzRN/YsSHtbmm6iTIsl++1ZYv2qt1cuS+7/IFO6nc9AbiLaPCPPkj
GfhWIUAiwfP5L3ZBQ9BaBZW9zMXTmgzMBXwHYQIBbN5RmGTaImEwAjV3AI9IKmUj
e2BXdIvbfwqG9026M1YpWqG6sAVasKQ4gTfywKtxBZF+EbhD1iBWuErbBomRULQq
cZBeWupJx+Huw1NUVk6RxKYReNW84LZQqEBolwnUVwaSvrPFJ9WzcBAjG05WhFK0
cGocQNEndTeurKPheEWJZOvYxGJb0ro50CY9wbOE06CHayHELqwv3OzzcnamyHeF
8pcazxSwP7gXHgmhLBTqt/rmVQrGQEos0BIlRzF/lDBu3quHrFNyG07BD+2fzwdy
jLwtQ2M6ANREPZqB4vWToCK/vi0Q9mTSBwhQGY5dQqTfIoFms9AC4rBBfjpCQIax
OAveMEQSZ7FrMiRSEua+vxUEz9gp3XFc+kyHfhtdH90KRaI6neJo8UbUG+lEaxVy
sR/jRVXPVSDjEYphOxo4DIa1Sh1hjY1TVeewA21KwXKx5jXMRAL67K+G9Yn5AJ4M
mOe9XYo76DIek8y2uZcL3sFtWpaWhs77z0QL7O3t0Igp0sZZLi3XHoBPzl05gPJB
l+0C1NMGAFQNEWlAwFFXcrFvVx4pBF1lEZt6FSGVLZ/9r2HFCLmfVF6sobn0tM2H
uFs4uD/tuDvsbKsA8kZyo0CEIvsgQ7KMBupUZ28IpEJ0tp8c8c0tMyfpzfXwqr1C
EXi6dVyGKBRkcmWmCMHpddx3GeY54juxzwN5sDCiuItrgcyeB1TwuFTJ7GEe4JN9
Uu5qcg530oPcjbn79ScqnpJ4UUWuaKcWRcH5DROyPwkMpbfIKQInSsen23Bbpdc7
5pvBn0dKuZClAUThR7R7VZkuZy/Oma9fG2JilvFWDH0BC+8mGelXZ0oA4HMMeeul
xJwnXOEJtp6l28IDua+E7gJufXovZYXwHhdsmnME6UaI5fzwSechjGHqUfE5c1rl
NopC7G7Gf2oBv5kyt42MVMWFkVL44/znvORWaMf4KOgIdOvIwIh1Wuy2SELdr1i7
LDwtIdnlDJnVpMp7xs11zUuoRvPvT38z5GFBd2SY0EIHNkfwGmtXen62gyziGsd8
6Otc+E5tF3guYaxbfuadtAV4eU+F32BPccf+YgEKz/w73oA/ur005EgOA1x6+NtV
QdUAlvTngQQIRmBfUUG8VlgJc9jD4SULGVBrr26eGriQkfNgWFi4bep7wGcYaz8y
Ip6sm1M72/DoDOOC9xlrnfC/nzQgXXiAz8D7ajmwM1WU3/O9BacAtS3K5L8U4JvB
/d6SdOniUw1uy6YIBCkC8dNVprCgJIK0ETe0Hob5DYoHBrTr5OwR0awlIhcfG661
P+AmliIb+kftG/Xe8Z080BLS6ha0TzRf6XCzrgePmhu0oZlsamvCI67iKEEaGCZr
aW4lwzp2vpq2dw9DnIpkErcSAsIfGos9O2spFlxcLTquCxGUAWIEBVxUXPkf0nme
6Sl2IxNrza0vLgmGGJygnMLJPJnTKXz/23G3oj9fx0ZEGMUai5+qymHxu2lHGi8A
Zu764KDshDfhE6sCZfedTyxOM8teNLAR6M7aj6nnjvtz0qgK+00eFsRoCYslH9IN
zldQSN+AUQmCPpi9FcNKi/gZ/IJrJtJGpzGZ7FfdOE5gD+Z6wHSjOOWek9FuMVpP
iR04QI962oYN0A1qsJTU7/PDkwVg0jPcEryE11aoWlA+vzFW2/1xxFE2vnkb543N
g+6yeRL9edjNTyFh4Sis/9DB+TZh9JUKzV7keBFA966RI178QoMgING9ztppA9Ej
MTJVNt+R9xKquVD2hcTCRcD82do+XL8/ioSnILlPt9oYLf3gSfM0wLr1i4CPqsD9
9otc0gVqHPpbauMFS2bq4BlmnabUYYwBEQ4WRCHs5LwRMWoFY+6y+tOuLOBfFCLe
thzkxP/gwHrh8seQnmGGvgFyYi+LJFPDibzr7yPBIGkdCHamPrYFGdLFDZsGPQR3
W59KiJn1nUqAL65mXzucxVcBv7NBuI/8DszcBEfBbkYKhXa/HgVc/HaaCeti06Yv
w70MivQFV9GyAVLv1kDwYN8EVGrsTyuQLFKtEn9FHl0Gu+wEZCvNSDMXQvs8ChMp
jadgKVRWBuLcH93io0pqFEsuBVYjeLFMv6I/HSx5amQyhMAfANWx+XoHeZgpexBd
+pp0t+H8Yx3qbtXcUwaGqVaaplED4IIL0g/looGIgN2IwL0LsRA68YXQqJjl+e4j
401fSemAfZdDrkGfNbc6Cl7qWZl7pngFJcX1Gc/y7Pi+eKzfRVuBXWISiTbWFIfI
n8LdLqwXaoJmzfIoRd+woXIjgONgQvwSIKJhX96ZLFHKxyylW+xqFvBiivEzqoay
oJmiyCNfIUapeUKgzr1NqSgAhVTfpvq7Ah823wucB61pAymybk9nvUtguqEUarnT
L2iGWTtaCwqdptfGNRwI13b/Zt6dh3Jx93zjDSw0L1WzeqGzqI6/9zF2WNDP/j+S
AFy4HhZndgW9VAHJeo6AlLs8KOkxb7EgB5aqzdpSpz/ZFBBT4Zwl8c0vdAF2V8ID
pXEvfpcMBuiB9H8X3Af0kn43nYrplmtQkFEQWjqmLFjLOt/4QFJx0XrSJUD6Nzut
baQQICw77pts4c1XJPsZFxoRNKo+4vlHdP4RgNgqjlih5ErNXUUFf9UOvoorBICS
FjCn1M3qPRQbdx0JiLt7tR8GNasxiww0lC3rr6RsU2oJ2nTtGobB+OSsTzZkUryl
tJxz5uso8ggmLS2nLn2HWJbACJDJm+6juDOZ7W2nvpw7q2b/lqhTBzfQnqsCs+ZA
ZlgwnXVoj3sMSne+VEGC5PUPXIvzH7l4+blUDt6vhwkkWugQwIsfTRsaF0cmdx66
2eMNhaTT5YuyNMIHIz0N7KfZBtSlokJjXLiUyzCp28j8/LJrE4ap3C329fiMWiVr
yy5xHmsOMCj4Bi+Ml6N2bXwEEfEXgXwKaINgyKpR8c5XEZenokaCRqzupH5ZmAgF
nDYTyutARS/X0AqeBGhUe2RyizifGkNQzVfOls7L3ZqbO7ZMzP80971PQRc8HDa1
crIovgwDpRDLG6M2qCVTLBGSqAmEdzaPlug8g/zekhrARtGgscQLaqnYCMZtaLPk
OBt4NYdIwoH6Z+YCP7RZAx32p6XznEdbqQc9ZXiYJ0DkEarwpJpOaj3vmrjPs6PM
zcQPbOsxZcVqByNGjjCBHuf/217kwTeoc70Suwyb8VMbu8/UnWo9XlN5kXXBsWNh
J6TC8FrBiNDRXZ4CEvPD+jLORNDOcpFdbYUOz3ClSlWAVUniPmWsvo4YEBA3kPKP
hnxZ0TZzmQRYK602b1WsoDuilO44+3KHmTb0njA2CucFRhpHbZIAzxBCd4BFzMos
4Pf68LDQBjuavBtDHRYhebe1+lWZQyA+aeOGDmlBQQyezOpxmB7+ab5JE598EOGX
pp6iX88EPaBlMva+TREoaJKutwa08qNtSTuqWoxGB6+DqsDyaLOj2f4GPubadRAZ
GeVdjTBHUncXxl9iP3FiABFUZWoFVPKsTmMeSufbEswhG3GAIj2NfXoV4JiIubxK
W3Uok+spa29UfRXYbZc4FqhhdD4YfaSKBvVjCYk3/wgDiqcbsWQp+oc2Dj+1JSYd
jO5UCGTlo2tkWjhoBkQ4JLqocpl75+XaeMje4Ix5JWzJm8zKQT1MkkPkVh+N2aJd
ydR4TzCBy7PhDLOslXbrNwcnYqwMhNzPzkdvQS1zujxcECOHB8Nss9XY1myS9Qkc
J6qfByKxP8r5RpbDPnHkwRmm2fmJeZNw6FJmKN0CLj3iHQzg2srogct+8KgrJyKO
lj7SZLnN4R15Y3ySzYncevgsrqngJMkRaXAvkCkHbGOR1Q4+OcRF5BxxfBZwJEo5
+NOBQJkFQi3ZP48uuUKQ1ndShnvAZJewXe1k72Ysu1rQbJaN7yq0/1qLbrBbCcjh
TwZbzkUYPjfTx9EzElXgM56fR6EuM7xbKa3DvtRWS2Yrdu6+meqrNtd+4r8Fq9fs
meW67jhNJHHMlJE9DcK75rf1lr6bND3oWUakG7FWcNuH2CkM9qvBqe49fAtzdNXk
HoAamaQEvrFivmuJxgGGQIc4+KpPKE9eGAkEJM6kUvz/QuB14ElnVpx4hmfebMxQ
h7aupG1U+CEu6FT7kSW4Iyto6SwjQo24Ad1vq1aOwSTpZO+dS2xYjACm+yu9oQiW
4GME+REXsehM6paU/Xp6FwZvllxlFcFn9Qf0NL5WUzcI3Mv36lHM2EVEwIvCoXLg
bv5U4Y2Y0zYbo7EaQvAIyxVfrIcxFSSh3JN/PsylPnpPGv6RK79+Gb4LodGKUOch
Jw2X0jv4ihmehf0dDNzjMgLAl1CcO2s5TQ0BNpRyRty1stx+N8JNuayYj0XQ+hhZ
POfXKK8zn72lu/pC0HUQOoK6H+1DZ0Bq6VP9hMp00+94wjGbOWUk6bC6jna+z0ey
zGOvJn7kveqm9a5T7WiTqhQfVdhtv7wbptkLd0UZrl62vJBdw3aWGC51WZC1GQ7U
/oxYL6RgpeECebl4jjk6jZ7RktTWyHTV2/WjeDYjgDlL2ir9taWLkZI83nvZDSi8
3U61OeiUMFor1DG9NC/iEGUPN+OSQB0q1SMBvt9SckRku03NBqneV89eUo0iI4Nn
PMssR6wmzlHTNiRNG35jBDEp5c7Me63M+WcO68y46TWqI62cS/+l9KUW14fbgizi
CJQkRDjOgcGRWndAMfVN69Kf6aOBWGV8zAfvi8KmNCAK0xNFs3tyQHVD3zBF+atQ
SfgsO2MumcsUK9FKFZcD9ySFGhwFmrPePlbeDcbJIbvOZHYxOyhLUM5BIQWuT7AM
0jmXZET/oa8mKg4yls/u3LR4ZzWR7aJJL9tr/QV5qveqb1W/BUfSmTl/DWbwBnLz
fjPv2mBuR123rNRQgSH09npwH88Bg85qQHkjRMkCCkgDTnc3uSj0stMZ3qm+rPof
qOcqkwpvxjIYfCSqCbl0LcZNpWAR9ZNSQ+auBitiJ9xNXPcxH5EYWu88MsuIKNf/
nena8bKZfJFMAxQGt9kaUWvgNwlX6IhchwCt8nN0Pcmn8UJsIZ/+VVA2RR1+4AXy
8IhPoRrSjUS8OZQoRBI2mBk1w3Zuo5w/YibJsKIX1YAwd3M58PLYEbowXkD6l4iD
pZsbDjHrM0j9+cMevm1npBcqGQdT/9HOkmst050tDWGAGXRddjANIOS2KVA0fa4V
WzKTMgrxrqptJeUesQ8ouAtTmuTUadm9D1aahmFhwafy+T43sVcv4NOUbGjAHne/
lmPOf+LdQlxDdTfDMY1Ruo3XWTDYRZVYYPTvxBI1wW0zIjxOW4nr4xZX/4FBSwyQ
ua4iZu0kLvr676Kqn5UHQmhqQdh1alJPusOYKHzQWdvLaUEbBRmCWYXf+MYfN5yR
QeP9KTB/WBloKeuOTxEmGIQdnPotN+2RP3Va5iW3XAoARWRPZpP278PFV399BEl2
AUSWLC5hRtmNXqO8CvqZlk9JYQxe5qnO3CfViMXoRgPY7SZa6FNbfaGgM6mguGUT
2tfu8emsLalpW2AGAB78+sDPCuwgcASVIDTVHv69q5zTb2NHIdg8RT8O2eTmpVfd
sUSC24YzSHU7OYFU8WKtGqKwmcb3W0WQnA7elrctpesCYKWseaU9cP1q5JXGk1cn
iZCZ+s+9JnCjuKBtnO12DjZnUhaJJhfix2ILmOAZ5ZhkYO4EkYCvTtJNoZBnOzHn
ddDRB74bZwnBrj/6TL1q071ECTXaRpmNRzfSp9wKdSu79ZF5N/7Sjw4ZehBaGKDc
EHh478jJdmSmcvqCq4QUdSKDFFtV05su8SvL2a9YPwhgx0zN/MQr8D9DHEdvslu+
wTeX/Z5Qop2v09wmUfDmXNOKkZzmh8n20v/RDmKBgd0tB76N2Z0/CQQS+LxbeqCE
RDZ7hUVPuWOTE+5sKqlX4KH4jWb6p9MN2HsxZ5E1sC4BE22SYJUs+kLZAA8vOzM5
Jrm0h3OWqUVuMheW34DaqkakozU97DhN0s7MD8XTQvvALav8UaUtiZzcnn8b56N3
5ZjtibYDEOhLkhXzQ3erNNxvkPDmKHhv0li6MTi3UtqyGTZba9F5Vu+TCU6Fwmvp
MVgN/C/+WIQFqdIEtxsTEfZCw7PCmhgR20O69Trh57rKpDA5LdhW9SGRoyxw0jYz
Nn7sRScLIaoVS80mYcuS3yKb/4o8L8yF3N3FmsoAp11YTACbvHWwMt0E0wx1zsNV
YAg+8OYeNGJydRy8Dk5cqlYA6HVBj5kopgec2KpDij3UWLiJgpjLOlFrFGgdBU4Z
bjzrG6YklaK6tyWpHG7NOQEcDXOwrOMo9Wh5OZRAGk8exRZhwJ1NDOc2E23wVr3b
asnja9luIMTgZscwzf3imq+41+sVW4eqZmLgzboTGSkuQOOhjDKU2fCDhKSmDkxV
vHV7S3kPgLHClXHKjUB/i2Zwf/0SNtHWoT22BJfmMeT0mx88nFs9nB6lY8ph+oMa
3IK325qvL7Y0+8osCIFGZpFnlEkkSYh5xSHRWcnGN3fv18IKrOaEp8ArZCvNtCGP
rzrMnxDB3JZDLu9g4iwLkDyXShrcMXEDP94J1QsoBMLdnV7U57gTCSwuyBhPhgtL
KS6cQM6tOH0SdJjsW7VUWfJrCXqN3kwmy3VDSCvQgc8RstGkzlOz4uSKfYeS4m3+
D9fWe2qF6X+zoC3nTKAoksU9/whzVBnJ8AnkrhAKN3uMUmq9Af+x8+2hANE5pN0B
x+F27gakI98jlIo/ndl+tGOqxGgxoePDgSTw+p5qX7fnHLlfO3/Ry0pIkIb4LFH3
cAfbccfD7EPU6Sxg6pnzP8oAecj+BYjSpWkxieEb/G2jIjQedxDHlWLdoYfkkasC
2Xv+0zCO5iQRaLceG8J8qrr7h0P6q0GMuR3nDXGItusHRwYM7NICzz+95RynHYvn
CdDLJ1ZB6QdpekWZmq9dUi36N+a0D9nBPLgoRmIwdaY7Tb0B9Q+G0P4erOs1FON/
sDMkJEBc/Q6uRhKeV3ZbYZe4qXrOLF3ap8tVtGDzaB+Ql5zjp7ozXnOMaNHeVky3
mP4WY032O6VrOZdOE3WJMe88FtRWB33bTYo15D9ANP6N2mMpjbNK2LnqQd0ejvQo
IpdqEJ9+fJnZSixRqFdImcsPHl9k/Jnr69LUpAJTozqYb2toeBTbTTKQzrGMRoLY
4E4KYRas0XQyelyyxTnKnExOxeleJLSc0riVUkxluh4+CTkNRbhvlxUHr/dfdfGf
W9qro6mcsW9nRizLFwMcGJ6yUGBA40by/FPVSFqcqmy6Kqap09hL0K6lSPFrxSfb
t4dKNUP7k1Pjss1YJOiBZWVpgXNKBSFxy7L+kXICHFiAdwP21eK+lAI0NYZaeGGf
zFUy2rUaExlB9dD7p0yYWAcMi8TY3947dG4Ka5zNbUFX8+sFei5vYRRPX2HonQDi
9scSy4jbueeld6SSOA985JFc1OVxcoXZoMnoGiaL7PLh4jQtXkpK/gMdjsTQt6Un
rSXyN6h4eswbCdfahvzajCy+EApTBMbiqRworqKfKrYS8KdrBF2C/9SYoJMfzgIK
OYlVYxFcUjg71JVbuNvDvMvcLPh3NQZRZUhGAHGIcAK8UpcdQOfOYUjJb57yMZhK
vXQnUp2PhqgSI/1zpIxZR8PO0qaLdM5hWuinMOo+xwaYv1IKbbkLMQ/EBTPBfX4U
4mAKZrYKF9BA9NMHXjgBO/AJq00MUkMa1QiVB05mM6ReXky0Zm2Xcw9NldrbvOP1
ZLbTxao4UvouNLAxwaXBGOJ3GF2GrmeC/Udncc22QlgExmYUQZuuw5miIthJdq+X
m0i64iRvyOz+xCl3AheLkXtCN9iRyAG6KPoAkIcCAVlAqOBTduz1H+W/9OoDvYAj
ewDGVAHbbxt41vVfoNng9gxsne7p7Sog5FMseOmNFDBuDbwZHnVaRm03H9Bc6ZwV
GTVUzVA0CyLng7WRl51eE0G5xRkwY+YZIChUphzTK/G0yWrLqZqdq91JL6jS3blG
CC4sbVC58pHKmPaziztfwLPjTeqq4N7XoHl10/DJ7DkiDYrWKGYGVUMrRUzaP/C5
4oCbU9itGqtQGPsB4lh21vckfeRXWI7O9Ly0onQK6Tgap9HImjtYd+wstPxjKfCR
ErCjjxqMoowoWJwAd5+tnhhJ62c/u/84ACbskx8AQmIfoOYzwPM2du9cpAJudBtg
Vx1m46X8b+9WMhTkEV/jT7Hug8sUeISYwOW8Y93qiCTTvOUUFJx//X+zdiO7YYKB
eOUAihk7lTBrefQT2YgarV5t1zG0z1VQ2gGjZNFtd7W3l1+TYiAWDBGoIvPm778Q
EjKU9V98IVt4eW7WIw/aXEctIcUotE3xGI2t5opGkWR9joB2Rx/+1t0TzFCxl12+
ZSdY8zBiTxPmRlRwFVyhLZHzmVGdj2P/ec79A+mu0qVnO5VeqS112XtgqC5jWbrn
DStNDZbNYRPiU1jM3fpACgcSCifM1LFdArCGtq7L3MjO+WTw9zMQgGo1GJSG3kQ3
jbtirpJ3rISe4Yp1bg4/n/e7sn8DasPKQgc+FKNNYaZ5s/jBRZKa2v4kHGNqlk/b
08XjAMb9ZjTlEqzBZjC79pgCbMY05tUY5X4T8oBQHVtXgGhQzI0TepaPJWw1/YcL
fvWvvqFD2zAqQ7z0JJ7lSIvdnPv3eJVoS6UTk2J6wEBx8Tx9JeNAcWH1OVUpIGF5
1R7pf0LVCAPdNB5jwxMOFkAEiCKUHLlr0nlv4dF2pls6mMOuQfoeMJVjAjT4WbiD
FxXcg//zSYgbeDfwlciv3CB7V0aq+zn9cay/P594PZHmiBk7baobhGxlAr2+OPn1
7IAT4JxCZ7QpT1VnPh0xRdtV+IzE42uxPFPGu5D+tmBOvu9GdpjKEBRIME/2nQcJ
rtDbK9ujrPnZjLLbSptnQ9kOdZZicPZvtx4Fo62WjzDUz1l0QP8LA3CEPtHX4oIY
L81trx14is+F4ZsdsJWd2Nfbn4GhF4Xq7K9pFpg6VzCsczeD7yLKbVAFIMYN5xjA
mIJspLr4dSdl5+VTepmT6kSDRIPwjZ2Ci9wCblUaGK5795ZCay/5LjlPuAS4VFYb
pnhnRvuoXCRLW/5FiZ3NYBij1/ciceGhWVIIxcPEkPWN68Ix0RLQDLmMvHaK+UOT
+HLIPr2h5wClXWtBwfEQmcjmTGlHH8M1L6iavfgwGoam4/X/oKeh0MqJiF/hKfvn
1pmA+AwU6iQAA/9Xnaba2s2EI5HsRiCaMuPPqcVMD8idK86ca/5rpl+mKVG3HVi6
1bDYOoJfYnm69OsBjR3n31U7qIOzlCXCvdAybJIhkR0PgEpzzvmWvzUr9pJBNmv5
7/w5G5UXQvpMSdT5qyXL5NWiXXBcluXwa/ViSa3mLHqUNn4WM3yl1Na6gL9c/sCj
MKO9jGXXSzF1We2DWub0pdt2J0IHu2S211p3HjaA75/M9Z/KSDUXAK5tqMmPoe1Y
nBKyWoroQjNIwnAjAGhz1iWef576kK37BPENVLNb2UTzIh7HeUFYfuEWkpsLpvVo
dgWHGrMlkh3hnqPG72Zrnc1EEddqBlxQpw7UWkm5cMKwQzB+ZwtoISZBYORBFayQ
/wv8MdxLmUaMWN+QdijP4DHIlM7y3sb2WCsrYLOFxbdA76eeHDtUK1C8s6pWHs2m
GImZIPWg0YtTHn+yAcqyipJWQvjk42Euxg1wlSZYx1Tbhp93yQToyBO/TyDNgajD
R8P8mxEyHoL79XkGqP0Iwb0V/YoU+4SnB6Kfhpjxl1URvUn9lBA/sXaDyj6PBd8x
g/fjnhimDeu596NdKSWqbQCZSgPCgURKOQgvlV2dTBvQbNQZXNtPTcUInBs3lXOW
CV9Jj4MqYh5e2hRHjcWIbbrQfT2/hZAfXHDF462icz5ej0GLCNAALpSiD6kmnRwj
9Pl1z981M62KGO51Vu+9wwg2HnhheACK8t+mvEuC5t78HZUD7QEonvbubnK9x5u2
DeN+R5ti3KmwtYIHaM7rbtQSRmIl/9BWY4z0pnriEQaX1HCgvN22AS5a8UuXqLTQ
fxhYOCjmo0glY84OCbBpShvFJAZQQpAVS+0Emz4jYXrrLqDtTTWyAdEL95wC1HbL
pTWzEW+7CjmeRJhSh90bu4ZH6I8gn65LLHZpIQexse98VxQz5gHHeZpfy5xboIb6
3pUab6pgoU1LnGEmI+915/nefIGPLzcCuCX80fHhAb1AW80mn0qoSEpdDqIUC1gs
ZdNRLV5Ov9q1WZIp1fVoVt5T9ztXenrb52+Wjtcss66akxCus1U8U9KdIp+Vz/4a
m6oQ8P7IEho8Y35Vs29szgIXnW4poawEfH72NH5h7fV3twfj1H7lN58xSN5HLwPl
PoRESOyJXwhowVf6RHQ4+lncZUw9SXZuLeq5VgvAsUts+XFklj7New5O6ejIvY0e
NX45yrxqJhoStWm+LCVwXNTZIl4ePL3WxeCrJ1xB5a4H7EHBh+pIdvT+Pror3tap
ezvnKORqLz88SjtGE7c8pElV33nEDplYar7wPiUsNLjr+Ycg9mLxbvakmahhsbjI
+uVeo0Mx+iek8GJmGV9KdzG7SLqlPM2b6oIuD9n6fhH+3fTaVYy9HuineDYDvt3H
pfl9slXPgqpjM/912Tp5wquoUz+u7tUbsXWtngN7ikL1QWm+SYgyEgJkPpBl4sPp
i0Y0LlnMZOaf9uY9OOIrXy/MjJ/UcB3BXHGsx5vrcacftzpPv3/NAJBTrMpoi98e
fkpLNv8j9HpunQwvKs/Ns/cNPLlPvgO/bx9hxgb8xqzcjlrdR17JYavNv0+utSr/
DeIOHW434q3dFyyrNjLaGyaJ/yfMUFLMe0DC24ko9cyEMe4UmEJ8+j8CBUzV0O62
O/fcSRBJIpAuVV4ULOsy9qeEKHGqbFWeqEzm0Mg8id9JFGpZvTUUPRRiS+tViiFa
28bT6WVx99AcTMvvKnrwuB81YGJy9gK3j2/EikrQ4ebRUt6hZUqmJSvGhjFBCWGS
hRUc52MvMF2kAX+TvpTNkfs6TQ8OToWEAmE4WDjZp4Xf0EUKNBPBrSJEf+jsdsph
Eegna1ZR2FSRQtlzLbyAxRu1c4XtZ615OJtC9EclypWbxb1sSB7GK+SNXnGLDujE
gX2Vbv55RlVCGOtG1Lz7nK37mhrPvDo+WWcGBowkZg0J7OmuqYYJD6b0WjinjsSg
OCZVzya52eYwErpUJyZyZGGBusIZPtZ5129cXLfbYA+ZpDbH/VNUmxxW+I0sfCN6
TWxEqeXPoDLx/g5L95dqqVFuhxwB+raccaOGdBQDfWRJ+iACS9koCdgf0gtNxHRD
43UFATA9p+t7VlDvkX5hNYWeYuIJSPaSVhayi5u/muBykajITUhLReJABNFPwK4E
vABNG5TGvl65gw3Mh59+QyrA/TQVUDPgsuSKw9G0CrkXRPSlrdmNOtYYevbHuFHb
MeweUA+5wI70SgSBeDeJZUSXP+0/7jIwlsdjbNOasIR6MVRFwez3V6+iwGfdkcDN
TTlGqHFiFI6D9Wtknn+wrMdwxFD/yH9ZITw67lXCkI7Rg8bZwiEqP4Q7FV9MnIbJ
+k7SUzWZ6uyP44J/olicR2wH67yAqtAqpT4bFCsdsHUZK1mHtyq4sx5GrSvKUvHN
5V+dAudeOSSMEwh8gTxxREwMR5gvaO15n1/FY4MSOf03Q6ZEMh9sTp1h8b4Rj9u6
W+k7H552RwmXK34SX7KXh6Kn57qntHqaGajgHYmzCUHOBBatPK83fw/Cg9BgZS5C
v+3RKHqp8cok9wmtdKS15nMvOhoYi8sCf65m/t975ljBaAjQelUuBSRscwgiWzZZ
4if0cECHKEwpnpQLZe5aYC/bgRebsCWLpBluY3n6+RH4lE3fJzhawYaCRl1i8Glh
TC1o1q0J5o3Ef2HXsqWrVosuqCyumx87Ft9aqdNxrC9hn3oy6Yp7gwrHKzi98gzn
Pw8rH20TuMMEcRPV4bvebZ8AoCBaahioEwrXg7MB76eXBAPCuqhY1td0Z3bZqqtp
D4j+KP967xw/LwFHLiOqvZ7Xutb4oTYzDdKaP2eeepZ3PI0V2H+er6GP6LVlnneI
Nr4qg6L1baJHVZ40rtDpvZYRn06a3bRqG+TVpJAnAq26xBbQRHebU9avCFjJ8pR/
6OKVUnR95z5O/Qe7Ze/5YTot4DXEVhgmj00UJ1y2kW+Jo25UHsgZwZV9BDPuftdm
4BJxU9ckTrp78LUH6Szk0JcYVDx7GdAT5+ZvYjKn/xXr/wJ5iHH5HdFXKghkNWCp
uD0npoEnGDXyAJU1pTtTweXlyZUi78R0J2Qcgo0PjEwKUB4Q73aJeh6o+lTpDrQU
31BO753b7wClO2/g9AFHTdVNAR4ucXTyrqs+t8LhXnJjCq39wha/1yKS5gxiqLFU
9sU4StRI4EA6Bv/Ej7cHrYVE1jxTdMjNyOzJoUHa6ulnFpamkV72BfwpJbhfhEDc
9Txq601ULFi0N4msk+PZpwy30hEfpSjTIWdWF7s1d6vU3mTgpaOhnKh3WGs/zMn3
7Pwkx9nOchr+AcgwAibxkc/xOkbY5Sa44jlEUSlP+UC48LVjN/2hL8pg/YPoxbgN
ydNapOzr0G5czXFBJWCPXr2lctP0Dcx8NOpSF4NJoct8rAU1z05aVYkpusFmPTFq
cyMkMDjxvNk2bYVM8+sM5GINx8T+UTbCHnitLdOvTPfxezoRAko2UOOotayUfDEl
scF5LFl7aP6rMOscgxIiIzqg60P0xeM4ediIeGPVGZIFN4Kqr5ptrYQ7vUtWF/FH
ZFj/l0YXQhSaYz7MGJuIs0S0ygHCCE8vSndQmKbYGT6hYbwRZCMMCHlk/xsG3+jN
lPFlAU2EE4wNTUuwpyLbUnachJz8//jfr6M6uT0j4oqrHm6s5puWXLh07eYCZKwm
Wmaz/Js5DwKl2ZWYJsed8cil9D+b8KXLtjXbmyqnG3ORG0SUdeKnLNVNOhv/lPn1
2Fier+FhMyqUJfm8zqAH3HPVzr3KbaqD3HP8J2ZJZka6P5/4DWeyoirlnocj9UqT
kJEh6TZ5iCBe83UKZcGxWCUKjyEX3skkHK671318aBXdnJ43gVJrSalGzXrbjLeu
gusRk94iuxup+ar4tAFawXAW3i9BF1pCoAxa9wJS6E8WMsvkq6yjEIzyJjeDlpFG
3S8Jn9m+9agR2jCuhcaTD/+Xmcnw0jC/YxB+ia1H5SeNdszuVMafHI4W0MzPzwcL
RKhbgIognnbEM0VmkMcstocUOynhGWsgMeOjs3TetKYO31qNpAkIQz4cUXbUjXvQ
p424YtNvE/jUc6F+AUsP+wrRckx0EMeN5nsgLR3Gdiv0W65mrXQK6hYcdqPT9MCc
J1ZsR5levxFAW57bDfQiO/mrMRhueMoee5K5znP/je68hzYgQ0/ETmSMCw+J6Xb7
duBmWRjXagy2EZkk7R4dA6DT/sB4Kwwhz0nX7QeblrDsGCHSSTCxds2kmZjGWIxO
bVlRFSnOoL1p3Y5dIO38PYutlnzFnCkIje9PPlF1AMxgp6SbSoliSEKf3roIth+A
Ko7w2xa09bc9lkmUb0eXvwGgn7NILXoj6ss8rMJRPMUiMSdLzX+jlU1Vw6E1gzeZ
ExGpmpIJ62LWsPD5sY/6znjNtV1+HuDNUmNf+OGEZmQZwTu9BElbMRbTxa7+cYgy
tCKU3h2B+dI6ayYhgfw6OfHC6sbMJDutpIEslkZqkRpe4bfjbEFLmW0oH1Fe6Ar+
//aV18GW5u1YN0drV/gAZlZ/5QPqgU56leSSpzKRD1Ntz24Se9jMTfLg13fvV2aY
Oweu1QYfSZg6+jKr6WeJn+NInUADqrxqvUMDQV0mpdgaBx0RDnvEVTEmzNWZVQYA
EqOQJl6gkPCUiksPjOr3U+O3qOcIFXQZfvgi9GwneSgCAaBylS7lg7iNPnjtisUm
8XVBUvQub9frHmTCptQSK9mj7BuFgmh9fozBk5oFQrsVgqLqHnTrzkbBb9p+3aXJ
7pLhQoTg5sOTKjZE+pzy2w/0popWLBLUlXusM6MhFiWff+mQMUbn7QMfQKCFGoDm
FDnV8SVgXVaCXgFNEuyeeEi+AD2TjdQBJriIlln6gBzGY2TbI+L7z+m5/r9ZWpRp
bc2Ml7lgRSPOvBf8q1HgTQUSNx+lwssy/VltoKjntpuBJWqHiWK6bUg1/YQ+N5IB
252Si2lMRafnk7/Evk5EdmiSoTccdlV26vPOTN7AF2hiT0saTjnbvXbpRoAQlhXZ
EPcjTNj3oPOZTaA6Az17IeuyNMBVGOIzCQyRf5mR0YT0HXGOW8cjrMOE8WJXtv/A
sK8MPJeMr/O6F/ZbPFtJVNqlCPhmFTW4+RugJpX50l5p04nTwxt3DZw3tygUbkuc
aShUMdOPgUo4Ug2H2fOPp984bcKchc9p6pEabKgEoKiBKPOiOec9MlWOzcqOoI1b
mNzn+fspw4bZVJOfTV3LY/sDroc2JFWR/4nzr4lK1eHEr5HFV4cCsupz+aN56Djm
WJpydSqvfsB+vHDrnM5bKvFq4GxCMAj+VDQtmqkr9iq3jC/1WynMgH0WTgp8sCqN
2RIehfDPaGsTIkxr07WjZCSzGK/1fxAs8gG9qqcp2bsIe1WJogPDDiEbEuOp6Dfc
+PcoFiYGc/xtCNBkU6ihasdtjcb350XswiYezn3OHZeTcu56//XdadWuf8oD5w8C
WsGtmIE/pP63N63TddKopvPK1c24spMD0Tjt505PWR/C6IfuVicZOzlUbJ2aVI72
71lqDsi0XwnSrIJCZ3hdFlh6agGtkbOAAKilldQpeoUESXdGzOQZtFPjgZdmzv3e
iWen5dxd1ZvVUMHC0ut/DUSwoUxcrj1NQzoV37HPjK8yYjmGa2om9Zud7+Kts6V9
jsiMgrUJb5VWYYDMU0XmSwU/Ln/jcsLYuYRnJRqfPmi7OiWMQyha38x5+AlLAXM8
voZ3dD8efULQdBvXii5sFhl4Uve2H2Kbc++Z42oif3+cdwtA9mWFW3IdsrgepcSR
JNRAAGkiVrS8u+LhRQ5CFkCkyCoV+1kU6xPJe/hhjGkqoSgqap8gG0E5FAgRSHQG
QrJ6AUIyYHBk2hNpYQXZRf/63Ke8PU4vstVFhSIkVJdFWa6LuSI1UZY4/3+0hPuG
CWgCJUmiPNnGI2dDz4TWMQce6vBgBbmVqSbWh1bSNAZwjGYtw8QoiSZtLDjshAKF
ruSrDAxQ8lhaw6c7z8T2Y2T+BQbaKECF465NpFFSeZgOqyAutHTL3gwpsjF74+Mx
4Lir9lqUY9OMgC+F5o0Tcxo7AkQm/Ev/mF5MB9VakhdFA/C4il+/MXKCeVwZdqp1
BeFKIPDCfuugLT2RDVvTb+tw8eoSFALALj0AfNLs2M74KQs1N7VhLT3XgJxzGIIu
PIMvPcH1m3+atdTUq+bQmlIi8lXM0eLCi+sNX0GIYM/5SpbGdObz/DZcDR0iuokS
S5HhD7MgTrQm4My9ZocNv2/wUixZPf6o8s8K/Tw7sUEHa2tDQzoEbzoyPAp8niKe
nL3nqjzWpbIEZM9QXP08iF7ivQw5KUJ/fEhI3GeO3OrVTi5HARj/NX3Wf4yfgwHm
0k1la/lBSymrdc01ximHJzv21AZTFG/HDGXykhGSs4PhzAEaKG65NAq4f7jNbvCm
1qwkkvwE8m/bmLt/x7gyQWIVQ23hmLQjoseEto6DcEQ34igsA+UImLY1EN7Urbvx
+gchzigBdHg4o31vB5PWY2gWB80RH4mzeRoULUFjG7dSKiG+SMJrFhtSQI9laxZx
qzeV5KyWPVCPgFbFbqvjs4jddRw6B0ek/V5iA4rZk8XxkszzrtjqT0zwzmnX9au4
1dgRNH7Dikq9ueROFxyW8E+no4bJbc9a6DnBcGeXoNhu6+LLjW/7coLwdy7IQa20
Mb9CJnQwTHIGKo2Mjn5wvBOPRrXuNBiJxrGSDl0LxriVnFLDoujGBKYh+cNtPdE1
wnen4xcoN4P70WBgqiOSv7+fvZzEtfL8146G2krTj9HQpONGTjpAmyNa6Pk0SVmQ
o8C8GVnCN1F0Du9uAVm+85jw8vCZeJ1WtHz/LFaWHb5k17e94eIJHwJAdlXrHxU7
/gD6bDbXkO+vtq6hsNFakTcufOKEuiOnfWBOxjRjY7gqo9rZY37eqHUvLSLq3vGR
mKsUmxgpQcUz28KsPgNQjlUbUxOLSrxJ9va4lxea/dsbNiJzwnFyZnIMouNEg6O4
9gVdhqkxt8Ezeg2SlNds3D7v75mb3pwid/BVfCKdXdfGt222x5USbDtJwef6aeP6
S0ADwrQ7+cKWI5Ro54BcaVlYRduiJv/YQ3piG5+XVwjRB8pILevOtYZ9M13TS7lk
ZmVms6GKWoNZ/q84KDeQg5JwDb+uVW7p3AH0Qyfn5GhOCMZFE3WtwUMdh22nzDqk
3/Q8fkvnJF9wesYn3YUEP9HgQfRwlL7Gm66NsIAsCwfcP2kN4SU4KgpZkd2I7FZX
FRh+2c44HWhhFCRLNSJBjIuSRKE0vkXGovu3Sfqr0OqdXyWa/H8LzAcHM03WVV9Y
pLz9ZsC28GOyj/slsnc/21Sm8zxLhfCOeyQB2FSnG2aqO2TsrskqbnTw2+ea3cMQ
rSa7dRcnfYqKoPk4dFKapgUudwuf6TPUGj/rvUEBpi+FYKrOO7O64HXfA+hxsO+w
d3wLjKKNBaDMJ0Cj9S0Chd5Xciw+mNlUSNP1A1Rw1OF3ift/ihcvGDgXgKLg1DEU
RcukJR+hr6L4Xl5DWyFSfLZWeUhsQqVOkVI74FMVYwSwJicESyWdLyHYgBxjJ5CR
yjIDrQthrPChHwFwMhtolvixHSPSVhhs1coRMKEGTj7+Fbnf3z/Tl836On3/LScl
jXxd6/YrGU0Ks5z8n8T3iKeYncY9w5pytw4uNQ6B/udEcPwpn2ZiHvQf+3YIAk7t
2fmw92cRFTg1VBRck7hNEBFmjQ+xBUy99tuHq7kq25MucDXSOuu9mus4CsRVckHj
+Al98zEKCQ87qsMWGJv4Ihw9rh51FWdkxMG95HB35rmuoHlsbqQ6hyPwWeZX3vU1
BQ0gEZUptiJpuO4b75IenUa7va1PyXIRuxeg7+SxXIeGwDCOzJ76aqGLTeF1zRiK
aJETgb9XYTr5gpjBdbdjKqPkHlZ31P+lCQxoWMTIGcc56IVPwTS1R/9RWACOYVel
OPJi1ScL0yIB22tcgrWtYGqAqc+DEYbGmJ0eoQa44XE08HpiPz7vgbgevPaxUR1T
ktJs00u+XxoZCILOkAAHUdRB+V71AZnpRNhimTjCJ4t7u5azcxNcchsW81igQeVW
ZtHQuacue9/ep5rJwRUgt+DxdeG22jBdcdYPe8RmnWIie7GFY9jybseDvB6Km35R
n11W/uiMDIQRi82sBhKqVda8d+To/VqsK6Q9RHK29f/O8rwgCUlWUMHrA42otenW
cUFpbRMbMUH5kC7FQNFPWTxJQ+D1W7dBrU27Hv6pOFMSeSBDskbPGKJnOyFd5T9H
ENxTSSP5U9xMn8+GOVwtOriO50Qsu4/A2ncuoyamRL6aNz7ytGS1iRTmISoRpeN2
Qg0YRMYvJAVTDltlYPKazvGIUZgE/TxGxqXfFW6igoyX8nRNgMw6eaUa34RV7q1N
jTYeBHrKa1IvjOcn+EEM3sjyBt5BrQgPSxvf0ftqw0ZpiDQAmmu56o6xJc6RtOAm
dNWh/6gg7pAOGQnHHIbxSosn3Hxg5eMADvaHqID0/AqxkzdA/pc28ZByCrAfm9Vn
l1eCrCbCQuHML4eowGPaW2q3ZR1G1GLeNPT5dfTIvk7ILkz2jQmDKOGwj0VfEfWo
a7HlcGfBHohaWhs5kwu9VI9opbkZr5BSjBKjKFS1rY102GuH0FXBVmI1Tz0jNJ7u
q64w0QMNltChiU56NUmxV9HNyd8usfgzPyEW+v8W9wkThHmu5Qu1+bkatI+W2zj5
Of57eSBTJEF5nqTvpnMRPp0ZuQNMcfiNC2eHQ3NbjY5t3y6MBkZElt1UttwSPtzB
e4dItAPwl5fveB5+nfewPtFh1Q3NoOKOwxytx3IU0TcYET+MRXCw9XGVeVzr+RSr
oMCjoHBs81d0oLzjwkl6vJUcsia3f0OyHCW98Xn+xgDuyrtLPs8RoFbe1XGEB6EU
d1wgHdwdGVXI2yB02T6AHEu3BiVFnuqH2WMKVEd7H9ZHrpCdbZmCs9Jq7Za/dxPz
DqXJ4LWuJYjNzQ80M0j6/h1XSiKv2SbeC1iYX0kYAd6ePFtLxDvErEdZ2gmQRlf+
Ia+6B1guURl6x67k6a4OhGsC864sB/RqcaNIsbSsUQM0IIK++Lk9g7Z4mqftY8Tk
J4h1k6M5FsIwDYMhSmMTdwW0dUmALyHCiPF7tnaelBrygSPw/smx/53ITGgLmnh5
xMOxYAXC5ylzdx2jknvYerENMIaprl8H/YQEgJF6EfmNjpc6v/suhsPuHFNg9rah
o1AThZ3+au+3rGf2NPR3f0Bb3BUVzWlki3eb3NjM5qg77zYUoWQb75+XEINPpcF9
VnVUC434Q+5wNosvg7pTYmi+/nTjQNa/nfSy5satKFDBkrWOTJaJtxGSf/ixcQFG
/pnmS8c9gbwSxf9WtzuVqRTdoyv4XdgXYnXTlpv2GxQ0hHV0EZ0dn/wiQukhWD0p
IIil7Gn9rwAi7HlHX4ldUeef34CeTDAXtzhrTbbPfE43njRbIfZTdNuazyyT2BV4
25cfiosGtCBlrl75MouqGLY24h1e/Et7PcKGDbI5oBWlwjMVARmv6EAOHMgWcTJf
rmWMpzOVYylF8plnXV6GaL9WOKJJfEbLGePXhiA2ep8s/n/YGkQtLZZUst0bmXr3
gsplmdvg/bkkA6HG4W6+Lz0scMQfRH3rVPj67vKyzhDHNhIYPu+Y6K7CvjMecQyO
nTY1zWzWKp1cTD6d2xQN8+gGCrdXFzjD2QepFG0P5t2eZV9PwuyCeUUX31XyPhlc
73EJQmKG0yJXEmS8gpH4sw2fQ6ykUuQMJXla7fzM1wqyt6rLH0PTBvChAuW04s1T
deu7Sgz4aIJf4yIBAMQ0s0SJ8I7hCo1MrgAO/jQ+9krhYNE2vwvcstAinKqHsVlE
Y1sKwMHdZVCI82W0HtZ5LmNQFitpAw6r45igopn67cEmL1kRVAe/4ulGe1vE2a++
BRGLmx8w80j7EPLTPxdN6eDy5tvRymTmzCF0QdG9qvHktL5EmV16ehJdetC7cZgg
nnVPJq1O5m1LxEHJSWWym5Ithg1GJ65drOGrBO1Choj+mECNzIWxhfoFKYs7Z/r2
ZV8uabFUPdlQw/0paroG9uBHS6U8HgXTpQiXpypiu1EeGmHWQtN4DtcK4pOIJVUV
5/P7jWjOCtncSEH/7K7FZ2CWc9NrFse701l7DLvuQHhbWsXeGFxfWv+ZiiFWOGX3
OJ5bfFFayQdPORXx+yUG8wzjXfedGuGW70Iyxopia2dRP+lH/TVc6c9EfUkO6eVJ
QVx5Yjmha4tV+SefwuvKPaYmVqSTaVCoCLJis5A3I+hk4GEPtzDP/iNniXbgHZXh
7HmNuqhLsIJtvL5F1lJ9dXDsaWSQvsJO/iLPuOkAYnpT/NIWGpfBnzIENopryCHi
qKwz6hFnLXqC0hc++7KsGd17+9mXbO4iUvjL80j/0S77KIg1uIM+nmjy6r+6AjDQ
hd6/iFl1nFmPArNXWMENKEKHA24L8rDed3gISjes4lOeWSdINDpy3n8nt+L+OAne
ajd7GM4p7bc1rNQ9I4rUym5wuREUvWG3ItXngaRKH51iV9f2E1d7MuU3t+XQ4oTy
hFf+NxD0nYWNrgsKOaFINl73XJR5sEPjaEoSfHcwfvguvCqjSaaYXcFRxjv1qxfI
pUjETfWjeUCdUS9TO8JY6SXxQ+gO59XFDXQr7MFb/HsjbjViE2vFfXkQuEUnWbGa
VfAbR+JWtnnogAP8Ejx6S+d/FbJ3n/l6FK9QmWdU/xceHzeXoA0exWWV8QQUke7O
dohYzUWrV3lW3Dlh26qsjA6nt42VfCSgIJ9Rsdi4jKt00KAH8TTfyPxESqu0FI1G
kFUFy+i3x6AlfChd2cx2QLxxisQ50jn+8s+HIXmde0NhLBDsCsyR4aDTOO9YPg7U
NYuv9J2E/hVReMrk7gu62paZG4Q68EdYyibiTqEmO09R+Xnh8L9iFn4O7YDVjz0A
DR8Vqv1HyLy+37AnXecx6cWTZ49j6f1vZZH+f7Yji4J9hUAeHcU5WYq1/qXJWskD
Hles2qnAvEgHqqesWI7sBi0/nk/mWbTrCjzPunpQrQf/3yxbJA/1cKYpum8ZXezI
ns9j/eNxPMp5R/DzfXPZYgU3a0+1h47b5aN2NCSbQFKtiN+DBZRrYDX9MXeDb32P
1fOAz36XA2ICZ4P8PYZQeLgjxrBpx97pH1UAtNoyCKfa0US0yVazxfFnIKfx3uQP
Asl3FmHsO7pFQ/KQow5ZYUSmna19iNz0VIU66Hy8hMQgmfB8PUaymvjQWiKsPN7U
gbVKAoZBCgj8L1BTayx7z7ChW0t/0Lb8HhbIHaFn8RlYLusHUpjfiKBKtsJrtZjp
I5VRk8eYorKIjNZMUEwmW65AIANtKReu2uE8KrGVsF9gdbUZ8fITuHqF86vXH/yZ
vG79wRMDSeUgJq9p2immRNwK1mHz7vSp0K6saxA7PC/FthIX6gkRYV8yFTdkOg+R
ymBL3vxIfpT3EVg4N6U5W4JIV4OhGfl350E0qKsia+dOwkaNxppzZY2o+QjU7kj8
A35PJUWaaTeg22sc/g82RqcdGt4QrvxKhHzGY4g17WuTXLme7dWV8imNtEGUEi+W
yoLH6Bl11L32VVdvxC1HwpkIQmeUOegnBaN9epsVOEGUP9tWgu/Eb63WKFbwijat
MVZpG/R2jpxSA88D+W0wgFZBWnRUrOI6+nGwNCDN5R2bajGC2sU3h2CO8yhM3qYb
ZMx9XRvimfDdOVcmL/ykI4LZgVE9ufrCSDQ/NCrn86I/8ZU3j9nIIM+fri+4dcbw
lS+Fmtx4AvapW72b2ciQT2Rm9xCo8H8pCVcRzQiAIuXjAzfxH4MxfUEjg3uf31IB
c7L16l6/7cFQMRGLmaAssqxN6WyAB3E12KaEJ3tpZ4mJNUzkGL0T3MnzjZsrY57i
Vf2PdYu49FX0+1EdEAUSTZL+8QzfmSyRuAJRxWGieLk+BTlxi3IOyIOLwQxUOM+9
iCoGxJ3o5X0367z2+wl0qMyuUg0zWPIVQPvY8SuzgGgwLCliJQE2VGJVzISglPAB
wK7L1Pz9grTIPrXeRe96cPsp2D46AfLyqyCibAvhvqXHuaaC5nptH/SkUuB8sydp
TUcr69zzzLHel0l+jEFNG3agMNPY4BfhpAqcdxx+c27yUnUTlhdvwi00NiG9f0yC
o2wJ/QPW6jgu/0cCeEHJJJ4De8SNAhUPURrTLkVRJriFju9R++iw6uGhIAaKGz59
PNY6ZKUxTTzatta6m8NME3tgLKWMPx6xQekSzviWFACwt3CxzIJZiFyuMxt/kvbt
vdbTcArEkUB2IStmsp4otVVtCOeav5tgZB94q1lNUlZsPnzoCxVIXrkjIrJ/J1w1
5TEyO27davsgrkUw78ImvAPpceaLvrDBCqNZxPxfOCKfDt+Ps0ucYq1nB373R271
c7+w0Khx/k1Rjg5471nsVGR3VPx8X4uHUlT3RQYiR3NMnKmJ6GT0xnFykEnoSOJ+
JQMdq0CJqKYg7Ps/ZxfaCK82YY1onWULDzpFsxDHKPiCCyxUazn409syLw+fwHgd
lPnRD1GonWwHGHwmfYuWl+cE0bDJ+mhZbWu4ymFNKvGiqktRytRVgPpkyysM50ue
eHTbOZLuTZQ7niEdYT5KGgKr0nDwkg1Y+LO7xcgSLHr8UYRIziht8dNq85ph+vg1
rxwbyI21/AS8l50S3kQHYuuHknpQyjVlePnEZjacO5AOX6B4xpbK+brqmef0o3md
4t/wfKgIxXW4k6SMBSaGzFWVdQicbwYCseIuxIMBr2s8ky/U/SPyB/31QfI2bVHz
1AwtW+qEvddyrgweLKhoO1MMI4Wq8pDDqWWaF4fHryZr/b9kADGLGaHRxC/HJe2J
GSX5lCu6+jnkkUjN20+u2Gsq9dbcViJ1aVgX6X0pzVVP1iE5jZmEAhOFHuHgjgfr
g09kRCECuv+GztM/RBfM2WHfLMkbJ44op+oumB6sw80TeDGwrsagVGHz0kJh765d
qGso/j9/RGySDcF4Fwr0Iw9uCC8IUwLQ0jHCAzIbYNYgjIbnJ55HCk4QpX7HJjLS
On1oejJIHI7q4Y13MLpbs+7a7idtapsNKR3SJk/JoZ8+dKu2i51qOseJkhB5zO3E
9n1NiKD847nSzz1ER28dBtT0oGC79XldaOdTzz4zDX2SsOv1IAZER8iHAGTpUqRX
6e/hmFVCZz8H7ZMEar2VXFRqXEx0fbgti3uaOVTmVZk0ViobS2RRNCZgLn4a2xG4
zS+Uma2swytCHr/DG3k5XREKhVtdQ+enMgj1SgN327gUJJOsUE4JahYs6WQ1tVkF
OdLiDv49/TWl0K6gJhgsVWtUZwr527PU5Ma5Q9Z0A+5rP6dsg5ULwJBGsT6sWaBV
8L1vB648vR81oubaWElIl4t4ZjFT4XyJeAUjQkeBzWENHfxlF31rSAWadqb867zn
CME9IuR4OhEhrsgtp5n7zNdKZfcss4z9KtLwtlWkUtZRqOStUB7Zg4Uzvc5yXjpo
Bvp6e8ZWpJoUiKS30ByT0ch9Q2b+0tDe8o5jpxg7Gsx5FgxHur2hca+lvPzcJb7L
FBA8V6gWVQerwapa0MQ/bIZYIWE9GKeYiLqa50g3nTsPfmiox6I7bpX3kpkk9pYX
YcAwRRTrGnNZ5kGLYigJI40ASRXRvU/2mIaAfMy/GNtKwUYPIprKwVaOSd3jhC9i
lq+PkKCV8yzccTP2TO2FedSZ6H78QzuEUR6tCLFRthGIGGXvCa4hr6mbeJz2hrB2
5G5g+LjVfub5dGX3djn3qbkhqXLhCkpJ+Y2HSTtu6/hHRx7sJikWxT6XdpqApdTv
jQnPEejOOMaUqjnuCQPKhlUbN82EbUIsYLcMwDKa+dHANj/5KDvRqPKGkSdBAevL
x/tHdCpuErhRIxvZ1HbQxy8SQdv1c9j4KohcL3tWG1XgtHTrBAuvKSJ6Gyl7ARgn
DD/YiPmIhR7gefDiW8ohjEhVTy8v5cbzQWTgS66z7YoPReHoxoDvtxGIMWbE97C7
jJ/bopz2Y0N2kw0iaeInzA2iTnze3K/PBRL/3Xf7d+ftwXAszuW9YAD+lnkdIPTg
2LjM7d8SLRJcBpVPItMPSY9U5MptHGwrweoZe0xjM16bHFB81BHQhLNi6aW8Wyjh
uiY/unWdnYtEsMsLAjW+nUszxnqmWQxOh9UAHLDoAcdJGFJjluj6qn76nSBu8cwB
5GY43T9qN1pDGmgnrsJ2j95chdySxd3k6JCzVjmLdb1b65V0/j9bVobGd5+5EIds
e4oxExj7eKcophMXIfp7mlkPBv08CKPMn044rmgAY2RUOsBXKB9N7nAsjtyljiTZ
y6Vu4nxf47+csxmYodL0qWEL30OXmI1/26rbD2nPfX7aiFDci4/yNn3usiA4vqDo
E59Zu5hgikERyX92aCTtjbS64t0CaEqClj3CtV3nLfv7NX2pOD7RpUSuDO+xOHQw
VqyfPbcJ8T6B1Ty3idt2BY6XBaMaL1+qXt+0J6d1cifPqIy04c3LaZG0QZVQhcMq
5mXP6QLPvdA41PcBRuo7fIRKOJVV2jvA9k+n6AQSEjB4Nbwec62l+pvfKaYSb50Z
3FdXQ4RWaYs8KnAPRRoyxyB3IYdbK/wuAAyHd5zHDzxwBBxxGxcuVZm05oiawJ8o
NZgXByM2OQhif6sPGN+jplgRXglJdHRL0da7DZzLgYByyDofGaBeDuidqo96JrJn
UMv9ST26ftRA5UNNvAt/92tABuLC+zrldXXqOklV+ot2PyqpN/y0puE1beeUos9/
CG9Gg69Ce6BTiaI3cx3iP9HJ+Z6wa4ckppUmt/aM8NQyh6gpXeaKVWOrWQ7114Rx
qrUKIjXWcPXZiahJ18R6lD1HFGCnuwKaX46sHwjDe0hSOM5H0AlbZ2Yd6wlx1u0H
4SJO2mNptoQLoGV3lPUzOuI1hdCW2DAze/SLzWzp/ZxucocW4tS2hl0v2fbUO1Xp
ZZKQlyiYwkam/d2Zltnn3DfaK83LG+Vx6ENgU5AXSK7AM18JiT63txAOBtH136Wb
J78RQH9jMr0numVF2eUVPvDR9oiIOLc5JVt42IW1clEn/FkXkOgTevYPrnnE+kef
0XNpM5ViTm3E/ozUKwkHUTanPO5WXBQUVi4puM0YZ3bVzrbdX2wV+DIRKhibCmym
aS3kXGadgXDEl1ipA0doPe3vuveN7AX+CrlT3aEts1ADO3KE2Knk0eMryGQWQ2lT
xx5ntRoBQEu9H5SXhSJW/1d6lIWbw+kWH+6KPBI1wlvxVbE+I74BSyGjxVdzIKao
56HMuoVKmAK033Yp1vS/jEAcVG8KJerjlDbLE6JyVPaMWRpPHUo2850c3rePnPkf
ITYgZvPbeGPJzZg/aKaD193FXfA7D8Hc/BFpGBg/uzSinIJP6gFYu/IWJGBZUUN/
G3TVWS9QTMdBRmdBglZtUWSrAP+yLTwsdrCqifLl4eD8ReaSOtXELq2wc5v2CRqQ
mcpo8v+a3LFHoNnk6q+VKeav9/HlCnu7OHATsFfwgTUMSkDePw5Lk7MIykd8A+Yc
pddmv4FzhqtvaRkqQchHHUAEw5wTKp0F504mzXSHbE3ua6OoPRGXnw/6sgFL/RUI
GSw2ooKxywjLp2txzKBAVUDx/+DXvjWJSoryPHbDmJ5ShYzc3zrysfN41gz0PYdP
O6p+5Ez7c9i1Tm8NF7uW+Ja9nyFI7Q3GeToG+ISH63P5KzNihxNZRsKbOnU+xJSZ
hT+0TwEUdw8qspq3n3BHpbI3Cdak7y4IgxxS5okoIrJUskNQkCHAfMKXdwouHGci
3eLsPhluv7PGvWWbXubi6aVBnPywWfq9w6ux8KrY1rOEmEv2NM7yQz66qWAMndT6
w9eNvqsHNRDT+EytvG9JphvdYbdHlaJ3VyfQn4DngdP0oj3k6h3kudsHVk0Tavjz
XWK5Fq3/rEhNF8OWvDftPvfSYWPAY/9Zb5+H2lrFZVvww+vjJfcLCAFVNL+zWNwi
IwoTZe2mSjfmf9eJ/j9jCS7CO4S9XWH+rsvI129/C8AB2J1ZrX8lzsH3YtrjpIJW
gEpKoqTsHXzp8g1JoTUN7zpWW4nSCYQeqeT4WR1zI4ZUgvkmOMTCSHqykjF+nBzN
Lkn5+zjr87PsNCobR2uSjtgIrvBUBylDxhLOnnqneeGqQ1SngzZDhiKy74K2cNL8
VwR4BeZuNfBlxtcbZq7lsowof6i9lUAJXFpyb0PvKPcQyNkpODKRlR8CvTjlJWpu
StgUgUogkuEAoprvUhfVxazpFkAYapma8W7bQcnzdU8AcvR27yZGTwbzBAx+Gkt/
rm9THWA1JUPnNx/Q96UNbirlV3WZbQwOv89CIDUhJy14843uppN8KcCDwsRkdgHC
VqzO3MS8odFk+HoqNiEeuiB8c8LDdBIcxdz5H1rgDP7QY2WgRfb7KFY7dcSel0iK
K44mrB6IXWjFn+vOOVeehzquNpU8WDAwOZnCvK4vv0kuoQs1u/+tNYqY+zDY1oQy
yhDy9eyifg1JIt1z3rJiSijZ9C3x37CsTI2Aql2oF2xcp8WVYUXRDlEkZf15jakc
jTMkEyATo/8HshyPoqK5AkXv3n8whOV1AK4HZrkuAg4cI7V5fLyYiYeMWq03r84l
3H34VaOYXDd2TlOQGVz4tXyZvogJoFmimusrkUoCM0EyoSxGE3aP4MIX0GP0/Cfw
X3GqComvOazqMZ6YkJIuaigy6rVhlEW++TYEFx84OmthuYvyoTP2ArtmW3dSk77l
/md/GHNifAgOr8mGM1HiyJIXLqGsNEEuy90xPGDxxq8vZpZtjltnP/UYDHf6oAXU
qP5KyqVcZNfa31SVjB5uFgotPG05apHs37ydgP1PaaZQcpe5yk1lCb2W8vNwzfj/
STxFQfCV1TJSNpBdx85/8pjq8cCLhYMTYkNJGhZrOuHL25ZfSu9LkgMIwGHU+hSp
k0Idk4wJ1fndhq7pUJUH+GFMebxvB42DM77XEHmzwlaXEPiaL8O18m+x12V3wKcO
nNocgBNTwMNRsQ3vBSSDJ467W4f4Qxcsie57GjNhxzZvZ9VyIn0R9MdxS3Rija05
JnylIzRJQR2nlfUSwa0cR7AuE8F//QK60wXHNdM0P8+1P8/f5X+1ov5Lx0IRVJsj
SaWRjl7r4RZSuGr0qd2v4iFBVQBdgsOddUG169kW/XyR/ZWU9avy6IBOBwvmUoVw
xxGt1ulKVFdqsrdQgz158QTRHMBfLpybfZXss/Mnveo2Lic/kZBAoQpXzmSJvr8y
VsFQC96XU+gLdKb9xsUR4DZkzixyJRdfB4jmzi3xcDDW5X4LBcxJRqx8RiHquFL/
587XA74EfNysKiUXpAqjPEIBnNz+GKDLGs61gfLFiGMJkE+PCOchjKoWnYckrWeE
eX+raw+aseLjkoXbsM+p/C1NT6tofQBzvbIkycZaEzzz6NgO9Pt2KrB0zeZWOB1m
1sWb8fV1+8hCYYjXRYPsWdSeUXlFeYMDUXZwoTvqQmY2zbDuAbj4ED7BKJFlG7Ah
5f+sooeVweeMFmNV5LtCCHiMGyfgavvMpqdGIvuyLNLbqnGulVTE4f9Qi4gq4c6B
gUXLu6RAEkrFuKWZRmyGQU/ecuN3gButEZnUl0klGI+U8oAN+46gtVey/4jmvwn7
zhKaFK3CWotxX/o9EIoNBztnth1h/rNCNmBty2KMoSV1/eAEo2OOGIOJ1es6VWcj
qlxQKxZ403t/yLoL8M62u75UIygPxNyqXCIDq4OyeK/u8cU1Zo70uZGbOEoY7mUI
BLnuYnPgCBFso00j5ieiGKGW8NzSsqpzWviSKYInymwCpu2bA8NpX9imwS5eZ8yU
q94yX30ItfZpb0oJwBTJ1SB11iEZctdcXJMHZHJgLJ/Yc2VAYJQ7cJI1h5W3brYu
xzl7ssRDe5/GZ9R04ek67rzkQmEhxTtzwFwZZrRinmKwOB8lyjXnFaLK8FIEjAkj
Laq5ltk2zAM8q9FZum91MR43cEl2xShRRAvq9BN0XkQQEru/Y6UaKIc3RRNxvsu7
cgW3MOVQLYKK0yLmATT5o8X7GYIDrqoNkuEzLPME4Y20eGep/zPaVCtEWySZZib8
hMgVw5V9nkkf4Wzm7hrw7u3QUm6hbUoA9vFpC2l6eljqWLY2ulGDT0YoGrqVjPkK
ylxTvhpcp3CLvMDNCLzHqjadaors4wd5gRSdKNDZyHhobvjeCyrcdLqtt7DBFDfR
bvnpZLOnXdtqmk6WEWlDvb4s3gma2ple9EUf8pIhMTN3rK+rDtNP3ZYRS33fF2zV
kIbg01OQEefLz10oinJ2FS/EnAKmllPmKrpqknoin4vAWNy5L9Jrz9jWrorazNGz
Up2SvrOTxpb4dA4cEK8v+0H1ImByI5XWgnkFJ8bJOxhHV+mk8/WDsyPosP97iq7I
6xKuYVOJTBF1ToxrLVyhHAVQLDna5fb2yWL+/rhpmIWE/IM1EeUtylwk1v6EMBt5
0AQpBHg/tCFKjiBAkgdHWd0RwuJJ9LpoJeZBYLBwSbTHrA3F9haHYKxJP4OMCGwB
jVWD4xUEboRgh6uNlzaSSQBSVY3gwZese/R9hG+tEuBaeCCrG+0OrWGef6alpVqb
ysy4tu1YNyJKLGRhMT13tID0HhehXWifmc1JtjMTNNp4zAHfR1TkPuoIWUmOlUai
6qYq3E1h0JzvcoywGD0LnkURjGyZf6oJGk+IK5CjZP/rcFDjHj4GfpTWB4Ok+Vfm
rfPuJb6lLKcTijp1x8T69arhyA/gWG97M4tXZ9FabS8d0DkxJRHSs6jLca1LrwiM
LufsAmsPWm+wkb9+ekfypJ2cPZ7WLoxmEES73Yu/WA5nn5nRBK8bsn1/FttSqgOk
Ev2exxip9KMmnXR3cV1OumFXgjbL09WMt43Gw/D1flNJ/xr04uT0J7lINjEVy7Je
858zzVoVV6mA/hMEyPgRKEXK2WV27T+drEMYz/2JyD/WiSwEgX4YFhQqiayNoCWF
jc84yqUA27uJqpNDvhYHoqpZkeEF+VZB4X6l7wPdNSTKJgwc3SZhem1Q88M7RGDN
9mjOGoMaAlR1hzel/0CbOaSszv+Y5qhSnllGyzg8QV0meQoyohIjFb4henDLoQxo
+/PGBXIH17pQX5Sn7B0OJdRuD77S3in9xNRD8cdt8/16ve0YAgdBMxugcZ/C0uA7
66tZHRo6hBev1125L3C7awZalieIzuZr8kGi5+/p7VkcDoASWYiBekQUkQrwKEYb
4AcTo55829LmtLavfbxSFHf6QMJdakXhvwbcHOOzkjXsdxlrmfe2d4DgFuBPlw6n
s1o8MBikrQi8fUEcnieYzsEh5fREKSPW55Hl+9TTUK1wj7HSatviKNLVlpir5mJV
QZ4MNPlhhoHN50wQjnWRbVF2W8YdMxhIkQrQORqszu2aBQCObGc8f5Aqa34oJNzX
fv9SNsbbaSRDIx5Ec3H8qBu1Im+E6s95wD0aPJA+4Xv94IUt6U6uWJ3ggJ+OvcxU
W6dGtigesnuCWWyUssWsph+dDj+rShfirdjG3NCA/g6DQ2gQ8aPIpjww3z7/xtVn
iEg+/lbDFLOudLtJZ1NO7jURnvTsxhopLGNn2GjHjtUgPc3hTu99H+EpiwlEFnw3
NynwqdbBC5lZjSZYQFOT309DMTqdlksAFvQn4WeLUsqX2xWnutKJ3vUYVq3wu3pu
Dn4gJG3lpGrNZaoSUOnHZ9wCwYM2dp7zn7caxnP3pw7stje1AFI9K2yoSql34wVs
HRtCX4mPsKi/MLVg0iQXZQIapEoIn37yecblwNHOdwye62ABOBsHqPUX9JmbyifP
oeb9CUNSRXC+CCgF6QFJBsKBXFA1Mm2M30IDVsFy/WXNlhZSJhKPThweuydFJlv9
Oj4OGhF23nMIMuKZDhF4jAmJ7SFi+EhcgRY8ZIoyhtwNAEIaRYDxtNlt/cAx9za9
lYfwjmhOxlttYg3yxZy+js2aVTRFKasJzsSZ4cv86U9jQPvYEoxz2kEvcubHXNHL
/+aEl96QvZC0eJyqhWr5SwSkTzy8sSrzrpxrO0OGEtwrzLh3ScpQ9gy4aJNxIyF7
Arjy7Rj12XVU54HBl/BoY7/cT0EOp3zy6nSFVi4TMduO4EQh7wfEoojaDKBK29Kq
zo/9kOMBRyvCutHD3zfER/Bdb6/3YEzfIwFH4DFV//w1gmia6VPQV7DwsM7DFJA8
S3idpzc6VZFsklUdw/TJhMwYXqk4CjiC/dqd72vZHGoj3s5yIysfmuEfbNJiXR/T
O6+rm4Cl5ufoEkH6xCEu3xMQUSE4QYCwylM7rddqWmCtkosHiXyXgxIA4nEpOQkI
koHaBbym7DigSb30+gkIAZ72hklA0xIqAHS0YgHMdEtv4jTM4ETd6pRgPsTrT6oQ
SZHDUDGEEHfj19l0teDpAH/KpLB46lfluoaYwBd96gNZ8u8EOxHc9UCq+rWi1FEn
aS5gTM75u7ALUTpTcxSjBHi3+2HP937UIG2KQz7IyoG9nH4QfEsyTWYumxs9FnKD
6Id0ZLfO3ElMuU2zTniiwFt73JVmcyEnOH2AWDvoTVS3aaZddZ1dUiNS0rrK0qyz
Ob6yMzr6ZYcy+9AJ6ISuuxrOLOv99ou4p92fquRc5kF42v+7PuNqBBh9EJ5zY7Cn
nlxiuSVbMhz4G17uNpWsv+DJBumNVkKYeEq2u/0iWlai+eQoeMi1TdIpfuq5TXuO
cFUBZDJ2DJ5SRbOAYS4R18TXXfUpm85oow4OhOqlWjbDStsfJnYJZHOoPvmhBlC+
Yctv5QFOHleh8c3wZblYmcUk1uSx2ye9+ypNlKwQxiqzdSuqAiILU6ZPyE5v/9b4
WIP3zUgAR2n3VY/ScHVZzQ6JkecUDZ8kobE30oIaezLsd/qV/odTeB+nG6sDeyof
mUTAPk54NaIuUQVVdE8GBO7duuXzp/8sptI31VvspOVU7q97G2TTzbPUT0CMmX7w
j0xpBYtaifetcsnFWx8St8gc4xVJBSv3wJvhzUp2fA5UhbhIwuwFExdKumEc7QM2
VrAGutrph1SjlZQtfmJ7WILwOEanlOrHS5BBFJl3i4iJAI1KlIkgJkBn/gtMdK7W
cDA7NnWNhibbVZfG+TtDRIvJUtHHb9rBFpfun9STMVOoxKKDNUBB/iRpzpRQ3lSa
XLuV2JD9ueD9KXJe58zNhl7IgHciP+9/PYnbb5Q0qTfBh+6sNp46M2X+tA9WsGL9
/xCvqfnU9Mn+x24XZHMeJtDbnP9aBq2wYX625lrn6scC099Q5EXPm4lTGXfR44vx
CwR8V1Nxpe1DK4BSzJzvfAY2GLc8CbFSXaxyAGwJu1JTBQoVVj7dCfwKupJBEkzx
tnuhShmgLyZHi7f+wDawqn2qjhKGDfAwnUz9psJFvg6ntSv8c+gQOSJM2MZMOJSn
KOsHojPDutVfY93rQstp43sOMCs4n9SmBuD7x8lUQ7/R1xecedX8uSQ4eYkh4lMS
9xC1dM5S8d4rdKQ8E0WVLC4xp6iuCf7Njx//L7dyiplMjXSy2wKLHURtxwbPBMVL
wv+ODxi5UlXIwCVhiQBsHqeh6qM8X48aJ9eEGbFlDYONvdbp7Xsp9uVbYhGJnKCN
8PB3dZPmlWdiMY/4C4mqu6jjXHlS3vzg8P3NaBqaP4uQZBunhn6EMw0pS1xSn2qa
EOJ+rxyNet8ZizhvSfnmmAa3Lqbc29H2Xa1nXkkdztpJ3NpsigVdQuxfyeE79T4R
ZiM7xM9AiouFgnRsxIEBR92DUiBueqEFATtpFaOsad2/jhF7D2XyiTtRFuIatKbQ
0gHVO32Iat3vN1hSmlp5pnis4mc+9QvJw9o/JmsZOiK+tI5GKh5jxc9lr1TycHAr
ueTUrAlxi0Vq9s4I7NVwjwKUEFYkeLb6oSUGclXvQGcJa4M+VtnbOCDSt5T2TjJg
VOjnuWMO112Qs/5mhtQDMBAOpEzXUTtcI4IiOxsSxE74R/ly0oZUyz7HhwB1fCAN
cx03ozTvbOTBtaTzFo5cXx1Ov2e4V0Mr77RtxtI4o015qQCPfAHUWncO0YP5RLcG
584G96LFvVJiSkBu4dsyD4DQPKXydfZ1SZpsuZqN1pY8j+mIQToh6v2p7ihKVt8Z
60ipWW4Rt1AbpI2KeZVI1jKj+b68vqrq18+Xjaq5R2/sXnEOfMs1MLK4KWUP2+Je
F+oT6b7AksbI46iwlh5tTts9hNBBnXdsjHdCLpX+SO2dh01FJ6jDVmp1CUJW4N5B
xODFTAs3QnNOZSqBNVQhK/WBnXhXTPVHohldPTp8GgKyqyXOXi2fLONdvapugMoq
qZEGWlN5e1WBG5MFGM8lZvEL2+E/cI6AK0T3nZDkW79CdNLLOvXE5K2DwFwm5Jkq
MbqeGDCBCyvSqoUVKiPeZlS4ep9Ydci+mZ4ocBNk/n/BHAcb7OW83NYZpFNirgDW
MGjShHw5+IPYZC/BhHN/u90nXaI6D05trioUTD2+uJY5bNY0yem51B7iAKyGZAPl
grgksevMIBsfIr/IXEECiofdDUAzttgz5zlf8StKmD4nA1TJbPaXjVlsZEYQdp1U
uoHLMqmiCBnCjwBIl7guMIo1K4XG0oibXyOA0u4I8otfc757SF8idSNqjUdeaAA/
y6qb71I28weJw+osswFO06LFBc41v8TPJyn+AAnSOd0CqozJBTx+73tjDNtSGGWU
Dse6XIhFSPusLQGBwE3ecpUC4F6SEq+WLXWiJj475ADdt1Fh7r9/aq826V4MTFDS
mJxd+z/r2AWYQqLRWt3s0AYkUa76bSI0NBsZaRraAyqBbl9HrCoh4haY1QZiLsrc
NtfSHSHpA1fECqQC4S1MGcwGWnMhN+8c73t7pdrOwnNVzcgGeg8jgEj1ybInQz90
7eOovTX2pKUc6mP0q5O004FN/7WBuJ3J2W8eOu0pbNzZWQ6csX/LsN2oVm3cPDEo
dS1vcRpfMN5DA+6WUKmt+m+GH26N+NzGzsY89yJWov/d1+88uxUZe9Oe1BbI0abk
sl9YOJ5w5+y2cSmyKOGsQ8GLzpzIHoFlAFQYyjOXcSqpCzFPu2aSp746XRIpEyGL
cta8wsDr6SX0VHX0rxL42ocSXzKOQbd876ORxTaN3Nc+xAR7avLMlYt4aHDmVP12
ZZlNQk37y19gk/3L7cOASzMB5hJ5GQQ0P5NVUEFbKwwON2xmQ35zb2w5QqBpvkOh
j5BtZLi27OEVQRxeNh9zQRGxsTrjakHGM0WPC/DA4fpfEuUqCKWt4upGcJUJYzhv
4qeETU4jUd5jJF6kagteUcySFIILvpq00sLGQ/j0+snT6sZtViiEdc1bCllAB8J/
XFF8K3xgxOGH7o3Qh0kZ2HgCn5avSeD5Cs9K9nBDScpRgcpxb6+gP3C/a2U1oGqH
qrirdlu7WE9lznC8a2u9U8ybDC03OQorJM0/Ycu7wmdZQTmag1DYqTUCfMPUZm65
FQs8r+o9EriSF24ifbyvF9h/lrxJcDVkXcoZcLyLpUeMZXGmcL1+efl4sBCCaMo6
VxsxK+8YyHVkuVQCHLG3EU/3kZvtlIO6s73pUzkOr/v+adlTar/BiJAEafyXgNlu
qDWg+GR47XJOiba8mAqXlUUJUtLpR94eTXgcDXeq7B902AzzgOlEMTRytsU0B9Ax
l4HBRaQMyXcvsRBgTdS7efydUhVcXp0Gs6ByeP7kjbgJYZvL1fbeNdyYHc3uHdVr
xOoIknQdx1nx3AY7dcApOgEymIy2x8pXqc6RrJ57/RDYppI50L4aT2v9okbhFrHQ
TnlzITqJcn9HqEuzL0lf7+YuzWtYLJTFuwUEPE4AgzdZETUwDqfGERlXTUAoJNkS
ewDwXNrn372FJ2HeZfASMNN+EAHiUD4+tVbB6u9P/Pje8Z3c5HlFjJ3ubFfioCiw
vOP3aMfPDfrZtNi4q5cjF45jZc33xHljQjOYeS/xpz0bMrzW5+6/jdtHU+NNsaiQ
ZRDY7m34ehmCUTwuh01fTyjpG+Hk1nJCXhFYtiHdA3PujmRIu+234HbYb8VWsasp
kNrN+/HOhridYdutVerX2kgtdokSBYdBB+hRIrYAZ3Bk23oVYeaxQ4arPQKQmian
2xdTEtyZwbsgMkmL4fnOVuRTjhlC79TiPDS7/a4TTvlYv/4ufpc0hpyKOom6T/E5
NGIiu5O3Vm0g5SlP3mzswwnNT8LkfPAC608iXQOjKAQOJfux0NIkbBJw1qW8UOmY
3Tua/RWasWnn/75RhVYzHm8A/cvFsIjfQNjMHaJ+EX6fYjeIoRETiyXr6fxsBZ/U
g64oN6pDYnXjCXdCfgwmVOHex3eGHpOfYISf/UvvkCZsEvt3Sdcc0awb2K7WvPPk
ZG14BD38R35XCliAqk4+3dn7s9z9ty5GYSDLhiW7OR4zAxlyfr0OWqogRkPxUmDr
kaHGwYaC/VqvvRUae4FAvl1gvAqeeGdXxIN3JdepnQAPZoa2U0zHEDqwhNXqyxc+
332ZwPSmwz0lAuxrVEyEsaK9zIK5YbpKqvMXy2c2g8yOv1ChdRkT7BKqg9HJWamP
TfwKA75DQQK3dLMFIAAJUBD/vz5ePa5Awup17J0PQXCsO5XHAADngez6JJhNXuVE
/S5L54Rb759hRYHHiTv9b01ALWGXmx0TerOMEa3NXc79zvZJ5lyp6ihJAj+4Ke9I
DTlbRwqNXhJn3ZXhhVja+YD0hEUskrzgwOYTqq7VuVYD9yGmfe4MmPrFxDnDmvGg
c8VYyXiSVtbtpXF0YyuJFkhstaLaZXRhh6PBavTkejRmD1aTlIt8ETQrYcfyZN+N
mmZHPmeafxukaRPM6RuEJ72YGUVj4lyI5xB4O9Fp52jMdmPG2Hsbc6EH+oRwpbPs
MsQEzc/Kuc0xwQeZjehTswkCdTYYBJq8XzkMEzOtulmYbgGKStPrXq867im3eELM
80Q3GGv3feZV6cwbDrxMFXJaSV3Rd3jaU7TqbA65EDkE9KV7Um7oZZMZOWDH3rlc
DD6flB0l+4QE+qrTVmG6wGsVtvmI8tyvLxEF3giqJyXaO+g74X0UP7Wm6YnBTqGh
800eJpfsacpETMKDNrnGdI+iMUw+e5BNQPvqbPMPJvS3VClxnsnama7dZYxlP1SL
fAfthqZDLYvust6M/aAdRhHEP6yiCVGd3xM2+9HLBhcuTs+7QR8LxCYM/3L+xpZA
35M51msIUmxj2yAyOvUKD4x16Zi+JWbG2JfDDZRJtCCSGBXP9BglvVgRvy339Sqo
GxFY30ed/l7XgjYK8eNC6mMbjrxXaF5vyrnZHD1E/H3ZeeQv3wCZ7cbKWRQoKdRT
+eIRlMd5c6y2wL/CFxfsbRAY/ki2TDcUcRFr1ta/DRZxnZ3qIJuwkgVZJviSqbR3
cXAQPawzxT8OA7gR+tbyvrBAiJN6/vBy9D9G2aAgrk9tPBSlFwbClSmrHyup1931
Vj0Rif7c+pLmOa0y8G/wx+c1b2PGTRstmZWJCLyTH3q1IF4ziKxSBgLPJ1LIpwyO
DWYVD3R6lkpfgMHIon0TG0iadHheUnoT1Xs3TM6znwG+mCIZTMTvwwABehLfFgSP
9BNUb88cP7nLIXycnw2/yFN9yl4GYgzNZPLbYQIseAszl7I55xZU8hMxVjqDTMLT
1Q/D9DTjvn5faoRdQOInVorhHSztyIJFcI4FL0cXtNq4gwcwj4PlOhUJMJ6IEv1/
ujsMUnji8ZhCRNIDjnTa6qr7+yI/Hb2x8zWzb20iCAj3raHwTRrrSZE0XKgwayv9
zz+MAKTUTxxCwBbOgjsa98uUAK6ZKTlykM7eyCfn7t0auWbT0T6Fq1s43PdPlPqf
Z7XYGSxhqGv9ZSJuijHmhpn3CLn7FpvbiP7USjuwzz69mttM3uVoCkPDwS63q0gB
wsOqBh6yr3qNHVpqffvpwW8ZO7oMf47R2hrLXI8ob5PafRsa0zsoVNGqHEqJaARB
agobMrZN6bGwN046eNutzaa5qefvva1uGcgtsVRnOVv8YptYfxKucKEFhkOj2Ulh
Zv9EZxkI3E0d3Z8wK1EGTMvKC9HlN4TkXw+YpILT1mHePPHuHtd6+u+B3oM8UAlL
33GzXpaGZL2x0fShq8FEhweTh7tyF8Jm2Sf5TfM6eX1jm2U4pJMTz77seuU9WEPq
QQdg2H4qP37sJ/av+g8MgWqQlBZ3wAxljzuCMxgW7uGBghaHKtGG7dk/TqWn9axV
xST0B/N1OAdBnm6HNQBQF+jdU/h4FWs0BEIAKw5PwFfrXO2n0YS67uCXt7DOpF72
Zg0r5Hnfag5iWozlcpq38mfFs7N52R290SBsYrfdUGfnATY7Z5+1AOvO6YR3vCEf
kiHYxDg3mqfEiP4KlU75viIQtpWl/BeNS3yusAqpQ0J96pyskmD/XOOfyFLSXa0g
PzBuAbgOzVjNVTgdPanJ3+uyCGsb/OXTJf1BCBxR4/f8bqa4TIUZp3CtLL0YRW8u
rBybdQ+kiILCr0fzVQIeI/7xNjE0/Fgolw4kPg4jscLiQ4RpvMYSlnble95HWHfc
aVNY6sZXJVcsOu0nRDuhP/qa/shFhH6ZQq5y+mO8zfvWclx7RmGh1iCs8rVbC1YP
LIrFi2A+CZUtHDTrE2U9palCJJows1Yd+zCdYXVh7YOVCKNB/fgfVJUozXzb1uLD
Im6B8sbD69WXZxLTQzfJi7D7o+10JwPs5kF9dCQxLepBhaE0U4skeGwybT/MA94v
8tZL6MSJnIkBtKr0I67TJV+vwIFdkQi6w/vG7DZ7D/z4gwXr2VXEylDQ/Xpop5RY
b3F/j7wbyMDg2JR4V8MY5X4BqdL6dUaTrkyoP4gfzYJmueuxmD55iiXrsGqdqxlK
hFNIYQbd6Ad/05+wAd8zXq4sNJOW6hoip0SHxo0Ovs+29bb+aDqLs53tA7cC7CZ1
eRWw/znEvWKeiDuDghuHj4PLkQMUd1RNDuRoQD+9MaypMxpjcPr6rswzlv2zdZMB
EJqRzIdNsANm0KLHhDl6O+M1d+MJzWncIqmYaO0rfL/nw3VbO9DWnwJGrwaNXZ4T
ookKuGnHHjNjtbKBooidjQSJqbvVh+pPBGySgEGdgK4SlZgXXA9RhOAoaOJA1ekD
vKpu6Zagol0WvdHMP+9uEu9N4ueSagUm5PJugegsJqXFcdaqYB5ro7ykwM8VupVR
5Zv6LlmptNWeukmb6bmpS2L5t47WJDYwovzK6+NyL3qBdBx4Jf9k4Xiv6xJpLYaO
cAm1xcFZ+P1/fRlF/U8XlczvZ8pjYSIk8mI06Ur51OZjQWtPUzwbnMIdUi4sR1Dv
DVQtAqL3KaTBjNbzxHdCCgTw6IsfuLvoCS1jpVAGkQfLsjUTqoFAa/cGOuDvaDAv
0buE7oqWroNfjmxmR8oX5nUBDrpO7/5tG2YBbaetq6ELuA1MxsmNJtlJIJSAKa1C
/ibXG0FIH6TM38sUuazTCsgGIGCZkdbOuE0xdCxfAKo60v0nWkGuVZzwIh30z+aS
21IXJACmocVQST2xYgtCN7VBcx656USg+FDMWM7CJs3LdjdU5xK3YB2LBDwVHVIg
ZvGvHAYh3Jf/13i1gM7i7OE/tLShGuM2YmzUWoNy+z+pmndPN9bSXCMCK835JI8W
lougaxoOXAis9UJUNNBr7hsUWHqG10Jk8zfiqG2IRQOVkt+2jK9zNLi4pbzAPDnA
3kR9CsLtYtFEdTjKemAntKKtBT3c5+nZuTRzfb9y9O4NTPpN5ERbcl1AopHG+5I/
IuMcUP3AOStR90eQsOWgccreMEmWNqw4juGcU/dITzGkfbD9ZawzWT1I/v/drH2M
6UQ5PPWytx2opJ5L6XXFS4x45HlKNwFSJpuzYENujccyQqaZ6qOYTRq3g5ZDdZZ8
f6KiudO06ihLTrD/lNzrlIYbGcLPAVq1zZqrVJlqBfcwu0Qb2ruJLOmp2WSh0eS8
8gEnz/Oyq30ozUTmxSE0L7MwQ6ZFJl3IVmnjtKZjS0KGYe/U9cbu7xbwG1oIPBnj
YbfkLkkVuxLO9/9ddBfS0+ZnUTNwQ98zx9p2n/LGhva7O0TAtYZibVVQhZALw+Gh
BpgY2CZcnnSrJhZwsbj2VPgJOmVj7Xype0Rt0vfz4Cu+ziu29thcEfQCuCcI6eHJ
dhbNDjiDNNNRP0zQHyu0E+eESRd2nSQsDxxd7Yqjv2rhU1ieSoF7gaqPBHMrd8Vp
KgScS0mm42uIkFeGNrbjT7eorsaKzV5MnpB4xuDGLCytCaCeSl7siRFe20JMutu/
utls+eOel159AzpWfyT46N1uVuT2XNeVEzVAlkiIeFdjWyAQEDIRT7tLCXNnO08q
Y55W3h1ofH33R2eZ7bQE6MWKuzHab6I+Y9raHU7/NrwxfoFJTBdV0xdpnREBrlwU
f1FucDFr29XC+p1I2UVz1Ys3m90OXUiItuLkjVyuqFlrCwnq5oX5vl6dW6HtLRM8
25q4Qr0ROKBxuA3ebMnY8N50mG68Ll66VBLFLvfsRB+qXvp+APnc+9AWUk5QsMem
VUixJQT0lWeZEIlVIuvnij/Jth17/WLWV1Y+4JGSb29TZ77SVstFi4JvoPvkC94u
r2grxSkjFzC/ooDKcaTJt6BvfJuti2I10S4vqe5vOY7GK7Ngye2Kgi8jAQEG6BMg
hhIOLjnZZvWjwU8oJIqxOZhvyCbywTocvJa4w687Il2WD29e7PgVBimFmRpzkajJ
NK2wyiGtvAjTRG+NZhJTzTxBKcrgYNKxl7zPyLwOx4927ZFVM/Kle7qSRCQdJpTz
cbgnIOqiRoSUtalFxdku8+mKdDHFwTK4H1a8AuZkqZ82NSMir+zpmA30BJXdRCOs
8G1yl6paffDSdxXENwKZandYHzwUozGOKGtclouIGrf8MZi6qakt3VNU7sgdJ1C5
R/JEQe8Zg1dKb+5GCDRGPvifZtW+McArI5x1ETlzQcpu/sDMqzHTeBmtl2x+7sY8
1Xjc18NUIaCvw8OqpaaMgKxmlNhlTS72cGpRmE4FwwR+fKLFbZbQlFI/bN5mljmH
WvRxiG8y4K9NmgLpMYn4oLYkNrx7TKZa+Hv1n/6b5eUkO0ZxzkomMNWjqaa50auv
YKjB1m0oxDPZB13o9z6ZNWUJ4WPNw52D3eDbtAq3P/Cj7ZtJOIdcdO870tRGtoO8
NL9sl5KR/u03q9dqhOZvuudERK1jS45TBCLIn6G8pazgWFjcxC04qVRKzxXw2Ukn
rygp7TK3AWtwq+LwXCriCxUV6BAEfRZc13LPvSVOGxE3Pq6BVN85mlvzMMprXlW2
FjTofyzFviptfeJB+ZiCDtGzfWdLQXby5FCHB3vIrFt2uChuZJZKY/9GFXZUiMTw
gQrfJdXdN7GszjX8FpkIkiv99frNxQy8N26VCPHnzUF2cRIUQs7fBwF49TK9UCuq
nywZ70B2QSM4nuGdyQltvrhc9oVZ3sKTN44vkTDVezlZ0VeilfceSk7z0cEzkh16
v4DRi2o1VzH7YmENZpvzhpf1IgvgeOxrn6I4kMP1mzF0yUerPioeF0iiuwm67J8c
kpZ4YgIr8rnxW/g7Q/NPdiIYvmen3MZe9HzbnFar8rY9vSYWbW32bgxtHGZZhAKI
T6tVWjGsEgdImPKjaOwBNa5zBFwUzkaPj357XaEZeKS3kkRAZ1A4Y0aCenpsL/VE
6uI3eJcb6P45gat1wtKyhMfH0yAN1ef+8eWvOLnE2/mTSayuYoYizSLeJbtU4a+m
11eqspqQRbFTlgx5mrNWSrBA7VijJwnq6QLT6wOCbDjV44fXUtQpQ1skCjyWhlif
ZaoOI0n4T1gxYW+XSZ/0bLif3cjfPie8P69r7KkWS5VBSTdbug0mkpYYI8fb3Ity
pKkOwzPHqCgI38k2q4NrJXloKpLpWuL4O1rNIyQcOrDLrowwUNeK1R4rM0S4Ha56
GY/jYsvYIDGKTdODOh/sfivPuSPZz27Iz3edaayyOB4vAFUoGVLgFeP5MzVjH/h2
VSj/ObBoJ5z/Ov34YT3Y8BmDR9kRr8RgIHVgwL4wlg4IgVtIZAP9SnXWYgyDx2Z4
2qbJEjWn1KkXDZ26ZPr29xCrS1nL1xcVSgnttP8l2bnC+0y93onnkiKzX99DLDG9
RbfFFT/PL007WSilHfc458G3JCMcOHO23TdMZFnhg9K+JJ7w0WSbWJ/e/shdoBhG
3naJ98/+Q8GApat6uTSMjg5uFXRQORX2wcEXXBTWo5feHsac1LfFIr0uvtpYRrcO
/5NTeOzCJaOv4RlWevFY4pMipDrQxngx9HRiS7Ymq9JRWE5GZAcfgneGQQDgN0+O
NZH/lj2AVvSjnkW/JIDLtHw5SnfGIddfqbU9VO9XcKcD2f5N9VXZkce/OlwY4tTW
vcXqUG5cygeYks57HSNpp0QJTCTIJccAgmlQjgBHTlg5POqbwS9gmRV+073KTb97
8PKMw2hw5HHXxfrNNLjkRwu1Ownd+eBLMUHGO3mHPwG1qCa+J19KL+Gm/jl/Cry0
tHNLcZ5QgmMTfF7sROJhNpXJiOFLXHbGK7YS8jHKkulKxaz0ssL48xc8imPeAzjn
bp+KPfAM54uFf4qDi+fIv4C2FxO9vp1anZ7p0Jd9+vQ5JLs2Q4cS8iejf+F5vqah
hn+oqp4iExIIY5cd/VLJDE14Ebxapf2vZiou3kJPq7oDTsvHbf9Jd90qAoT50A6a
zFVJLUUMk1E+Deu9JTHsqqbpgfUQGqnwbIEbL7euAuV8lJGxeG2yFsRxwFQCuLC/
I0QnFo+FF9mc7YWSg5HikSZMOw0EeUS9gTvMUkAl6q2hlCNIrUstsyPsljnJzvHp
JU/IvEcOmBzgzxOH+MDL8H8hLRcSBUYhMkwP1mrpkreFs47xvIATATXRcDiT3ZjA
4Mrg9h18AynYQ6qVICtistqXTTcNYpg7EiAqj1x2dBET59H3+q8G8qkwoTOmiZ0s
pZ0b0MKajEO/ns8noAc9g0aEFYV+ZHURAGUo2u5D6h8WGfPpfa7aCByDc4oSaXiB
sT3wW8FdfnbEy2LZpSecuI7bwDpoRvD7r4WJ2Kog5nN5j5Rr+pchOzwazCSxcFgH
pyhvhOVbvi3NGQ74yjFMS2zMHTTUReRDK2WjScPyb18zaknK2tLhNRvf4wgWJOqV
XwZYqSRH7XrDtoJxxdJu2B7ZL0YuunIYgC2+fs94Upl0z/KHL4yoNXTYh4BUaT3l
4UUqoQU2Qi8eacVSzctb+AFBG7aK3XJ5W7kTjz+7NchWMmvXwiNd6dWVq01MLakf
bvAB/aeMVay+xX4PYQSD3uASlUMHQml2vVAfS+d3puaA9FESCJO92bp6Yg46o3ME
euumIOj2GTjWMCxiUZBH1fKvw07VGL7hk8yKdBIYZHNmQ9J4LxbuWjCJ6RQ71Atp
FQtU69Ma81Cs5ZDbhP9l3vOd8Wc1OnkJOntZfYkK3x/yodVlzjUsoyIRBHE+LYsN
EZ47nabG4VnOPa2/UEIDc13vnpXjkCf7YfWx9RnvkG1WhVxRNV3rP33P0zHQakoM
5uiDb6qrxXHI5uyqXPh7G5gRazYJAZrarODmnEkGEexWNQjOsMfURP8PPpRwpT9z
2QnDZVTv1PUus8IwWvaFM7FUbE7CcxTWql1sBdLShjsEiJDV9XzifGRV0cMbdqSv
71gu4ErElA+9pJpAatyuLN/InPX2NzLHSBduCysrOMvvu7PQznU//bA0zw5z7zCS
WriwOglgmYWe7NErN9GexfelwoIqiC/Qn8AmZGn06G5GBj3JCELh1A+i4Tglluy8
zIYmEnisLCMjnDXR1OuyvghwvbWurH/yYnY9I9mLXt6nKUq90ATXP70XN2LGhAfn
0S7ui/xhOFaaAJxLLK6UZCxHoJUEoEMO6Y2dKbZoGWUsc+OJKg2V9/K+6Ut77/7C
DwQU/5vyT3LiYl8Dptf2Aym2MUF7ZoeenQ2sLpdZ0GHU2z9cnoGM5PgzYfXQe9H5
5lXl9lrIBF5k4bft9F8WwB+23k0f/Z/Eh+VWwBnBJ2E3yHC2HY+k8WWpyWAqrYVX
zW07aU3GO/HSeve83q4OKlkGrccDUGNSU/WqIdb7YT0aMvW9m4Q6nWWC4NrI38l0
Q7qqSf5rnRnryyFrI8an//O3qBvGUr7FSlL5SJOgL9aB9oMYa8HRy7gsXMGCwUc+
yFdt4ao63XMeWrZfYricDgv5EEzocezL1RtulBmUP40gXXMDv/On1DNMgrg+DYw5
3AnrZarMgBW+xOn1JBUm+fuPnnjJcaKqnn/Fvo69Jr/U3EAvuWKv3L7h+imzxSBI
nho1WIf01IGJmXm6exBnLD+zcgZkd5UPgG+6Mf+zUDcndfUJ6RecRtPEQrmr9SMe
vI2zvWvYDtMHQeknLdZkJzU/K+I5W1kCi85zmF/WHyevipub6ADWneRXWLdeYKgR
U/uaGCubfpd20keYz7ShssrIGDlCnfSucO40qaHRK5UAOh4ALpYfT0M+rzOD9//j
ZWwCk4KKilag62KlKHlM6y89pX1C+ySGqb2VuWfDgdj9yOZH3ghimWSGLsCwnKAd
IEOXB0tXaTtVIZvbfgZbSaFnzk7K+DBUbSUZ66lvrB5HpS7NCIIeIdx939SSn9JB
jODwu5oP/7hZOlISqKrBttuwPXxfEyY/YX1hq2+ajJBKzPw7FzDlbDv6CN8C7cf/
cGsNdkKkxvRWwPPt9mRY8lnoUrVYeLPicHROS3mizh/Y5G+KyRTfeRDAua2gm3ZX
rMLfkQHgPwKBhjGuVC6540NHPJioA1Lx1czJdsaXCF3SABnIZJSIcP0wkJpkLX6N
uDcFRKF8MwpCHJR5cbZEUifZ40SVSAYxE3tMy+249jx4JaqT0ZjzRvl5XRLA+zhV
v+ewTueWOD9eQP7L8Q9gL+JX7PZW7Ykb251OfwE6kPtwQcd2oNzSbxTaXt8Tpw7M
R0vOq4Wdl4eXSKLtvSRDlsZ4gdS05h91n9qA6XVmgYmni+O75uuOIMKBgiWHwmwR
UUdyDZhrNiLjrp6l2rGVjWInDeEW/UNwa2i5qjqzFqEk8QkJ+3yP3n7bC3cQnH9x
kzFlr1Uu4B4sQRLVIqfDnAjqkCk1UgdUCl0T52CQZ2ug+qMd72j2acEw/kHLHTr1
MuMeIuGH2xMb9ctS8ngLdH/zXg9DQrno56StpeePaZl0hKh8/qsHcKLNYBAdrZcj
8jaRIMJrU/GNERJJwsYWdwEWqkaVtEsa6P3jgZqTgdG/YgagXZK/o1BP+hwHQaB4
xps0los5NdH/kHKwjfe2spLbVt59J1wP0kRlViPSX/328QdYV+m6uCOk8FlMtGE3
nV2F1IeG4kzC8jx8ZT4cKLg7GyGaS4zMpF5jQW9bjocdNwgnWhzgeMANzlcqBOCy
YQGkswU8TpyAlWhunLm5st9HfIBbdPnnF+uM3xL1XQKDO4Jpvt4+HKuo4zUFbgcC
gtYCnwJoFORcq6FGBGqtDez+Q6MC2LzUgNkDS2/2Hhql/yAQt7FJaOeLrSP76pJ+
LDxmtfGhcQbnG6h6gQ+R+hIf2r9JXksYeFTkZFethtxC7esvuo2/cfpoQdK5TAfS
gmczkRkAhz3MD622XCR3myKeo1B4MwXEfKazOxoPeG5ZeQPPRbjz/JJQky/OErwR
eSlij/dESkey5RKjzLF+9pYspWV7jGoZ0/iEyc4guXe7vmBktsWNWEvMeTDRB2fx
N9QUGyp9UPSdkI3yMu/B/fDoR+/v4zkzjLKUFevSLQ9UP9bp8QGCfoA4zEBBwL93
99h8EuMgBz/qg+w07UTpYDht96U4Q/+zjMwNAQLe4oNG7c12QSx1KuzmnSSaHvPA
wJUHpczTuCaZvYtZU1cYLdyWDl/eCBjdZ/09vkhcDHi5c+Br6u7NMDRPutbZN3cC
PwmKj8pw3nVx+FB410ecw2KmOyZkghXlijEVqv3yPZfAnd/Leu1Tw231BUUJFEsB
cs/Skpi6R31HswwW9QmERowlHyuolNZW50f/vrxTqOufvZC4lBIlxNli/ykPcb9N
WwWVN+pZu/jxq5BGwIAF98/Gzsjfg4vJjP8zFPvP1hkH+Ijze8R4bKVQm375KWrF
DaPj7U+GZpqAnY95PM2f7CuuUYSR8CqOIHPPZL5Jn+6wRbwMpDgwyypisoeUU5cE
+Yn8olpu/qRqO/LVPdvJduTTpUZW+KUe3t1U6fmgi/7v357ALmykfKIgozn2pVCq
tOLL7FRQXWZVSg8nK6AVeA3yy4U3+QWv5kgBizRN6u5G4Srvdhi5JLdY00917FGl
kTSBp6HpoiOzFCCok1r0SMoTnqap26OvQ50yQbdNLe0OYGshuIUS5s5GIXEHLSME
BO8NJQVFejL/wFLSqYoubuDxajrpZ6VtGDYlO8XaiZb9MezHOKiXqSAw0tP7acAp
D/MwOBtTOo1dunn7DCvKt1ZjdyMT/Sbr6Ja+UHl9lTjYjxW6VpxnBSaHkBqwWJN3
A2R9lyaqO1wscq+hV5KoXFWQ1ZwfE9TBopuksj5QE8/GCPpejNQXdIm/x2g4tQzE
ZzgZWhizqC4TPKGzgpdgp1uHJymNVhLpAZ4vw7gsLUovMbHnHCNNKwXuYYqG+C5M
mlmSBuCa0yAKTmfCYszKpMCxSTftDO9vo1+f3ram8gCDvRy+4hpMi2SaVHNuRHrb
n8BqXMYsb6d3lBa5T8c0mM5f4GEjSSAHC9uy1PEmykOr0C/jM0PqD9/dIS0qF3xb
g1Ooip60YCG8rCYivXCX/l6NL+rMJl2qB7PyzB5aLL+jftlTr3k0mvwnaxyN6ONh
7/nqE9hNwIFK0mRqNdKiuG0aMCKL8xU/EXJn1Bo4iGF2Bi0lhwwy6/EeW3ZWtjEC
vNo5AFh86xJVFS6l4cuFatWTn9jymFfDbzG1rLUSzuTVv4/0PIJiAzcBc1nLVXXH
2/V+yk6AsihxG9/0dbAE44oWEGUlsckf9EYXWHyKxZ4Y+qMjKs2/1YuUC8n8+DVe
en6pr5RnrM5AWypBklO3aXm2WV+q+M6fMnMHWT5VpDtQKoNNB62+6s25YFe+v21Z
YP7mEzpjZR4dLhnadVfkKO/scHMZWlPF444R5Hsa1OpMdIMsX3gYGKHF3qJbPhW1
auhx1q9sKuN7VIPAo25FSXeUiQg5wRbjNvFiuzORnArPVpG6BI64x7boo8S3Tgj2
Tz285VE03K9ETxtHC8o+SEU3j1OAbc5WdmMbn2MqRG+CKKuQrKuBACsPpWFEPUN7
DYQ5dOSZB0GYJDKYiakQNQk2dah3nGEKajMj0wdH7gSUzjyLCK+jCksh2YfIKhO+
lBX56EreTrenwPVQSE1htFDtiv3C63euBobQ1vbvILo/8CSukrgJpFak1GboDPze
HiOrv9oF/UaDXap0Oaz3ZCnLJMQWwctwwTtaojU+V5nGE1zgkti+8BQ6XqY+tRe9
8fjYcBFiGu2PkykrglSnjyQuIBJ9NvB2lmNfyADCPuoIxMwNrl2llrH1bcK6wquY
mQJCquClSDW7TOIvtapvxtBRJNFvpm0PQeWKSfJpJI37VwV0bdc5Vm68wkKGkOKX
XJg/dKWQV0apUt0uzRT95+1ya5W6xu+Y5CNhCBHiNMDdSKhATBb2tE3wZxT27gD3
iWCwk6nhHp9KX0p3ZAb4dv3Fq5WwEuLjDvXZFkhR2s/dP4qbV70AH9olTGH9A8Cy
a4TfX1emYm5AzHplNKZtkTVHXwkiWqMrv9s5c442hYkLV3tWMYQr5e114bI+2Ewk
7TJKt4daVWpMEc3877F6ju3y2n0DNN+/rxWgR4msPJbnKTURBNnejd1r9R/48/sD
4MbDR+IWQfXqOWDOef8fNK9vCVPefnaYimM9YaO5xyhC0LbnSsjIxIzA8vIVOA0/
HBm4F9VhhcIrPVadQGfHqN9XuY4mM7Fh2Rz0iAkmU8g0VkmEYzC+JBAt9nAj/ad3
dbi2F11F8Br9/FuvlNqMQImlVSzaqdkH7jAVBQl7YfhYNAK/U/bpMKXdMYBOIizr
tSNPREzrnoKXv54MjSvH0TmJDvdGi4X/ZVaYlgYeCLoXb08JeJpHxVgYSAeghIGA
WSsjbp8PUFnoIbwJn5QnYTKqQxLhyKjTungDccrxVvkp5SAKcFrwD2vclF0PlG+q
luLZ0CXNJePnagvyY2zcSPe6dOhVeB4qLmDMbLBwaKsqER+zlIqLM8+zEoe5s/Im
DF7jZGOnLp8zYHCL51tmPXly/sH8+nqTnkoHsEjyvZg2+iDCfWEZMkBMmEUxHnBa
LJ7c2A6kXs39z1sLZSfu23WbfOmAGupLpN/BkF6Dp/9jG2gCcTrQWSGOK0B8eUdQ
wtD+avZ2Jo6NHgHIA2ARvmhK+S47DoRkqSFZgbYWCh/izBMmvZLFCtXKgRHFlzMX
LbGm1mVWunhaAknM/jXB0MCHsSgq4AjZo+PzoQO6dDNQrsF2wXcGjZbm5foMJRCB
prbXdGOZoXhEs5Hqi/pKfnHOO7MVe+4cgvxNRwpDFibx9XCypJSIn58LBRWJaHDi
lvdPtes23paDv3qzzNwZmFzpOvHMbmypwwwZGABXcgYAlBdmprpPFvMBwAAa/KNJ
XYrNqW0ulVgAiUopnFR+jI3FSR6jOlQmnW1ko237Yn5B03VxMi5x0uxb6nsJxF4H
pYdhTfGAZl8arQK1dKPvgN09StH5RrodD2UnD76QrxnNOAZo051aUOzgcQ20JV6I
OeHO+LVlL/uaDfz22r8hlIn4axpoyOfa7ilFegXNTwDYLA4NsJV09jxV6Q58GNBF
/PQmwDheWujZvyrnER+JylIZXZiJ8g+yAgLHliSTHYuTID7Z1PgkJ2gVakzbdV0n
Doa+/49iiZN+23rjWhCiJuRhI3MK9eNg3pt+8BJEcDmVdW6GrlQJ8rBsxOI8rL3m
fcUDxcFtLZQsvWIr0XvdNvly6yMysj2tNmfQthoc0HUtMq+KGRz7qTjyfFGWdekm
WxXlzojHof6wI6xN1Yw7oshK+gu1BSothkxNjkqieCpjBYcGjRxDlxn2mC8V3wV5
+uAWyhWbuBWD3VagiG5kKjeA2Qf5r2Mw7qgMAWHQ2OL17606OJiI4ZFlYpmrY71P
TYQcK2m5Wc7AsUmOC4u3Y2TdSa1kWBanVu7DiYB5KoDlLFp4JiomF5jZ0iYlYU3E
My3rmlhAZc7J3uB+2SPkj4l5nGCEb9T1D5CqOi3SwsO3H/cAoubBNrUeDuQM0H1C
4jxBxYmUtpqk0NaogaulsOBm7TgyFrfBMqyAgHwvlMgJ8QMJpUmi9UmTdQGblEFR
vIo+uKDE5CVthR0M6SSEeiN+8pP5Ulg1yRV6ZJ1daMmvXB5xUb4VgnnMTLRozTY9
lXUndjF0CI8Ocik0YURtRnXrfXEdUFHmQOLgepUOa4LnJxkRGtPNqCDI6YRaTqTz
FFGhkgnDGOX1ZYXkj8pRPq89zBw9yi3cnsqSP9Mxdv7u8H3dZm1IIKvsqUtYG4Ti
unhM0asRDLm9756rcOKYTUgaGnRAS8JEEvhzUEj2usqIjs/fxTc5a21Kvp72H3bv
4IxBOQRRLWQx9W6b8QjkYEMGElnbYELRcmWIf1PhBUgAzzLpJrk48OQQmJJA1Xrm
MjnWZzJ0P7cBVBTdMHftm2SZz998kU1AHLiE3LD/AeqZdcPPRYME/2L8FpnMyxHW
Ck+oLPtSqoYmnmOeJODkNT9aTvTJvyDF9UGuf/aDdSWLRJBKfG1Dp5iRfbPENyXh
EJ1vO+A09xCIRgliWediTi9egxdl1kdTuWAfLyZ9xNLHZXm4OnY0SFeep5zO5AZy
d77lypR3b5oLtnuQVCr1au1PAIiGheZAyx2rN0ldM/MAvC5RftXNV9fkj1rMlzQn
2rbm0RwoYDTM1WQ+unKOMJUpafhh/EZbInBxteu+VAb5VW+IV+4HMGmBnbrFPP7t
KZGQxBGDYJodxrrTXfy6YNEoxjXS8vqUMjKPHlGGgJ3D2evi0a4OY9SRvlJS7NBj
2kQhXFtXETDvcCCSlefBLBhMD2NpQbo+jUNXIG3/dIzLq53MOBbfZ2wxdY2lBajn
DSRQ41Pg3EmDuOuphWICIaq3LCpnci4SgAi0JlwVQ7swam2VIjnIYeZjX/kuwk9K
d9hFf8YKSC7iqbozU0SEPB7sMJ+lDxlE7CLszS5bfzWzFReOCr0JkGy8bsYiSe5c
PLZyYRnnPCoMXBE6Y1POOq9bx+Tko/iea91zkXNUfsWE00DirrknFr6sJeCvPLHZ
UAGcVWGSnP1xskghbqzSqnvxcslXsMaQ+MaJN7k8AZ+RGpQqgKV444e/WN+//BTH
IblsmFMNboyNQq4b1R3cFuNj7bpdtGc8ZQuDNaHHkWFJc3CAr2SuAm+EcRRyTWbf
K3L9rBO1zF+EjQLCUPCf1JGIQ/Kc3+WtxZcQtoD8IxHKMPDAHxmdSIoiZr3jngFG
yMFZe/OScIcGAI+kWDtPoNBPwyEaULPvsxpmtt1ofhRw+cOn+zJLoDUFI7gD/DVk
JtuSpBA4g4B74I5+fvR+2qVZtI6G9L6eGQD5/Y1UiwPhalzKig5xMlXJoNX3hMS8
AOXTH13tAqvIWETHV3A/ZFm+49BJnAG0kL2XQHXbqj+yzmWrMe8dXtTdhMMLkDlb
8Jc24JuaSEgJb11CTTDOGWZn29mpcpq22P97usJ+3jnvCoEc1VvmSd7017/Y745n
22iMKjA9gmdd7KEIf0mJdEiKMWGpkv8BdN7h215Mi4EYWkRNWuBIDgXombpvr+Oz
y+XUugdCqd6yzfNolb9kqvCg9Ofa0F15adVd8cpDn0ITubOm/B+Ss6ysIz0xHISH
FEsDDjKLYtgrWaC+NQi/6wXOcs1Tu/Ef06iSLwxZ9rM0mFbVAnyGTE2uy/MGrLf8
Gw8+J5a6KlSK9PgwfqWZyrt3vYBtpE3eeLKkqx+yLQw9C28pbACuAa2bhN4P2WtS
zrcJuemhD4nhh8+cZzWqBRXBlPfFWSbSjsK8c5puZqh0vdb9QwVTQZah91IpNEbF
GPuK3fcgbEDe2O0PA8zIglZ+N2FMJqTNWAOXLZ/ph6rRiPLlGKgunIqzysewESLK
CBBXjDghbJ2x0d8SUBYa6QHfCI00k2viRc6PL66Xz9uyUE6zeYnazWOfJY8hw+eq
ADMO6as0QV5EVsnRoecfW4g2XmJtnXSv9ThAgtQ/5+HQNM+ShATRjPYLQnsxTMZ3
x2MwrfuLpTnNXTTvolyU53dK7Joazi8crOWxBJ0Cu8kV+mUqUti5LeR5UHhtYg5F
EQBOJ+uii36cUwknemJueuAmovlqDTY0DFqWglOhSMP9nyoFmCTT0HBWM22ALk9F
a9IV4j3B8OG5RTVjhxrjW5Mz4iUV+I4SvfshBL3MMWfYhTLcjtolC1vpCgTWX3S3
/wK9sEVncdIStP+UWpsNVfukD6wHf6lKWSj8q7Rr+MQ5xK9pGLjiOD7Ltaw5/cLj
uLEjVEwej11HtvjwT4MfKdju5IJRjYLGMG6I4M8hwUkxajRO+WBmtpkVUhpRNpvI
wWUGlleMNCh35s8r1dI7YwWP7X+3/K0l1X/v0PEiTpl/0c4VwDxbNqPhCJd9Mj0E
QUA2SfnM76NZEfBZ/HoNJGkUFDyGnkD/Z+CAbGnNkh7pjT9oC0b8cZS2yuVewGlc
pQE1qs9D8hN5r3kw66SsphfnSXkruLZ4MRfHQwTUyBCo3/JiFHsHWXjjS/h6wx6x
WitVmpvi01qLU190PHwbQ1tES8mjDCwUHv1hx2L1afzW05kUXT07LuLhGgiJIZBu
XtZjj0wSkrM5nN0VSE6M9vBS2Q0mZU+HmWaYH7HA6R1TRcUYsASfdYF5GMwhpr6w
+ZZeYnn/quouYLuqj5OIBufwXM4BDmN37vhv+B8es3MH9xkBDcdSykjZGDZic8rW
l3P9uwhW8whWw9zwOxCzwx5EreOf0CadAEhRNfhRYKQy1ZO7/RBoo5WilH+AksTs
SsLExyGbk56HZ5EorSp7XA45cvf7e5B5XCW3gktl5/Y3Fk0Y0Wh1mFFmoQ8FBQJp
edGClbrOfOwFG0Sis3yTVojH99uUMNbGcJEJobaupW1k26r/ZlyqGG0eTuXuPCdN
tINKv8gWIoVWISlEd7T0b8mw0U1TI7ouLPMnylFVsXYG0yRGo7haUxA592eaxbpJ
9yLN91bueg495vK8mjUDOpnCqJpYxVfjkivRuIUSVZlJMh9KlwuYm4MqbTY97vZ4
ALa44GMtHgPEbbog/B/jhQeWUnqorV1a74gAj/RlLREKkDHwVceAVKYU6s57GRIG
KeYDR2W7pyaFiOcLL4O4xTlocEtv28j3ZJ5Q2lCUb2MMzMb4UWngyMkywg/EhA1+
nNUsPA7hQex9iJ+26p+8MaFKf8BEiK7+B9766BaZTmPOHJsHm9LfWAGqUv8NS2gR
K9NVpj6pGzwI6sV9NZXn3JQQgmF9aWhxjG20QTNy3UrAVroAEBqeCj8OdNEr+Edp
MNdNDssGfAWoSeFwM2tFikko7pvHhWK/eQRlD+NOAMbv6DvZvZZjBQgu4gjAUMZZ
NyLB4sv3A+gPLUeM2GLohJSdTkvb2jyIJLYbQUu/AEsHAxXbeIqoFV+GOdEFOKDK
xHfgLJ8uwvJe40mI/n+FBbVv8c18TBuf4YJC1C767b5SUT9Mwf4eJxTRAqFUDPwW
OwyqoT8dyAxFVkj4/TllxQ/xSeAq7YZ33dkghzX1VZtmJ668BasqjCiOIq0qBATo
q/nQib8DILhpRuAwpQ6OuIFRqS7tpgl4Giq0+mCbMa/zrKSZpJ3Hjo+AHIMXdoA6
lAWsz2/YBfrI8GkDuhKZ5ZGV5tto2iCfmkvpW4U/RpBql8ybwNpN2eat+eKQgE74
pxbstWo58E+WDbdrJJ8hc8Oz+qfiISSSQpOoywcERXIfuslEU4c/j6SvLQw9pJSi
czlFi4qbDNCKpQGYcbpTARUvwwER8GoTnJJjfWEl8eSstbF5M59suZqQRyPQCPjv
/wFZDTk2n0wgnvPuYRI7+EyH6RQM1I24eS2ucL+rhrAfZticj1yp+vV1IhToiGeX
LSsItt8ywQTW/TY9Tr2aU7ANJlrbo7WUyuyhITOuNY1BXQQ2n31wxYTE7iRdXp1T
EHfIDfrZfG0IBbAtCF/VYnY5DrTm19lkFnCC1fQgreCb52PRrHGxWSFw41dbdwzt
LdbLQxiK9rBX1DXPTcw3w6w0c1Fm0bK11BV7Mp7CEebkMY24Q41XQFWBTquQY7SV
/BOyB1DVRtRmBfqZnrmFQMi6dNX3/AvyLcoFl+aBuuAzjsBSXQc85lf2CcdBnXAH
xTK3/+hxmvcFym/LUrRnKduVPK4KWB91Zp+dQHCWi7oUzcPviTChvpYYVmH0OzLJ
zp+VNegSlFQelIjf+oaYtRr0HGJ/sLfEJTTm2R3pK42feRLqNlUyWRemrUtAfXIL
VLqNngvJO0l3epSNBiTI1mfYejwKDNIQTiyJI/TlDU0KGmLqtKXzemVp5jaRA+XB
JGKb77hxMYBBRLLOn4Jtg2kdeXlE58/18tNBFEdIKumzqIVPYs4m0D2Ets8pD4tr
P1h48qeAi93YoNyZzdm3UXXy2Mhz/kRutOvrX8VwbNc9CQcX+yr4xMQUHrjNHyQT
0Y9cId8+/6qEvjHPSVs6eShNedPb0GBfEz0eFPtctCwoPi9oate6zZvYEw2BQY5d
tWnUc8/VKBghzrV1FDM/uT2Mc59efNY+Cpk8uwRIcdAxka7VcRnjxwqlQWYSMBx0
tMF4pE6p3Ynezt8yoiBvNX2nlO1RjpWByvnSAUOJYL2Lg3+410S7mRaUY0+y7jNd
cnHdLXj+7tidyw1jP4JXLabdn2Ie0tUh9Zlux/WbDbr94YQ12ok0PEARsMhfR2ab
Hs7MaCm5myaOyizsfJc0BjoEIGbDKkWX5E8+X8f4UIl/TXvBxekvAaknA/nxvhsF
SN4QbCmSvbQlsSxfpCS7Q0AOl7nwAzgGOS71B9yXPyNzHrhGZ+KmEVLpCEybZkMm
Sr4yYtHX6E5sTGp76LcQYzOgJqM7d95EYRa0rM/yIXnq6IQNmNpTZJXv7P1BM3PD
f7avJJPTm7w12x2VObCsisqiBSWPpAvijaj6G+k0oAkI/deZBLXKcKP50bMGXeKg
xBipJHYMppiEHq3/dpa03tDbTm7RnwmX0CNs+lk8IybyqAStniZbCGqHIWaFfvdi
TXPMsICKTJoQN4V35fTP70wYJHUiu6gXyrWXLCMDxRYp0hR8J+EZL3i8DT0AhlZo
/4jC1lY1vuss6xrosIbCEW0JaYbLmwg78x2fb2p3Ebns2HPMVOOwvkuEo9oCo938
sQNTXGmrpK8ztFteMfSsaFFD/0IYnzcdbfFTaOE9o52qf/niquOoWc1p9Xf8IX/r
DIY/2q0Y21TTg/mD/eZirrDAw35ayotblbyjWNTXLbTvQFiN5Y47eXuG5GW/IWia
jKF2vmlVfJjm1KLXedWvpZQZBjCbgoZPVF1ITXEBksNw8cT+GMGcg8GASD4cInW1
SbgoohueEwxIRgxxHBNgpFUcsrEBbM5m7oGCyXbNlziN6o5Ajxapv7t7HF+rk/aC
B0LBU80SNtlWhrHP3n6koky8PvHCNpGK8GbAFGWl85kkmofbpeODfQAudtzHr3BU
152lT57ag0dIgtEVll/YUu/Mg5fXir+V3qnscRBpc3IzQpLBdINqB9kqqgShu9M7
0jpiEnsG8QgOygl8U2tfvvy87A5i2DcO6VN1/qnmFR8/4lxyrUiziJG8hXcn+EWc
weVBbJP/Ys4rMvaVCAvESRodfQDxZ0PtdLX/VFObLtZNQjR8fqQlT3+CW3x2DD1o
Y53auKiv6TyqYU9GjSD0KAwmkT93Yn6QOB2s3P6efu3000xy1IckLwkBFdEcUzYc
9QVjwcCZ66cgmJVw2KNGZpZvqtMs36CCvIX6MQPa8GmfYBVB2cocZbXmm1mxDaZP
+Xsrn2i2Kh81J417APerDO4IGDaAWHLiEKMl6hMoxagi6avfIWIZhVnNdCzS9zRH
Obz+3vUDYW9ySjug0dnnHyfrXaIAzU45E8638psNCe0lhPllGOBDBq2z0CXXq2ub
TYP9TOeR0QEdzjk4aqswO72NT6M+yE7tKbHdLIapcFiHjD0h3p4MU2MrqkjZHMXf
piOFkptewuBR8glYjbRYqjItYrtOttlF7Lozn1Ch1c/k0NnAgjq1MOQMv3dcuKCJ
A74kocQ01EAiugBDfwPExo5d0aXFsayH1LS5Vmib2TWjVxoJsVe0+ANN8VkspMSj
iTX8G2N/A3pi8a0gHzcX/KPryHWdc3CZjdbtNbuTr2YxmfBxwAcXfxsCxS+Og+Dl
CR1K/VqNIHw7NnT2T2D4sSTPVhJ5gJP1MEkos5bPA79ZydsxWX8Z79ECepmyJITw
7M274O3FTeNlPGnUbVziyDLWwYGpnjHeOdGqET0Al3a9NmbrTWndOcs3HqceVEU1
zaZHtDLgwzMwcs1sP6poO46o3CJe1besy60E/xgLY0MGhCah7X78qtD+pv4OsnPj
MUjO+Ko5ehr/00ReVbXUovEtG5IZTIJyj4e6AjQznQDD9FfkrPfa0rOy7I+MJpIP
JlQvCyF+iMXmQAQIk2ljbxGN7q4v+71k6xvXV3gMGRvmafBB9hB4Zv1CgCMpTO8j
6TL58/6PdFfkEWiiVOOqxMhmw9WX3w2wygS2ciZrMpwnVAMoAWOmn5y2Ui7QXn7B
50KwFIlILDj+A6Pz9muoN09MW5kOeIM5pqhFl/JkJ62fXzzxCbuc+BnkzFOx5V21
uyF9Pj+3fmXzHua8HDoCcDTlx3p8zmRRea39ZnD4sD0Sr/A4SgGkMchRUXuklhTn
6EYat12m62ScxQIp0onpZv9sSwbxcJwEZFr3KvVklljoXE73UB26aPpArMaSWpFR
EZgp9zlAk/v1BJ0LRejOD5YB8kzmYK7DuLa2v9y+AP0xZTkOPdFwyITXZhT3UDaQ
tlPjWvhw2Rvtj8nidPc5stluf7A955a6mtf/TomBPSxJgx0lBcKJbTSd3spuL32A
Ybkjv8yW3DQ+2d9UfQxSGiSRFw25fHfJa7gVMSW9rqHnPQBOpKNakaWwql2tlc7b
IePBGQkUQSP8S3rsxZSWhMRXddUaGtmfcse3aiqfGld8SWHTuA0iRv8Bt5ktPHEx
6V1Hg59j/5SMimBdvMz7e6NehHB+KSknwI4xwCNswulyXpLMb0OHHgMieooBmgkY
i0k6CZCwQUBLZeuRvFC+0rjUdMF3jq/VVx+sFQFsABbNDoC/tqR6JTG11oBIX5Ho
gY9Ki6MuOT8oO/i583NMZOGJ3AsSXtPHkMuCyiuUTo8Sbk1soQMAOuWpmOAuLDJf
v2uywcxg7IeobTCUT/twVNAHpIruY4b1qp6Jo6abJhQjNImzl8AFZHz4+rleTnUW
JAPjtvHg/hQ+optwHjn0RHq6rfDoHw0i0iSweVddsbPH2l0NFbfqQXj1Mfg2gjYs
/he2SMJ/pzcOcJEsamk4ENOXrPl26nmfIsmo/jSGWfCiW0sm8/VzAcV/4t5PuBN3
zVX6HMj/Yk839C9VQgGb1ZjDXKmS3oa146tDdto8ROK1a4p1AVUxNFN8UwUaQfbP
JAnzQdkIIbucj66TBg6l3eGlJL/+ZkXDEWTuPWTxeMD7meufQ6hvTw4+hmN64oyg
2llU3r1/W0R5paEkRbKQRow3b7jHyu8eHJmjYFz5NkgSsLKBiACCakhWoSYcDSe0
nVyaruzClh6l9VL+fXgMlg1PDgwH9AxGdQwWU5lereF7+KZdgBXh4MjdBKu4F77m
wMr6Wjc2V6VA1ivOD8CwAjaSE064DUUvdbIt2GOS12h4TrAs8APuj6wG5HJZIbtK
BmI7qI/q6rKuP1PzfKngzvx7fihiJJGSr2Ib+t66QU8iaMDYhxFZVpgN5qTwRKqG
nQuY9BS4Vg1TGRrjwE8ZcYqn6min4Rpl7NdYH+ye/406S9f1riDgtOQ2ot9+4UVq
OHsewOnEbhP2awPEDtwJSX+2B/hy+nOQOc6wZaCMShl+/GNMYczsR7DdjZ3mnZDm
KUGbfCTggSpdw9RNvFCb4JY3NJ6V9TY7jyTk8sCgBnoH+lhsCMMWBs2egC8+TlhF
WBA62MItCHa+QKVbOIsBo7tVhuDck2LthXdVaBpnp8XSRLiVLXN+k44d3XQ7GrOW
jgYVADjLhcmKBFXJ0ufdjeeW/LwGAEGkN/rqqLqD7Oatq6Jeghyi5/WbOtmW0vaV
E96ce5wh5xqfD3wiGYPySo0BoMSOmBrhWut3oSrDQovvBB9Qn/xr7eO3eFf69ucv
equaQ43zi0hnnuQH4xJkg3QcZAu3MWKTNSjcGBPfxky5BPv2cX6qkdxYI34adyuW
idRFMRJw/4fApXXs40xsUBx2YoMdx4ycJy4fM+65Z5WIHYuaJpdxQ1wP2c1WxjL/
iy0xc8iMlLvQWe4HL/MxKulHExUpnORjh/S0ZGlUMSKPxjkLEApT20Q/F/bjZU7C
dyu4f1nFimKfjKvlfKryaewg0HcTpQNO7RiKsSeLnrtGGzAG0L11K6aD7/TRtt3p
S+FOPLB2RyIN6+CE9owINh0IOkRxliocu6npIiLhkIg5Ia8j143uhDI//D5P+n3M
6Lx2CSmLS2VtrjL36R+ilXJ4YgGcLlbLu3pAyefqjRs20E4p5Qqxr2yYPwZnVJCx
VQ2rp+0OIN+V9KdShmP+/sNASqmbYgHM3by0sCoAnnFsU8c7U144JGK27adVEJfl
qm6JsIBodiOqSg8rmCdiitGOZRYwpLGF7mjQ1NszZKJ+B9XgxHiqp6szs4CtJy7c
i9k25ezANVSc2Me2jwcdnpmZtwgyDs72qRGS2jKIRCcTrCCSiCPeOl0TBOb74Gyy
GrRtnTYlJh7KqhcjFfXji/Wcddf0Gf5fyfEOUNyiYxpRN2rIEzn4bcppP9Nwnqy2
zlBAPJb4JRhPILu7NqYcoDJS3W6OHFTkUkVp/oABR8ty2EnXjPSjCaM4OAdyKmam
2h9pLirT75zuMEfxEIRTRoKlEmihVnjmR+3YegnPJZRGcWkdFlJ2j2ZEpUwMJdhm
hv5JKao/NSTtjqMjyCMyVtON381T0xB2Nd1Nigr3BMzhz6DeJM7VDUrwYwz8Euxq
xNeHm2iVpq3Avpj8Wzpsl2m+oTAA/aIiFIl0/wPo2P0xLmztMkXQUtzLAjUhqvtD
Zoq0W3tWSQuixck/3K+t/U9jwCtKvUrPE8eLinoEHFaLzggufwaGMMYCwJJ7p4/a
+q6gqZqysBt58ElP0wYEfDhVoY+mAzwD/qi4ZYw+K6S3Pr+6lL0GScF0jE2O1gpr
z4aCl+dZq5IOUtOhSHo1F77oG53o71K7y8XZygGcWVP2z5S9pcW+a6oXFcvoZII/
4x4foI7uwW4qA5Ab2J6X5pGze50MRkCqKVd5cMP/TCRw6JceLR2LzFP4wAye2uAD
EpGEsJMseTox4+OAdU+hP3o30IjWWqvDvV1r3vNwxJyBrZ+61/9rS4DN3TOg3qnB
oND310KW3px+9CvYnn7pROxYvoeEttULn94eqHbCioI0C29ml5AeBjhJhfvlTPoO
erbO+V/YzZGAJG+sAxEt+S84JjdfU+BTSUiBTZWMA3llnngL1/6R2gty8GrMArJl
gOYxxiCM4L7KgC4zwb5o9IelB1Ym6euqaN7w0IjbXbh4vYEQ5fkLIAO81O31rOKw
GTR8TiAulKwDSMAJ9v2fRR6xBE44iVlw2lEF6OvGrVJ2zuTvj8hc7VH8dOmJh573
UmN9FXQqXIFxjkzdmaiZetKOdptHoFGwWw8zErryR37veV0h3z5dYDBRPUbP+m5H
8TbZqUpEllpqvAPfwNYRqWPiqDW4s5IKRbIO8gs5KSWBF+yUOAZW/rCEacyXb+R6
fxYbGBOazwKRcDvs3Q4CwScQTpjN63WkTT+PNFFrv/cLjTaNxfjTG40Kl3fJx6jv
NktOSPg0relN+igY6RgXVV8V4tAxRmJcYxB2U7b6gQCZBMSENc8gJVG5BVotGvFg
f5EAdbs2NFx+gyu2F3jrOqIIZ6Ub3mppkkubQjRmNuzYTzM8hnWpzJpFsKp5wrAu
c8LPxrC7CphKlpyCmeQ8dsGeF7T4Z7/9JDfUEub5jFyYBRNqsMJi8Tj4SAQN+pqw
Dl/zem+VFTJlEmsvS5I39JjTJqMK1h0PmemIVjpXg0Bog+9Nr2AEBsI+VHGt1PTg
OU+QPrPG5W/7IW1qjqb4bWaZL2owN6z45/OVN/j4JLj4ynr7vxOzJrchDDdR74ZD
eQUtxb2bUgD8bjyLl701OL1PKx3+gLIEmU932LrqJnIL/b4nM7dNx6LEs7JasVMs
Z55ivBzdy6vwrlUiNfbWdgPDs94TLGTpao/7HRqj9hb6eB+iDLd1ka0dPdxbyk2C
Siw4ictVBINe35e98lo6b/G+vM85IWLVyCe3E/8VLWUE2yyLUx08liHLp2sX3/WH
NMe63MMVu4iBSGOVRsnQrS8D8G1vwSQ2BBZfKT8VVwiq8OC/i/9N6chNWNmzEjvN
dQIXVKBLdPUtuqtCHKMdt/MXa1pTLvZvdgNRI+CBBWSahBGTmk+YIkNIKdAkiqM9
Csw3nWFhCiqEuN7vdyYY/+QW8OVaPjI/P9QKkAoPeOFACQc209/x/y7SmA8xGW7V
QvI40gVWMcK+LmSyHxUXPl31IH7KeF8lLGSzn99/recaLFkMXvIB55S33cfs1Mee
Gk9YSt+pNN3MrsjBGM2eKMZVZPnyiqIRIqT48wXC5KLhyWc9hPWCydQYhJNLV+ay
oQnODpYQWpKJS18u8MMhY4X6qGa/z3YgWwk+GdSbdDirUaNbbhNdcD4WgLy4s6ts
Fk0mV9KjXXqwIdigHSRmmJee6KwtqzZHpl0gxjDoWip+SZXH2GMyg6pURViAhe8i
VzQ5iFoomyuUI87xy0T4iEGbjSyBzxiHyosm6gUTlSOVzVYEVq+3w7nibO0i7SBA
feHV2U/1fMT4/QaDKbRStP2UFzl10TyNqQ8F4h+6uo6A9yNgsWup2S6tGxRY7rXW
KDBtfuczLWCSVht5OzRIldGEgcUravnGqz6OmMBvVyPcBu+0axiycIWigL10P5r3
6ufV37wmUFGDoyByY0sT4a39l7qVLVvdqvGbk6eI+SZ+Ybr1L3khd5tCtlizzNSv
woDuS8LxsBTcAEcyNWUqDylGQv3lQKC4zhtTL6pplvSVm9cKc5jd2lH2vKDdCPDv
5xfjB9PE2154zERfsHjbvcbUr2uIIWXsx1hkgk7ViGExW/USrgWdwswDZDC1guQ7
Ols0bS9rxgZrS+7+l0L+CGE5Q4nMByVrpTXVaT91CVOEHT2MrHp2Lh5Tv/eWYPEw
uzHtcTQrgt+vRod+eo/PmsrfPLzjQ6qe6Z7jDGMbvQGKRwruv40T77PR2rSxCwIU
RO+0dgoNiq/m41c/LFIPKMUdXv+yMPHwlNAn3YjsUydYIgMfsuHL8pksNJ4f65L9
8jvcuGjNkCKA1jtCqdBTDVQbDg6BeiTeGIWF7VHz1AJeOVwIceJWzNpBlQOLEVlh
9nQISYUqYCX6qW3eef+jS7g8yqJP2lQeFXIW3V+B8qVaAusTO0iDdycy5L7oxVvb
iPvOdLB5zAyIKqd5/PAfKNGPqqv/Ph30MwjteQlf+BgP69CdtvgtLVsTdrYKZOZC
7qJIxM1A5cu6Z0pYefl+wPuz4mxTUyYVaDKcP9EqK60tSlxktmM5ax9R+6aSMD51
hy/kpgQMGtIWyO5niWSM++ICKs0BsfPnEAMzbb2rY83tdqQAmdI8jw4ZgwKXuz+K
jFhZQl1OJvQK/GOu5Boew5dVQKmOuGz5KSmk3zu+iVPiMylP6kw/OPzfrVsQzca/
D/8p6y4SPMtSeUrL1Rj67tZxAY6u5RyWiBSuyY8VRUVBeVRng2f/URUIDjrtK/BX
nEGPRIF73sjJlmrvre/J1cj2VkNrxNO2d+Cflg2vcYUe9Atci/3D/Rwz/7EqluC+
bOsd7N3eLAJASXE4Kn+E7QbGoUUIowuWtLsJfNrj1T3P/v91al3TWJxXzbLsh4om
vb/jXX9xWt0bGE4qdSBS2Lx+0od9GZ4OBkev38RQ3VzswRHNXyDyiY31U8VxkSnA
FKnAkfVA0fVZyXgEhyCA3GqBnJEh6L1XONtFGe5MPZOFqA7Ee1Nl5IneKYHh64uN
b3Oi4ZJTSNccoNhT9YzSZQOFdiwu1MQ4bSbXug/Tbns9N7l4QdYXNMD7DpBNt9fc
clSUOUfinteTZC/77z39RsnGRJiupVvuzpkWD+5ejgDAgmiKn/5FByF6CPHvp3Gb
GwXKspXPV3RkSnKmBMhRwALn+j3ZoKsslg1UP7ve4coasuQIiLQeoHWFld+GGpv7
jR5Z4g7zPBqqnviE8XmW6pF+vtMQBQ0bgl4muNvjzz8NRgyBHNk2ElQU/dZ1DFSu
6MR0+NZ2Q9WRRwYXA116EfH9yeEaQ967ZZugfDWipsSCwsxNcx+cEjOkW/E0AKBY
Hmxt7EofBLqvNqKyR197uZlubJwSW/N8S4tgvZyZryv84sYHEp9smQLMJevHk4m9
DeSaR2gStjwkwHl6DZPI1fv7eSLNtNQLC+RK9fHpI9hAm7Pc+ZTnafUWJab9Ivau
DEeFUY6mJtiu9hT6W6lU5wjgpPTF1NJp0IJnSnzNKgVGlE3XhFq1xsdQaSZ5DTrL
XM9cM1gN0Sbprt1CdNsNDTkBcrsgdGq2EaatONhJAdA5rPvszRRuhsFQ3ys9xlHf
54FkjQxtZf4hd37Go8tNF1mXUBzsIlLtQxCKvbs2YKYjuKK9DXZ9y8yePpd9h9JP
ZYlyjxoNh3ZqNhRUapCcdO44T1ID22sMiryuWRQBAu5Fdi2/WvOCDj99L3kzO3C1
RlAqdSLPSUfrHLGyyRsJ2nFYWq572TtK2MUUbLc7TSDmLjHWFDCDn1rk97gV6V26
oBX8AvZCKqhg0Ng5pkPCqDYGb+H2qNiLS3F5L6n/IHwO8qNMSbtD9ZVrxJzkFhck
axyAHf0x7U0KGeIaKW/y19au16fxBisYOuBlyAOsqwMrc108mWYD0bYRwyQe0LAC
8gzX+s3lGwNCN7VvYQRGBYb3IwIDNS7GdUV+vqJIRrMhRnjKxjbT8HyOhfr3yKCE
HXf8xwgZmOqpjsV9knP+NVcXej/sGUnZiagfE8/9bb69cub/wMVB/jovaVkNYG6A
7IMCj7WKyKLvCvKXpaHBzb4GAYy7S4DCgZ85qLG2aOGQkviwJCIeR7wTvs3TB9Nt
NUi/8FAnFu4aT12/nO8xs/BVriwHlm5vivP3fLoDHUQ0xb8VmGGdid6ePmwxR7J3
+R46Y0T7VZVGq9ZV/0LLi+UsQJew0pdShz9QEeWfWl0toPEY2zP6HU/1kploZiSr
xbC25uXE6aMy+va6QsxhmaMcy/lHUoqd6dLPJkkJgfd5OP+uYVQX+iJpNmlVRo6K
Y1Cp2bs/vCaKrTvA64QsA/yoKCTcLnyDdlhakVE2EPwaen30kEwoOs9SVOuDt23S
s3VDab+5MUL5rUeU9XNGu7t9hpO4KomYbtmfFdFF3IbznJZfOlw4xesUj9W0l1Vz
OIa7wFm0uV5dt5fbvZgaRvOu9qcc4ueC8d/8gCQGitUjfb/IgsXmn+OVC7ZJOM4/
lQw1M4vB6pxpale0yJh6wfUMEZuYetQOhk7Ndp74cJ5UGtNzOBf0wMs7Um0VhRP1
X/n56j85TFbAmqIKAofwmX4wH46doZJdgpiXodANB2/wwZVNYLD7Zk0kVZNio9lv
JF+cMEE3PEP+hb3kcmhEGiyeWYHoLWWJW62NAQqZDtZJaw28TzEzgUfa+UU0K9BH
aRcdUXYKhnyVaalkw9gDauBz0JsiWkDAPdhRyp63U+0uSa5W4LSJ3UCIB9QjdfA7
/+FyEfRfxT2nrIRW/PvkwxZ+8K7aD1aLIsFtEUpRULnFpk9pDsWGTsaMUgHMkkJ6
H+rGOEjmSUFLCv61ji+cBHXL86B0b4v+IGc4TSzPH/osd34hoLWE22Jvp+ld5M4i
Uol8Ic7E+b3m/4fS3XXUJAXgVv5btHvfsxZUIXl83X+JcwQehuNVLQVmQGddYo16
0XJN0dxmb/+SL9TD8lj2WkJNW/bZYRQUMLNSqBNJ5TwVO26FWwSEynqSisoaOXIZ
OmukFbZTkarMmHD4UgcfK2+0w9RWZet5wu0Z21Sihf684SYdPmGfvEA2Hlb1OKa4
v8zwTjWT6gfej24zRC0AdVRig2GT3pKqfhRFL9yJDaAhsQkf6qCmTKE3aJlqsYWQ
eU2gM+U62h57sI9IXD1HD/QTnR4FwGJFHW5l03JG29uzr//VzJgCxIHNjb16EjCZ
A5cO5ykEgONrHuwniyBk9WJu0jGKJd+vmE0vBRxugnSqYcyPcDMPnGypMyaNyc4c
gkfNT7ICOZbJeU8WkxgfO/1U3ZxxoMwh81iYJRrAOPt4lb0CpQvws3AjrvjhEVt3
SQVv5yzQX5bMK+nqYNVp4X/d2nzLqtgsvClVYaVtF1N+CrVU1RJiBCChkqEJy/ik
Gqgajf/FqkoaLzh8hDq3fyQrsQ8KRCUaPTPP/LuQR6QEBNNa2WeqrY0mb4bzQfKZ
iwQU4siVvia2ZURqJjcUAgKpdHAS8OJWPndv9qRP9+qUMfPkE3+/Oe9W2J0kmwxE
z4WjG+o1afz3OZbP7eH5WVxhhe8BShmN1mVsbnBKoxeGAqg2mwrYGvDX0j/VRz+y
yNdVLGoAAdlvREQIr3Am/rd8VqpRji3i9YDY4h2MhlHo5ag2P4IVmtZFdGA5/L4k
V4YLjTpglybxz9hFdqqFNUydu5ED9GblS5gefa/24q5el6dhfqV3X+lbl9VZfDo9
Ief+QIXfBBqcqKChxnPFeR9HBT0EgBVREWbpp6PAwm4u+e6QbSSL6TMZY3WfHnKf
V7JRfxb10UX2e2IK32AiyienEq6otxIbP92wWwZQFE6flxnkjTFvkA2uPe0kIvCX
VIcLflrMnKDYhk0kQFbB6sxfPNCLQWISuHLsl1OhBAQ6uCzIU8HSkyqbq4QXp1pJ
2PqRuLRdbOQ1vjkkvXRDeBh9S8+AHebBBWV2FuweNgwqoZVdkjqdwNxvtGS07bNh
YN+sV4tLRGf1nhqRWGFj3baejvCPS3JaFMGXPKa53N6cFKpNut53oEBcJYYGXYUW
GuGQ/sZqA0gH0VocMyJwpQ52x6aVrHp8yMHSOGi1yQ+Jv8WCoMXkdSj3ZQhQKwpt
SGFNM/JzuaChgITDpbE7twmvFDpOSynYVKBGheDClkMe6PwiQ6G2X5JtZ4W2lv56
B3WBKpJVoRFxOcQ00ID/i2MegdaWhVEOJshhA5vhRaKqf4EruLgg23JGElTZv55P
dQJZU3L2TeIhxwmkC5hour7dGACXrPK0lPioMP0/3Z3TO6hGaCv2vaKO1hWDNAaJ
xsQbdOuwupo7nHE7dFIp6jVna9MS69gvLNl9RNPHNT1NpVo/28txUKufB0coOaLS
QbTyXwIAVAh7xf8rCB1t93TdTkJtMYHXoiB6LzN/za6SM8Vt0D7E3hZKqdKJXYic
giUoexPrfxF4hgVyelxmm41V4Ls4Boz8KOfeFN7FhMU7zps4q1YzIaeOvZlu7VJL
WRKNdZLqjLLOhZSY13D9FX9NGmNopWkHkGwwFQwEfkF26tq2hidch/57zoV1elhf
T/7O1ycD8whcA1F0ISRAni76IBeKmwODK4Yggib5/mfVNRIeZ6H0c0hpPCr1tG16
4S6VqyHwiwWK45USB8/jJwTjy12vLbhSD5eGI2lXW5aj0P4m7eeZDsfXt21w9iFg
dX5X2CqWf2Gwx9XVMuaSFJzipisyVpyCdX6tI0ezereHH3JAdabVEOupvH4Gq5Ig
y18zs8frcYk/pb3qokqhDX04ommIdBvfmp+XDyP0u1WpNTm++q4rGoMM9hK2bkyZ
P2mxR0cTbxFHZggVLfbPa/pg6mZQxN0WH+TejFA+x+rgAXzRXEWpsBoV+oYRsHk8
+SY+3B9xUzl2rW40E7xSsfP5TfzGXmQcYQY9cZnfTXiIMhI6PL7+QA/TyJIy7lXq
kNCpp2FjqtCTg45QNWZoWtCxj29Jx8mamY4Ka1WUiITXjViWejvpePKUznLiDVLM
VD9psZnmv0I60RJvUkuOn9aqDEmrtV4UgUwuxnoWUinqw+ONHQjselTLt3CzeL3V
/Q72MCOWH/kUSLFcuGZNIhkobI6ihA/wfjl1z/u5p4LdALaSckscT8+7dxHz77S4
PB7lyPyBwVyN99eJj8zeaQoobl7zYzXhU7DB9H5++Ou0Qj2isbXmcQU8XgduAupZ
9mtp7ycYxoMcfXt8ULQ+rIL+FlOldSdX0UufkpW8VdDPVNGQb12nOASgoP4G1i8q
dNrtZT9XEoxY7EruDKZjMby+wbyfcw3UZb6OHIhqenKjpoINolPBv/yFb5gdVORF
Wt56v8s/WhZZXAEXS0wkZ3y0resm1mbwBZY6ianBwtpPTvAuyoRDQsv86mzFEREh
V7RdXpXvr1PtJ56Eua904Z4qX7rwlT+uY2iL/kmDbhMX8rK7utAIB3njolZUOwjZ
g2gm0Mw77NmnpUWuibPXn5ZJuhrdngPaYbPiy6UimZwkxyyUoeMSzJ1G71YIYBq4
2r2OFvREOzV0dvYQ05/7FKgF0M/XnUnzQUsdQ6pnlNk3hRvR8Cg4xirp3vzggVOs
KP+Yn6mUKQLykmQKPdfNNBPIcd94xf/rjJfUJRCqaUVnqF52UPXWqDQY6k+jvxlw
Hh3/hr+skKgxALOI2rB9iCokXiiS+BIveyeyHKh7PfEUvzQV5W0y2TbEfVBjX9f/
fjYV9ZzIcAIWKsOXE4oLvbb3peBlwu0QBCAxdEr80hmUfNk6MOWUIef+Re3JbxMd
TnMoZsdCLgQl1JUDmYO8AZpFYDVhLDIe6PpmuAH4ykpxuO83NkyM73fdumR7VBlQ
MhbW4kgeLNC9HjeIFbP35oeL4uDVEDkgoYltcrb8Z02OFZZU/F2+I8x1n7qL3+j/
fsw3Zm1bmGSfiDQG6QSO03Hpso1dkVORxFhXrKwAEquDNoJuDL/KiomvVy5qm9YE
4/uCOCEGXO5P1nD+BShgOQypdbfyuvOoGVwLjNXlITVXMR3CdUFMFaPVOzwQx5+v
jg3IZsZ3OCOx9MFIW1NwT8ypymndYYBSi3OQqR7gX+hWY+OhvmkBFVjKTLesNCmp
ZRFeOONAFUdvfoFC3vHRkD/Tpy+Zn33b8XAgrtSfTY9J4MxcaCMElpfTZRJsgtlv
Hkrpp9nqwhkjboFC4Xappm3y0QUqH5lvDztVjb9qvZmL1EH0gF0EcRbAZVtoT70Q
1KomCT6QjfUthY5P3fcyuQbBfVz1uF6QL038YhW5i13vFQzs5WRRSBcoanSNX7yz
NU73mwkgs+mVskH+cN+4usDmgTxz9DoAGXTATgYc9/HpkmKYFxjKSBFvb48N2YeF
2e0fYW7YX/mxCcTLfq6J+3Vggd9g9r39/xhCzrsfZO9X5CmhIv6Ul0Lrlj9knvqg
+wYBmMvhQh+1ZafZKdbvJ0oib1ozLji+0zaiP62fcLT+khsrS4RtmBUWLdOrYLb9
0Elp9OxPZF1Ywluh9yYgyfNcmMXPNCL/zeorqKE9mADQoXAD3RfleXJE4F8ohmNO
9yt8714/MRyRe947pdHPokfzjNoDtuhRY5N4ebeGpipwZwVuTj4imfQEWE8caTYf
qrkXym/64m7lpFSAXhCYOtFhYSIWpGCkh9uQOLhXYN6CuvbiIBqs7AJE2nin2TLZ
q0fzUOhM/tsV5cfdqgj/uVn9uUjnRxhnvRuJbP+huTJnRwqvMn8Wmk6z4sG+vZIT
qBU06ofbz0AFi2OGscapiruWxH1RhagTrekaWrBGfv/2SpxqdDyz+luvWLKbj9Zc
PZSRUQzytGEIY/CU6lRYrcHhlmwJ3bf30p+zdQFR3wzFQ/s6J5ZGnvGdNIv+sunJ
Vm0KuhBu7DLLTIvPbjN+4KEvAJQ4NaeEyB5gQ0FN8Mg6BGwwNaDC2fmI9Q/nxC+p
uG3G+XWgj9ujs64i1RWVyeMlb8zmkcnSjVjr76pjIEifIwD5K9Xi5alKJJX2TPWB
5vGCMXerrQq5G5EqrY7IRROa/zLZ2wZvo9x2DrDApdbSCj8umc9R2l1z2Ym9nqRj
cNoUn1f/Bj1V9AY4A4tDp2A5DPH3x8UEa/DBmbnKlEYwZD6C1fDC2oF5EGrRPHd1
6xT3yFrBmo5eJ619FSDng4A+xdQySmm75YI9HMgT8WLCZl26gU6+qpzh4/QE4Ohg
0G29uEoUqqrMt7ydGjqQimq8jdjPbCxE/fekajBA/4DERdL9ygqwy6JsugmASZN+
TSA/4KiedTRHmp4xZ17fEsQmo+jyGly8lHalnfSotJfVz95pW1BPv/+gBfsnw7V7
wE5p8J4c7VKwlhIxk2HXypNMphrqtV8pqE8qhIMiWR1ov6v/mod7fk83JoapZPaA
Hnm+Pf1FfzWtjq7aQT2PXqrT3ZoI/IuS7sSl3ZVHnRAV+QCkP2nY3kYXIApkOG1o
2kc0ntSAFcFE0h+/wZVMGdzR83K/dyyUhsuEUOG+4HDYHP46wULvHcHmn/+MwfdG
3TCqWOsTMiXVtQWRK4fA9TiDygY8OcbjAkRm3XWy3+ACUFc6psR6DUlMO2JHo3WQ
voVbloZdkgsI0fBwntuRg2pHW9wDoEl74ZRwL4sAwTWXq6+3Dpx6mR2Q3Gt6P37/
0td4fSdM2elGJKJ76TobkQLUeCkDvSpQl7WFeFqB6SgmRoqdw0CEerVR1y89qD9h
danbPy6u+xC7b+87a9pmPrKYuQyve+C5S7XMSYP4LucWsPIqiM/nAph7/n6JnivL
JrtXahSZJ5b0Zrd2k6OXQd9DEod17k9tU6m1Y6XrBWLLr700wHW+ga0eSmfhqZ5G
QveCvcQ55vcpEHZCw6FBLan4DqTgbU42tMKM27bF9MoD0wqZ+Vq/VeOVdMuHf6Je
yzsHDbA5hJDS5VZGTSFxVpeJ6ayWu6oXp95l704RYIVcJwgo2rrfBCcDLdEcqNWe
7bja1sTbyZYGFOkrpe9KR8419xGrp4COWmT40mI5+NJjdLC0XSKCYo2C3Bvj+e6z
vV9ltesF3NVmUeK1CLttOwjo9R8h8hgS7YpshwLPfnzf2y8pdYjYSDx3jw+b9prL
h715oZWfb/o4IJmFWTrFlowVn5dz9vpH2rziIK/pO/YYnoteeLrN8g98KIZ9yAiG
eu5iT/LZyZ2lQmd+rMWSc1BRP5cnl8FOOT4XZa2orFy/mMoUovdoOStIuIkol9lK
cdhhhD+PPjWAVLg3QAQMxgsZMhFdjCFKDCCW6VlCTy0twAVUnKgFvhltvlzdG1qD
NR+88liG8agAmoV8MtqxZgC0dcHmwGHbdkdulEzwuEXqP72O41QQ8nJO/PloL+Wd
uk7esARN8bAeI6BO5eynEzToeC91X7fEKm1f3l6kIXfZ8FHsE3uysye0p7VCQqXY
PlL7K5PDW35yNAxtYAV8XyttWrv4XgbPB3lNvcME4mZrlyGS1eWVoxg7y9BmbPUC
xJ31YvMIMAQ55ZJezjds1DH+gVJ4DcZLHh84A3wqnu0cHeYOxNIL0NoeWMM1FEfA
tOJxw8sPh5D69rKiDKTDUKL7Hqi2syK19boF6wT5r+05tVp6WaNgrFl7peBJP8pu
eKiZ/peJwmD+3XQWmNc8E+UA4xLoM6s46+PWLvrqzefVFrEtrmRAAayhF4W1Y1h8
6jWMtUv2Eaq1rnWFfgTl00lhJTxLekfnqMn6EsW8fA0miy+EWgs0v9GRMe3KUFRW
gMc2FV9mbD/fTonk8uG/h1bOzTJ6vChZ9Yt4Tt/DcCUKfW3PStBlH/7GL6B4P2h3
iVQcqkV2613Dz0ji/tcaftMBcz+bb17PmXeCJFE811pJ8nFrFUEFkOSff8UDGhBL
Y4v3QtmN5jovpZ7XHbzUbaLKAUt1oMlQh3nxy6wJmVoPjygQPBLkiTFeQIyoLR5J
nUpRoJaeIZ1tMRv7dTUvfrASr0dLepPr14O9bfJ7zykjcUli++7kSHoIs7b5XVmE
lwOji2Zl4meKnexL/5Zas4zxdABM+vWW8YLULyaKX8qkEGcHByVapui0CwY8SHAY
FnUuhepw7x+TwEqqPNbV64/7gmuu3Uz9RHGLciZlHHupgeKr8OPVFlU12DhpWzL4
bBYDPgZqOC2nDyg1qvnoHdw3bNaMSBqbbyPclugPhbF0fHLP63bib4LZNriZnAL6
sr0Z1GCXEGEpCauAhJMCk/5S7HrSPuEPkd7hS3IJTp5oARK2KkFGu8vIcsTJ6YZg
sVilkkujOXts+I1WPCEkemgMawlq+PMlhrxxrVjRgmt0AL+Q+sF3p5W5c5GLHLGE
Y7vhk3yPkZueJB0EHIl6aQsYkWvFdysKi+DT43CvF3qXOxZuMG82w7dhFNbhZnbZ
7klABHoLyS6+oGyUw/+jh/zWlUMKFE5hg3YKysPGnQejWvpu0kV/Nf3H2esOzsum
LuqdzKA9XAEFJlYNWe1m+8TvpLWluXV9bfWZikniL5TgmPGeakUkMPP1BhFTBUG7
Y77j9UUjcHMMC1a+D0mFQeupWN0GiNlAfmfJh+f7UvtA7kw1qbDNv06f3fgoWoMW
kLcMiphL25EkBL9Uhwdo21wxBsWAB8nwQs63f20QqDKBQSi/SRHX2vZZEPCZWfRQ
2YSpEjosivhMvP0zDlUF5Q1Ditd7g7pTmOusfIddXlNIgrBh3GZFOGKsfIiJg1gW
voXjPJW0tWv7zjWeNr19fw/B9MooYss4veNP4xZqzSWndhKDQC8MX28r0kDdjKLw
doPogG106s74wyMAuvAmYPTb0gSJmsOsDj+IDpMw0kLyFT1UoiAde1mo9PuTatYb
HB0XLMhJSpuvoi/L/vmTRR7PJSlEHdGbHnW+HpJAt4x3hv1KAI0e46nmA+3mgMq6
h6ycpHNh149pr1Qrgrb4tUyT1lG6E8yCXbRGrr4xrq+6MmM6qvdmcFVR56vR4xpw
f2QHOf25C3JNeCPY6Z0WHY7DC2QJEsMhyXK11fyHeUz22X4wW6M8pbAKkB9DhbpJ
PXAz4cMpmOVKwtM9XHCYLAVu0WbuPibt8KBdhE1AhVrjz85mTGPLX45l/5qwvacs
RcsPevh9hI2HySQV6mZkCzAazPd/CuKCBI71GfrAuQaeL1gT3DQq0aola49hirLj
xK1z0P0od6pYfG4TwQr9FaXyUafjOXTuzep9cTUtvkUOo+adstMA0IyRy+F7i8HI
tTt31Z4G8dbYnngZBXFoj9YsvFQmVYW3ynSGYAk/OO01wxNZ/RgGXbIdWoqv0ynt
MN8cFeZSZBgWjbMF8l/5fe61S+Ew2DC+hW3vPUB1xfm2uj+wDi+w5EbrIGqtxfdg
8E1wo/UQkh+LUF9jHxKWUoyxdCs9ohkwjjVKMN7RX0CfGCBkk4aTpZ1Icv6QvZFn
4p+o4hbieK3F47hNLnwpewYGSnSTFA4pHjV6f0eaHORlAkR3HDAM9vIh5Ek7zqnG
Sngbq3Ym+p4J/kQcbXbELmO4ip5x+OG4lYbtu+h/fUj0N4nX/KJe5dARx6hMfEv9
vP19RTyJfchWQX/6zV4Tj8jnMOA+C/7yLeSuIu30ZjskJbT40TlI2uuY/yhkkgxZ
DgZKWUJUbeM/RM8JIdj/8eJHfaTJVGNuJ/74jb4AvXs1JoYw77FgpNUEEY2vn7G1
6NOf/M9/7JbDj02iC57TEjEp4czT7At2GvTacMYnWzx4LR5EDvYFey/CmAkM4Su4
+JQKdzwwqEAthSowPZQPZJoc6ehIqlV7LgFjzQUqkfC/Xu/qXVlDtqIrkoklKA/O
3n6dUTI1MPKcBX/2EhP00THQN2Si6zMRfk17a6HIjusejLsYP1nFyu7lexOAFj09
+4OVHnGz1xAYY6E5rGbG/ecWPqttbBuggp7MkyIc0U9U14e+A2JpQ+cLuOmA2ife
Z66FaxohSzBI8FbGhKq05WtYqHBIAoM4WXn8KUPKVrpUQCKXVeuDtTs8/o2w330o
LVW/pO7hwcCwpzOKY+Aw9H4r9ic0U65/YSWqpGx8bpYHDZ5YMtZaDnTsJlVGcf4H
bqnCc16/ITYIuX9Q3/CtmSzuSmL1l6LsTjFiHGF7ORJvcVc2UHd8HNJiZiwWxVbk
JZwMjA6edncbiUDrFrG989vTn7PyVecHv86hritLQ+N+5PzrdANQYTGF0YMg0Cri
K7GDfP0xtHMwXCIPUuLUg9ybCro8KEYbd8sbwXQLLtm1CXWt+OcwvIJXAasxgwRb
/8QbdX+A7niUsDU01tZU13BTfD3bEZzLYooIO10j/Vpmc/83pM87oWsyKa06LOf9
L45+iHKtqGv7taK2PMuXmlfot81jWrjah9ZxUoz5PpG3/nUvKjcfJRML048dEeVr
vNBcna4HK9z+mX2+1b/dp5ol8uGysbWh02I2dtT6DffVkQruZU4dHDq2WO+rVHN9
BoKngqxFqoDl5rwn62h+uPEl6HY/Cx29kSJh2DPWxHFMVvz/7oGe+y5T5fX7aWjz
JD5UlRiJSg33DgBskyTbkUv85uZBR6ZQ1Q6THp6YfQMuCNguy3aun69SnkFPDbJT
kFp4R0euhztP5uqSVjTEw/F6Lg6lftaPxHI1kgrBX4QQuV7dhxTXwMUs8IpcJ4ep
AgCxkIO7xOBPU593PEjqfsAAGWQUZLOlNlyHHmcN1gqbSIiZ07MBd12HQSBVutr9
Yq9MR6WE0w9PV4YONBpv7YxQXxuxcjljwTGWuwBvKWHuPIOyYpCJWk9YnFSe7K71
ni7pGL7myneKhVcf919Y6s8WAKTRiV11TrsaAodytJKzA7v9gBIndxQDWysmQH1P
ZLXBPWLcYS3oMtjf9hXK9ULg5Ko35dOSTL66eys+j77YvtryYyTLmwExzHpHIxr1
dWvh/9GZHTkbUTToIReFCpErsBMnvWXZt1V+Dy40U6Q9NAvxtxRg0HA35g0RYzZa
T2Z2Q9FpxlouPgqKKEBzTZoox54GS3DwCvqmYZD0HnoTl2IfTLllDUXIV5phEC+c
X5MYPdBJAhqjW6OiA0BNCn+xfIn/rzHOe/GeYu/nNXSzCEpFe2qFnYR/e0uu3cGP
iFdhNks5ScdER2OKXXLVJdM4QKYuELtCpCXH8fsABFoll9AZUhUROx8gQj4c9fm3
A2DYcBhD7dB8pAlWnCJNEl+/7xk83gvJKGI711HIVPBDB67fB5rTMqbbYNXbzekF
K7cS6R64a3pMhsz+VN0XH7A/+B/JFDEIj1qg2RReJxQgXtTMYETnlzUp4QerFU/F
fF+tDwtQR+zX/zqKUnubY3bTFGHNWRZHmGw64TVRrfdZAEANf8bS7ifxCmm7kzbD
RF3NWASVRcyO8ezORnudJN5zVsixs3+g2l99Dbz4dJPincD35/O4GwrSIOTX4Chk
OGa2HBlFUjp5WFUgAfgaMeP260DNExSCmVWivVpx7BhYVSpI8vDlrjCiRCGZ9QmL
zfmWOlJ4LhqODptOED+FAcB0KIFCpU+rQhhvlGkSNSeE8AHCyULq4aPKRXpmpCT3
dD9R3EfKfoHcCBW/fwp5KicaI/f1mCdZxZfluEh8vPgkBBxDpG/KLwBLVPH0Cj4R
UDv5Ha5Hebayi9TwSCEPiLpYv/HroO6W9juDNYK/YN/tBprlIA7e2V8zpDFOcplO
GEmKxN5VAtal6HvjEc/sEpTTNG0C322/++lo4SlId+UUzCpcyCfh4l5CnKaZPupA
yzIsvHnqc++jQN7oE/DJCRtI9kQRD92MhGzucmnnr9HiWJ56L1m1TWdUecfF8Ze6
0E1L84hkeNsLTNRozcYeek7soETMe+zsQmkldLMdhxwYNLW01WDzid/odc9ftojb
UzHSpg/QZPXzezt2wmqIZVzqOZn1J4uhNX3/g8cL5ELSSOWYX1bMxI0QITX7yd2R
wyhps87lBuEeT6bls1Xq9uMkQWA2dfdUrvKSLDLwtyN1MRN4+TJWS4+zS2XR3CjL
lZW3A+BNv4OrlZgQaxyz77te0z0QP5v9G3kxnGINJUm2WWbhuoxgqtDAt6V2lXBY
8eBqrWQp5OQaW8Ks0I97dEHuhOoE+ToexbuoXLJjA/M2Oph8rOAojQY7z583i+80
CT1X63Zdm0IjdQ78nGcBqOGQjG++x7+PnE+9xOgO9H9+CLb2Z2C30/TMYcwgkMBo
nhcy/RIbHYAoEoKPvDsnvue8b4apZrtuKKG39OxMMgSUBG4p+lDbbRaSu2YHVnne
YtbvMbkMc7sLe/wMv63SGiwH294wMqR4J0RondvCBPIKhMgxmz7KiDcsMRJSyZQe
IIJlGagoWVevLmaB8t7RsIDZ9ZKWVUyWbn7ESn86jcaZyg2SxaASzgXUs3Lghfsb
H2Eq7fb+iaO3aDqCqMwcwf5qGSuEWZl/El+ZvxvwGTagD8cxBMK5lNudqoRsemNR
5iESnICrROsBv124L7HVBh8/pbIuN/cllccYznYcI/3Ri3jXnmhB/7t/Mjg6WAfv
lj67t9LZegQs4e51hXk/SvR1/XUNHBsiY8cKcFXDlpgx/Ju+b7Uubu4bRRZT5DpM
RnTrgLjQiROZ8BMrd1P/DQFs7F0a3+1fxCpIel/qxm3C7PrOrZMaryuk0U4rLEWY
TECfYXcMWeJXUFBdEEahBZs47a0OJW9jge4DN2d0FZcXVzJFASeWAckOd/r9Znuu
w8/TCbiAC19sYXOV7f610/yMKn6/va5LyMKux7SmPOzgpRaTmI7LXsjTny8d2stL
FAnVrUK04mqPy9xEoYEo5c/w0oF/CeBQCSyFdgPtuSmHY1xKzf0Tw/yIdwrLwKHl
cBuyslRWdvL4MeWgCNuUaJr2aY85K/L4DZM+OKGuCKAgsJXwjHqWafpi8hDMpzBU
lxBCqcUjSkq9wjE0Um9KQoTgdHw4flqnl7YHf9agj1TKI0VTiN4cCAv2EzfJfood
onJk58MTmhKT+GL2BlZO6td9ttcBzFyTYbw7FOr0jd9Ynpy9cWST9EvlKtJkgjzW
mPGK/p+ERMgifgjt1HO2Tl1XpwklTcxZ5vSQNIAECsg6HtdPYIx7k3YjMR0xSD82
sIqgS0sWrPozXXM/Pa80DkMcV3vcSsqvOe8qssxLJso3ijUf6kaHy0+0SHEa7wxz
uQoP1Gma7tN5W/HAYLI49MHh35qwq0o8NZW4fCtiDlUIvRFJcDVCk0g7Qkjj4fgu
TOwm50hLlerZ2dPrKlQNK1XSygRVSN9oxtHZBQWgqTkmd02sPg0S5iIIaIlZABhg
wivOCQWYax3D+Z0y3kiCo4/SXRfEVsMwQhqQjjHU0bOvEraR9sS1C0g2UDo5ZvhL
tW3nRubxJYjCm/xjmBdDHpl922VJeNMnAsNkxqCUzeK0FI8IQYPZFhKcM6z8ZVlb
qzrEBsQRHN2dT4cx1Fpyk38O+6tnAB+jR4dFzsnNa1F4Fe5GZF3h2JgZuV5teufk
mvyNLkvgGYc2MhWd/3+MKkbTMojIhyehYCPNmCoGwnHFtl3U92KEtffSEByB3DLU
zTUDSDBZOingv5mWCK8/l4gnkIxX47d/0m3V+5N6A9dBhC1Njb/pwPJ6i8XS6KQl
yqM/I7bcAt+4LXd56cvQIrx0UkH2uNrFd4CLymJlyr6xcw1MDMxhEOD1h4lkVfT4
b5OBIIbaq3WnyTzABNPrPtiBh8S9KZPXErJ1Q0kW3NFD8KzUGzYYlXr3IimZCkwq
aZa3fzz94add1VNKrkeEWUkZnaPkJA12WSVGvRMrSElGr7vDXl7wXscIPmigN7cV
UNstxjGf42uxAzMYAbrPP4b71HyZyQguBp6B3uud/5ubRXfK2YUF4PLixKYb+2C5
oEheML2XfWkjaoDt2IOjXZEz0NRSLyjFzIvmBpV+wTCRMooB+MeZ6YlvddIx2Jnj
toq1jDg+RW6ewbdHHdWmWGS0oepFMCQmjHhbz4hHWw2fp/+GV2d/6y7TaBW/WrpF
CuQxRtlcFG1CF/ZEhOh9VP7Wppxi0a1Nd2AdtgxTK74N+iLfTy485TSivk/yfyeW
1SRM3I8xQLS1O/Du4SFO+1p3scUSpf0YxecT2Ffj96nn1mWLL9299v7KuQLNEMRc
e/kDA5+oM+BfHyGdQOYm1Si3VnZ7GD9mPz1Zk4lJ1YGb6iJWUhOWPldcqPu80PvL
onuGe8E6g3u0FYAHCSYt9uR2UIxp2UQjr1xoYhZciWzt4LlYwm4+UqekPKx9ljy6
bE6oQljBuwSI+CkQE9zDg92GyPOHelbddryD+u4mn2LXbaeXfl4i9oxAs5P7AR7D
1QJiJ9rST+jif75tdXLOzsSp3Gu+VPgl2/sSvuz+xwDtAPfcCtg86HJrued8b9pV
ByO3Gotm+jEFqMtSq5tnu/Hr8ibBmV4ZXHWN4vHSTmwzANsaon5hxnc1CylmKgd0
MASNjTo3mctWL1HKIbD6+luSTCgxgJ+NDpYts+epxpkSRn/YbirhRPEuHUVww65Z
gwpkaMCu56pFx2KfXwDE9QpGzeW91hzZjB20bui7alrFh7qEMih/+diIfiEsfR3m
l7pEUMK0WLjZtKKSshEaG+qKFTmiyQ/2shKejqbhYjNRGHLU2nB9diErkEjAaj8M
fTyQ49n/Pewx9XGzqluGLHRQW0wkoKpcSdJgX44FITChKIlFSYurGRcI+nqG7zqs
FuWZsZsCiJQgbEaLJ+MajL8+GoGw6N4tYODDzQbpLuQwLDy3eq6sgPw5bnocIHlV
+zfOyE3KQLbS1r6n+fOnNubiLQkurfFuQkxol+7fgpqstmPJed5zd3TIfimFGil3
Xwo+TnpFPTLOuAiwZuYA1hyB5wBp8pl1Dg3SXzZGUWP6BFZS1OHXCUAUTMwDqwaY
nFajWB72Eq3vpH/bhFnExGVke/R9VeADKlb/JTMnQ9QQachCEocI8rHDX2R0911o
napWgX1PMsC2EInAhF4lZdHklq4HBbkdtynBoWyhtg+HuBh1ahUnTSdTDUJUcmUk
GPsJOaSSMFkckyZwX3TMaEdn9E/rOE3lTRONXMLTbOI2CAFy2a/neHbt5AVMC3ci
LnRxM0RWCgV1y2zJyeqgyOWIpuoj9xTl50jsm582KpdNUkwxQzEkoreWyW3/ZHb9
VjHkqSMetICnwuQykTAlf1V5NU7VWAC3Uku0mYNOx9h+epVgDYxz62WcxDUiI3oF
c5cfHEyLUo9oLx4M6ZurUolfn3viwgQUY+SQF9fRiHq72BEUPk5KF47XdjUFfwCo
+4SLtb/Nbz8RcyZsp5FrZ3k6raFVXvEM272mi2vQwsb7tkRnVgOf9Gkx/LrBiDc4
jiHyo7QAD5G3WJn2dimLoaEcOUU0awe6JsopRM/AtTsyv8SowPyOov6KgV9eLnqJ
4636L+dPFbBpU3v5ijX/t5ySxycKXQKws2BU7PoUVfFFkd3g56JSCQmDSxmQLvu4
Dt6fw51ZI2vO/O6GtQ5Uf3od7Aybo5rCw8MglA0OjN81XS5heWyGHaXYxtEZxhOy
S2slxRnmPAUac5ZCEVFLxC3ZptMfEzR8dWx3rP7/eyyaU7v5u9g16MP+tn50MiAl
wENB+Yz7WZeSmmgKZaOD63YYlAqsih2Cgx7R/6vvlkrCoWNi4QKq+qP33+XhFg4u
PI36Fn82aJyc0qpJyGLdnBfrLO20gGP3urZMpOeIkkhX1KHhdXCg+Rhp7A9U8ZZe
41QlV/28+BFdhWSliL3uAEv8ZMjUMZ14aPAYR2KYcl9Q8F+tgC0Nn24I7vs85obk
vOB/utrjHrFYzqzYIapdc4jSWvh0VQdXBGBW/9B9rcqJCnT2giobOJjnC5g2feRv
s6pSzF6/UWKEAeJgaxKjQTel3s3TLRmYVlq+PpKSrsug/hRAqrqQC+3qQAp63W1n
qaoOxGqOG0/OQJlCK/ejI5YTEp/iHXCLw10xVKH5JwbBK9PAg8zUnd3obDByZsli
59na/MOMvJ/GSlmSHWfSvV9Rv/lHwCOnPzDzwDISK8wO9J56qw33NKHiWAoRACHu
pxIWGFrBvKF/96F86E89ThCdPC5g9GdIbmUtK4uhMvwOaTtFH0mpljnzmi0Cqzf6
RWoOeTxxbp1eurmaa51nwrck1pOkfDSfIo9cb2EqI4A3J9+3Li67qsJjfEIcDRQj
t8aoudDmSXR+41L0gyTXC1T6o1qc+//eke/8bN1Q8I4Kv/SeMX7ecAbb2y8xpSaB
2TpxgbmKHxeIAV6lIQrOIm3zCHRCWwMt//cdxtooW9OVsDeWsiMuqzhMmmsj6Idz
YDMJnHHKLR7zyBu1+Po1EwgMZ5OIH2+Pk55n0lgdX/CnHx61Ga5G5upISaWStl0e
NEBaYs2a2BDUVzkGfvuv5SGxdxC7xph42p3ve4nZ1gJ6by+JOt/Y+dEJxZ6ARJod
yfhVEI7qrDBZUXGPwftJeHCBpUrApmY7y1Jg9NA1XNVKjyaZSg1Kukp69tR827QU
Vwd88MBlDNfStbqS2ay3F4f0/wNGRPAv8GZ1uCA3PGMlXWd1XXO/caueJBpNmY+b
60Bxmpy39T7epbh8PCqAor/JxM8dOmCIaYbROnt1W9hwcEksb3cPyj5LH4xNivZH
T+eOHIUT51b/lPlSLCsG1dyEQT0un6mk/ZT6e3Qdu+440C9sXIsEhJfTGlJHytMl
8ULjNBADA5OnwtHU9yNOCMMsUoHqG1QooOq1JHZHMkVNauLNQv4J8I2au6NshaUk
1Rm315jbLeWUTmSPJ+UEGkjCOLNn/M39e7H7IKYtYX89eKFy/prP6uHm5s3av88H
0Cx8PelUoOTtB1cU5a9xW/StV9Pl6mhvf4sdFjDl51kv4/eCfoHL3lFYL4wU9Rj4
UmCoOhvBmzi8SgoU0R+f5SDszteAiy5NW5+xVofhOYZQE8X4OOAANgx8UBP5QcuP
dXXwblx1Fjxn8K2qMCMD64/wXl9yAQ0E7zyzUZBNmLyL1FGZTiATaPAxWubTZk4C
3mtFVfCNOZ5vluvr8byXZowLUE3tKb6Qfw5xe3notN0qH1arWQpNbUhFwx9KsgLd
S7q3yBizLT4/TqMbTtbFmUzfJ7oa13SZ/RGGsZKRc8xj1skaACPF9sMrHbAKXrD8
0kI33LIy4Hr9cFjO4VOhGoya1RUNVH/YwaAdbrGODB3x30CRj9acR95Dh+lYCRHa
xmhbUtRNoUGCK8t010IeJf7+xxjfCqOXNSzLzkbGPyki6Szvw06l1bQ4a6uqWJw0
x5m5pLq4SVUlioXE2sdd2J8LHQO+fUXBpdflRKu9QP7NwPOc2NBSlzOq+EHpl966
W0HYVaR4QTAp5qmdg9njE0DC470vbMKLlTu2vxWzHJj1XtoEApcUtCDbUMhVofSm
NylBbMb+S6V1BIP8wkM7ol2yjNN+Mm7izd4hHFRwBJwlRtsiyx4HDicdGT67sOUx
oRv0/n1PHgxT6hRvNudZEe3L9LFf3PwpkMyuHpkht+bWlKpfGhG5KGSLvgO+o6Ko
77ptDix9YYbwVckTuqQC9VP2gP27Q4KBuTnxBpK2Vlge+Z/YhSmV8WgAI4/WiMFY
/vlMJiCgy8ZM968SLNUu/P6UPNwZ2EH/WYXo2dF2zmQPqQvCK+k3kBpUkxXlOmxS
60IBtsirNc+VuPLR95yJuOz2mhMtlejnoc7CBHsN9kGJot3dwnf8maTZG30NK6Lg
FS1fYeoa36lY5kBh36vLdEFLTTC8g1KNnRzLHgl3vGuRuS/+zR8qUwQJn1MQLRUx
Gfc9/tIubgyYmTcVI3gYQK/aMV753K9rexV/5Jux407tMqzTNdxzXoPUzZxsf8uw
ZXCrf/oOeKkA7HhLPXFjYcRXZr0xMguHgoeSu8KKmG1n70dWyOntnWuX8ANw/mfK
PQcCd/hMQe651x++CHs5Bki9++EcDx63PhXLGBnjoF46VqmzLqXtzWAisn7d0/Eq
sepDTrPKwL/qw2fAU2xmcS4fcETPm2e5GtKf8aIKC4SIzfkesEmKR/tMQNhSKKPW
L93XpFEAB8fZY+9jxW4DSkb73S4y9UdMJTI05ecYhFJaHL3Kje/cYT05/PW+2Wus
yYyLSSC830/jlR4TWeLiXl7YxJlz2uRkKR3p8ljPAtlG1zva79YCJHvDBexJrmNO
DYln5FuCp5kKVxE3wndwHszNK/pzpj9Ks2F4KbFtZr5HxfYqNFltgmt8BbRWtWQv
5DKDYQobYcRxeFtb9GGiliRfN5227aqbEQPPKJH/OBX50qmcAB7tuZj62AiYfUyy
WiXdHJYeGsC0P1DzpKHutMXHepdifKxdoHbcRjluNQNymARV/pHi1AEIDu+CSxl7
1d9L5crp905VO515bfGpsy0CKI5opmYm6Glo8dl5NPs4Xbzc9M9Tz/mOPRMw9Yzo
vGVVaYp3otWzxcLZ2yXDZ+dpTRyGxY5+rDMO3Vsld+kWqIZx2qkcNvB4lO633zF3
m1vicdOHtA4vUkxjcYchdC9I9LD2bGWt+MOwbX/M1ImaxA1k14WjA9NRrItnrL0/
O0qVL35dq5g8SOPwJJsBWFNu9/nqAsGt6DOfFTrLOupGEidVxa2igEw+cvC7aCZn
xsC7QivHw2St+0G5mBkRB+4b5bduDGWguQEGkUCilOYAW81mPxgDhGu6ul4vGyij
rXxOJ6TWJsr6zbJvblla0t0t/t66Bso1EJ1ArKXVoGSm1VgbY80XMkKoC8qKO5qI
30JQFnel6dKIAUMupVdVxF/JZF4giQ3KTDBCliy2WCN50BgdJoxCwvw1NUAK7Zbj
C6OjeSokhOwtPOJmhVcPd/foKLvbc37auoA+eJrXop4A0I5z/0gCL1ZYm8UxyKr4
HSc5K9IlDtsfHFopmmNwJ9LMjyxjFNYARSzZ4HtTFFQZlny3w3JNU04bJO01W+5Q
22GP0/v9YcJ5rA34R4ZsFT7eS0nFYU+d4/vdVsjFBLEFlZRN/Lz/F+/4j7+5sMxj
Zzx1+fh9QQHxFAj2yEic0W+sfG0w6lySO0V6MQANnlkxkwxwb24RJc2X1O6turEh
F8KCif6rAaDRVX1HszMhgl8CBpdeP4+MxPAyhX8T5HrW5qeKDXdoHQGxHSjWc5C+
AKXjy7fp6ABLIcaJrY6Z4wL2h61xcjzTyNFr0IcN+tc0r2xo+QgIXsrLqWLI81oy
C7PEpr0bVXAf82Ge2YIpz9lbT9JD/GDAjFFYS/BS+uGyUEsNZ21o4ixTh7xj8dwB
Ix0euBK0rVfaL5xMT0Ox6XRVlnefwhjSKhVEH8q0GYaENMSj/KXwsubucXdOWA+K
z9L7Vnyz7BU7UCXYA60BKrdZzWG7w8uMmgxM518dOJBQpnHendgT+tCCzIIzysfA
KzkcbudR807CVeEBEu0Z/nAq+zsJMauUwCf0/7tKhhhDXVc6g45All4xb7v41Is5
IhOnnv48fw8O5XIMgWrOL9wn8P9008skJRlbD2E/eVRXxEXl14yogT6r5ag90EYK
wRHXyHUIOE0bfx0YfOLp876Bzbqf73vv4TcmB9sBLUWGj0YsCM01RkPbnf7GOOCu
nwOrzjWlBtJaVrS3PxLTFN65nd++g3dFQh+rA8DYwR6Y1KBoFWVsD5v4aXpz+2Sm
HLVzF00ephT3wEhcw5XCqR+VIp1xybIkEAYSsjIksChT0nmCpp7SYDxPwJBmxdmc
Q0ioRAsGxFuvbs/pdcIiOa4HdAZ2npcS4usELgNVL8NaxAEMpQKjnPMlFBH9slzg
kBYlaJZXHskWYK+qfGKLzTfzCixKt1JfAEkrl4mE5NogTTZhw/ZjDBHZjpjiAZ8I
C6wPOeJ4CRIhSh5ZIuFrPXkDcWEFLgs0RW35MN9xtyKnGJoDour1IB2GRb6EC2v+
K2F5uh7CQwcI1usZbqrQHDd7iQsLSG8+16MyZReYveYdTi2QFxszQ3aSborxo4s9
qq6LKHV3bUrolxox0W//vgwqfVOeBUHGPZqXtw2SoEn6sz+ZNF2sEP4QVyUN/fjB
7TGkDymnMfe24oQGffNjIb3UL7WJNSViBUA2vvlOKDss43A8KrmdjJpNsCITo3ru
CzNSverz5agcJX3yns1RclVnEexHBkg3MfmR45yNAfGVBIp1wgQmBY4b06dnwgzQ
nFQgKdXgPfBKg4XTa7aSmQugSZb3H1AJEW7g41s3CCHsQj23CKimh724UPaKn+bQ
FnLh+//MMVvoUxaqXcKG2mbDu6GyDAXu3E95dtEiZAl46IXCWGOBIkgFaA3AeE7l
xKU1A2g4PWvwxV8Bx98nZZQsCeejRm90twMoVmJjaFKbE4NFUruIqkaYcRbbJUcI
DrJfAhbBZKRgQMqN/q8afj/sRNgd7XXf2ScJaK9NfSut1U4e7/ZLAQ6XF1/wh30o
dn+/z1poIQ7dbGeFqMZ2lpUkmGGEJQRiuxjoYJxt5uW2V8XDMemfIZfEn7HlslEK
xwD8sa8211AGt7yec35XvOFuIXdelcgs2tH8nd0MdwQAf+V54iUl/NY0PjKkzKss
J7bOpijQxIC9i+35wg1IwFoHiiyBlVpEdiDLJjNHVIRzEaK7CWI79cBKWxnxeF91
s/4efvRELTKGB2XspWbxzdU326kKTAQ/bTc/NxJ8FaR2aDIrPA9L5kcMsj1/NUlv
/8kfEj2KoTohBuBcIYEBznAg/MHRa+oCORrwmmrW/GHOse7fp/ux7qidxG5R7gQi
IHa2MdzrAysTWA30c+7d+8oQIlgf+iDZVm9xKDVIH9zTOzEc/BtGtiQ81eGRj7eK
uJpeJVTg/RgM+GB86lZU/yg1omZn+kXO+irtjtPOcJ6CPgwTK9yAJKyRVTQDUUF/
sgi8FllAZ4laWQqs7CPe+p52XresOW8Zek5qHCis4ZccGh4PbO10GOv78+rTlzOU
Csj574nExktgVc1Ogyt9AqrXf7t3v4UFO9VLUlmfBAvgftYO5XbpUVzC6+Do2Hle
6Gm8PRhtCBG4Pj152L6hcFCgyJGonfWyDAWJA6jKEI2sYobULbGJNzpIVP7DjY8/
PqoLb0xQP+7Irz+Kew2bhWYIIkrdQ/mEtYwnNTmCjkQCnrP1LXsXoaAHybhcv0q/
qGXUbj1hO/YKu3aYboVHkxpC+AhjPvDIUEnLqPDpHkb9Tk1JbXSHijVPMn63SQx0
zTbhBmptTzvUlPoU9Xb9l2v6XYSkSCqNySUuBMRnAV6BrqrNBlc9QuECsrPt/Pm+
M8ZpoQ77YZa39ytbZJGQm/7zkcpAUqYVPjrMjxOQed0OOFW8ja96gCZ5shIG5Yt+
8nPmVXOXrllqcVsFxUDiVGDGrEBpg5+lmZBrJ7t9Dvy9CSEXguyba9XEcxM6lUam
13zO+mUqlzlk8ibe4EKyrGxDHaNhE7YJCSidcjxQDWAwJl5sBVgcZYpKvHqsgukk
0b2PMiligmctt1t6hEA378hiKaOf/TESJGyzTCvHDDxL1u+6SncNCGZITn/FjBy3
jsi9vqm5cxF5tJbanIuZhRuXfz+ImO20IbLvJQ2Vwp/IKpi3iPnNuZXTQA7FUbqd
KqJEP92Pc/G8pvXQXnXdUm3lgoFoArdbA1yLsj0xN9Ec+85YbVthRmaeTi3Y5umK
WAPBbVs5PbwzaGdPh6ib6JTaWdwcvrRuemnXKbZUM9LqwJ99PpAxI5AxjW2nQ/jc
MhrlhvFMvwYvikV5czNbqkCt5me7lXMLIsZNHZHSAngGdvCY0wEJ1MIo2L4/GEns
MXg38NrbmfyrcO2ofkSXvXGGZIil3jjPNtzE0LHI6OooWuq3pZXP4/CWniXBs0X2
8RbAoqDTmPA4Nu+q35KGbZChugMCSP6TIaWwPpuBDeOhf0EBxiWwF+J+imi+RxPm
FJsZe5iz7isePmwO7Wl64jAcKyaXDxFCxZwAZCbCHd6OK4VwLhQrxZpYMjpuDz2z
GqYqNiRopbcoZAX7yrdP2DN5NbJVxaJB4t8tAbPdddJdFxf7CyIosWD1icOIAhjn
kyrmyx6VZXDmfe5fW6N8lda4wSiR+EtmVnTleeSo5ZjxVkLJD7g0rKBv7LJslmft
7Mb8GbUpoyfic7DOFoyTklz0Vg5fnPr7ek65WLHFp1QYN9n0hCL0rHEOXYYdmLhP
3v3WTH50wl1PRCKQp9xTfe64dBKLjDx9xnFjL7rRwVfk1wIs3iwCLwznqcfAABEB
B9d3N5KHqUvMO5EeZMRkUnpnJQdkCrTOiTUums8rSuUnBaDUAMu9+se7++QcbWkZ
HZyi5jk2qbjMbu95Riy5BTHXwWE+Hh4pP62IDe3PPNT3nbSuJ0F2fj76VbMcSitu
cLt21CoswwTT5nYIXR46zkL2NWJG9HdTJZH9M87ewvpT9yMUzx2EayTrnOv+qv4f
Q9HlBSwf5MvNGu2c+M6mk9I4WUCYIuMdxFMeOZq3et5X2s6IIqzqDve2JTQG4MBI
zXAdb81lzHtNTzzxSseIsoBojlpfzWfJuPGxnMUUHmn1NgtaT+bQgFaTmq1GJIOU
gVivUrdiy1vDJ0KEvxQpjxbW9ujymVUEjJsdLUBf7toqUR+hfUUhogelhpEPGLUE
8ScJKf3etrtClVAqDxaWaTAj0/EvBNI6oaGoUptxoQAS9xjonpLSPQlabfNGA8B2
zRuFt1yhIRszo7g/+vL+DCKTqw3LzqP4wJKWsv+VyqBr0cs8SCcbOmT3ZLy9Q4hx
f2ZDryhKZ7EiND8GZa9lfm+C4Auj+ODNfN4CQmq499MFFG73qef8NgeH2vzf895N
g8klZAH9GJCmkA8afoMKb/5xGMbHZYXSdYagNAmU4dJbkFg8oPYvXdgoVLaQCF4N
iyVx75L+dkNabtIi6zEUemDkeMV9hAJ+Sc8DtjrhrEWB5el5cNtMd3U//rXwe1vi
S2j5qYXbGV2F7Ae4Z/vPJKD2o4Q3VTUEuaBdIySb+iCRCjpr7vxTQOweV0nONnhS
z+0MIJE/hSixsKSdscJTd9CYKKv4DY26DT4Heoxz9vh+Ed5su44gd0DlO3a0JbKZ
6CY4sbmHTCmGls+yR4QfmTECtPeS2cFAuWqFteQd/NFfzEyPnNpmo547393KFNSL
CINa0qCnn/Xaw2OgBkDSmUu2xWnWJXqTHi/GO+lqkp31IPY0x30QDUYgGiLqdFX0
egh2Y6T2e9JqVhRVwPvsOXBvpu+BsxpJ2ZTOPpqCYRaSXjgbY4hD3w1ABNl0TYJC
folJODVZNpRXUhYESs6GjcbPk6v9UU21DwzpyDTt8lNrSZMuVHkdc3vt7EVds1Lu
yX3aXr6/DvvHNTSO675nJuAklcfGjUC8SWs8K7Xq312+TCwf473EypcNLPflGuJu
JyrbwE3xczGOUDx6Vb6cGKLJIv94hah6kLcUF1U6ik0xnYkGajbnLyixvIQ0YQKO
Al40tl6tq8NC4mStA+KWGsMXjrK1dk/duz6hz85567jMulDFyll+TXNAvW4qjM6U
ZAQNi5BXKYG/K1s7lxImBhg5agLptATDGijrOceZSdVZcVlOuIChrYEmjPUUZz2X
Bp/MqjayyyUOObwFjWS5t0atvW1f35JKUId1srmZE/k6nRI1nM+bNXTNCtEZlhyn
swqdZwIA2t/A3L19ouVcqoanpDlMs0Z99YMJMDqwdKm2C716c5WnWKfI5WXI2wO8
KunBddzOIQtJ4ImUeOBQPUyOc9njFQGIQo379fdy6gMPTYUEElpF9+3lkXPipYYi
kqSnS/NjVgQQKBfJC/jWdD8psyLSRRp3s3UegCpqJ68KYpF3Wq00BDkRVqG9ys/p
ahYsWna1EWshj75S2uHlVdWibcAg1J+0RWLjRTJn5ugLhw0xh0BZ5Mdvu5aY80MP
3OQQzJcMlIjMrsN+io0ax+EmFEHyW/3WtjQ1ruU4ZcDqONC78cr8XeGGWyt641JB
vdT3yZeuA6LwoLjLZAkubcy+ApAZqNTl1O1Cr/dXUi/+yYz5rmi7rKQokNsTCj+J
krfpwD0CzDUAkIDkdjUluADBzajv72DtaQBJZxDVWuY9yXSX8sBKVmdiZ+8x2s5P
SSeqi3iZcijELnnE0QwyoqL5y5UWQc1S7i9NAl20xIgu2oR+U1IH2e5TqjY2Cl0Y
ducPxAct1ENqE0vA5GZw2wxDnmVUjxuqJXHcMMHDmdpevu6BPk0/qjpl5LLIK9NI
aE+xx82lSP55b8ISEyx6VZmOnDIugKhxnEyAWhm3AxkyZmnBpyZx3hxa82vdUnZ3
MKCF9GgM2Sn3x8rFc36N2WYYfLf8CQ1jeNXZT3oKwpqJ94GJt/KH0ypSNBF9HZtp
/mI7v8CFFMWVNpI1DVGMbtS8Peec6HZOiy5k5xEmWIR7xnnhffB0IpAJkdC92To6
3Sz3jc9f+IsLjFeFleg9htrFwpRRuEafqtuxoW/sKSMFnR7N9y6NYYzK7l2vdEFC
0jrzZ/wdcjAIPQOCt5ci/LjR2hPdSwiL0y43Wo7dJnJb6JwJggU4FJYmi3gcBjuY
0p4uE3RJ4QzkwsRbRShIhE1nyWNxu1T0aH7XaptWr7gSphjVui3Y0uUYTtQuFbVB
DPjrN6jjGL5olRBdYEdF4ezhJS9Qm9UmgvV0PPP7ZciE+6k864LFItVL1fQqds58
FrOXvdbh1G8S+xPLMyinVMzwQ6apGWA3Gj3toM+Aw55eQEekjf6F27DqHklWK/lp
kS9oQI+1qFubzsJ3+CfdbaB2rq9ojI/Yl/a0UaXG+i+kB0ifCnBwAgUwGJgm0ymo
gyQp2FxqR/3nsnJDOqHhz5LNg64DvATt8fOmM5gYJIuwg5qheNhRoDlcMgwlUvjP
b5CYkIst4RfbLh+/L1Tpl1Cn6YgcDBLxtGYsWSSGMcHwG3vmXTFU1sj67sUbyvPi
rHXx+BO23EABLTiuG8ptBkm0w4fL6kv2ZYsSj9cK+ZNF0u8CCQ76f7qfRXah3BPa
2iBER8UOmn7coBMP4s7ilRlLaA8b8FDEIVScY2Dt0i+PEV45uBOk4kQmi1LajNaX
Md0u2QCWIcEYEQH9OD6vcjM4g/av6ujVfr0jBdzZBEyFlyCCut74ONLC3oHUgaeE
9oNuPz0cDLhtjF5O9mvsbLfKD6NBm4a/qsEvkW0ZfpJr3QWruYCtSpPyy3C3VhfN
aC+Y2Qoaj2EMEVweycfNrXv5r54hwlK1GqrgPg1OwPjXUhqJqVmTy1EaP/hFJvEX
3atJQ0lgL1XNew2rrMfNUgBjF3RyF4nhCeTQL+z0a1BbIEPneI8l7WgNhGzdEafS
J8a5E9yTPtF6bd77JT63eQCDGBuvz6MUitVCtdk+rKNMmUu6vsuWNJSkOCyp9dHR
zb9Hz+SKuFdrp/cwP9cPVa13UArAg/cRPod0/3+GSUY2kLrPM/Wiw+OvIdi5+JMM
PSDHfz5n1GoI/8+mNMAa+eKfsqS79sgfCoEdhh2tJwwxmK26oubY7+BD5HptqM4K
TizRXt+cRcMwWpi7GikMMRb7xycSUlX4Hto3VC9zJeAvriYLVRf9og/H884marPt
uDW6VFGOoM3KPzFKTAX1rvdIyxIK+aqxC8sGVcTvhAl2rg39V8CcYFmoqnKYjwbO
DOvWFjjy/zhkmjAluraH2Pa6IxGhWRvy2n3SxZuiz0CUJc3l7FEhjyMLCknR/ynT
t0EheOp5jVdncOuL2qdUfTewgEnw3WMpwngSt2ojrIBWXQdidoXEqVN5wYVySHtg
aCKTZpqtomeCHxzLuHkqKbgEQSqop9DRJqS0R7q7kzU07ylTo3I+oJCiV4A1zMNC
nsJj3WkN5jkMoJqPal63zxTE8rUXGK5ltW6yokA1hDCxc1ut01j8/OLbob5T0C2p
WKoBrsPt1pWmOynee5SnvXbtVh/bENGHTDsBattHRyLx76wPb1NwBrzxVZtzzDl5
5Li5M5UlxAoZp3Yc3N/DXrkYxR8YExS3gW5sHdmPpLh0aBXAfQREEsAJHp3nrJRi
na9ujAA7lSm1Tu1xVrIIhj2aRUPiGO7b0UKKP+RB7HYdVFUMHU0BScOCJRllRCzI
og1CY1ggNxKWfueRjEFnfjh33G0LQ4ODFTVA3B4dxqEl76lmt3OKjWRnAchMHVPB
AICQAHycKLs6FFYqKTRr3hjURlNgFTZ8qf1jI1ULhmzu8Yy7nD4TJecwo+snnaVR
ExS4VqNPwdlgfYQ3O0IPvi9z7EvQUwbH8dyyYxWrVuxOnVHHYo12mVPGnYK8vKBF
8AT3Utlg6PEU7suLXbvOlKFdJBgOamMWj1sVEGfxThnN2BfHW+pJo4zw1C27Hpdv
+z7DbjzPASPyLbBdJT3hrEF1wrNCo9ued1MOhEj08bFPsEutTgKjw4GdGz3yATKN
SPm4fEK03CUpWnxUvHgzDoytsKoW/ZHBCTy6Knixtb10T5k4R3BQ7Cyr4Z0Irb04
CkS9h+ugvSZL2TsfDmkoUdE+tYEoEEDIiBULyT+vlHhCRzQ/6dKe9J+uf3P4QuJw
ECm+2ACVIS9P163tjfiz4bGgkXGgNOx4xkJpaaQF2vLoWZ3qezRKVse15iyKhkNj
ML0Vgd99Sd0usebpMOdRs+FuxBpL6Dqhe5owe6AiDV+enfEL/rOJNYKjvCSiVHO0
tSEpoBCaqkOlFuE1/z3YRdTaNAaPEuWup2NibrPt2diLZ765Y9cDw6iD0boBI2p/
cGftAqX3SEMk3O7cIHvUI2pFA1dbw3nKAwP1h8JxodJJNMHPxbR25UO6vee7V+y0
Q8/8Jkktvnc9A2XZFn6viwd/opHtl1ndV6HFtBBQAzF7TvCyWjpShsqpvLNMocdh
3ZrXJeIq3HB08d0thYWN0wUzCt+rWIYHtie4gXtEu+7yMj+eoIjhGJIHSTkRmU0m
w28oY7Yg/GQwwRu3+/0n5slZaNb0aahsyGQzu4TToBzb+qyyuyKKpdulf3OJWd9f
3jveBcpsFSkxoWNgmbaHV4gaEPRYMrwJTSlLcBRTpkgw8YgxXhUX1VHm9nNvTCM7
sPJd6jf/gIw4BcWI1u8GGmcTf9fC4OXgYBOYxUYkXJuRgsOPjq8eR50SPzUJvF+4
4kpeNj0bd2RcxlVgEjSYdcAp12m8RgZt9JJ3Zdvaf0M71xvO+Ay59Yx+IsNJ1wYH
N1ZJpI2C/gR6eSZ9tfz/CiCnk5hyY+jz2bzAz43iomADhr/je3VKI/JM2pW5pzkc
H6pzcMOy8wNKD4h60Hn2u3w7rx1JL2libTRdUNqb0LaM7yjYbMGPXe0nP3P7Z4rI
ojlUUAkWFw4PkxkcLvTlDpSnY3/nPPIbDs8u2tL1D4zYXVc/y+tNCnno14C7NZex
gTtfEd12+clpcnPIPVSNyrjSyuygKYneuc4cCN5YkqtzDCHyy11Xh4U0Fo8kK+6i
xtB3F2qimmFNwrDcYq4ULH1QetGfL6nf/vOmJnIVpVHAxLr8w4czgoBuKhFKNJ5+
8MlTPy9pikVuvgK8RBFyTpygX0czIEF06IXwoEfb1BGcWa0lfaYDnGks7QeP6ehm
Af9hDaxSpGCh0JIAhynCISDSpPfpj1dplTTEJcKKnJWvlVd6X5AWDFvABSLaRtWc
TBXa9XeE9gm0eySeFQpGeEy0E7hX3ufaJ3eNYPmMzIae/BmNU362JMA8y03wJMGD
2HBBC+C8OZE0OfUwUF0R96djpFOEw/1Juk1Ir8IfPH3Jff1P3P6Sdx/qgIal05S3
G7GN5bF8ReVCjb7fXhXxhPFbiFyGlLFEjYez04yNwHhQA7FKAM66UlavJbmfLf6I
QVaZ63Hivodv2Pt5QQ3N7FNQlJLl2HDuzhElaVRbsZGbJoKD4Kpqn0EX/GZYgRZP
I1gUSnjxSfotHkA7fAJuOWl4Se3QG3/tZTl/6BglcSZie9n1v6cN1fDZxrKmjpY1
ypQYNhHycUKE8YUktr4WSRSdXyKuokf70phQ49NnX76aGK0le9IwCcskvdVQ0yr2
P2bdv9iDBvon5dbpMdVJfBfllGi9QBzwTzhNU7B5MyrjJYO7wWgM9mevDRdyCAHx
rtEnZLE8kjBAX4HYHqf1YF6ZoO6E10oXvOV2wu9utHlD4A5PUtRZh1OCyEm/Rat7
0JWWgJbf3reRIUrSVBvnUep9SHAN8bzJ9wAHwRtiNOqLJOJpvsbQ+7Bw+cYagSaU
KtlPoQHxCc/0SqJLXE+dw572l/B7zuLlizZ8oKph8UNtMccWzmpZu5fTNNTlsyab
m9x1Qn4Wy8e6ujdtkSqftwMmJwdoLiAidBB3PCZOb/PcE4hl5kNln1KvPvjpZ3gL
QMIjGuO/PK2OcuCSdiHjkKVZxZzzpoZynXN5GNXvw6JDawhHiIeS3S8CMMX43EqH
UR9im6frq6yP/tm3HF9K2lf5kuN3AJJoVracHk/1+AOKsJUrBzftTWOmcSqkGBmM
45eRB6Rv2FPv0zF23PwDiDhEetwyKy9ZLtXjBE2ZUYc/XQfXF5QjjL/7PV/vCpeP
LldjJQ8NdLRQmMt0/ZIB2sZq30l/c/5f63jpSg73qhpoTW+MIP4fuvIYxaPz6+Uc
gg8bdw3P1KGAzOhv7mIbaz5TTd9NZY6vpqnyUaiK6OuVPUpo7GTIYApTS3Ldmpov
qEDOkEMC5syvniAMhzdVrsyLjyJueakZSg9rd0bXqdM+gHFoD85TZDUI4r9j6m+Q
HB5Y4GU/AA9iH3mBcVYA6RGfZkwLaXikDL6+zesbx5fkOUzDHExL5zfI1rONcvGO
Ed+N7flB9/cHptmFltNIXX4wZ/WgIZoxqB+0AEruLxCTjorThu16cGf3mozmj79m
Aup0LZq0rp8N+OTeUZjqBn36tX84HNftJ+7NHftn4bxHpuh/6DAuRrciwiQxI9Jz
fjqFgPdIDHWSLDpx5gX9lko6u+WNTKjK8Z2pc2L/MP8JmZmI1lX5lhHKI7ea5ExP
EQwGyPU/7/7h82N5DwUzLoy1UXUggC0g+0XRaStXGghw2BTzQ8yKbY8czsmKBGBH
K+BCOVfMxORGsDZlaufrplVQpIqykID5S63U3yp6VZ5MagYdSF4+Lq09lrNgz2KJ
rqQv9gAQCHaciiU6Ge4ul86RL+Rl7smxxLVOzspFj1Zow+3bKXakdwoTcFKAecxn
NN0CEhfuDLfoli5Cssl/Wl19qxSsWJe6EfcFTtF1HhPA15oM25ME8h2o40snrS62
ZiB4eoPELdTBxvZIWsvKbgi2cZkoxr0peNZfewzOwrz1x8cqt/rLqA29knMl3mud
vGSlkApbeb5Y4wmd7Iy2+FOKAWBlVzckgDRH/jLMdpNpowr4+ncig5NR63TO2R1c
F/WWSmCYD60rQN/uVu8va3C2izIs2etYIZtH3kirRhoCjF5EkUexbaQxGwMW46wB
vu8auVurGvY85La/TRNfuQuxTrIFHYix5Ib4+ggb9LsoZeCYjfrne4dwKcovenED
5s3HXQ+YFFg1CrPSncXpGJZDc9y+YlYNzoFMnxxldyQBun6obMjnjj5TxOjWef1n
aKVtEcVPG8PN+iG8pkCRaIAQmO+PwYL7QIhO0Bsi+OyWBWIW0rNgHfYyCFYoUHve
r93VEmqha201/BOQwOz7fXtOurL6bicW+ZD80nk88cs5QT4SJxU8kNo9YYpDdc2h
nCSXiHNuBrV6WghFLb4ihPq8RPicrwH8ZszFLK0fBxBEcCuSgZd786dn+iHiP9Ck
XBlLyEXBEtJ80cxhMvLODZJiTZ4LMW7UTXWihj7Ua8b1pZmBZZLEHLa7PNL2Pbzr
Iha4aEtgLt0m4CzVk17elTdGMg566Iwl191rZm6eFYzOmDzGtyAqUir0/SeGCwkM
OGusTPtZIbSAQ3OsNf+DUv+uTrulkwWvhXkwmgKauTU4Tcd0KtrUxYeJ8LC1GwEy
phxlkwpG2zG0DBBBCdtc/NffTFUKKzeQ8qK4saWquSg52VxlVywlp8W48BsqoRsG
hIuMXRaxJ6m64v1JmJTc2RjJbPVzNYhiyPlr/Fj5RWnphNOyipLB36lrmhFF7c6V
acAAwH+X5/qo2lR73OzXsO24rYrnf0THFgAqHR+JkHLANZMLohM9I7PhFeiQMsoZ
2Owx/kED7j+jxjHPwDN5ZyqaE7e2KLJsfbxdipdYlkE4y/256XFuCwTU3Z2qFp62
txcCJ3fDZXipQT7+HniWihBIKDEXYuLrmMCBnHRm5ovjDdlryfcXUrP1oDrL2Z0d
B/qquHWPjNM9QTFv2FMi7CYgi0V8zkSlGWK+LY0O0b3KgbQiGGQ+FNdSrhCRnKbq
yUYTTDF4EdK3B3RuI2No0niHHyTjDOVqK8O7kpfqzd86KvgyLCe8lcIPnTKxdxIs
PfvM9GzhsB6a9ok1GwQtPyVAZrI5+VBjK2LbBhDXABLbzytCA20fCegM5yfApMlW
xfR2xlmn2x1NK7F4ekGqEgr6ijlJzZ/1Z21ofPAS81ysMOjgEIbEOO1ItWx8cuze
kBSCXdazDxDvEp5oFt3F/THM+Om6M4cvR9N5hBTqCrX8CqwVfgNw1KkTeT7pROlB
+0Rws635+Hrj2IIgc+aeBUmVIa1iY0zcCmPHDwrNFImKicibw7IzYDN9cgvStN1i
YFkgrtb3xaBVzrPw+lKr14jY0C8RumhGej9t4eHkyc9K2lCh202utLWIaxRtppA7
xkacW13stkVQAPI40zong6Z7YNSvJPVhu6iMGOFJyz4XDAr+puwE2LoKZg5A3bMT
qGje4sXh+aGtn/leVnqB0ITnWyJTaCr7mniCYfzz+WqzyniQroQ1NRWbpM6/Ja0S
CgycMMRvCUmaPEE5O+WQTQCJg7hJ2kadfkuZvv4Az91IIZinqFZmHI51jN3GQdTi
/Kjvqf04DpiWoi+4a/5DskrC+V0WJPGvXf33zvjJjJLLQM5Tni5UDcb3oOx63jtB
kuzr9+T8iVW5nG9IzDgcO7kKIu4clYkOej5E9dzRYtkMk5Ap18V2H0TYeCCIo3sr
PLfYJ+w4ztVOvTs7psDpjrbQex+sLuNoXGHmPK8t+MT4YcmXNb/NsDAVuaELt7Wz
E766Ci2+3DBXC+xZcqLl77XTq7IyYlXHe78U+9nTRtbndGtvcodnl+j0LgRR/tsw
Gbg+BADO9tBaAexUTwTTFcECgGs7yDCM+YW/zjhK6LXMg8YORGwZ208iQNIcCkkq
D9PVBZbtikQB6CeMLeGr/XpsDyfJ8YGrC6orAMNfu9Ko7xVqLHrmBTLcBASbt6Pd
crqn4Ibs+DZ8WPFyg81Z+q0ChmVtFdy+TQLCacJWGIX/9msULXmbL7lKUGhTu5dX
vyfeRG+Ji2OjchofBts1JwYij77ZrcjzMiF/YR1a4/neQcGA98oz2HFhDTaulS2W
DAFUYuECX+MzqIKBXGIz/W5zzm8YRNWfMetikr39+n3wGs/mOxyDJsMvKqaMnUd2
cD+I2HKtjaQDE9W7aHjN1oI0ta4zkygItweATspLS66M/otaFpDeROeNTS9ravMH
v9+b9CAkT5TPt17g7lj8/g2PvN2WGndvvHnGuffXoR3PRsevZSssIt7HgAAtB2jE
pQLZSt/qVVdcH9zANzmEqPzf54VgtoDuePcq6QkYPndmXCQ2+NPpucx5dokWUyUH
KWmTqbeZ5CTzXCnsPGKJdcLBlP0s57cyeCOptGX4L3KEbndGeNnjtKgeFmKuSfoa
eGAsq+fIXxOcqs+KfnIdk0oAUpiqP9w7W0bDd45OmOwUVIr/9e0YewbqgH/363BX
lVB6v3BG1oDRE0AFMLXfhmnOz5Dz6xl8lprr/I9fFq61RXg1YOsBb5zi3URgemuf
1yThhwUWyzfHf8brAtTQ+VGpKnPudtUR+j2Kf/jNc/h9wNT1+L8T91qrGdoa8O19
yjIeCxIQp4kf1bgphWDYEn65Tqvow0hn66nFr1Cbr1NJEvCVGo0e/UR9p5i6KHOB
A0yq153V79f6nzvTLRNfmac4IJlMdYP8r/Cq45/paBxnE9m7ms9ew76lzpsXiPC2
JrLj4rwAK5i77bpFx4K/VxLbM1aylohGmRurZ7Io4hELdRb0vYCff14w+sbD9/jW
v27KAbkeRy2MN/NPAGJwyVsEWGYrGTFflKfwKjJrBgejOhztJhc5BdPX7ziuoNta
zMQ4Ou93U8sQPNaH1KZ4lL2vok8p6xK9ngW4mR8CFnbizTvZH5lDOXnxQ8Fumd5W
H0fZmpHp6np8Y8kQOdp8x+9RrkBLtbpcGP+85LtFJFFY/h00DIAC8+BDBIkE/3OK
GbUobH7GW5kOw09blgasmRCUz/vqOq4k1/YpBBxLAMsKMj+WthtsWbknGqTB4vNh
7jzxrLNXVkCiPwbEbDGPJUTaC0UV7LJk9iJgG16NxKxN/2Tn0z20QZEBrEBEevC3
8pnhNWZrES0yKhaNQzJIDjOzxkoLbnvOF+9g/umzzIjDOSMFnu3hDbIfRycP6KMf
7S8eVxHbDLQEJHuhiQaSgU9C8FW/C0ltJi0jtYEln0AwP6wR250T7FPCGUSBQMc0
TiVtuA6Slb5CIQRF/42S2izHyJSTPdYTfqX/tPfL/MGQuKSMjjiCOVccXkZn4+j0
cQ8X9dAqLR+HwUAup+TC858vEb/bmTtKGDNl3Av4XxG0X+o4tULTvKLe0o35QXnU
hMV9WSBtJd48Xl1T/rTwAaRusaeQvorPR4DeDsLONupf9GF/bBBmDCJaQPr3kh3J
5RgbLYKiy9m0HVD0mXWvhAv9+tnGsOHO/PMgAkm/d60Mns7lp/2LJgIoGleJ5R4K
fXtxAt+dNVVazOPW8BEE8fWB/08C5Nci0eQGmTO35hlK04SyThhqDxXITrKrfz8f
jD9cOu3goZQgOQ7YOIAqAf+Yue1u2LvIDlo6zXWr/N2Y+030kE/L9/WyAwucUpHh
AWQdvgnBvydlYn4Jm9EMuXniyHjVhPlluLXlqxldYx9rWKEZfJWe2l0ugc+2ilWo
UZMdzR+XGVG7h6q7gtF+UiWriztfOsJ68tCquHnfRDgjoVf59bmF74ybKPXDzSh+
rDHLhaopnGwFtCK4aqsaDvOrHVgCjc67Kse3bTdxGpx2/pBJWn8eTwydOLZRV0Pn
y2nVgdeoRJxlCprZwtXLXWwWw+4nI85deFt15xqRihcUb536K2G9ZtZdJY7gjs4R
14KAsZp0ywzEVxb7O1YAydXK6ELaDvFfv7ZQp7DZtVST5fynCEieRqCtaPxJeUeX
uEtoA5Kdt7mY0nz/1BouMchbzC9geu0qZpwav/eLtEpfzji/kyFS96PzpVCdMXE8
WFq3VWu06MJiU2sB0a+36cuJU5Hx6Yaqpo7prYYtOoFCLuQuWKazyo6gPLiPYrx8
t9Sst/CnpG1WWsaV02hJXIeS6QSlnht9yOompVOhblz8CC2bM30AYMZcnAEKWaKR
0a5RwH73Mwvqvcv2XbHrLAbXglLPZkJNPwYXfTiMlkvfis1AAtHokJS6nYaz8N+S
dp7vfQkElxjUJOdsJ1bm5mfXTde/3p90wsMrOutqZHvJNYRoG/DeyDtaStFYgY+X
y7LmxQ8WwUmnM3pwosf0MSAGXE7kzfdvr1W1+drTtDw94RrdETROMV2pD0pdXC2c
WwGGMQbv6+CTEkjBzvHr4mAnDEnFHQqADy1b9d2a/5dnNXgGrTunaQlFMq6f0cXt
ouNVLbiSWRsF0+8ZZZQk238ZzjnKnWorG2fvzClw/Lv6Mt4uPIzMsiywxsBBynKD
mxP7lDLwRrqRtIGPtB4zC8KM5IOz5L6vylbHmuiT0vf6OMbucZXbsH/YpQialp0l
uXw4i/Z+8gdHTkWRpJwQVP7h0nQ5LCfYGVA6o7YvRStNwtl0oxPK8alDpUysoh/I
9FrDVB1deIshIsa9DaqkQuRNHd/7dcDX7NRDm1WXHW6i+l7YEYlYyBzdSfhYZ8EF
E5oegMdiDmkuQ8lo3olvQNFraHIFsDrdVRKlYm8ssEN8Yzm4Ycz+Y5UUqPhkR8TG
i06YB6KjPgxbf/CD4vVxwyutuU+SO4aTFsPRSZJCSUbf7MFb/KAkQX3xW6sjmO/P
9iFs1xsHqoGXurVsXS2byWB5IUvJFIlfig4ApIkKOQLeoksYg0F7F/Rq/1N4X4Ua
slQtHkFMD0uNOXGbwVkIzmmATLc+t/o817gSAtMp+/ul/3BKLwwC8S+5U6jbb5A7
otX4PQp4sFnA4NfWj1E3CAAF8bClzBVeqoFLG70/1xlFh8yZkdCXvbkm/3s/auEA
a9sqUUPzh9dtZe1uvA2e2KE3dc25DS5RZzl7rR4SQoD/GSNPgO0dezwW4mvCW9Ef
EC6acQNnhxFwGDETPK2wY4PT9hkV/sCqFZn6S+TEV4uiBrEqRzTa3jqWPPJl55qg
G0esDHP+zF0LIKcJz0om8IaiOzgfocu9/wzrR3T/k8AYl17dBvCLDsvam1a72Pmy
CFXOyjLml45Ywrrb6eqJ+a6o/amq3tAg5PYcUwPdYhVG1TUPdHUhSI6RpuHBJ6b7
rBM1N2bKV6qhYAlqjXO4RhNwRWBhOLUpG6n9Zejy0UE0AeOkn171OEyM4aeRXGW8
H4rNwJdvpcYTMy5/gbV5NLKNp6z4LXOrKpfKOmsciPoODbVXP3x0cFiBEl29WgKe
qVL79wl+QBSaLlDlnZE3B2AcffvHGetUBFczG9OqWBdNnLQNmx4K2p629ZY/Ct88
jFqAigU6eyJrO1r96z/6uVped1m1v00tS/fSXRpZcm/w23dtB+fUUaglxVnReBWy
9JvcDw3GlMf5tATZQmBzdKtF7NHVA+BI2USaOHd6eDOSXRFW3+OIy3BZk1M3GLPU
Mcgj3FZxBbgj12jQisFOTxw6sK6luVmaU3kTqIM6qgPxt1acZntUKPoaRSBiFXpC
O8gXznJoNGkSvic4kbuVYtCeLXbNT6dJwdKT/mYJZRl5E2IXJmoliSvrCMUmqhK5
EIQCCswEKN36tJMD0d8zCyG/sJz1PveSGs+bZJfHROv5larPRKNQjRO30XmOR8y1
u88lad5NOs2Z41//Zti2YGr+SaVKLBL4oqVXeGtd50aztoqR28fhyMzAspio7Wlp
ChlkVL0IK2H5snT4cz9PecP1g+q/QADqm9pj3wNkhMTVKRs2PoW58vt4RnYm3Lz5
a/wclG1XLMKGbzabD7IcJqt+sK+7aZDCzP+N5NiGb6Y94QoygIaFoA1Q6WAy0qIE
CU4QbQXpVE7Or3GDfNJ65VZTSCR5MBg81PFQpZ/lEWZCdYbhDEAe8rAwcOwHG3iI
zw9TtZej0W3LJwYm4kxHt//tDt5fpVeTYiSxypVvOHHPCGZ2WXIObsp1qzjLsEkb
kY5UnApqGuKadlSU4phY858pYjPd0FogTyt740YMYKdYEy0pE2iyFxwblXrJqoxH
4bDbaIeD/t2eD1ftGgnRGUOc7t7R/UptRcmDhbb/2XaUf35Mci/Toh9Jfk4UwzTM
nGX5WAu8ovIS5I6TK4ByoRsPj15rRoy1zu798k2ehIdyU+CFy1uR5QD5RSaCz4Gp
vayASOARo60VDhLCqMviHBjDKbSazIO4FXuil2KHSQJ7rg+nuviabcv8gVWdBzhv
945op/PjewWsV7L/8//XIUTLuz9WqIsZaz7g6B1GYfqygZNkvsC6XpP7zuNUScbw
LC7y4Zsz86X3FWONOa4w8tND3Xkl9huD6vE6TAfucO1NveOKNft/Ms/BzTrgDkeY
CHZ6p31mQT+4SA/0AYQSjhFdHFyAnwwyAqsRai3pw9eVOdsvIpkUioBAWxoDvUrg
kw1P2sdtT1fCqmCzgxaVLiVY90nO9/SOg5+HZWNo8YucvddDIfBc6buiQpqURei8
C826qr22ed6ng7rK+FU2/yrFHs/subxT8MIh9c2q5CTCR6CczYnZfksN3s8dkCLQ
djJW+o+XdCyAcOOeF2Dvl0ZuKhyjZ9/YWIHaIsLGXEE/xeTvkA5hAk2Nr2ckXiJi
z3/Py6ENGkLSUabBLNBznjJKbZKpND2eZQTyuQeCmqzPuMqyek6j4IBXgplRnNx1
aO/jVTM65K/L+JQ+6LYIPaWpYhd9K+yK9OamUSU6BnHCjl2x+1DSoSJy4xL2bUMM
MwodnzVAoj6Spx0wRGfZjhEp7QC4HxteAP2h2ZdIonD81G3gXgZARf2BoHEFzEwA
EMCuMT7xV/anzVFC1pKI9RePH6UYQAH8vXvWljz7nD0vqFP6VnQq/mCE24YotuTP
0l0J1CkzrBeq0D9GrZsDQYWHJQFn+gbGrnwbfxrRsduUbE4cMCygPE1C9mEGflIG
ylJTIdve43qwkecJU/QLxMpp/WE2owCoL7DamFwHinr2qTELdz/t4MSuWE7n//9O
WH/esIT6SJUfIJp/9H8My4uPeCYaK5LGcKaOCx/jmV0Zj/3B2So3ifDMvbLw/mAO
iwoAhbelzUgiiRs1nZks3nRhnMZnWjunAvnfcYDjrpVy9A9aQ7gdkI5psxc+Ympt
cwDSKn7xeIRzNNGsPe4FPbUu7elpiyDLrdnqVPNe8EWCpluCni0CjckGbicTChbR
6TiowRQQ00N4EchqeNW+807kzSGtajijS52Dufx2/Elz2iAX8QzWw98LrfOV9Ecf
WxHePdXfNhmoGUuFex4rIVPRtQ52KgIE6gLrSFJJvXmIS6UNszRTlC/72yMuetpH
4pi5Bdv5tnMT0R8+BohQEzVQxUDKZhbLmSR0z203Dp6Sn6RmLH8h7ax0ehO6JKu6
n6ziqPhqka1e5vXYdo67ve7sgN5rGCnzq07ECkrN2MUInJ37xViGPTtRod+m1zu3
KeUnm9dW5rP8pl0u7FByq8gmRxCamrVNAkk0we+G8rRcpyfOpxzA+Mp836cpQn8P
p0sLVUSWp7KEFUBGzCigUB4ZxR0SIMyXd2rNNJbjwlfMPjq3qjm9R9PE4tu0oHIa
pDFgZUAvwM75lKdC9iWlsDOR3UvoabdHkNoBKoLp0Lx7d61Av7wX5tKC307lDMDk
nSKzMT1udWWaIN5bO46sztZAZM6SJ9XAhOI1fjm45oVh9fXyVPBEU7qmjN8MilH0
f5WHela5S2DQwevr0R4Q8K2rk+/+SksauU6+kPh8UoP4QXu6RcKoDIazQxfGnCE6
4ZqnTFb4ShwRjEHuXXnSNhXdIIXs5ktiggRqP/LMDuV9gCWmDlo9ks4LBPlO+aSo
f/cs0WTCL90i/R5yZXL7H3/q1YUxm92eqeNLfcY36kK3U59zVuqOx3T3MNZNmo7g
Mc634NTE3oIGMN4agGoq6WMDBYSINH/BZu+GhpC4z2AUpYq8fiNx3HW8EnSDDhS1
HcGMfhIko8hixsSoF2jrppLaAQBoy4Qupa/DP8C0qeO9pnbChsSA5yzUv4dUJNdC
Iot5dhxp78oqL1xZQHEaK/VIotaWDyD1P+RqeQ8IJlI41YfQQcnkHxUB91aH/l8i
SceknqymHOCFIXKfxFVJNpqlfTPFBPh3fwEdhvSQaJ0NEDcLwhufclxIrlzx0N3m
V4JRiTPDbP0hgFg4+3QtqgX0H/synsJdIuKLD8YQmZytUxOhfOfcu9NUFwUNa4Gz
MoQ2BJB+xmMr/TTEO1/XMsaGv2awGV7rPp66kmXuTW5cDZo+XWeVGHphcSI3xWyP
PE/rpzH1l+F7Azh4YqlvP4VnJbdusIPK78sAiMhmzurX9kCv16hpebeX7sNoLJjQ
jW1L8UCCfMmpIhYZd/9ZDDEL29qBqr6CClXFZvpXl6xYxLjsfKPN8+WkjZJvzxNQ
Ycp4WHo/BBhbO0C7+35Tkbi9CDxrPD3Ocg3QpKepnWjeHISGwsXhYPJGSk7UkJY1
uQrKgBh0CWyNFUTAE2vP2JDMoasJ+aBkThqhH2ihVyYsTTWiIDm8qYCB0S4pI4XV
jkflWKk00sdyP71H48bhnQFEpLRWTMqIU4Z9GLhByRIgcZnI6OvJp158BR+Z8Oz7
bbU1uyzprTYEF9JJxRKmgITNK8uRAcbxK79IDciCy9rD+UUuYb0Hh+3wYGCYl3B9
+jwZjVwRP9bSSf+jl87+nnkGoEW/GSQ1MyzB7uawKfqEPVmuGrnVvJMg6gYPTzdX
FhiXISc2rSakDTNecsP8mlQhUKKA0gGLECyBZ7lI/+Qjjd+5v48SnDRq+lYxf9YU
7k1uvRGcVSznrMOIpNN4xk3BoxncNjv+hK4WdKLZ5W/Ru2EH+pe/qdOHn3IQfjH1
K+wbKgc41pSGqxRKjRopZy/7FxN72/+aAX8QFnCVa68SHsDwMowJu0T/ybQmK8BU
DcaeozUEowNI3QJX2g9NdwZ0LYdh7i0pxd71OSaiAl09M5V3zeZ7GaqZ8OhPlCEB
bWoo1CGLW4EeRAxOQLsS4L6N1yJYEOz2sBE0ujSDPYqfJsKF1xMLaNdKSqLnHBis
CbtH9jV1h/8VxPRfiAWMbX+DduCPZnPvyVKCd/uHxpyD6nSJJQhKSvUcCpqwaBoJ
7vjzDmzeLFtgqqFcp5E6/tYMeAyPAau6Wd6tICzcDv1e7je4jrcxyUFOkRJjXfi3
6pS/Tk4oDQXzRhvpOF5HvZ+a0SvuMUs/41M71qUGMnhY4Xl4nD9w6s87JmmJ8vGY
Q95zAMfmvTF4whjSzTAb3jdKx7J7JPEiX2mxO8zfyi4iOdUGWpKFYlVD0Aa2Kq3F
1CWvPWxshux727Gfip7yUUVHOt5AFvveuD5TTYCG7Gu4af5706y3yOwuhicA/iar
cPqzcS1TMGhMbYVLnsuvL0fTWSvoTVb9ul2hVT/g6ioeFyACruWUmWmwYMA4q1LF
Dzs36QGEuAY6pUzV1oBx1WJFY/Ybw349AQnSnb+Y4iRYsa6mJO1+tA7r5v+WonDQ
qPoVjZjHGTid1QVfu+BNeYv8r+lEdsu/X/VmhxA+mWKbqHgiUnh6E/5hUFHc6LyH
0F1lKOZKPQ4cTB6Mzly1NJwU1mehCg1ViFu8vDPkY/bSyT9smBMU72t5vsK4O2yw
ryMf3BQiqS2TYbTv1/XPpr6pw+RNI9AiXxMp/ARZbSHXfnA2dSYhlYg+XYRc34yM
qLfvdRFXYoCeEtVHye3DCQEeNtifgH6157bUZ6H+1sxCknR2J+L0BfUNyw/qCI+R
K0bagyB0OcxE2oOcU4jDOY3rOyiRpyd7uvoFK8OPqpvunRXzWHAO2A27zZ1Zw0fx
U09M7bwNiGaYHCC/0LJ5p8mQtOBR/qmvXCo2bJmYCkVbuT5rP/n6cIG8zA8xJleb
wqbLRXJI5ReZ3pmkxQzm+pE9cpQEcnbkm/L0Ek7RT75P4FbRPbM38uIZIAa/qNIs
sq/ufJF6096NRjLeIYH7dI1dXI71LurMz6z9QPqqLfIxJRLZQZwQ9Z9c0Yplgw6i
mRG2WgC6N05qRlBgBpdYqZrbQby8EhEiSzw/cCCRUfVa/ghkaG82J4qkEu2IDqkY
zPwZIcZKjtDl+3wVVChu8S8624AEgpdih1zHMXFBjnU4qMaLLSS7JhbZuy6EboGR
dK95H9DXha6gFyhahEWsLD0rEPnt1lvS+koxSfIVZQz2i6CRIsYlAYbfCGNWiSYI
iI3LFl3uDhOFn6USl3JdtTXk7FIPff4T4KhtY+RFbRTYmg/UNC65YG2LtbUSAkio
po7Or+BbSmtVecmrEciiVkCcyTtThmbR3OdJEAuCxDc6OnnLROjekFORNEp0mlQw
nSZaZRXvtv2cJdmXl7IyiK3tkRJVKsGQK2ii0o8E/d2OqRWdcjHHbsgrC89/F2cS
78IdaA8CGzk+f60hzCtxWJ7hEEz290qE9iLK7v4JweFrcmWLs4gyrShq7DfSy+GY
TrHfroclNLXxF9LXrMOMJh1u/U5EIDduR2J8pApe2KZWQgcqpqmsH2Ry8GqMYeY9
8trXyVID4S/VLNKpXQDsZdMA9JE1Ih5T+aWceElUYZ7g3FQ+PTB+l+ljKmvy3mTQ
Y7KPkgo96xLXweEDHQbGua5qIB3OyTU1QQE9d7q2dxa8rlDAJkDzeEKAMp3HBfKb
GG4Rr4GMD2kU+VNUMBj9mQovLj3EfafdnhvzGSltUejlR6pN0EkYVSfgfDlENEds
BtRvZs8LxpE/GMTXJV+s1nBLTqa6yGvhVK1iC2pAky5WCzSGmmI2Cnf1lbeyWoat
z1Kv6j5dwIKKlciBWkl3IXex68rfQmeNn4fpHu0UZugA35jqxSr/gqcgdHfBywzI
KSFO9u4CzBkOz8rhN0FuNEJnmd+U+6F1V0hrJDnB5n+fgKISJi1/Lr6/UG9rx3CP
IZy3RELjti5Cy5w5A5WUpGWvMqY70KGUjAtp+LUy0/Ia+V7dFhE1wsiUAW0/JoPn
ysZjzZa9BHOEwzhSvE8/OCwNB8dD8/I7S4NMyvV9Hj078+0rJSUuX015+OOTwIl0
NNYLKGmM7Luq2Z2SuZ1F5YDp7+DBdSO8pF6o6PPxK0RIw6XHRsk6q3PTkcD8/Xrh
qf5yuTWZhLwJWe4VNUZ2BOcyvZACfH3kUXD9coCtoPdPTRQE3RFAaiumvdi/ew8I
zLStncq7ORHnzjHVhwEQ5C3xI3NwzNXD7+sNf+6/XyAMwr9jGrdTaEnrAwcDoKfU
nOX2gfISkHA0ogk2v1B0Yw9sAj1QDvQo61JMuXFktKnONQFJIVgO2SWU/RsCIiPJ
ULb6KR24Qx8JlK69geIj2CKTneVy7yruy+1Q2Z1GEsDRp6an+upKQeaZb2D+MN3O
iUajiRjruYVSbad2U9Dgv9rv754Vbok3rT8czX09w2QYne4l5x3kcIn8O2mwE2+E
EEj7gDArrYVBBBTbzWRLGfh4Tr6NSjHRnosMRlcJHC+I7ThQQlSuhil7x4odcQpF
n1XGdhRnhqsIQ3EBLrEaiRuJgS84RLXAOJir1EKp6AlAplM2pBHrrGEujc7CB1hS
5akdO8JlhjCPUJFY7JXxjRspR/ThzeMPwhT1h8+9pniff/k58gsJD4/c0LOu4+Ax
RwWL5Mx3JzkT5OCeKbdRg09Ln8iNqxhp8CaRRYRklYg14I/PgGDmmTl5Akac+dye
PTTw9GIDTveZ071v7Cxt2lrMCqFDXkLOQioQ2YJG6DDiWih6mlQfrvdolqRJRFAi
/bDGMxVFpFjBzOozbakig3wWek+IskA0qfReDRQtn+22g38/tXP0CS9TXZG7uljZ
yYQk/b6r0B1yF0Z1E4/rDrYILEbrjYB/q7RO3pY5K/HgcqCvE7dYaD1piYJaWMZo
gEokpBqqem+5HzwM3TjVk8EbHfiYshoty+WoUQZQQgEGLSKCaNJ+Q6Tna2lRnpxa
idiYXJQcypotxFJWKpPNVsCHo0XjMve7R3WS15cb0pEX55pljgaeDCRguRUiObiS
AldWrHxX52FWW0rKpGOl5a0B+ETQfpAzclaqgVvpeTPe1PZk1SzGOOufrDYIHQLO
663osn7H+htNbgrOkzFA9QwnGQUdQh2zd/Q7xIFLIVJEwVbaMaIr6jL5zq9K1P5k
D7/2BILtOF9XOZNrS2YDwC3eJBva9mQqSEZ+xk0K+i4UNCcDsuJIiyG+0KYbhxyF
IwRuSixR93s89o70E1uEuB5yIzu5S3oUCtQmwDbUfKGi62sZeoGG//u3/vhEaMw8
TKPoid6njY8+8GR8oH30Oqc6pVpJL7uF8yc5YGe7H2weapl/tx4KTsGW0Jt5H4F0
6J4Qa6gZhu9AL1MdIhJSRWAlgaxXK6f0Hd4dPcjfZAXkF8ZyzC88QzVEgxClYb+O
xjmZWqQMWGxwpnqE2+doCRnkZrxgrDQEeQ3n5vXBij5aontBg83SkZEkjtyZQNMk
2xwccG5fQ00UIgFGUn1n49RAwIMlFXsFO38KHS9rIjsgUkakHsLt7kZYihU21MET
95GzXEN31z3oze/uxvyYOYlXN5WydNu/ooTJKPmvyDAPXvyC2inssf5ayBrUzO+6
7cMl9WY3U9P8sZdWbVkmaR6INgCRos7LvetPvgGKuQNO3i9jCNj9f59Bmy5LgO6l
L3RsaTfcotR5G/ULOr6YY+KM+3UqLVBThBl4kqoNNOTs/UJYFddYu5Y7QcW7TO9d
7DI00hR2L7d1cUzT0CCleI23pRlqgHaKckI9eHw9ntoLUmILfuT/S27mkotQDCya
NaCbpyQuVC5S4MhTFiiPhcU+gOqCa1oZePRrOHp9SpHZMOc4a0otTtcJEO7tVZ2V
nNEGTssDCKlYbqapsppEb/TuHShwomvUuQzvu2HzyYlR00F3SMRsl0PCKBveg7Jq
H1G+OjCNXjPjEYGQ7C+b8IrWwQgr9WnCs77F/mVZUXQIL7psigmn48Ss/jpGwByM
sFYrMqjes/sKF2J6antQUmfr3nDCGq81IO1+hLYWQF5ZrB9q4qlV1R2TQFFRAi6p
gyQ6BV8k0LVq2rWLQk0XXfoYyNT82zq1Wy7ZQ9skc0xdjr3LnGuacKf7Mjhpwr+x
0eZUNg9jCTqUcIP4P/T//heAY2w02Xo6kpwqsmFhJg0B04GaAHDdM9cBUenO4/UR
4a1JJAJ3Frv/rdiSrrRpNJhSTsuyslpO+MtTsTsmLUbte9zzmSgKQ86G4je6Dl3s
1PBkd3lRnHlMcccQJPxqVsLgq3KjH0fsLY//ZESWux3xeR1RpHpoxS2nJ+7qPCsy
RJuLwSvn/rYQOTWJLOlrBhmawlDct01V711KFdDJvTXZc52sW2Xw1LpapChC9okN
InRGF9BZl4wH0BhmecJmKz+M6Jn3u4m/agRJE/L3w57V65n4AXgs/wydFcn6eWUt
HEH5zA7TymxwR4gkvKw7vjMeUcfbyA4/9x4DqS8Dk8K/YDWm5xa8ZtvCS4WPNl51
08sQkrCNkJ96hF5123iJNraHWaKoROqZ6QYOWH6RFrwQ/ji0xMuKVbuki0gaIJPr
xB7yKmU0dtnodXtHDu8RccMEeq31PNWHqNTteEuMgFuSzkMCGLfd441rQ7E8HRB0
mb22ToBnJf73IcqJOlvyvDERyBLes1E+01ROUp+E2KmlSET06th0JNQgQ2jiP2fQ
y6gf1Kgg/e6dtQTxjYexWIR1NkxIkMOKWJJ1VUpieXjnalR5+sZDjDpDLxMHDmwH
g2UvxV+/lfD0Nz05Bdf8SoO7yo0sju6kYb0gg8tzrBuEWuJsaKM7ChRr/2EiTxIH
/pPanNkWsjvi/OJM0LsN01rVePMMNAfR/3mxTne3xapVSXvYTrDV1hEIU72J9M/P
5ZCpCHFS0qr5PGmVLKrkMN+WJ3c1m1VY2wGkiZU+ooITn0EAigH+vvl/EcHYBsdh
yGno/xl8gVCe9cNzW0paZ6cALpVaD37zCrDr4rsLa7Jq+2jK7eQzJMETshG4ef9I
jeUsmDEOBZzDsQ3cDWLzHdoNrYXXGv+x0OsxxYycEUayQi9/ecpMmpObNKA0RIm0
Kmcyu1gTzOznaHlkrcfn4Bk7TL/1UGbDMbKTnedbUNqg8CrL7v6xB6tuzSH5ugdv
zpYa7I9CkR/dT402IGkbJEnEgEhNOb2dP2GjxUl/RXFLpGFfJeZISYmAG0P895cj
3TvDjTBpKZEnG9jmLh4lkxquf7CFDWRzIn3eNMOdftqewG6NcO4CCaURtaR+3WsX
2wLK0LweSF0Siim4CZM+6finSbElKJdVUcyLoZoHVasBVaP4e251wmH9yLYc98T9
cnAq5nZCQk/CAmwfwahLjC2vAQHD9CnwTE2huVeQt6+qYrJN5n6PE6DNaquMzoN2
cqO6HMbuIVYtlD5InALsYpx1RRTMDQM4kaXNS+9MCoqrWvOms7/8Y8hYzqBi8tng
SsWIXnA/dqQh6cF+9kbhguBNED6Gr1tetQQa2S70in3l8xv8YiM3Nu2tr8pOsyNa
4gufhfNhLe1JEuBUqiCNlkIbuTrdBCKX1JKTKBC9BKQs4RRc6nXC3vhj7P0T7XGi
XZ7iMsSRh3wLM8ksDYGeUgsJuIZ0HrQbLG6tMcLTQP28TlAk1uhIdT4HdJtqD1uL
CB1UHIKRbUdwn0juKboxCnXJZKhNX7ZV5654vNMAoJ0gdEY7YL+m44SkP8u7mZJE
Diykfl4+prYH35gfahzH4QKCktPTPVaZYTVGfZ6UpOHHmrMSj4otCClxRC0Kf/c1
jr1/vgr9tVXfhlssvi9n6PWVpHwLAYZ4/q9xpc/8b9NBArnxv+BXR/ztfm6UFpKd
u7h18LukGE0cazrGjLVAxCtTfBtOElARB6p/rI35e0ZnuPbPvrVM3ATEBToWZFUr
XCw3Ijc98UqwjX0rHoV82Rxi3EstQd5minmPsAAejCpxO2ETZO8goGJOioWU9lPi
rJFFts4EnVhCezkxRSI4kQ0zu2D69H3C2LaLu4YkVZDVqqYpp20278q+PMXaJT1N
h+YO+g/4BoaPiF3NmGPS4aBtctJXg/NXrVtMI2Q4qgAHlJBtKVnKngAS/3iDQkT4
zIXfz17Wc2PFCNElDgjE4Dx8pbvDICPXUFUI3DFQSkBeYkottsdHrbS79kZRQs7T
jzwA3VWQ+W+jk7nxvToumnziBVGsi6sd0iMHmZwzQxmFVcNmIv0pZuQU5nKlDXWy
Oc7BtLqj0DBu0+fxMNxYviDUCHOCTXPfQ6hQIfnLosRJsxkDFE40DWM0kWQf0zrf
T4m/ngFX280CqOxOrJJOKZLxF7SfWC2eOB3hc3+IYfO3SEKrakLiHxTaHu/vTz87
1/zIdgex9VEOFad2QnuKP+rE/mf5AY6Z3ETVSB0oexNo5ElUvDKuig3YGz2353Hg
KCjdBvpua9powoICrpJW/YAHjacoBcT61FCvxFeXsq0REs9mFtdIpXcydeLJDps4
X3xL9zTpEnjY7FvDidx1s4klx9R4B+Wt7x2K+kSzZBwYIuTKh9E6gqrzugc9F0qe
Gpq0jUv474gt9TmZ01ot43FapIOJeFu0oW1TSWNU5JtiH+an0q/PiEjY7sS33Mq3
t+Lyyoqw7pASkqFA4zCS6NohNiLzJTSALHi8hN0N0BGRsFeSgGEQtlVh/yI+f2ML
CreTD462ApzFnVflgX7QfFmEaAxdVD8fnhQFteFnYTyBOiufUhBzvM51STT1uB8p
E3hreGYO2vEYL1/DTuJrzVqIPlPWrvAtC7RuCcFJCQiFtGT+0liM/K7oUcd0rbMw
QjvpriqfeOhgrZzLv5zFHNnBe6qVxtcBZl7wdixITblez2W9ENTqJ7MuXmuqjmJb
zy8V0x2PWhYppdeb6Apg1C2/oYvN2RTaVK8k1IdGSiL/eNtxfvf1ZPBVfyIgtYKj
1rqfgBKAc2dWwN1MCRzumMEUX2+7ScsiHazluRWCXjgQUwUH9N+TIsNxSIzVx9fv
c+HD04+/jTFg1e8CG1daht4CWjWHRqNOd0321wiNvA/P4cvP2wlNhkW+24vYHQPQ
UeFFjAjotTC8cyYTsr8vplji8bbMWFSZhadHP9fzzZ0km1exZhYVWBEmiHHChrMU
FIpdBIJw+d6lgiAuC1+xyqHwaYhJfwxtaeEkg0q8BGed2zEpEFRmRc5aErJMvpkT
AkuVOhMN3Wgt59n+Oez5bWG5rVMabkhQBEmIj4s8jl63a2IdrEdGnK1xQDS4SJRT
GnCUZPb7I6ScIn8uDppCLdzWTCOXKuTkugemNQuQMlilJouxrgDDlacMb0VwmCRA
gDZ1u+dS4cCFxgvjlMuBTzu2mdLxpNngpFz7Mg4BI8VTm5rTAZ6lu8SJxiZDXXcm
dHtNqQq5WWt82ibSd72MTos6/W2VagWJ6lqnwqhucsvRc5HjBncJFppgg9+alcmd
/zApnN5ZNguObxyjZWfvDnmRNCiUTP0jzf5IeS/n+UQntSSDaeNtHs4uavR8138K
ubdd9LlElWjbWBNpLyKMgBfOKcgghDZJP4ib8xMy2g/twr002yrMG25UGX0vuPq9
ZcmPgHZ+xlak2o2S/ozxllPAoBF0C/g3ZUARBMw/EndCJC8X2Sg5Ix3AH+LX5+Ie
SYC008gs6pGfQb2DYjJUh6V6SbtLdMT5CM4golx5a1LySxNj+loTXEpEpPyVEWgK
KDorv+gnuPtRozdXCI0X015wFuLzYW8/Zoy1VNJ2gzEJ/vvlVscDF/WqNkEkWz3K
Y+5dFAalxOhrh/s5iiKLxQyi5pafcEYi5Sr5ihOzu4CkspL4J3s+nzJqVEOGFfiE
cBARAtNVd+QRfXYoAx3G7MCdKIaEebT2nN+lSz+LKl7vDfxGdTdEse4voxbMcaAH
b1+JGlTdBClkLK+kxeer5khCOp9aPrWAlPzhHwHIgDZ4RKIaUhT6r+1h8jfepfBF
mnKHUuA/niaLavo9wwnelMJ1J8wdBgDVfOtqdgezwCg4kojH6wiUv8W+vEyqbtEF
Gc/wWDChhJvym4ecUP1EVaQTpRdNZV0NMT9I1gk+hbt0m/wAXNdoX2ZJqZ1wcNWK
KAoEkcdFINS6mHL5wNDv25ZxvGCvNek/oDhDdmzA/8K9O/VFcfOoAhkk8TNMNTs/
VS03LcMNT4KixAEcUUteJTA17GZ6FBy+S6tmRLb4bXsrakDunUtt2cjafmR1zKT2
1dO4kHBZp1icpl90+bGoQYTMEUPzeXQDBIeBNCfBPma+jIXWhLq/hGTgYR6Y9XQU
xuQ62PLDs8eqqM4qtRB1ly5nL61CmEBEYKTAUUvzoIOI/JElgkEPOeYROe+rEW1p
uLcdKe+atDU31bv0ST4Uj0UOBbNB41UZtCSziuKE+kkTCXKi42egxbbr2wGPOQ2r
bS9npXfalRiImuM6bcSEamqaG6yFjGtl6W188/B+QAh14EXNl28pnTm3CG9pT2Jp
ALw8+kmgfqw6aiZ2MFSRtPAVKOqNZmR//9Z+JAvPVHG2O/SQNG3CE9bvYxF7uzcd
pihOXmaBLIrV3tKrc462RcHm9gL7cYcs6L08bm9PxGF8BgRVKk6MohyOI3AFSM4A
exHbJxTCiDmCc4HK7VyepM5x4N+EgdwjWZal7+mzvA/3cJfCHCogwkH8Ilc8kjiD
RjD15++1SqdzE7rMU4nk5Y5Ec4Jwr9ZR+CkoLOtCm/0wq/e7uECivXBbbVoYY61J
Fv+wmfC8p+D0HGa12DCgk5lcLcprpUccfBlK+STjVzyj9B0xoIngho/0RoHq7Iab
Cx1rWk2wtPAY/juKZ3hSJGI4eIW9t1as7WHjaiXIHvtSprZgjumCIEW/NRtK5DfJ
ZHUHUiHtvSvzo0H2uqpWT9J31jprCRvfUVXtVUuPvS+dQKRRZtm2ilBHIy2lvFw0
hfjWfJc4m3o8xmd7hnq2SAB9jEzI/Pt4PEWNMf6HsW8WBFJxi2MDHsS2/RHdu6XU
33xkDvD7S3iNu7XhxVJ644edWIWEXsY8GSmiXHnzviJhPTb84zNVOtUXhBJge2k4
NCEm65OO8r6+SNLud8r6R9PLJ1r/L+k6/WGR6aVTb9MVe4T95rhZM0HLbDKInQ7a
8UVBQwgwnW+Mg4Set2pV1ygktAWJGtHvukC72QNLEPYUYC1yuk+ZwE0iBe0pulW+
9MK6R3O77tWeoVy4v8fxMcI99tc52IZkEKA+UUO9MAu7WHTYTaeMzMgEZqwynWLU
bJq9W1r+JX8Ae7LT7rbceFYWANBfFSEr+L3EWPDvDXxG2RN/lHhKjzK9igwodSWX
tFdZ0QVYGFwaecqpkIZfszTb7N/dm1KHsYW4HSkHm8mHQtP1sTyJPRTng5f6NnDm
y+v32iXR9MGhZDs3l/DGcbkve9Spwv2kZnzssxSg9JBnoNZzqrllnDV76sHPMhj5
D9BgVRngOmwO7hRDWamlzVy2ZNbGt4W6lS/0l31OAynxB/dWfK/xp2GcISxYHuuQ
87idrtrJJS4MNNfXp3YfE9ViG1Kroy1utBk7XgPuNtWXU3ezct9BcVbU5HFLOoFM
FBrdqO0FG0om/2gBqQC8F8UbC0rK40RAFzaAcpO433JQiwQeb2uJ04ACKgKa8EYh
39CpcB6p79Se3pTUcQX6NvzoJAnt+opv930voKitllwnI5EaGzuW+hp9BoTd62qD
cQX++QoTuuuaNS4EM2RaeV97xauChrqjRSuDu6agRSSzPvkQwjr5gbaOeB1DFxU1
LzFkmPljkEctT8m9m01Da9qXqSHoE9Lu/ZfYtdjD72baVkXfuZkX+MmGAHG01rTT
9jUv0OzX/lAta5ie1VaYdHWUyS/tFNsIL8jLq0F6UgkkcKJfLp0JZhJBStN+i+zZ
CiohUasR5oWti+khy0cHO5qQUV37wlh2DCGsjG5gGpKUAJ86SOlBbJfPNQ0oUR6c
iCkKcGm3fNkFSFDkyszF3uuTZeiZwLt6eqEtP5USMDMw/rOd8GjOBT1QhigYEhHM
kYo9IMwf/LmYF7dJF3E8yhhdYwwAhD+DKv4QwNmMmCPkJjCYeRt6jbxUy8W/qHnf
uY0sgt4ilW8aMoFYAO75eVDeENjz8aTdo9IFCCarp44cGK5R8OdK9HZhOb5iB/uq
RqabocT0q5EvX80WElWgKv2YyUPRZSSWr2XHchr3/SzfSiIw/pQqmuO3MCPy9XU8
ztwHjd9CfVH1RFdcVk9xPU+nhTeA9UwXFp8trmZozEm35ZrehBhSYNAnMlt5NjWY
YXVD9WAefQkTf5dym28wcsLGn9xVKaq4hztL/jUezjerm44F7M58dJ4SV0IklGwm
eTAeS0DTYCeQGDlGR7SYbcv1fixxV32X3GRk3HKCQ+OPi7Hz9ZTzhZ8iViIPSlBG
uttWxqS6ZTVR5GNo4mWl2rQNpCC1+uVAF1aRYkHl0vUqouEpJwEwNTht0CgI0Zw1
hebNhXgIiuoGId1XZCI8oASTykMrad0Kz2lfew917gc3+V7A9jhWq1H1EXBTFvxY
YjBacmFd6KEmkF4jhlEi+DOYAdeInvxa6P0wZuemaBv02x+ErnrxWx9/newsiFdE
53IUARxuAGg04dgJnTdT/lqBrHd2kQwQ81OdbRpyD+Lze9EH+qYbXl0XI4JX0+RV
37NkqH8a7LbkDLBHbc9PTBFf0EKURD/uQ6nk1f02TVdQ7/hiYhgFGJ7pDAiPcaL7
K6l8jnvwmQ5jQGD6Fh8MYMqABllJCATetQ5CIfsHMPgBITFzPA5suRTTzs4U3/gl
k9KnRhg2C5bFAkMzwenVMEE09rC/J3MK5uouxOrLloaavrUw+P5TnBXvBSIRkUtF
gRoNuaEnnmt8Q678lo0qibiznBeLO0OVfnkwVpWv7G47L7mrguRKxVdrRmM+U6CT
XEH+7FuCs1T8SU5OEDuvYHg9vHg6sbHN64hvvJa5aEO0Q0t2qMF2hSERQWRBTARP
I68QQzhy6OABMoRggA1/s+u/+RBAGvVctD6UBWvKp2AKNYhD2PRcRCv4E+f9lMO4
g5odVozpuR0+w+KqrCNxShBBloT68OfzW0uLwEGnnaH7iXTB++FZUxr9m2M/sLU7
5iyVuEz0oSvUbPwc92akQnsEjLYR8Ycj+gPeotZ2Pi6ena1cw6aG2I9z77Ca2VI/
zuxXZ19RqlcGJWlJkjEg7XpdHOQqpMY72JatoA45WlmiHO/0K1mzDPqCvSFs8d+r
wnQm7SepYb7Kie5WAm4JI74De8UraEsnUQVAicD+efL9UU8FJnjQTGTDysGVZLBq
1jWs+3EtPEU6fOIWiZ7joIOSUSYUZqfNU3XReR0JmYXwwlG2ag2x2lfgQLOng/OC
yiaThQ3fm8BsuZeKas8iPyyjwfJ7ZuWonQG/Dl5glIZfuGtOE3JOnIlCZxZCMZNE
Z8zUhtoMIe18mC/XSCyqXn8h2q6XKfh8QkQ9L01A+9bs+QpEE/yLpiSzPUUwQCHl
Du/DAtGFhwWDJVw24FbXxYwV9FcFmryWdtYQUun14Yq9h+XDSo9LfQ6vLjQQ1orm
a0y6hgB+WHQl16nSynfGrCjqX7zWuIJLCv+4kYeL+y9qou88t/nIlJo1imWz4P3S
wx/Uf8xekgh9fy52GLKlgNqloi0Cjh9F6iG4jKuuFMqxLtSh/aHJB1uLjv7+DE55
ly5rM0ja6jvmF3DYapf+v8AEN4zVBYIS+H8k0/sJWNmROvhk5GXmAwDgwTYOqI4a
Nbt/xq61QYYc5I3egIOtF3BpqU4xwWpyBVQyU2J2Yb3FFscovDygDXXq8OJkxYBe
JRCEMVxZRw//H/hbqoR2B8oQf+sHFd3ZDZocXFK/vY77lOkLo5wNd+PASTqXSKXx
bBPFb1aE0Opfco2USLMqgHzNSfSakh0Pz2GCXuOVA8NtyBixDHVneBWwON9uDBs9
s4nTwxgMJrPR23SR1MYgC+V9nbAt+ACi1QnxPNM54g+d48xbvA6fEwnWoD0xO/+J
9NglalLtMkXxfECTi5/Vs1OtHvuOZ4YxmSBmkOiUX1UFYz35Kt9BbuAy0xPko6c2
eg2hzYV80qsYlcMXLZiv5W7t9JQ4chziROtGz6dNNhClzuxilrMFM6RzUc0FY+g1
E4DYAK9BvDg+Uky5eRj1VDjbfUkOkpqyfKlnRgRQIOnsxmEEKGHOVfG7TipDaKJF
wXrhEk4LA4jNPPrFkeoHRcIOuepltupCKhk6+fR/vUAzGccKm8PRytskgBOhKIRG
1rFnZ+QgNEuo9Rj0oUfkD3swLG39FiDwUenq6DkQpEMDSdbldGgc9Hgy+sATyyCS
erFMw+pfCWeozq3eAB9lk4gVUDDI38reB6WTJhROGmdJKhqDcdA6PAFqqySBTeNs
qIZKqthOuXx30XG3kENEXuEig1vzVISFB28YhWV+kQwVyZrUv1Jv5bLhG3IqGOBw
f/WwiVvaNXL9fJ+Vzxvo2jrKvm4TjDY8AHvoLF3y63g7NGV0Rg6oAmZ6C4tWeOdG
6SHWRcfp372Kg8jq1xdm118+LK9o07Z5jL6+AMOOax3/+JNCtuegP9k5XU7OuFRN
PSBzONyMR2LFlawMzwhGfTBZ7V2OuBHzX5vkXmve0jW/6mfv7KcF+gDuGXzD112Z
+wGxCpSbi0Kumi8N5MFCoYkCOdxco41XEtIzuxGPIbWsdKhWiPyltJ0udXvrbJGL
/oXXQ7Othj0NsvNGRtArZ22zZdXvw5MRU48PTUGH+M5KS2ob6siHH/PUyQRgPEF2
zxaj1xl8IyB2fI05yirIxy4JXh3fgDBqAI24m9xkxvzT5NffcQabukTjDSff60EQ
1NVZjJSd+ZZmfbgMKfIMsx/LzIirE2GZFRgIVaAVl4dpzLpr70mjpDoEwqDdbbHQ
hVSia+n4jnpCy0cViN3zABfK3yabZIwQvWD7atmEEzmzN7CTJVHk9u6Gi/zRSSqJ
pLddnKB9j+eF8f1AGaboYc+6Q62Ej+UOdaHJsE8RhRkLMiIEoL6E2i02iln4uP1w
WrjVDNCGaGHCtoAOI/+k7bm0VVnWHib9C3swjjD1J3UAO1ajT9lqv/minO22ByBz
lNfWCF3r7MMoOYuMZPgdzJav86+SaJuWcmyaNyZ+UXDg3snBEQ4wX2MUTsN9WY7Q
CcxndeJmMMjIirDv8zclEX6tv76/M+B3LgeMs0xC7hNEZIKV6KefPPirTUR7AMv0
eB3e1hQjSC74r/whletHLSI0Z5DYtaihOmNDN72tLnqjAK9/CN1DnR9lnvCAeQ0N
k1GnZoD0CS50dgGfiQc+FS982NruMSzWfOvGuihPCyTQNcjyo7WsCuFZC3iZ1TPP
AAWhL9lc8yYxPnxbVILfW6BXHU8ptuNn3IGo9YNjmKtCQV2AP1sYaVxjvebdkkHl
dFB11CVNT7P2QctKnvmVGQ3rnkWhuIFC1PbkZp0JQV1CdpTLa4Vh5uQah4bsApRk
yV5u7J4GtbtwZzjtrAV9IINCChIGYSzZIxlM8qkEn6hUlwKcQGjuxJf6IVBC/3G3
Ik/YVboBRBMukjV2jw9+ktG8smj+eprFsLr/sqff4DBt/Zw449BB7LB3pXi863uO
NtLC7nFlR0Hy98Eom5kT9j+gV0WAs9nQrzbfK1vU27/Fg9wnn2o1g6YWKLIDqJ3E
4hZZ4x5TN52P+fVcoFF0RrPpjyo5fxWUm3dhN9nd9FQ+UD5HrEt6Q7G2nX4xV9SX
XT4BxCld4EgPa+mLlDCN2I5U66QvkUAShj3WLBQLUEkc6rJjTHpVXQ2SXjLV/rKf
dwDIf7uho4Wh7nCAp4JhxGAmY8LHvm56jSmF3BuqSKNV38Xp8Zut2cRTxgxDMU+K
H1A5fJx1KoQwufXYxI+IS8qa1Y6TECiHwtniusRRngzsFuAd/9tdq6HVml/wvu+q
ddYra8+hlC6ovZazOP2AQF6YSkQcGHtSMSv2wJy5ohusvIijaZVOCM/9q/K34Sdf
b5cWGVEJe9ydqRlltG176rHkGJ1HXCzKedLhpuQNa3wglm17QLlEnaK0/a33frd/
iPdSDAXMb3WYSx65Pgl7w+3iZsxmKG8h5rTHDEnzrBiqaxzZjqqJret6ela9XApo
57Oeu4EZ3TeB9guFdwlnwZbn5qsj+saQhKgoIybG148rA9VmsjqgbYY5oR3MUSFP
N2zSKNAA2NSihvLQq9h7eakIskvNYV+dov8TwPgOtIPgWluQCJ0ZY0v+xU2ffIyb
WXH8LpaJQ6qIOqEqn5n0gslNLhcNnvpCWahQpcdlSdyeaQdd09gW21CvOSMGQEdc
vKyaTeD+2ZA2nPLQ/CdODRL9/XAO4g1xiMzq/XvNeUxbwSB1xoUC2HrIn6v5Y4Np
46bA7P2VsVz1p2+3WiRvYbG5d2EtG1TMpTkjX5dRUxXtvex36voUEhSDMUu7FTk+
GuZRY82p8Jk7U8h+5eFAjqBkIMObNn8sgcuuaM1SatbJwnIZJrAsAnmgRw2CzLjR
5VuduX0YoJxS88Wz82XYcQGlA+hgtB7XdAqYRWDqo0Hy2fXzYkRqV5hdP7JwDkHb
+O5i3FfOvWgHdV9cztgkIvMAnqo1IjaKE+VvWLilXOTL1mhTo8hDdu7YYJIO9q9M
lYas/f/FBCf/B98td9SZmftGDtKVkCh+6B0cbbynVffFbZ1U6Sxle4GeHCqHwMAf
uBc2QJd+ks63CwSmqihr1Sw/9yqjBKsONgsLZIOY5qoREYHr8OLXwcwpqFo3exEJ
9ar9U6Y4cxzDe6+tU8td7YKGW4AwRZk7mAMYqRgp8A0suBWZOVbX268KwHVtoAOn
rrTghGVzeOp/ggjvvqb3gqrV/OgzagiXsMoZAtfqfebpXuPkQGma9/nKGCy5TxcA
vFZJ+IjgTAXSaqszXKx9y4CwtXx+b6J8F5qLa8JPFZACkORc/07N7QNX2EWSi8ZH
EqTXVVlzzuTS0fYfwtiVPO8RoqrvA7deEhf1zP22X9EXBrk0FV5OG2IMFSXG2n8d
NZorTn3rWBMPRsyYWFoNqNjNp6L2GU2srGBkKhmk6alF7WgsFqR/LWjCEN6YxmPM
b8LGHVYdKhTfDatI1iuWSkrz08MWUkUwguYL9hurtQcD3Ztv5iQ1WmVV8zfyJ6I1
81Kcuo4kylmM+yQYJcliz7Xl6ExNTlPd194qO3J6ziZtPgCDefeHeMBIAt8Cu9+o
7XOYBb6pOERkwK+PNVkLD8Sn+0zkrPVsaHmP+RUFWVBDEHAEtjj1IKsTt+RHvw1P
gcDBMveLkyE26xGAF73usOrJfL7qLLpc9TpUxH/UsZpOF3K1QAFidCseYPtgDniV
QwklylFi/LQm24K2gTGmP6CDXb9MASy5PVpLYYyf8OHb7qq/AqSIVO2BPlPNL0Zf
fLOo0xvjX1LwVRrMbY31B4Hxp/L+1tA3him4sD4iur8pBFdOW55og/ZLfUKgRv+J
QAk9W+9jIa6kdLhik3K1XxKCkbBWw3Oe/cxdeApO8HtNLUhgWd9IcW5DINVd4phf
wUV9M2+ZjTUYY02JRwZ2Ux1xRVSsWxYhOEnqL9l5EMLmDWnnZlTCvsEb1UXEPWJi
b5urgbnOO8N5b5OlYgyKvIJ1hAPjabQJ71j3LP96yLmMwKl9kSl96sPz3mouNnzn
ERKbPOUpy+pyYLnPAqXi9HGDOmWNsEuFuht2A6p5cxT3JBsux+Kjfp+g9M8Ag6bR
Bwq8jAbiLwksgY12oz6loheMb+Ges/llIEfu+68fjo2ySFch8QE+oWfep8pr0O2c
sJVyH7a03SyD9wU8p2WQXbewFRSovfLCtcFxqDvqD41ThkrKvI9Ye6SPR5p1jekJ
bw/yNOH6/KCC1OJpcJ4KfbsOsmJcP86MMSN/xTmhWcYgKDgyk0HuIixhh8rPNsK3
4BWnp001Ui5i9wv9ZzNl8mA2yxweV9LvoznQPu2k9cmrTnvwYQHpIFlodbYD9lkl
0tutWUfis7Y8SywMru7dJUK07HD8r72usEOdybqKyTUEGFheO5w97EsfafQISfAw
rEi7J01SlsjeieZXD3p1VFuklEz2jam+FdAAjLO/LEL8D6gyMVpUbQaNv0VUM1tC
wQBL0k0ypVj6EbXE61nzvVEY4G/JBxnyHAi+f1uJRs2WFOzYDqgeObijt8NR+AKj
yKMcv9bdsjntPBxMo0o4vzdtM6603PHrSlceUpf8jjzRopG0pYhLdAgT4Sipb4Ji
GkmR74k0+JMQEshGxe+9d9pqE/dui9+o1BopQjX19hKvhBRfWu/s3CDO1NDvwe5j
7S5rmx0LW+jG+JQyNeaqIVnhP9y8XxN6vwHOFBev65Bw4ItYtBFnfgo0KWHaByiG
Mu2GPqQ5DKNZ+OrKt54LFeF78NYRNK/N0gyyF0IKchlyH4mbmJMXm4UxVCaw+pyh
ZwiV2jzVHpZ3PSD3UAv8/xy+w9Zzp2t1Ad076AHxNUoyd/nfuzNVqUmp6W6kvRDC
S1e0/JhQ31UzPtOhCdOvWXvqyXe5KZR82YjY+DFyiQ2/s3jaA+6vmcZpMBOzAgGK
KmKVsxI1EsVWEktyBQI3oUiRL5tYrvH4ci/3x5tfENmYjOPEXd1cuC7cizYprMeB
G6aPeZOvnl5CqCjBR3NZQvrd0VA7jGjwApdCLkhI1rpoleQPtCgkojkCaIK+TKAw
iJf4hpbIHBEgjOdWwPWIv9DCrbXrXGgVAckHviKIQygiva72Whm13Zu9tSAgRJt7
QVwbExszk9pTcbUXghuXpNvfAvXCSIuXrNUyf7+KZcadW73ZMq88Md6UPV2E4TXJ
iAzzHzMtIzSQEToMA05wrmVgrB94vTbh4wuGena34FKFI9/445Ly7pYb2GIyoqbg
Qac+h/i3RIoUwc1Mi6ZpIYUlnhNEoj7NYSdFkUJVrdXGK9hn7x4h7ELwHLVLIV50
SwJHHEI9owNihoIKwlQkzaXFiP1TBsb3q2mEv51PYgfzeXIzL2zMh18CPgp1MdyP
lRYo5RUuuuBJyOExYeh5PGGmpDolO88QN+zv4Ekr9wfoiJ/f3ivu2NOrNP1N/Kz9
SFm0sGw7Izu2rYQmYa814huqBaBJS5nuCaQdf40QfLrXSIlvo7yPmKGNq6+4YDpH
3b4eypTYZ7cRvdbkEqDwc0c4AoBpuTqR+x54uvE8iQfY3Fejh7JkysV78hzK8Kes
VHjQJTvW9VOKk/zulSJMQ9HlLapAWUhR0Gz87heNoXTRXTRl7kPgUSYMr2fc+adK
wLfGaddMGDRoZS0qxISsgQzllbt+fKOA2HqP2n9d++TIGOoUx4KPp8d/8OxzXLBx
ynkcjONHbjqcrpE9CcUFLgxG4XQkvJYzi5pWqlEJ7C5avUewX+j80/HFs9jELI5q
ZNf0dSoaJXeXL2nLYHLWOAZp38WsZbK0Gdy/DrfaIp0tWghzQ/eGpLS4PPrGV3k5
aR1hpH9IB3xPimeK0wl/8ZvNEPUBoi1JySV1vZXKRy8KfZW8XOUktKC4iDsHKQMa
7jxv39JM9l4AobtFNs1MqKyQiElQ7GyELCIXBIC2xrDj6YIFG0HmsOM89GpY6Uaa
yDAlfav+PMsEd2oArklCBg90g41hJTBVLISvSkgClddV7A97UuH386pbJSFJVJh2
hniMusA1s6RFNj0OWBUo5lYmtyQnr1BktlKCtbQQSQjpe5J9jwC+gS9c/IL8YlXY
NM1tdlHubJACziksjoxtOgvwwICFyN76yKMfaPzP6Om0/ZsvxqR4aYlxqYWylOQg
O7LShVIAaA4KocYOgQCuhJY5VoWPpixs7mgi+NBXJVmPgYvzrhqIMyknSPebLGFo
4mzOGqFwbwwGaQMRG3WIJYM5dlr6Ceo7BcW533nq0CADzeLqNZCpyCsv3C3uGWf4
YsKHhfYs6ZOhkRoGWeasyK8ZoSZfTauolvzaBT7u8sKXPCQWr+rid9mgivxTuoMN
7KBGEs8HmmP9WrCQ2bz4QjjDyWSobiyQbB8+aDfKt+qO8w8RlUl7qxrODYbqIcXK
op60PMpTQsX6yt65mlvajdyqs6eEGvmTmvq2VqLRjjiZYDI3cCIRrDTZ1D7KS1Ny
8sG5/zfBLWi/70noL8cq/JHA7U+ks32ssdmQSobHqzcEVzEQDSekrPvwOdgDgx9L
G45KCQL9sj/1cLRwRA6eNp3FeT3980gZXY/Fi9jIpXUPGGRxslOixApvqimBHxBm
sOBlbDLEUPS6Jkri65eY4aj5Lx6H5lAOHsx5gKNoJfOzI3I0X/2u3Zf4OZXuMjpN
fyU162viECsPMToe5XEwpRoG2wcUaNQWVUZsGAGw2mkqFGMtxuCuL1lson1cGZ+o
yijlha2071VOc3Q8tahWc2rn0aDkex3WZXytYpGjFH8ZurSnVctsgYidxnRjCsvx
POnOyygTndJwBDCHrd4X+La6S2zPXFjywqdWO+77OmKEBg+fiVflTZJttITOsRKp
1YJn9YXm3aFH4QFhEk0peeRXW+k9iCmv90BQVaWyY5q1CTbkWVabEHOL+ZDpjoJ7
4Q1m7i8s0aFvnBNjsS7HDdIvk1uXYqgEbHn3AI1W25BZ+sqRBsF1nvDI+uHisly4
d8nsJYqqBmGNBAPUE5aDDoVH6w1nlZWmZ4LedTInae5acrJfjJnSXvbdztYBbYkI
FRIBv1/8cILON+gxVPKm/qDEo9ly1ec0QqNQl2lhOWhBmHnOJ6QxWY13zo+EaXLG
A6e5RgOI3RPtA/e/ruMNSKtxteU9t9vHtIeCOCRSqeD4pf/o5hSIrYq70iP6tuMG
sh6TBu+wGlQfHqNzA+3HgdxtbpPl3Ue4SwW6UXg3P7GXuz2EDqZCjI+ceDevLqoA
fkNj5mWoSUy3r3H4SMtCu7hbcfWZonlRI0LTavIldg1w1ufaOIe/8fKMQbN6+wXK
8v2HMYsc8iDHdpUHpwhBcD4JuLbcd/GlrytU6uWwmW8W36JGhyRCdtKCDcZ7/2wt
IWgoFK7bvD7ZDTX7AmhybrosFAqpHZmEM7YC40ataCwqtpvuwQOjUUB9i8L5qUgo
ZIANVhPtTcwbU7Y2//ua8X6+JTXsj83h4t407ZL/z7rhRHWi/h8IkZLFH2GvDxyE
3WCt9Fp3GP5WZq2aCrpkjUVRU4uTsdYk7Oxx/D58/Bayp1lhB+RJMuYydLw88VVP
2CEweTkgteapO+wb6wHadWtv3vUBXwSNVMWcKCCMjKX7I0qtn32b8BoPpfwxKFPY
7qJffOxPuUjzmDiEtoS4MjsNiGWIWJFiaOIY+bE5OzJ44hqwjNubRGe/TH0ppU6t
xfr45XlNvVA2D+NTSgIy9ql7wutaXXM/+5ytcEukXbrRRGuozJ/FtImdPfzAlaun
Aezlz/jH10X5H2qcw/DxXW1shbbiBZjz5s4q7RnzOXZsYhCVmPUp94x3xxmZsPwL
aPLsIuktYkAzOKCKJVYnM8WENJdkm1DlriMefQ0c44xlr/k8XjJRmX+IdmanYWn/
QoHB41WwFE/s3yw2Ki6Tn0wyizSw2PRBcAFc2Fo4HSUbqXJkquB7z1XsNYTWmQzP
OeKB1B0hjJeTobAnnEzH8hGT8frYgYJU2Mz9u8JZnrHfebp63xkLW8UER2r2pcZT
XoUKAngsOmezEEu9Onbcd7XKQwdS+SqMR6hLX6zMLlMvDsTUQbwSsFpUtjffvYGn
fZepZVanJEKgkLQiqkIvzxLt874VFSlNb8o25nM9Cg9HE3/IGmUSy3jYxoWp6G2O
0pBSYpqrJW0yJz93JdkHaIMXJKSwieZmEHowaL4q5t4WgNEGXq8Md2ENZLL8z90W
GcHaO9X9tFRDcynB8FZ9ts4lZrmEX1DwT55a8RjZqeQaaqRFPqh57hctnu9WayDS
/By/OnVrQyIRa3gBUyfk9kw769wzGegKc6LgtFNqJHHTJE/M9SkqRQRgyuWn/mWq
l/Sw4Wl3V1vh6yoZj8+BvF1MWpTrHDilWSPU1Xsr6Yq54Wudhy2zC24lnFdNMAfd
M1X3nibeveUVKKnX5anDA6L5yQwWECEvzV2UbnJmlRm36FgE9p9XfRRUinWdDMIf
Pw7TQO2gpZ8PQQlUq3o9NRXuotav0Q/7s/XBReHg/iJ1lmF3l22F0K5cfhEBJ+zy
NaOK8A5vPFNJoU2+EFHKJvJO4stOQr7jU5eF18oDg05cQuM9YtqSIDQt4iWoDRcx
xNUoS6FM+TKWoDBFc/kRSXvLudGRjxyq93lCWgMrdvnSdqHZbOWlln2OHnHvbeC0
rn/muSynJZKMG566x1nzn//H1DDWinGdF7Y/Bgx135dw8oqvvrpAze+2RgXocXcM
NevCCIzXzhGxnI24o+xFe/N45G+dUNjRnVFrCYYt7p0ujz3QGkkhIeA9iWp5W+i3
QdaGO0qO4pHKWqkP5oS0Veiglholglon+jQlMoJegrrIIktVzDj2y2di/ch+cfhS
GJEjfD4u3XGU7DnVbV4byPxR2Rnid7n2JaPhSv8nlPpnnqmCPHXRS4gQsxJmGziE
gZpE6O1prQVBHSHLN8WUqsNlUia2S9iSGoRfwCPkK1kUh71H801BccjSej98OY6C
EeZdEZ+RoUxmQmJXPQnBe9/viTAeBJ63UCY+bbUlRocYT2S5jum1z08Tkha/4jIJ
lqBsCYk6jcmvlq/kj/waBv43AMxfgWUcPAIpTtBom5GzqWpg4kDVkiyfP//u0Tmz
xXzb81VVkVDwzJBmtn3UdKhB4ewzO7HmEro9btGDc/ytgOOXYtQLZQnxkWQZLqRs
kIbD90Y2OoTlRt7qnu4rTA2TuriB7W8OXVMSyxQ10wZ0s2LO/zvWI2HAPCccwDer
nu6ivgHXUDFIP19N0a1ne1CXBoa2LeIUv1qw9UtvWPD06aFookccMFnq6gjhsbDe
4roOmUEpwVmu3H5wGcqWNI76Khjca0UZfFguOBZfWctgQ3G6ZRlPwDcF7B8i5BaT
PsdYM6Tu5wnuqBRscciP5o6+TDYAFFLgLSIXs7GVpU+WVih6fu8Kzxi5viF9n97z
qiPckC4IOMi7HjUgFGuvdUTgYtK/GadDuKZ53UZnfBt0LmAfhAXsRI0SgAJVUhSN
ibFqiQaeeUVI2xL/E2jwRDjg2+Q9ND1p3a2gwjQJnbsOWMDlxtbNmSWAxJbxqSUC
uQetdiIRwqg6ywIRmOvqTE/WvZYVMamxPxtc+FStckbhBdg3yHhgnDkgEDZ+4eUJ
tStR28sHLDiEx4HfZtlFqBYm0sTV5kaZtNqbLKYHUjCa1llDtiYI7GMR/bM7d/S4
+o0IG4KdMLMp8/SlxzfoZKv46fxiz8A+5DOJGWsVIImCpnrRVc8KsYwD92OgoSHG
IRD75p3PiDQMHk9iHM/BeUdJZFWA9pJcwDW1lqj9pU2HfB6RRydYkYrzlk55Wt7Y
mMNqe+qSg/gj2pQCrqJFgeBEL5iP1YJi/0S20Umr0HpUxJuQqSG9W2eEKFi5AlAu
ppRoHgxcwtfVCIsQ+ZnrXXfQGp0Zqf2GZiw2MN3iDWX0M8JNAKzptD4fNgEwvbDK
5oN2yU9nM9NkqKK42PVpf1B/ik//673VZl8Duo2PFeucXE24w7jsi2pE+NwecpV9
sDkcAdZloll4RKwmhcIbDJ7KZ4PL+ZrSAuLHTn+TcpP/D32FBpP3ldzun4QexMPK
I1aZZaSknUyJTM4XBUetkBYP96argFWP9Lps/Oc2MWZZ5WQKgF5Au7OPPwXV/l7N
64/ogf2vNxsHgzrvYre6ruUvql0ajUh/CHxANcUApKdd00CM12PnH2Qr52Wepyge
iZ8t9Z4S0+ZZhUiIOvXFAL9xHBmebnMVpzzNarwPKats11cY6yYmyXJO9JxL2GPJ
BTtC6AJPdSlTZB+VUYcnFXQxdIlC8ao8mKD9URiO4wiLwfrZ3/PVzzdVqprsIvvi
IFPb/2G6WFHw/VkDogaEMb0Rb+zc8YCWXm7IrHfelrNd6flHHO4A9XmL1mugABHG
WOnhUTdER/gAbV7yBNly0AnVvstLpv1bKduIwsdZSd+St2lAn1sApAko2d5QDBVV
vOs2DvqOoI/DT+YvYR10pGPEEVn/F2t5qsNu/OOpcUVFoNLY9Mus5F0MWlqZ2qfg
s8D3Rgx8mINTxEyhfLPydNukGC4fHlwRq/RMneSSgq6HgIsGcKiF/Ax0MsS8PtRB
zgt/CMDeH0ubdD90+uAfj3vA3Ah3CRc/ttG4QEj7FBIsD/IjphlzDLzZ26kVraYM
FSvPOzYhRR+BJ9HnpZNfmjkHZ2PV7SjgX73DVIt347wRoP9g++P/fp2Oo298KNoj
23pwwhzOju+CNGDpomg114u3BJda2XSdOYD33WLttyaaqj0JfgdOrQ23wWZ3XPUh
rx3bzRFs7l0JImokuHcgBMFbpbJoExgWWleO+d6PMPohdo7eWojcPyb90EJkeDLA
9RKG+4y/+t87KJ9wmWsHe9MDHgJ9yzi5X//unUAltgknj6UkSfB4FNGFpzwONXi6
E20gDGfbf09ay1NJjff+dRJ/WRVF7V84ihMWbxmG0zQf2SmtxfjB4Jb10pM0uU03
lTLoJOX5l/XR85LnoRXPVsVohOCWOjgbmvkup9t6B1xQRgYsA3qLdcM52O76WKuT
YZmQ5uEYjHkghUu2AyOoiiuujm3Y3UyD6JlIptOkUvrVWDfTsSPL1L9PRnvQNfcP
IV8hyV1qJvTTtV5TFkeGn3IvHZFaE1H6FH+i0T0B1DtPuR737hylmoc/zRoawOB8
CfAq6X8fRYqVHZteRYJNxaBp8tAxCgCPjmSnGzDdcHmqnoWEzLonx9XV1Pe5YsIA
SELoFeCZWhNuCWXr5bBb6VjqbGoyRp0ekxoWbLH6OfScNwJiIJyVVHsNhEmBDdtt
1+bKTvZXIigWTN5erJTywSKQoT0GmmaHsJPfI05FYMBZbHxww71q6GWNM+8xBwBQ
BiPKbWo79ET1wslSh1t4s1PGeS1m3pvVhVfsb23IC6Qn4036chBUOUl2dDKU7WbW
FCzJaJbc8lOgISht07iPt06I7OEVF/QnJ26OvS8D3pHVAgpMBEX5mWLZcLRLGcNJ
CyPpm/6D+gOcfWcn8pP/1KrkKeN65eMhzk5JDEI99XZ4APn9hdY5Fldbc44EnAUC
4l6owIGRg1tb4V9aINV4a8PR2z4eWuh9cFVGrWB8D7M3lxAn8y0T0vdaazVhBekX
LN2QVme8GDisfXjLeyPlLxa6kvu/9Koe/n7J8FPhSn651+39M3hYMZt8L8g8EQ+f
Xc0KmiNNfqM48kTG7SrC2UmsJCZ+Hw47OdcwL7KjEU6ovTAPhLu5+fSEdPKeyGcJ
9UHEtD4Fl5NVvBCEJY/3OwQ9lifmTuKsCtXdzYQi+0VZV+ibmqXZn7MQVieLQRfd
Hrvby4+qw2QYRghqLX8383o3X5p++JO8HHv0val4XG8gp0c7axaEZPbrAz3PHRBE
2I3MN4/24STkRGWIuFLR0alTlJUWKG4+JD9I0C4f4UxL89/x5TDqtYYsce/DNlHh
ee9BlCBLU2Uxbwkw/JJAF6SytBX0QB5mpCq2g0ktqnAKBHL3LOdZwoDqrL6F1DTX
bbeiKRNqhTY+fyp87okFt8lZVzxNENeYjO17n3+aMTMkJrB5pAl6vD7Afw2vf8tx
wXRM58wSunDiiqsuOwdUfXWIbvw6N9hmss/lvEuTWjsc/re8D3YrBMkULXKPdJQm
pGnMEamkMt8eFmlAAGfI2QOnRad6zeki2UKIG+zmi6WMRyD2HsbpM0v7z78gMiw8
9S/Ba9WCvTgq1O7bUIWjyjXsR1InzLn6XJJPCbf1RXQ3bf0NxwAUPORn4JspYvq8
bdDaYF8inGumPxEhezclnxINsurIAgjXGu57y8Nn2SgppMcjNX3lIcuywMWh/gsW
9gtAwTK9A02wfOJWIJNk4lPeisVpQdT+zD3O/7huX9UmW/jQjPOqf/W+l5XZJQHw
WAeZRiNemeeheznhaFYb9DkQZz5C9OJ63qUVHFjwRfmmGwKpyrBdP18wJwT1bgr2
X8ltcZIhfc1LG1vCdo9eZ2j4a7mH3JjBPq0sFK2TxdVTSq5Hq1HmfppOn6S6vLRa
keIvtsaHXBnH4o4rmZ5BlMgw8ueyoRz+1N6ce8gAW3n2OWH1/bRUdNhppF0YkOY8
2Yq/Tg3pdSBS+U91O4u4PJABvTjWwhQ4gr37jxTb5s37jjRrK3fJCU5XLx8lZJg/
5Qdsfig87ln/eok6N9zdknGC7P5gXaBD2Ui8qbMZKwsxr4BET+SfCpFHNNjpOlcy
s45KM4y5JbhR17Z+E4J2Dg37Fq9WZeulqVg9ZqT7k7SBsLCupGbbleI4lusF1eeI
MJQftvS7TAx2u3/NouHIb/OfVq6LlSpVljxPRyiUuG1m3kjFXyOMEy7o8DDTOkJt
2P+D0fMamylJgFoIV5r767hl7IBg6UQvLTnMEod02l0WyTbjMikIJp1ts6a6kudI
7wVywqAYcyIpRXxCfMscgVA2Rh5Aw2CfRCFvNsx0dDULGP1RGiaL6LQ0zFbALChS
tvPJLqxj1yM4O9v7jn1SOY7Jsb+yPED5K21X+KBUzhjmUpuH9F8/wiAUf6bVuK1f
8eZak9ffldOq3bUgvdtdBHIepEI59QMkLrYEIYF+yZ1DN+NlLMzdOV95Da7O1jpK
llRdVTEuWSI9J9HxClAxOr5OXhcU2NxY5MSjkqRZSvcniLh7N9m5Bm+h0RTDVTcm
6d0mXiExqOqd8ULKadZeQMgo66cUl9PAb+aoHVw/D66JYmFqRHFw8O02AZsKqOtD
PXCZQ/Kl3Jpf4MS1XFOlh69cqSXm2Xv9gwRX/qu3x7yoRFRhfn8dYiyPdcp5qNt3
kOrD37PFNtJCP2gMhZpUPQXFsqoNkUSlXXOUxmQfJeUMYH5hdEQzZdm7kI31XYFY
NmeOPa/L9kVfoSkOxUAnnh2+cphCqD7efTQG7iMMK9ZnAeBfUQZ6ReUqz7LfrrJK
bxoRaMDHvTYWxtZlGVktYf56MnhVjjUOAH+8kqAw2z1pdCU19uMEEdjLd13naUYT
Gxf/zgVmFLVDR8UgEYShb1+kYyGjg0ASMi3CsBfoqmE9aMBWzyvrqfQS5OUv+L1W
Rkg7W06XqMtT8T3Jjn57PgWShIKgfY+heepCoFcwFX77nhXfDiyorDcGsimVA1X5
PM62exjSj5w04M/wIxWMVDqzXfViqzZwSrbFsTpwAoy8CXEEzjeC4zdp4X327/Kr
EQT7CL+HRP4bHP7/sxuoVvLS/6BGOfOcB64sZaAwKq8NUDSTeBPGI2sevgKVh3lL
S84Z5MpLwjCv1r4qS4rZTsv5PotV6sAkImPiTefpAz+p3y1h89bmt2rxfB/8qpKE
gUr5SyST4pLrEq9XVQk9RMs4pH3pv51jmZ68L0zN40UOyCtyXZTGKG2io1Y0S6Pk
G/1IvAaDNlh6fqr7Px9hrHZEOwJm8ujU2HSThpHbJaCeH6Pwz6mbTMWUSJX/VMC+
2j77JKeBe33SZpwARsFuSMdAjE29kGcOPv7UdxphvrDniI+cT4D0kIT4X5W+UaJD
Qv1BdHFH8fWqvRVeDYnosVnxweLpmqKZhrq3ydHBWBSFC3yJ7Ww/mgFziO2gMnlj
gKf6nacBxmrRBWzRDmOF0ev9FQSBGG6oBtuvSe3w+BUQzpPp+zCbUQYqTTeIXkTW
GixOPk0t5uIqZjwcxOgrJehkhUTAfXuZCqUm5r/ohFDfdGfxZRxw99lMMGhNj8q4
piHG8c0a/8xxUYjo+a+Y7QvcPIUenSqG8jwTdk0qLcQQnRa5u4iWJL98+XUB8A57
cVLMG+WwX3Wm30tXkUth13q0LCE0yFFCKQu5IjSYB2Fl/+XSgvlZBB4tOG4Ve1xs
C5tbvR1nJAV0QHZ/a+vE6ch1+9hUjBAhjEJqwPNwEbZdXMJJNB+9CwWoXIy/NTOx
LFFyic4FzDTvNyOG8actraGwBQf+1Djo2+pl+FkZooK1Our+oHZDCwZ8OhezwXgj
HHf6TBUcRvU8hIZLZkPgOe2ggYdflETyILlItnKgwjHpeh6syeReqD4QSnQv2sxL
9KvxeGZxQ3VtNsAeBBjPjGapeBZJR2zr0BGVvhuT6Wf9P0hcKxrYd2w8aIJUvISv
5+9uNGV+ng7saiZBNk1/3bnCwzPI3WvVBYoUHz5JMgIHqxjf42OUj1RYW8m7tsuI
eLjiATPxIXD5rIo0mMyYTfO47D3XLgIWgpvb2Z6eF9Xbt/tdr9HR63UF65oVeiri
jYxTCc455N3ei+2KRIKhUK2n8eeWQ7ZFfZ/MDdQebvLXkblzkJ93UOfcm5GPXuP3
NZKoMWtmIOlBvHRDLB9VFTwW2UVyedUtN26fBc/BFNe6DVHg+RQNifGVrqq9yYtl
Ezq1PvFOpaRqbIDZTfEJFV+MeHV5uIgd0rHmg5jaM4Yztk31OgVuMIkPI/SNLTZl
gjCkl98R1W2Q69fjBif4G5FE36GiNCBXmmH6R5bbsQmj40UvRywUw5aS3WRcLNRL
vNFNR8w3We7jN+uRM2xcsFSyC55hku2RLOPv4svY4hNw/EEgrdp3qAPfCr2KGODi
dnHVpYQNaHqVvc0wO7kGCm1twMvWI9YpKZozLZLP3VgVU4q82tKp81MG2JYWjDEm
GKrHqrwkSAopN7gi0X+kn95BUKWw4MGPSw2KCGel8Gn/vNb5lk20oASAMXfI7DpS
Fwh0g9UkeL3JhIbTqRvIVgIvXuzFvnw0QdVTU33zC4bwAGP/XMsgMGBCFq0yHc0S
/Oo02KX8lIisggsy/8Cp84/5DU7BuMUyUlPI8/SE+l9N04/IhNUykxYWPSMm0BCI
bf5usL4Y8taj3boamiczZqXwA5fEXxJwu5n70zH1/XTI45J3MDB6QOvIINhCz/zM
r2xyKsE1fjGgaryZfhGWzop+igBQWXyZQVEVeVQFv9YMl5fSjqF/wYmRmX7BBf1v
QSo3C+cwigl8DQuyagjBfUIlzfULNujtvu6277fFWtPJG8MkxV3ktYfQv6bs3nEn
0D8Q+4P1xk+Ul06oRI/dCOckajnZi2jLANXAsTYnGaqjp+Jfm/TW0w/Y+WDjAs87
4v64zGcvL9S1mxg5oy48BGfe5O2/l0BpkBH/p8joWqntsfOsaIRnPUE5tJ/udgck
0obOv1R+7NxgwNN+5oq93t0ZHPcvML+J/MChM/lmUdtyanPXTVmBfYRsib3elwWR
JUUsYt9oS6hWfnWgEXlN2bx8srzUzIOiQ2XI0vsl/rWtkwCEQliPq1SdHSYiZoV/
+8MRB017r2IL3JCVeHi3ebGxu1SJya8UzMYmJzpTCIe+bWr702RleFnp3YwA+UK7
ZQ/sXhcdjmyzG8aSXlNuVjbhnfikqqlwRIQGYLHdVYFrhOhFvp50EjJCpF5jtftz
1O1Tj6seFUF60q//9G1pneq4qSs2pOSMCqdtNx3KB6u1wSTf2iRxW8vVxY0+OYz7
zWWce1QXkLdajiUkPVMSPYH/A/Tz10P4B4Ki6fnjYZvOON3NyUYXc88oDKpmo+qz
sawaLYWVf2OzgQrDrjuTdRql64cRxC0YYgMJFav9ZuYrMTVALXV/DSODUOpDsGbY
uf7SCHHy3X0PX6EHsi5fv/q+D49Dx4c8CPMf5WeLc7zM9qq14PWXQQsdRfdqgloN
v6bq1Kgtq4NsoiHjZs37bkmg5e0x97VK0H6L0pUiuwDyKDqxwTXcPKNZdC3YCuuL
iaDJWYMscMc66qxO/tx7bFRy9fm3Krsok3Kcu7f07locfmZFuE6flYWeVxNitIsu
toQ92Nb6NoUGXoVGfVqx5SPii1zM+7hJW9N5WpTjslEsPYR/qlYMD51118sr9iYD
MfP3G+pMysKjieMPjKDHVlqBqpLo9x56CwKvgrXpyk1H9GYanBbmkXvb1KMzwKV4
2o3EFLYa1Qy8W1ZIT2f5uYlLgx4OwM2E57MwocTxNCtdhImUwoNJpW3oAz1kHPHN
16WZUjYT/47Q4JYFiLfIA8MhtBPfc6zCxLi9w8+e7g+W6nEpoTSb9Q69Nuq1r5Vq
+qbhYCF5FBsjNy3K8Ckf/Luq5KCO56IIi4YfA3qu2Juuh0bhbnoH1pf6Yytp8klT
Anzt7cXXUCorA0RW4DC97PT0HlhR77oORkgNZ/2JW/zvnRpAjR8SUJbOKloh///c
J/qLiqsWtZ1RJN/G8NJpc9eaf+gxrhwayALyUgGoyCsRwDeFdOQAZMopB6sgU7XP
uqHOwxBHgxW49wmvF0CjySH1z53ejx6yAidsz0cNueOfZeDUFgDVnL9+dSu3HYdB
bLpgvAkwLFyHNn2OgqGNmKCC3PQiokRNb2ZKpwhdzVbjfsW1ReFpFk/wpWEvXdNo
8MNpc5Hsi6fmK+4Y8xnBS1IJfczEOOY00c4SktEO1+Veqbzh1namXTLI0W2mRAEV
Y9BG5p9+Q/P91KO/Gy89i5hW+Z4JVsQtHWHt7QTCYg0XJFQ/dr2E0IA66X/7JGaV
4/kJiVqTACi24bUx8fVs8Iiddb2XCjz87y5K3oIIckknjlxiznLPwdOtcKu6eLD9
PUShvigOYACiVQbJDsiBNNKKAFxwJCEj0d0McgNYM57c/lqw37nZj9fpcxmrfBjc
gpKYmRpBd7J0vkFXNK4L73kAsXECKeP9Df7PnjGExutYm6ASwq/UpvpdiI9sszMm
BJbvoZ4BnC6LzfIqkgk4HtIqmIa2dsDqqbQv+/BzKNy3Tgz5O6lLsVLHVgoZ8j7y
45BBsjrZMRaTEaMwqThj0O5+oHkzMxNsrulLSOcqhn+zHYnNolZWnowgHb/oIoiz
Z0npdvhgtJtHvnitrMuTPONak+ek8AIdJoNJtB8I1RTyeNL2xCAKj2TDlUA/N/H9
PKGnkVd7sol0+UKmEuaKL0wgPgZ2AdgaqmlwD4BI/hjMTf+HXY5PwLSGgRQTAMUx
akB8udo407ZniIoKnhLUUxjSHzFuntr1PHJ+yx29XUu2BtzITDfWRlPmnHLkavps
7MjNtkFm1kjrKLXamM2nf5HGcBBU55IVWNTeh4jP6IKpD9Pb/M9ffkJ40rIy323w
qsYUvq8dvyTHGrNbHW5UaF8fvXncqzikIY3qyuhnLiy81V90oKDsD4yGhxUisp0L
aF0JHkrHaGpHbYMl83YU6Fcy2BpRBflDM/3ikYGhZ3TUtpTiWa92OtZ5Tv65g1fi
KkUoHaKVfu+/tMFtEy5aEQtimtoCAPkIIDRjstRTg+Y+5OCUYTahQ9TvntQSO0H4
8H8TPpnwMrFF8h0rdnTKg5GO5AIshhXi9LrmfHlB52rAjmcjL2RFOt+6wrmrfCER
qzHxC1xojv8VpzKTk5DFsMDZB0ONLZ5GlrfrmlGr/EKxQFnluw7axX1fMXjx3wdH
vayqcEhvRIamde5iSeC0LG6nIVGCsFebsintwxFOxx1R4/YLEzzmxdoSMaPMake4
iankb6OFjsGwh+q62riGDs/tLWo4MVGPvCU6rgiA1nLnL8Na8cen3LfNRbP1Qeee
HaamnRE6boCebDAo8msSVIZ0Nhn594q266rscac6ndcl5AaIw06l3ESDVzMre2R/
zp23AV6KLJgokV2OusHaPsJDI5LnW3U06a6VIlZcTu7PndD1mSuydPQLkJifn8Yv
cXEBLzi6m4q5Io8j0a3/4eTaUYWKl8tv1AGWPYKyafxALB1Mv1RwaMvbM7AP+LgZ
uquoS8jf/qU5i21XskvYsghd8SoQlnqIlH0HL5suc5E2bEYY9WM03Mw0xEO/0G0r
p2tXYt5Nkas3ZU8m2HGT7I4uZG2NYzXJxeowQKK61t2YmV1M3g2uC1cGvZuosYY4
kvzfLjGHF1IEKzLC7XHo+G7FW9KBalwOtY/dqQhsSi6sUxZEXnOsS8aIuwylZWfj
DbL9+GBmnrVByv7jP6oyRceTa9xGdEKVEyRB8e8PuuyBlNeAqSCvavCiHETGKqbE
qyYEPnGoF+QkfZJX1dN67Ep5wGJEOtSpA9Jdb+wsN4sxL1bM/78Ujtz1YmRKfUYm
UUOMFTQ2J3A9LFmnFScKkLFXgPQqIVfXUDiG0dMtsD2dWrX7WICMs8P2yGjUMfUC
9+kvUiJmZs8uYWDes7lzLhcmpbjqaYIE7ly/OEME/asKbpFDoKKic4yjku3itFwn
bhGwfS3rp/HqJz2/KmyTAYRzmUXg2Kg7adAmMy7TwoMfjos2V/bwrHfFbuU6omg4
+5jNgQWu9oYGQFislVQChdikT7WFMILd5hEP7aG17kxNgGg0Y5bcIpV4yX6rq1+2
3mTAbH3Sk9NlByL7AtBkfwJekI/nE7Aj6msixB9CFoWEXlXUbtk1jPjQl+UgIJKg
G9//Prz4tbBABpxN5vRvi+m/g1iF0qFO2Svi+ID6RjENFk3gXPEVLaS6zvXL4l4p
vCbmjAFO+XeK8Hx715S33/3ql4yhRWd4aSAPOFbM/PJ0eLTHdJfltnfrlV5uKd5l
rFRwjRhtRwsdLbByTbUu+MWaW7vsp5KO4FNncCzPxakDXSDQaXHPOAf2LowG1XZ2
Le/3DLA6Jx1zuI9EFbEf+Rk7zpeWdUZg2s4a8OgYiKf5ni8GHLQQXBmoO6DLljkQ
AUNxL2/zwMRIZ033nXWNAC6yl2brYMEPUd0FDHqLC/OHqNuwzu63aklggC+Dg3De
vLu3DAa05Hyhh5DbsUFdTnRreqFw9Tk31PaULfQauNnUO1N6rezYgocs7Ba19OwX
zSIZvM38m4w3W8xX6HhWhocs82rApuCXyNN8Gs3KNJnTvxqGC3mFVvgNvSD11kz4
/t7ozf2DR1G5XYv9w9EFaILnt4xVkmLIjwi1ZMsKoi+6J3qz0MdzCrk79s5klxzH
RJW0pg3r3D3A1Wmet5eDihvb/cCdD1ori2BGuJlz2DWBZYzV1hPrBMOY9gZCbrET
LYD3CvPI8eub8wQZ6wX/+0ZzSSxTWgyYA8YEua6pSV8h9FMJVzd6K//lSrY0t0TL
Zgv0GwKH/UzTs3YMu1SkUDdiJJRHp8oJ1BHC2hr89+GbLMdOOy9VHOr9IcW8sBEb
UhhJtxuLiQoXiiRlBiUzkvRqjiz5HHgRp5REayNdNryMbDZDRPtAhygfVE2OyU/J
RlJ3obEVHM7iUYpiwtXTQG1ntjhegfEO8mfB1CNRtkqzBV3ZUvNNNtMFzfWJcYwr
j3gSCX7AYl+OA/OV6LaDCILDP8fEZ3E3HwplkWrqSXXKDhtUBSPXEJ9EQt6CUQCN
MLP1/TsUJgsB5rCvu5KDUn6J5Kt0PrafCsdGwx+1pVK8nEFV4DXu7AAFxUPNFYeg
cHzk+vtAnhKpShsxT+8B7Pu6sGpLnIj+CO/Zn813PqAE1miLoMC9fLBM2hrZNDDe
jrhtT58hoi34HHx7GEfx0f+3ed2l32Lv2Y77S0Eon0ibbR68XDxcGDhVr78fOCEC
H8lw0scH1mly7g3eY3aABIih6SI4JrwLMVkMgWpSKUBxG7UTHziR7iTNzHO9meLQ
LgosrKmNzqd5FxxZxWB6T2qfYCTOYHEKGsd/2MezfQVCWi+kcIF8CohrgP45Xcbr
uRK64Ug/QaRb1CBNv53Rg8P4DvBSA2RRyodkuTQAK4Kz8hhB5bxmtG50jbLEHKz/
zXWFUaWisFMwak62NJyKlfNG4m902V1xSb4RbYEuu0FoVmON2MiPf4xGoGy3xYgr
8nFQ92peedKDfq7DNVciXXuMB4HKBOkKY8fR1CPBKXw/zb6+mW++soYTqaqUtzdG
BCkpvVdElZFNq3mRYA7oFfvV+6nVudn3tvyvC/PLVOnQAy5YzCyVVY1W321nw0n1
mTHwwgnRQowQ7R9xDMgJMu7ULuW+R1H1ZogqYvdrnEvAa9dirVCllgsh25wlD647
WWAOk9LHeM7TeW4AH77QK+VJpdp9W5UNYVVjCxkcHTmimWUYqnVMAhZ0iE61vV+v
feUyEbbrL8n6tHGLncwBlydHJl5tgOUCn+bP/bNfD1Cz3o7cKg57Dyf4BsW5Hshc
6VUJqFmQO4b3GCAZeEvsK+MRw82mzipga5XGTHVYCoKi2c7RP4S+EjW5KpBQKWe7
hVKVKeeUEeXQAR0SMKEXem+eKpBp/PyefIC/4bj7GgGt6ERqA8hfPfBLebCvjSUw
lx7D1rsbpdCEbwiulAjlFdlEBTUReY9bWSQkJHwj7v+jwHIHOFSw+mYWu+cvh1bo
kb5r/n4KSRCJNvBoWXRvu4bMSFYGLkICAWp/L3vVOI4RhcvcR/noXUFQ6InOGlE2
hHv61IOWX1x6vaCwE5QzKpjx4pdY52TKqMVvzo2n2qahUdTuB+TtzsoA5oJXGrsU
ez69G93OcIrA5yV2yqimUfipMqRSiyJc3ulJPY5BscesqRZp7qag+TPMx6msbjlL
zoK+LugB+1YzkWmEBNuIWa3hIq9w/9kEObx4/B6TcIyYp6LepPNzQbVmU8OAbC5v
WbLckSBn9IJpUkjaA2r/XTjLmpHFlL4HkzjFGOxO9siuJb93SEM0JKfJgXV3/9Zn
kFN4w/HKuVBDluA/9YjMTAYpfBvHJcQAtUdGzSXxGcQdhie6uTWY9N9qTavcUPTk
KcrdwYzYRDdTZjlv0ntwGxmnu51oXSv8dpAIadp24wbQlN0ocGYImDWnafCBjrwr
13/VsfAwu+R99xuHqiuzVw3gkgqATiOj6sKJJvPhIOZ3rFneXeMH/40kpGKfhcr8
vKwM5Ufv3p+I9yhNh+aDWKJ2GrSpH5plZswsfL+Te6sXiZMnOAhD8/mFW98fiVgn
1bY0e/Rx3pUaXqwH9GO16iF+z/B2gBKqM0o4QUN0E5eadOVzAlYXkIvg9vuavTDr
dyApa+ONRxBv8duDsTrrMSle37gtp0LbM1TQbpMuMzZ/hypvoWBQxtHR0V5v78hR
wKkaK25FOMDZOo5Chyei00WsBXZqBjjsGI/KpewEZr9vm137t6pngDwa3gp3i82l
INCSgY04RBTSYcXlC0koLkHR6AbcYKhhnOqqXDbrcGTIpZJlHlf5EsNPYbC7kK/s
I7HiooOblZVjRaEEeCMPQ1T1rbfQiJ2ReMvVVmXtV2GKw2Y/48Az4coRbE79icRa
l52N5w133wruwi0cjcwOwD5ARmJf01c8rp5JSgOpLN0vHCc6T0TJalYcdCr7jhqE
9p1jI7etZXDy1wg2QAsfKoyD/W/ScKB8k4SzLmUdIvKWTCiYM2q4gLvgJ2Q6urUW
wIPn1SBue1TKwbldaHOnobpivN4isgXqzgoGCPCn1v2f4DnC+YbW1UXScxi+hNQ5
bZYV3/YPWwL1xYtprZQO35gyXFAmahZ8IM+zjMDRk2ia3l8fPx+m4V8OZIu7t/oN
Jt+YGscXxDcH+PQ3/d5UvIUcMVsnqisaucyJ0HiPUiNhcFTQwzIQ4oNiVoUPpSuq
Awl9eLyQpUMt8sD6WBXFjRmSs9F4SuguCbaZ6yKxOaIBbH+DbxHozSbEN71eHCRY
L0lWvEY5uBKtD5bP4vSmxAv6e/SuKF/aR8vY5NV0jiUgQ61uZXv11IH4E03Kplro
uLn/g0mN9ugxv3obkeYty/WegiIAHwSWxBetYP0JObafQyolB5JLttcZjH5SKnrW
NfK5HpMevogfq4whTP0LJJgdy7jSUj5QqAI4w9VnvKSvawV4IzHl6ypnpKPdZOIs
dx22jYKKgh9gqO8S58Ry3X6CJUsVh6hrP6ZTFzwRFOox6YfHtPVKgkSv2bje9ufu
gjsV53tYejhJlOPi+v/6f7Efj4TfmJ6tEFuNwq7sBxvaTaF6UJsRmCctijdAJPHo
E3/Ai4VG6Blo9g3G0PbeB5kR0T+P1RT9jA5UTn4X60To8bQnOYwUruCwySg8bVkC
7J1Hcyu/IQ1E4jVwffjk7hsGz6yYbqFJN0x6G2jlK8+qOOO7Xu8UlDYQHD0/I1Nm
n3fTcChEhD1kp2kiX6R77z0STIjUTnWnD2kUtLz/SPOY3tiwK6fhX4UjsiRX4grV
wpXR2qDVUC5V9Tey670fIRU1KS5CMQ8BQRlaUQpECgMIGzj0kcKDu2V1EaYWbYzl
dL3K5VnhopW9Y7cO8CosIbtKZTNaD9VN9k/sS0cS1VZGrz5Bi7PWOt1qXssRl3ri
GLAz6YO4uUQcZ09CqEpG9Jgs0NDF1UvbokueRtTwGiZByNNiwxQG2j773zsa/sXH
uOcOLp2yO79x1HSpBZiDMkyU64VDOsf2z5wwmQ9GpzahVox8meZscAlo2evHXOca
l0VVmIjIzc3Ctfd9WQJkhJBHNRqoKKEGXtjmbcmiL65dQ9qRTCn1nyuiMtZKxlhU
r8Wb7p5MvYgXkaRjnmhbf6AE6z8dEGeHGyAcZzlu0UZx+6uBABDqS/3RAMd/nH/v
RleRtxaPFHjLO55Wd8oOs7mL1BBwWG2JiMTQBEID7O2mkWx7WRaf4LXCt0sMrasY
k/sV9LA/jF9VCoCxEVv1RnZErZxO43kOU9geLErPS5AtJg/z+KpqJqg+w1/Zl++T
pwmYWhEHbQbZdcQAagxExWsNKhWn39iFFb0A3JMpX/bxWtyDVXColKQCkpz4ISxW
aY91MlaLp2V/jUT4hzt55QCk3Y9vYQiq8g0FpWGxAQZDuSUDKSnGK5LSgUTdFv5+
/Yj+PgErcYDfS6Jvt/1/Odd+WLzzFRi5WUnTk/QH7VEfcfE5o9TD9QmP/j11HqxN
Tnt1wG3pAySaWiAr37zV0MmvJ9Gi+zqzLJFLzLtnCwudNMqjon7qQ9tcZ5gAwZoX
P4risEmwHdQO76FdCiCJGfiW5LP3ZCwyd2DPtLSRPjpy0pLtxzI0gThMi/isAmcl
s0Q7mnFRgRoJUIJJE58AdznQtoggfvxXTZfVThA0qnTedqoFrz7B0aDaEsZ/R9oe
ecIz79rZjsnij9A0ZVwuxKEz7IGe7GCvU7DlHAe9q/07X+H8nDdXLHwaxPQzS/1S
IW1koObWaFNB3GcoD++CWtFXvXQRoFUBa0AouzqchE0JzW/Psutwr+4CkDdl7VNW
O4u0KGwKhqZMnF4eRRsxiOt1ylazBCE0z0hiWwwV1CrWJ/GXGdOtNS6W01pPovsX
u8UMrYnidVSz0GTs7bWM/kHfY4xQsv+9H9J3mfHHB/VOi3vNbIBCfce5sisxZsvd
hhUhjGUtkgXkRyAie0rpClkpzO0UzxFyie5HhjwhaZjo24P0FuQvvEDCDbuIWblF
bAKRaVCQdIP0+2CY+AkooUW1J5/t8VUOliIlMX/ERMNVdNns+0zOET/6zWL16EMH
v9WxgEbTzDTxm724MdPmanvHV7s/A0SwOfFlgXmTiL5rysLEEI3/IWuEa3xumXkC
9Qa39XlXegLj/wy238HFE1oe3T+eZ3bOihMCal5GA2jsJnjd/Q6K8EcVoJh+TWW/
vscloBmeIT5kx0x1+Tdm9g6ML6XohFVuXggpT8mOSPFtph1GhijY16H37wu7N8dZ
KgyhU15WAwH6xnrrpKys+lXWtKkPpNi+bk0FA2cVURaA3jx83fUOEZknod0Ow/8m
NcrtgrxsWOfh0oNYZph2lPvHV86zhHsh/sbWyXqsoolxMVQYsffJki9AYS05jCom
bq6cdh0SxatpWpUSuxriEs6mjT9VisUYpo3CqRG31du060niQUtAfXxfPiKgVt2v
Gohy2NU3yhOEqzG21J6CUFogw3r8rL4BSwtDuPwFgRecaADbcvwv0RbNlntL+oOl
PNr1FZhMBDAu67zY5+5mkaIwem+ltY4laAqifoqsQ1h8AAy3UuM2QeUuPW8i16cA
JMZ3GH8blyq40dq97gu1Bal0tKjwG1PSLXRdjjAcTkyn5DOIOO2kRqgVqaP/p8ia
jYgg5RzZs5+Pt801Nm2dDxSvglYCdufiY/pqx6uSgYA+MiA35XBBC1p4MCOP4c7s
gpxhLlvpAbU7NUoUN8e8VRekhDH2qysgTX6EvJVypueXWLbPJATXWoUYaSae7yPr
vQIuUoDJl/za9CVYzRzCfz0AlQSxJGf3OAtSQRNuiY7WbUa7GRzqXN7HfgAdFWXj
KpN8jlXTIyhGEgR53JT0zUNRd8FytIjx43Ss5wV4vvrcjXDaYc/JepxLPKfnhaAU
gz0gVaUrIXH8l+RvXAsdAaabhTm8ReZHmzXW9oQOijxuQJmigdZZ5thw+EXQo5vP
EH4scEdFbE+eClrs/T4nmUSCcT2V/TT/TUD2WzgrG0oOM8EBQcKWSQ+QITkq/Xnf
ECH8VuXAgN6HvBy+CFM3y7CCtPd+s0VMudbxXcC9frxCNmJgIy62Ryvx3COicoyQ
TzqyU871d2DOdq9GCPYwwcnZNTKHp7zkv3MW9sqZhYFr4JNWr4zaxQfRfMjjM1mC
h7Fqmkd7zaER6uQIJirNJS5+U90BCSNCAWqAxsrz2IR7jBU3ntkTDRYVbzq+Jk46
0fUxwWURWn0ckN1klD3oDZhCoxpGpO2BRlVhidEZFT1HGEMjn0vtfjaUw8tYRykg
M36jsm75kjGxCQfOK+qujdwIr9Ln29+klleKDgB/GAG5B0GT2STLcnX00avJ5n16
G7hyzkRVWlgEektTeHQcXTR1+DEz7/pjGZUfo3CT4+dsLuxQHxSfoJd9EGmN6n2v
X8IiAfrYi+zlBlOPFxltMhebeOQGTTZI+UipzujH5DbyNC4ADIcseMW9Zjm7URN0
bsal5GHcPkW9oGZeO8hXJCXM7xmtGvX3dKTD/MQc2DqAnBejRqwbRtvARRvmGNeK
wuOiWHN74Ng3z04Dv2+AxNTUXwrP0Aq83aLuXStiTUP/F4K6ntrAors8NDi+fLVk
/3PVH34jy+y9sdLJ1qQd6NQCmjm37/bZGmhOffX618I2yDldqthZ19JybQT/dCBe
Xh2mkXT25BDAkf0g8SscM4by86sub4FyO+GBaAHL8+NGMZzU5XYLfyVIcRdHshX9
XsX09KaUmQIDRyKt/UaL1zy3hdgCj190HNOFbWqIyLxIZSI+DdHufDsoOg5Dp+8X
EeWYD8RJYMNGy6aHGAi27FKnBX5FEWxVP+S4YiBbFa9DfbgFsb2LQjWSdZ8OcpJJ
zwRRbHSpP5vVvRPaEQM6VdXafhT03N0YtGyUkdIrtMdIGJkA6csmca5sqdiY3fHi
BUSRGS87hQCsDDf1gCAuAv+WLCnRlAFzi32sjsfolI+vDNoLwuZZquCczaUKaEnn
5ogYDMs40iH/4t1fQJWvDWLF8r+iPdG1rBO+tklmT2WcOXaJ+PSpmUoMCHwcNscL
qgWoPrvCiIM6GUFSIs+wjIG9gOFWpAfzj6mJXPA7shISAcEH35BW6/3A3RGv7cNI
5mDPW0pCAkEONxjNU2+MQurTlp+YGdTPh+LAiNrCQevf/BRIiT5NN2u6SohSM7FO
9tLnHJNwO/VubTc1A3AsM7hfK8sDDbi571C5vhfCjOfUoCuKYgfUKt927srCPdmU
LACtvxI3RIdObdxKRkG3J3vmjcdl7urMlpK2YmKuWvui+HJA8VEQSw2r7E9JB2vL
NGsbkDYw6YrL4d66cTJz8eiKl2jN8/N7D1yOfX2etGBwRLgZRqR6pvnaGKRNHDuS
HQmICX3Kn0gRhSynsugfQDaFViiENapTBSuXEaUIWu74HSJtckfiA6y/xRx4iGc2
kIQT57YMOed52O632kLN8JndoNbDZ0nqoCP6NJZZkECTSj3PhHTsCCcIoRuZbEEe
UtKA77SCcpwlOyO1lrGMfB2gBFY34kOkPXQhbb9tEI1KkTbUz456zmIPY0DPU5pX
JjiNvjmCWmeH904F3iWBWDe8Xu8nNAzR+eE9m13u/pT54ftzJhlhl4bpYR5hJ6nF
IOmhu3nQaYKMXpuITzYhKhxIyOu0qPOfW3eCWr7gGRn3aYQEji+JX/nrifisY7YQ
wmH1hqcdUsegKysMP2RXOPjgXT0fLj5v3+w+eUM418J+HKkevJFOkHgZi8VcWBhV
6/wheK+izV4hTyzh0Q04IRTooYkqnDGG5VLpAPRh8cN7uV5q7p/+Eajt6gDCg78M
P9aLOuxrH1gNCswsxF4xIKSvXbJpX1FrE7N5e/jO1Kah8CNkdb5qz9FwgGqdVwMr
iNkyHuRQfLYKv/kt/hJJlLcxHp69DELLliQKq4W4oteu0PwtWol43n+ZGqcFTJJX
z6SXHH+qwcklqC+F2Fe83Ysel9UMvsKKo+xKIzp0+Z+58RKV3t35Kir86z9pWz6r
8InPWO+E9dM4OQifc9jO7tNOhfV6GN64fuOwlLAgxsTiuRKxp1uPLP2pLa4SXUuG
EhLgLD1Z6Lg2VYjl0ck+Tpy7uyO9AXB4JZtn4BmcQ0dgYECJ5UZz51MSm+U5rwpw
42N+DE8JqCldJvpbZtZO2MGj1S3EIHQW55x98MRic3Es7S7DCmISbiTqwjaz15qX
PQ9TdYT1BBdfTyImzAx5uZnJu8AVeHUErmYDcAyvi8DYraJDOiKaA5kUJ8N7+/iW
OihmUMN4niTiZLPuQ2t2j//3zz71Rhz5PHR7T7akILXTkyUsEO6Q0aA2yvnOIW/+
3JJ/A8gF3ifnZIH1IbPCxuk37bAjJ7W8a8pBMwo3x2VyWGWkniKTZ+q7krHyy3LN
nBfE57UhiTksfET8GZ7Gu/KOmCZsM+Yx9z1vTWwxKdQcvFjjDMjJD9+/UcSfXoNv
mxbiJkI5W65jbr+zE0F6XEjSzttelupPhZQVZahCj4xb9uSoUuzskp2QqzNG+4ut
++9bgzo5b5pUDuXoNN2xmY93i4phMQd8Ng3ZK1lfDn5NfgENmvz8NpZCEd46SBlg
4LUqULoWHc3kNEUPp9YRbLQPArL5jADf7M8iB4HJVp2R/xIIZ0wzY9z1crpA0mWQ
C7G8chJKf2uWtV0BAQlnBpQbMZXfn7Ud8ctTPLXj84jjDP26hJYxkO2qXYrX57wC
pCOb21wKd/WE5OTREwzUkuIDGAPVUmriFrtVUhu3CMWQucMcj9fX99NvJCdikG8f
QnXjEmrxbEP9sQ4CWntbDc0rhhzgWuaIJYfUZwI/tEJ8w1wEum5JqTg6DNlgYkpk
KuIVCfPwPh5Bl0vSg83kFADKvRFpl1VP+dXwWJpjxd+3kunCWwkwVJNSMeS01LBK
y7jZVpG77pOTCPLe23oNOjNJJx/iqaYN088BDVNVSM6b3Be20nL7PcOR0MhvXb7n
dDNXuWZF3rA6DvO9d04MCgUc4nU743+JONgDlenCtDIcvnLRg8B+fN0Rx7HnoZP3
c5gm+DI4zZ+Wh3gLrvoEN9WJsCy9w3lo31cPd8bG9JyFltawGQfC78Es7M5uT13S
vbC9XdhSSHBqZZghvskE2xSvZPxf4euA4W5J4GM5ybFwyfHT3wXL4wkD/DX8qNPr
YBWHc7wXO10sCdLH89pnylNeUHft0p7pvskAmJSnILvM/9x8juPnmJ3PDKwjm0CN
kdj4ssnzZTX1H2cqCudd6QHVvp/LEzphwgPDBMF8FAruUGMvrELOAuSQ0CBd+gad
NBW9BI5yHEn4uC72gyy8m1F1z05HwlSWoeJEbOhfI7hstwHnBWl+n4kMu3U8JFr5
LnycA9Vk8hzcwv9Ss74VT1ZgYUXHUIISJ5M9DqI2i1H/pGublz3ttiFh+mI7LGNF
bGUVKvL+5IbU7+seEyAkgP9imz3yvQwyKD6NZdYybcVCX5BupbVtYGP3lZ/UWHz5
KX5dwTqbtSkKu9/pS739LbqcX2kp+UGAZS5nHv/ITCkjbi4o9PVC8IME4If/gNTE
XuSSM6yKEsTa8NoNEZXRSBL34/a57jKBuevkWQfYLTlStBzCqV71fhxOuhH6CXsb
PO6Z8AKmHPm26Vrx6JSi3dPeRalKI52NMqYIg+HxLqONr1o+kM17M/OpXTO/qWfs
I6hgUTNwLUXvpCQqTt8Td0xCL5Jlq5x3XH4yH8qjG0t3+/V5ZmKKwSBkafRjlmim
YMIECNZpa/wi2QeNPb1bB4SWWN6+UVXOMgXcRpovG1hE8BoYxUMMoSMDxYzt7fOY
bh+9W9BKFi5lEreP5ajbOO5rz2uwPRSjmIOmDO+ZoLpiA753YcVmcm1ksi+2aZsI
zgH+cW2XZ342j10fNaIwnNP2oJUD5GEjr33Eedj9Dwa0FMM6IUenFyv3cPg8jQJb
SFf5wWMgK/8H+DGTwugH4QLPZqJGJy9i7mRTUx3PtAw7hni4k9ZA/99Trm7H+j2D
E6q006uVEc+L7jlgXDigoKDSdwOnf96NXZMa0h+mdkj24pPvbbiJKhUL5p+ukMvt
UbHejlCUaqJFj1Z3RshWVMTQeoUlq8UyWtcHcP6fi7JbDocywF/ympa35cO8ekCz
omgG+2QJy+PTCupToAqpbRjQmGDdkaizxOYXaQkPdnzj6pXh7/2wCaKzn5vb+qkq
vgDW6+gqIKM9l0wObA5Xotul03fbPRR1WZZFWA51zXA7NOUOxtfYDgKtsmwjugAw
H1xf/Lk9pWZqN64Y0IWXq+fOlR44UZW5FECMMpI7xyVwW70Iam0/LRDcR/AezGrS
iK8gHYikxkQuSLCwsBusiySen/Loft5KvRFfp+niG1fXJDNJApBfwO8S1bfUvObr
ekpbL9u/pskHN9TZj7x4HRy++tQIKmHZH3bgbF4Sr3Su51HKtcmlQPyJ3zZhKX0i
r7fx3xqMTGuTs1dTfqzsbLI8voaSURCSTNTOCGUa7cjqdiPx2Mq8qHNjrWDEz8cy
EtmPEUbhojSx0CfnYI5MmzVlqbthSHpS5cHX6HYRH01Wngs0pHtNLGdFwuVOkiaT
EL+jNKt0UxV0XGnytSvTt1bQXyZsCqfF5rh7LKnNCJw+NbcpRvqIT9lVzKqb+ZD5
fmfr7SxihVQS97YMwJKEoBpdX4mb9ve2UYvQe4TIuHt1vTS5nItfLk2wfzbDhbVf
HaJ1Ou0z4YP4tMB4cyburil31Es1ugf+3nhyiTjNp47VpOlhuQSrVv7g9ZbJPKOr
KllPyGAKJWWjPH5jxUlAe1wQ/qA0KypyucFEp7ujQemHLTUOWEA/yaxu3oHNXLwJ
HjaP7ZzJ8scUMnhRrbBKMN1fTjNL2hIifSDNNtJrmywgUpyijMw1FOV0ujTn3fvo
PVKky8rJbjldAG+oGBNDslJWr7ch9jAuXOrar9jhzllMCQWz7Fcd3RrK8zQG1sOh
mm0/k/lm0TUuW6sq1so1s3clnKOxor7G/V+IaO/CXs+61uZUD62Z8lT4lQMhIS5S
ieXlLOa3V9MEQ27ieEyTYHwWZugOisP0EPqkXWLbcoZQVJiIAZr3Def+L24uOpFi
e74A3aJxb9eX0DMNLirgE28eBSA8spd7M154dCpT1swhE/hlvh4t7QcUqNC+ytdl
TxPZ/N5PI3WEqB7rtrvB14EF81WEjoPDHI+PiiIkVdPwWrlt/w5OVa3CUAnKM3bK
fht4wtWCzkEcq/w7hYAqYq/M7qIyoWDQ1JWBBZD2/MGSqCIWFWKtzygq3kXFa/VS
5YHXFb2/gk4Oe/Cfv3ons4uQuKcohegx/QuUXmW3uFZLmSNHMbdWPi372Rsg4WYm
u0FBTcSzVUZpE2/vGYESG06xwdzkpp0ceBhEjcbMt2nfMQhGdVXB3eBs3X4/Gq/K
i01pkxNs0opZCAQlPX4okT+JZiDSEJQhsSP5TUOF0ETNXG0Ic41kSMVhp19FzFKh
tBngVXOpu6wamrjAtpRiUBUBhOwYxaPmrCNVe0LZ0dc57JA1eaCL6St+hEZWY4vW
lBe+BLcWKgyERSKSt2JYyutuwYNL7qgcMXqQPC5KpflcmCn+euL1vhBh2WnWo1ks
tBIuv9u+PUedTC6YBtearCtMIFGPHlc20j0veOnLi0AHaZX3JXy+z1TeqOKs4wwk
hhYUV04imu9O6Q+dAYBl/qjMK0QlBY3p58vLvEUqYprb47ayGwp8KPe0JWnxc/cL
eiiB4M6xGJ8w+5TZTXYGi15N3pvNZXIXtR03Fhr57UNo1/oyU4CGQ/8K1U2+LPo7
/Sie4chenMwwOesHSVCTPRjZ1WHs9lUIO9BUbobDlbE3LdUrU9ALwJFyWYW1iaS1
H2hAau9BVwebCkvL9+B9bJN+JZyF7Nva8qUcNrclT2hPhixJqo7nc6cWf/FrvJMy
8QEMTE5oBt+SFsZPijZrVfeGPZ/Jt4PqIpxXWc54Tw6CBqJIHULIeA3AJYrEueXp
yNVOXbwIWfLsbOT70RlExiAr4yV6Ke+8Mqi0qrFWiI1cGvrHgiu6CJqfIWNDtq6j
yGgA+Kzt1wPEM1I7t3r5mYbGPEmG+3lySK0M55wa6l5wUVxLlM1euC7vs2YGxcTk
EG6Ec8VryIx4eE+oCuJkKG9ROMmG8oZtQigj8nlovnFQR1YRzgkfUw5kU2KVirPh
X5xe2JEyKny5RuXGTvVnmH9jFHB4VKRPEpPFS8Tk8KPMnQZ71+fBRYM3ivoSZwhf
IxfM9OMKcHt9F0NTzzBSTUiQZAUOmT5vi+vy0Pt9NWCjUAsldPmwhGfDNffywYes
dPzZkQcPawFOLN9TmtCbs2Hfn7AXErrRP4JWhjej1VdYdTptMnI5PCkL+GPBf94w
AqhYkwgVI5xufHetMBapYlDfRoYS/zknyLjabDRksB32gVtjqUjO8+uP/4aJW+tY
+kR/rMpqSVVXgAmOipdGKSwGUcKSZMoaw1HnaZzliucReLmMasYp2Tn5nZ7+NT0h
dO1sQtTRMQkub4Fh4J2i4257ieosdVyxN+wYNBKxid6E0hFyzCvtemP4//6102Em
7uHF8DGe3YdVfh9CIqhgpKZjkAUxIh3gyaMyYgG+jlNfLa9G2sNUlehBbb51DAu3
u84okKnydlQPEjCKbSlJQODFGNwA+DX1zI9zrXo/WCFZzxrDjRKpXH4G8Qld5j8K
elEv2y3sukBdp6qE9BSodRrUSou/uYEqqRlGHROzgx0eaGe/ILeY31nKY3e47gD2
XUmFDiN4UKE2G2sVvfrFHVkPga3k+jaE2FYD4Wxh0Br5a6Kve6sYnz7riIhfyVbR
5tAaakMdkQ3S9y1HiEbNMv3S/IPbZQHfaptViaiNywCsG7EIAp2nVIgGtd74B+X/
+x40Cu3BlQVdaN3NVW8sGA+C9xnRyM5s2e19sLv+KYPptr8TP1OQbSsyjp2wK26v
BG0eX+NGB5vATWULSPS9VdMtptQdRk5a9mzcW5CXZUMiOjsmLXarptKS85Tr4MvC
PBh8PJ1bfE9cHfZkXaGEDtyMR6QLnM9z+7J3H9cYmQ1hsV7uBc2dpvlPiaPzrGK2
7Ey0w0SAtunI3uVXw9SBbRk4AfnOzSRIojkwsy519bKCfAbC1Aj0cBEzddweH017
A53VJY5oCB/Uy8ZjjW3V1andHYBL285xYmjlvqnTQGuZ9tE/xt2QbUdCyZjMC/dJ
CJqmuMAELwZ+jivbgp8sDuddkfRhSr4Al1q5c1gUnRo+Ylq8fLjFaL0/iFdjR1fw
pzx6FI9gOWbUlPgZVz1GvAWBo8/DOXEXnKr18OBbGDgUmH0YvoSGxkXVt1Qf87aW
uKnW+8TOj2q7mPU4yS4vQYp8rWQFzmyvxebOfmns9FhyTrFxtK4dgEevDciTrTQX
kiLW6udSuPKTaXIuBXKCHfOU8d7K8o5PPwq1iqTsadKNlFZkji4FHeh6d4aYkLtI
wwSEUSdeV4yJvRob7Jy9zLv4RN/1y6ddg4dmhH/y9VGqJZyhhGzGGLdW1aetfGnS
tVUlrZaQz4V6Nslbnrl1vBW6vluPf88/1Ep+z8YXlABUjecfBzzfbByAzWa7U4iH
Ac+11YtNXZJD4A5iuyzruCZTgOVDjoY6967odq5+RjWuxcZQ/+MXN98KTb5BFdPB
yqolaYDITdJ07j9Io8RaAz6KAfv2qOwcXKejZi9DSRyL8vo2u85eTi8TzjkeUQam
EHzH6SalRtjiO5WEn8HtstKfvqQgYzEb9Og9LeP2tabPtf/nOxOTrD1rRVui18dR
+e/j7QECPwZv/EXHoEGubNH00kJ3SAyjQtZ4NBuH0FvkW5mjJIqjRXwliLmDOQer
w8NhyGKLsvndetZjY4vX/oWUlRXhrX1Yih/mKyVkT60n7GqpTiqC06F+8AIkjaVS
E0G8AomWpfzk+1tRc3exlM2WOcI1Yp5ZDIL/lWYn+DPEbLaRQfSSWJpSDhbdFfjA
iMNzEg+SvcCq283yR35Lca1kNngU+AxiqBOoXHqWMxTxrn7ulfnv+XPfEmqEZNk8
5TashGjDJj+AVuqxVDtN6kG+Y5NViVg++2rBh04kV8yjkU3xrnBX3PzPUedSBqLv
byy5c3jn1P6G4ljAJiAoAMxm1mMPih7B8gvB6ApRvCBpNoHsFnGpJONgBO7w8j3W
kk3REPkNrS5yAjBqKj3E79vn0UajdV7E9UmCKiR6VIMuQCA2K+1/VU5C1hi4aPml
LM4wLCUZjcOUTwsBKRvltwCwv7ZjBob4z1qqtNy0C6kUEypf2W77f2roJEzDObXa
61O90g3Xo20X0nTQvkiPdwUzxfUHYmcpkiCdfBZywXkve7zE4kiZdLtBXEwY/XMF
u0KHZvFANENlwYVUiJfowfZji8PrY8+j9iSp5sR7ZyExSJOslY9bb31mORVFjqVa
KwjcvSBHfmXlnG7b/1ZA8rdak0s6d4frwYad9e4gOTJ9R71KbanI85+sMtNFkXTh
1FzT2iDu2tKyN8D1P8CtNLfn2nz9/zihxAH421TAhd/WAawMUg+KYOMSQ2kydMHb
zFIMzhNZ3OPc8QSpvXP4hqasUuaxsBYf2M4cYlRklNtpOqgXJ4mB39ir4p1alchS
zuilIGEF4AxXoVYnA7ZE1bdbT8Cs8ZiOM1P1azt4FAIpjIXtp6yM5BibQ/FTyXiU
iEwp1QjI6uxNinr4HWTcRg+2+ZN84GKBKpF1Xa3FeP0t/Wg7i1JnWKHEzO6fC5Kr
69vsu9BpVb8PnWGdcuPgtbEJu6TvoAbVm9UwqmNgJY6FOhElFIygDEdKtnex/FOk
TDyipXpyIl0T1fcCStoImtM3VAK3mvBLiwUHeJJnBshYVQUFGaUpz5Cmo7NsnId8
vOeV4WggA72JZzDWapoMCT+kcm47IUedCU2DLQ8rX02I+x9haahahe65n8JsspxG
SkJm7jz5uYRDex0lcLGZIdsZoKCrE1gbrAvSMMMVX+Vhl6CG/Yk57GrwDOffZ0zh
3asSNXNSHr0ip5PeXFsoPJpF2S5yVW43p47NFMRj13oSXMsp4IvqfQymivKG2Cm+
E5k877FCp5vCRLyPob7dRXbhUbKYu0x4nXTozG7SwBUEnMDpqGYLoQfXbnayloh7
SXbJBEYmPMxB+vXy2vW41nJND5Vlgbwl/yq417kQLRo2mYLwe6x5kckGXYN1hwKn
NB6s9lOsi/HyJPyq7m5qMsactUkVRHFWkstqn1g1te22+SApAgu54B5seIW6sQdX
PN27+z7SLSpiN9UWPnHQ/gKJ///abmLw5joOvNH+R/nJxD0pthFrKxTqbuqk4/DP
AVTvLbo8yO+hvRFD6tjPucNG2ulk6oEP6I3wiHcnzN+NJ4uxWZ6jV7tgN2+lEvsL
U+PXUTluc7Sk5MqGQ5UvCWBk+bAWnlSX695/Zkjs+khhHgH8b3np6Mi3ERM2j/qw
IxGXbTbU7YuqwhZDdhIbF1ePCpJ5aTobv5zOUWKaCUGflw/8Ixi8XccLAuXF8Pjy
mcUyTLLqWcf+f2WzviMmVgowiQI4lekIz/Aj4DGxO3iugrCmUOEcHBNn3XvF7fmI
alKuqoDaeUoY4/dJXiu6JLZZXETwjRFK1qH88Hw+o0MG4dlQBCAWIjo1WX83VfuZ
DqWMufE6tLREj8n9OD3DwgExdgtX9iC/g0e1RMdKwvmadBK72nDw45Cq9FeMXq5C
0W0BIkiI/AUVpS/FeEXk3RE4iZvfB8PUsGZnW5Q6gm+kruHyg70BbAPv2uRVvHDj
KQwu3V7YE78oN20UfFW3Lty9c8uJfXjv/L58iHdRylH2a0N4i5bwHfn9aikzVgNA
XMPDktYnqBFFMxxWodL56G2DJ0+/D+dh6S9RkoaOT9NBk5ZNV8ODMZ/FnTi33N6y
h+EKRT9QInHcVwTL9GbunCv1ECK/rVoBHvISbcXxniwgICcJVzu5G6Rn9Vwql4DY
e09pKe3qlHD5zbzpHUjsYT7qUV76kWIzecMa3vNgjtfRvL0KdEsqoN3AiFFfyPWA
q5P1b8s0+o670JC0XfgdUmVsrpdIzWc0bpqdUCkKmN4JbDJxYKUoq8Gob+PSi58Q
XsiyYa9soi7R/MaOdsOyZ4KxUOIvYnn89XxR7BuLmRGmtdMzdWMoraMiSU9ZXo8S
n6bL+I7t4XAryIM9XTqlIUi/0/VQWYWwjJmAWsV1FRJYGdQNHiMCaH5ORCfJfAMu
cs11LmD5iuO6nf30P8b8ul44Qg9grsWp3swNDVKTCDvSEhMkA/B0wfOs/SRehWvf
ewJCDPoMq8wGL87NMcSpKpewU1UDCpndryUXI0ytqnTh9r6ffOUVFxIviKSSO/W0
HZNeSzgJjXPXL2eoBF0XLdAgTlrhxOQJQ9Xa4V0NFzyyLFoEAqwo9HGz5M2Winbr
+lgQvyEr2CJBaEwbFRX3hIcNuwDNxjCyf7QcY93NoDUriU34n05V6DGMhPSuo+oX
7xpbrUMGLoD7ZPztm8vTwDQ1Htte0ybPQ8HNJhMaiG0lBJdkmdkpXNpNVZa+ZoE5
Ryd9UhbhX4hUnsjiHBHsteBDd4h9l5N8eJg0BbTo4bPvps1vynl7i2rojEDdxmtO
Sdq2tqq5sEatkPH63a4q1S8y3QQnGe7uzLT4kYMBVtKZKpKww3IjYhLfpu0Fsq49
nyxlLILJ4Qzzc7YvLVrf3mLEVVCnMZyGzeKlyHhN11/rc/5AjhgL800gbOkohQxL
YGDS6/GSCMg1ANw+jfVwE9Y5Zt2yEQIhkoThbFobEXS6/AvBLzBWliRj3/UWnqcY
NQvAcxgpJfScg0r7uTqjuRIAg5FrjNhWQxNnUvNErbzw/0WsEsSqlMjJxXJB3LTx
8vTJpBViFWlTyh9WQC2sN92kmPG4Afgnsoqb7Bz2CbDsRcs0UZ7Hlp2mirtfU8KK
kktfdfpEFtfdk/GTcbzoHPQWwqjldPxm2WWuX0WPXutO7c3XLCFT6D3Kl7E0Fbg0
9AvLfOiQ2jq9IBmZV5VP54xRyvt1H83KXPvET0fxPRknXj0JD3FKps1G8X+9giV3
apKA1xXh+SjS2pzYcUK8ufZONB6mTsGhm294nVw8wSTmT47odA0ZTkMgYdMec7pj
eTPh3VSuyPW7PS5hJTqqmvOqS5RYL780co926n90dZysoAR6iRypV/zW/qbRTG9G
zUnDIWNjl4L5+O5IfBJrmNCSB5t0TbDjAp2jgW8rwlj/5VyBMnqHUym2XCkzyXBr
4wbCCsdFU+uz4UmXnumCZdjSC3lummMaRtGAHTrlTFzANJ3AjAb6OSAeo9D6OieG
c9GohN9jKrdvZTN/XwYC8gc+R5cfybWZLwtX92tLT7YZCurXs1Bo6kAckMmSlbtS
s7/F3pjJHgahQN7PwJBzDlxdmCewgR6DMbosaP56pYV9PwMnplENM9QiLvd7rO7Y
eR1dqN1wJGAcZOarEIpZBN6MFR0m5dlABBDoVrtQeWKlzeRJZY5vzJ7Iza6skP79
xVrynydpfd8+lhI5IRTw6CNCPgP1g7jScWPbUGA34VA2MOBdEBMXTHRpdpHkB1Av
Irdqc6eyOuW1PQg1vKI/Q8CwVRXlq0cWri4SjOda9QARqhrICh+KNWXstl5LRfrJ
X6lIR5+7W16uPyruM22pCYVyNl7xBHNpqmGhR5Oye1taER2futNdVv4k5H3PWZWe
3aHpa93w8esSyPtppGPbC1a3+k00PUnf5PSN9+W1Sb4BodcV0ag9RXb8OLcZKsBk
Aqk9uWdqHYy4YRTpB0/bDB0jD8M6jI4lEAzoHu/DKSRWJEjbFcAz/K27rZpzFJHS
3D4+iaCKY1eIwDGkiOOXDi1zniVzgmGLGIhBRDOKkaMH3V413ZeFacJtmtLvTvGA
y+oYMgOQEDkQId6f46iA5K07SxyUBM4XPlma6P0+em/5CXt1oXRM+igOAB4LJfxv
HZPJXQ3WOz7JMKaovnEDwC32nGf5lcDN3SX96TBaMo7RbtyXisV0bFzigRV5uWIT
CMm6qJONiEjHROKiIuWNrjHojqJOQN+92wWUxFIACABkWpoBoWgq3yO6Mh39NTja
l6tf40iHUZX2FRFHixOGT/xHs6JF7bcucAI8HXh119D0d1P4r/ANtd48jnz8kogR
GAkhDsFvZ1yFGD14it3x2FhXK3O74ZsK4WGGjFxbrHJhQA6YfSle59zu62622Mde
J8h9INlyqntMY5jDXMfHgu+UAHFna0gL+6/tThw2LAgx2L+2lLpQlgTQFWi36JIa
kNnp6rh/TuMWjc27qV3yNX412lP/ZV2PAh4LAovbgbA/TNCddcvxyFSL+erw6aZ8
Aj4AABblceCd+f9HGZ+TK8CZXVHIs7HaC8jn6WB88GhNw2HydQZM3fptN4X11Kiy
ELE2w3vUS9c49DEvar3zMFiVhZWUrVY32QvMeut8ILF4Xiyj+qGIhkXyMKqymWXt
Q/uPX6gDGpN73BoVZ6iWfPuojuefiTleklcWD92Yq6F0tU1v5AIHdbcsx4bfHCzY
Y5uEpi8bKFceUJ9IDo+mn1V2Im8pmQ1IiarGkMupyZffQNiFkuuLpLNkyaOyEceU
LE0vs4WHekDQTWqkNJ/T5G6nk6xT4ipB460t7HtV33Ps6k16sdQZFts5JontXtjA
gkfBLSSm0ZLLpGmMVHIJsJegUQj3FRPB9O3MfbRHJblvdxubtuBEMZ2YKJdXS4RL
7A5AiMfM/OcX/Tf6+islMeQFpX6XuemZ+hQw54lUWPwpVVbCLR0uwve91BZdA+ek
NezqbJW0bE0USt7xDKrIv7lEfW6ZUp0Dg5IkE24ybHF20JEE8p5U9waJNN3FJTI0
IPXZkBRyTR0j5iWBAxQ82TJTF7Fgt1/zv2YqD3BdVJ7O6AzaTdEmt7SlNwYutM5B
i2K0/jf1b0YcxoGLoXNwxz6f5fv7Uag+nPS5itKaAuOreQb9h4140AN8OLH1uyBB
f0yo7UC3N9UJD2VEhW0zqOwI7CeGcSfDUuCzkBBQ+M5XugciVDmITjl0mvP88SDv
6aVGfKOCoXy5Jn6FQRbVKMSZd8ErNl7uyLE+fGu6JAdxJYyeBQhnCgM5YPGZ6fSK
iie+9l8qrG/YvXXFHFYxHEfNAIA9uF4eAOxp+AkHnjqmOta5qgPfdVDsfzEPXXg/
D9wYjH85IHkIXMTKYEJQopKITPRi9aUnu3wOhAz9Me8rZePzuAFf1FxNEemFeV+i
BkLffLH1if62h6kDmT4Mg/y7BZzdS0je2RuV+TDsmuvkeCe5mo75NkoMBV1XT4oN
JCuX7r05UeQmLX0nfXtQaeFMEKhZokyadM3AggFtJwoy8ORP8UkDNYLsCvIJfvc0
ct77ckK+wQlbppegmZnCco6br4npJ/mqjmLcU4mziR8eIYdz0MvUuJc2ylUH1nXc
+GdD2ddZCgmcWqqmkajCExm0PvK5CUB5o9Hnr5vKblanQ6DADI0ySzXzJSGqIVkX
NY7iJD/vWronxAxMvFkUEoDj30pJyt7KbpYV4Jf/1sMzk8mKc5H7cunCL9NuGjI5
RLDNtoBqapplNJJzT/2hhzYy9nHebKHZZo02BL4bhBJwcnhIeP+0oNaBSog+oZPZ
rYzC3Kmz6TOVYt+vZKEk7797g0mn3/g7jPVsTW6fdXOYK2fhheuS0FbQPHZ56XK5
+B37pCfs98o5sCZJluKjbsPTwuBTjBPvJt5WKf0knTuJTd166bE4kxtH8NQ+YPFk
+0R7e5+63h9Y5SK0VeX9TQJxsWxY9h4A+uXEWBoSkD7jrmDU/lN7osHGHXc+FZth
cryAWpP7uZLRjKuDrkDJ0djoO6CN9ltqGhjO8Ah2rPaChmZno+LaP5oifXeFMaT3
ay5r67Kp4NCTu13WmHZhBGNXfJqyUKBUCaw44DzgoPml+eRZUFtzFcbFKCoXsiiW
neSRqt1MZFAh+PRUiSfSm9e6aHrHg8nXOIsup4q3hnUesmRiVGzYODS5v3dtiGW8
BDd7I+TMk8Ioir/AJI6AqtUem71jbpaDNhND8j4DBlFBCoe4Vr4e50IMbaCbZaMq
2nveyCoim/nLdWlxVr9Nc3gBdFtOs1PHrpznZGQw3q/C9ctAiPEfB/sFD0ONoife
fRhdwqKlq0aEwVlu2CAwxsa1Zcap5jKZ4Yh5aVsXBQJQQT2YhX0L9wCR9sFcd0HH
3W85P9rebcWWQGq23KbvcDpr4RxEgbPrjqI4SiQzXhnepxVoSiEQHw8q0W6kwQ47
LxOZalpjB+aIyfoUbMtrt+jZVAa/0Eg3YrT9yjbW6K3gStIqNulE9wS1jJ6mrXJN
eQg2veU6FeK0JgvG77XBa4DQJpfdKZEPrtRG4E1IqKNa56RdWCGmHBUYQvSqzosp
jMKKdoMEqaszz+BQqX0dlpSMTqDRN2kjnD8fHnbyyA1x8bEIum5vo9Qii/U3C7qm
unwhpD1oWUDpt58T5xooPQa16BC28qSW5NGa9NgyQrdUhw/DB4Is2rNOMPtBVoBl
ieLIMYjm8ZIC58XD/oPxqBYFYtIbMaS1g1IumaMU2bRWXAWcxhLBgaXxv7uImNCc
y3KibI5iX6WpbuzauZLHRqKU6elkdvYE82cMHSWkeANUGEUSOzUwzuiGnOdwla0f
qzxGub8DsAUZmALUTTMusLmevj7oo6pTf8pXf1yHeTT7tbSCEPbw9zDqnJoCIE37
d4Smah18w3EzoxJZ989rUQ4qRKBrpvyph8/mGyDFw+p53564PuCvwDTAcOT3Qtbl
th6vX7lsjofVcXNDTh2m5S3smEvE0yF+LpFD475O1SqncntSjVGEBgeuLuX3gSf4
HIWPXf+2WfAoqK7ioDGCuULW8sKEjr9PthTo35k90XQX9Q78vl+rOU6S2G5uIA2r
E7krDvY0u3tQy7ffy3p9Zeqe056fNqteLeYEnb6ri2fGTbMK2ndL2E1rNcad9XcJ
OykTQ3UObr0uQpFv1be26j/N3uYQiW4MoeG+Y9g/aXWhOc7fKuaFr9k8O2Cz1rQo
Fbguc+gnhZtyRe4mperK9hB7DuS3LglQO2V/PyHwgZbp/QOwpyM7c+EUf9TyZt0M
YS1o7qqlyRZFxKSXXkQNcsbgOHhu9VurWFT9eO9+VOuSuBmSmMVpAOT2W706YM9p
ehX3E9iETWHlsOFp2zAqQYz3Rmm1CFZMMao878S48fcdf2ME+ZgnUTnqiJlzFr7a
qn1qMtxkKpfM5Am3uKxc6bAnaXrujd7RW6KG6iuLUD9c0QpU9+LxwHTvjMpm/b3Z
K0k3Uw+noRl+/swzCyO7OxuOyIqfCn/A01WKAA1iOirm2H7uS8nzDiQpatNeD6xW
IUWkypX+KfZnIMFI+jo1zD09xvUl+zS4FqWcw9MRi6gnSAYIBfj47RtaziIS66W7
743Sit5sB9EPBKzngwLeHzpE2zARvGXponotvzez/JS25GgSxYeXseEZTEsSond+
MWo5lDc2KpX4FmOW4ZciL3s23Opehv2ZFRjbXmLGDRr7U89nW7/ULWV6LKptN8la
lGvz2qXdXqk79oFQWal57CkcxVqsflcibnuxoEftIgJetHrfOdHZ9ykHuur0ZvvF
aDqIAgwI0oI1JnmleAibuhhASJySwghd+py7dy94ZmOTzEbqbaisbUIcgM0Pm496
j3vJ1nvAtUIP5I3DWVy4dTM+05Doz8E7n3Q2pz2szOGc+r0hXZcbstSNSiDTDia7
HlhjkO1WCRQpO0leZ9WjS4oU78e9Kk5rQB6/Jaz3kaP+iFNPDS2VkvjjQ5bapkFw
9fBYBvFlOOpZyP8hHWMgu2nmO/iJqu7QTX4c7GjebaBrQdsHRFX5hdIVAjbJdbS7
48QkOmTUOd/DqsXJoAOId2nTItOadGH4/1EbI3V3n5b1xD6DvIKSOQsJ5KSpQSB7
6/FnOElwJuGh5LZlitBTFSuW2zI6THxhSSd2FNptOjMWdoyd2ko5CcgDtBUTMcVG
TqbTZuJtTfXNoZNp0ogALFMYnqQDc34f6DXwPEML4BDyq3valWx3X7Z4A+wqyPvH
gz+NwD2lVR9IBfY6t2fnJaOsQnSpil/2qWYFXPUmaJRULMu2x1MrEN4MmZaNCckF
vYYCkpXZ6BpH3UjxYYTBgCMJXWJBl9+g1SgdUeDVGzSssKOAcW9YgWJJlt95Jn1i
JE1HwrMcwLDo9wVOJA0vg9QQvkLSVVg/liLBXhDdCuTxB6zEJ4vJMQ2UbKXPQiDZ
DsqB+4IKIwhu+yiiJtVztD5j1fa/eg91yEl/0oIFAeL6ZVISyzRDi7PfJTg7PESf
1igRHhjDaVWEqruArokI0R56jVh9RPYyZchcA9H0MOR+2vPqe24yBGevIByvDaBD
X/HqFyiB6bFwZvldllJjuujVgLzpKaqR+g8mYIeamLhauexe4M0iiSDKXjC+L6ZF
X+/JnfjxCatb3zG0LTFpU52JJxojSlY/5QJvzpIa1xUWgAHX0GhRRXLsOe3+yt+I
e90FJ7WLr8laklYW6otm/VcjhK/rt5R5ZLJsBfthay8NwIlf2OSt9URSPaBTVWw/
7ODP6RTRZbuFcAv/SuqTjGS6MUmPGAZLVev1ugSiTyBNIMt0CmdLh9bC5N1AnLtU
MiM4ZlmyO0NCVAGbID4LyHXbZU9ZABFaEu6WHCEgaWwUpwOd9suFYfJyhBWVoe0N
TgmlCUW8GUSVoZG1MknO1vxGdpxOGkrz1RGZXEp5BVfQme0AGjOvyeaS0tJwfo9s
O8kgvNrKQ0N47XhpIPUBacqfZ4fMUyqwlSq38PdEXXhHWVJN3VOKvujrfWVR2wdU
GYZe+KKYeUsLHc4gGmN2tw6wGMVSmoeqca5owYlgXfagk2tvIFgjsEq0l4LF62DN
BpjASlPA6AcsgomTjHAUzEbY3M/lmMgG9FDlOq/pT6UaHlwUOIquYmwiYMnDQyqd
kphzFGa7EEvT0yjKBkdUP3LzzmVqcrKpzvJjHXPhu9lg2AIGWsXRhmuIL6nPV3X3
ZO8eBOVka9Q2dxuQYFFoczvSe0L8uCFqVOb4uQPQKUTiHCj8zRD9A7BOJscRuCvw
n+qx0g4Izub3B8WdZzO9ZiOL8B4vVgWVeovUf72BcT4ujgoOOxXBVLvO+QkIhATE
9iqsPWO90MGOgXUl8A983wImWm6kiLxo4ShdYMgusNLZsXeE+csJaHEYLI5ZGsBD
`pragma protect end_protected
