// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
sQjla0qHTMtw79X7W2Fn7rQgkFO8L/tclnClJjtFJW8nW6oLrIvH9LrAwzVC3GwG
0pShtWaG9azXPbHNH5h2L4NiOo0S/8J96vBuwj8K7PtI0YjYiwohW2oU8Oaa31F2
e0N6IcHozL+IxnjJnKJ+ErjY18G7k9GZY1/V2FL6mPc=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13968)
aHrEvbhlmeTV+1h1CxpTEliY0BwUEADO7mg8PIyrSNsLG8teSLZHOpwGil/0Ochb
NCvvGRrxrS+Av9jngJaVNpCpN7PWbf0rn2k8iZhmYvNXY2KDOwqjolhTwQvUpiYb
VD4U8sUATRC+AdnHadR145LDkU3ClqwzIkNKoQamEbwu55BG7CDzvq4qpVOmnth/
L4+OIgj0r7Gf6+mcSQo9Rb2Kfyjup4UeZZkZXlVxFJGdACDx/LoN5DH+dDqdlK+D
58gV8sLMiaRVZoezoGsjxv+Z6GQ3jF1aDdyWKMVO+liE6IIFkyOhBC9r3GO9QXal
b6vjULDpMAGuhYA/MBc+w/Uh52JMdtMQvXxYA2NxHWYpxx9s7lmq31xy7kWqvbf2
Tuq85uJTyDFdY66KAU0E09r34gRhFV/eYK+FOA2gHwczAZmIzYlrv7FwOvmKnuGY
c0XGobTIybTC53HOCo1qAbtRG8cTObSOFhj1idH3IxYNQDNUH0kzC5hqlSOn6syU
qjrs9i3TbpMYpTgzbu7j4VIPzuwbr/p871EUbsBa1cNH/cS9kEN1zM8NZxpXEhmZ
6nnzqO8rXm5g0PR+k7ZAcESpQOGGcdhrrHambuh2LtqKyI/r+LRWKwdAfeD09Dwi
L2v0eYnGZH+CTBtVgrnrlWZiikmtoTceslqyk/X4PD6ir9GKKzDOEoAF76MFHBxT
qY2r2iJs4JLJ3hkIjkmpOkRGeQYshbKFy3+g5K2T6ga7I1ztvK4DbmyerQfLti9l
zVaUgI2s0Wx5ZsunKEUgaSsbi2T+xmuruxQttSSWCjn/u6vOxbU1+eX5FBTP/Mmf
MoWLhoivfZkQBFw5aHGd55PjX/r4fzhb+6WxOJC1/RqGDs8Eeenr/vm5aP2uTHc+
CPwwiDkpcsf9R1a2KR7I5ZeOFqciCC+tIDXx3aXD0uZJVHwy1Fk/xq1fUUyZojQq
KUb0w58i3vocpaakbP0L0jBHJJ/699Uay2StRp7bBzEEcaDgYzkHdWi05pBFRFJ7
wRotdwjpB02xJIK4LwZ6FMlzeZbtQy2HIjZXevnlVipQSM0rMI9k24GaDt7Th1SU
1oQ2u1akxdJSJ6P0ye+68vfnr2EIdDsS/U7n4l+ZcCT5BdC56xSgUf+dmDNQBO1q
LdYrWjJq3rCAKyefsOa7kv0IdqAaG9V5LMJz97Yc2q1lOkp3mlf06ox8elE95sFS
Rh+Wjt4AI5Y+cP8paasyj3C/D7XYjRLnB6F/TgWTq+QA2GXMFAQPD8VVZfJlOFuP
N3Poj6tleVobw/MX5/XkWgQaYeaj6seR5eciSGp1x6l/7mClFP6RHbqJxFIcvd52
oK6JR/chB4R8JFTiA8HwbZY5t7pPCShR8NX+h+I7kQklyn9D4p46K4RvLseZD+An
ueON2VFUm3NFsh5+nqKYhr9+Wzgi7ns2wnkJt0OkueSB0DGVR7Mn8AGAhRS+EBkc
WxbLZWAsCAk/IXg48BYpIxrDjN/N2IZtfU9y5yyUc8TeoCG8QCANAs9NjTQE4wxw
b6oe8yst7C4qlWFibBI3HVKZj7VCxfcpsBanUPD9mrn4Yz7XUfxZ5IyAxIJ178Kg
Q7XzH5FQ5+uD7M+WgMxrfVw1emR5JufR5sUo8KnLl6umGCbNwk2OYFSrpE0mSaPR
Sp2zTNg0069ArggFT2rKnMxCRRE625/MTPW7oAuD3RibuVdpxmG4md9qc5NwrxpN
zJJz9dTV4ZCt7Zdv8/byHKNIn6ElVx3bGIJI7tvoVhFxhgPB8UlzkRhlF4wurKUm
6i/f2Uh+bR2jkBAYmihv1+0wBLcQw8xnsFHHrBdZmEtAn6JSQkYQBWnMl9Lo0XVB
bYQwCzFD7A8m9hWebTvgB+jipMm9AB2sshF+M5r+Rv61Zw6EJyyW+5G/XBqJcpzZ
G9BmJ0OUH3jQhyAwV+ET96j6ZhWIbOPdZlptZp3Xsrl0I0hywQiVZiX1gHBj/t0c
E5DmR4RQVgXT8Ure1IVfN8HU4QL20nzu9ClFvhCuUSaMZqWqM32Q+jM4uPlJPKG0
8pTrjPn9SSSo66f5DcfgiROXVSSbgYtAAcwA8CLdnl8hSaRo2EhAMpSA/k345iP2
CGEG911JjewP+B7+pA9PJds0fgt+nPU47VbBCEJO7whJ8boNpIxY0awUL5BR4buX
CSx4ARpnfgpGSp750VMJuWFoWRLWP3DNmb61wF6Y+JSAbv3TlFsDATvBnA84J+Oy
jgUSY28XZYPkeaVLuHrEzKcK3G9bpeJQNYjgmN6XoabTCi7UoKq94wi1EIiAnTKo
aZsB2/e4PLYdCqYmFXLp7Vez9e0HtEijPsNd1ECopxsviPlJyerPdaZuSMyBLj/x
nwyD3O8mp/dq1nE49aMXW76vRcY4T4+GlOLJYe8shYxmAKQZEyNgK1wI/DG/0PLT
Fgw8aicFvwjPKibquQloNTTt03O6RlZXMYlZS97nefItUUwB8ge26BCD174rM6H9
1TAywHGncSuhdDfuku5TCquCJwG4eWxR6tk1pTERwRnbatQIDJ6pRNcXTSv2xl4V
biG+y2K1zKdMD1/+nojW59XvtB23o8OZPwkQGoGjHMWaL/ec2TrLcyMn+Yidg30O
L7U9w1A6lmVL4BBPiWWVv+ZdAv6bVHlSdsuwdmp4OLMZpwGYD0e0FQ0RkuW6offq
pKqdjzoaBu6srH7THZSdD+5hqIQSQym6PQZSq2WTh4Gy4IQ+iBsrVbdMMnogIEy5
h0bpgLwWwm8HdEermpL7sXkomHppbJn4unXdFfuRp1gjO6CWRJm6p2Uh8OHbrPLe
SDUQrTK0fV5S2BPrjczJm93nvLHi7BdkVsUtr3g52TNwMpgErKZ/Q+n/yLpLGO3O
Ark0HWPC1RLqITZmVlbQzLaXhtFn7F5YPUVqRUX2greGD7WeU5M/LE4IfwKZ1nsN
cORLK17ztRVwDXvMr4dLmiboorc0vLMQeS6HdZs5xbgtlc94KcuSIpdUzaZbjIuL
h3+rZOs3PYKdKVwAOa1thg2Kpntq9C0diDbeSCljCj01sGlVEiOJO9WQRDt4zRNR
x3bKYKhmya08ht6wuJqR5Y3EXcM+8Piv63US+aQmKmS1/EWGxq3uc9oruPti2831
zzfF1RFo8hUpmWTKfwQQ0BDgZQgtxAuSnIU/OqjxsE5IxyUIAoX+TxusP4eXxnma
z1d3g69wgyIVv+m1yNjlA3HvQTB6vszrbvX6IiYcK+YOkw4N+0MWY3GuMcISuHfz
uOWz04sLushQE812ovx2s//D26eoGRX6u/ooR+G/8IlGxT1SoyOfe4I+0VuiyNN7
Xmkv7mAagRC+Zs0JJepld0jT03LzpEpAHyWBXnaVUlXJBA2eGtMef/TSfT4K5yq6
/yY1NuGrAupD1am7BfRRzSVOoRsLuWF+gJhOXCw0sR31ezgvvYNt0P/gJoYTkGIh
Idvo6cu8ecWusj400Wrjq8mrW+IZG1e1yEzynWHf2MPhqjffX8GU+nkdrGhEQdlF
UA1M+olcw3ilOZQz+ibMyxLPaHm+IOSa615BS4WhFRt5SxB6TNUCmSbjbT5DI598
1jqCsr4EoH90jLowoYcV3hfb1wkoXHRC1bNVkE/OfTbHeAIdPvkVm7GuF/zjfICe
UhVIPYj0GBwfVvu2oy0Y5a1rBFJhwkg3b/HbEg0WG5YX1b2cZfOkm/5F7JuouQ7y
rGSZNMfaUovXFpCJ+87dViWxj6mNco05uNNrHlUohCzFw72iFSaFTlHMsTTLo1Pi
FSFqzbDZzzHXKmfu2ekjBqygaRkakC8HeqZfxsmr5F93yXNunNRbg1h3c7GJS/+4
M9ta5kW6hrxxJGrJLAtZJfH38zsGCifoLINA2kWtEXspwb25MLYLnwgj6XhMch4e
Ut+0lAj6uxtHheZdzG5XLEzNhVjuEny3aK6MBTB7S887DKHUMxqLQaWWQwz9SBLo
ioA5dhD6BNNAg7/SE37rIWYLfC2hQTVPvjXtEafBG7MX01whV6PWE85PRdPoT+H5
C3d2Wfj07Fcp1Erx3TDq+AyttGWBMlwS3TL79DpwdRflf5J8AQuHF+WFgkS0LwhC
ywPj8mfAnvX0DTwu2ldT3N5h7LSV3x90DjpsVUWNsI6UaHhDc9pEmnW8qNhaqWkW
X/ksZRcjUH48TH2kNLszjWTe1NvRBzGJfwa6KEPq2ahFVSggdJgsSnIBylRTrFtO
amOzLJOkWF0yoKQHB0EOEklMMeYA22thO0nZr4n3UpShEj4bnk6GPTIgchXfjjYR
zHTmdz07s0kfkUOBYhDsyxNjIjO8eikkeb3Uu781CqjBYhRNfdx4sf6NP5FIDfWC
lbSFyi0GqyhGB4psTmXHNgvDqj7NFJf4v1niXr2ZCg7uESrMfyen5y3p60H+kLyg
iUqGDVPFRviuGydvaydeXKlLXJAZMh1c63aTgO60f8rmMd/baMqRd4qJrWk4M22I
t45s/uZH/fFx23MA2sK31ldNzX+RzeLA89YUaf5gFH4MjezSrHlYzmTlLzw5zGyu
xDGBTM5lG0P6+w39fidt5kAUMVv2OsS8ZPI38EhKDDxOK5BuuaJCxgWV/mbrRb3j
Agw4o9OE1OoBHk0zQv9NoyG0xGneHtahqE/ZzvOEQNYEEuso6MilBrecrObXDmuj
ApUDVWSde5Gzocu/uXyk+6vQkeR19OrCyjefN7ve5Q5Vw4dNAB+jCmkTys4aq6m2
RoxTRnjZpdGGSibGHVxo89x0Q5CdYbrMhgs8Arwe+6980fy29bRvvAKAp48nCSKC
o+jOumVQF8FrBt+R6iladozH4soQZ8ET5yadmnYJoACW8LwNjVYUSoYggJKXUwWK
INEeMwNU1KRPP8z69jkBFF1+Gaaf78aNP+PHQbbBfUGKZuqeo6K/fCZ9qe7zzc5W
VtoSw1WgL/cDaHwqo+L8EzykTw59YqEzQDuwHierGpXqwotNmGJwg6L9t+IpGjbv
V+vYjSMfhwJq5l48ELCFE9rEMdsO4NQbYT6e+9wTaSjlpY9Ka1+4m9ffn50QUThL
keqkkB2lA5akKAl4GETUMnmK1IlKapPQGm6I4lLRR1EEEHSai9ngRbdxT2cq+Ma2
zP7kYcMe5XXI3ZpwMEajsG8H2PTfTOG6HEkW4DoeYI9kw7PI1pI8uD32B2kE6+7P
XrRcCvDt9HQgJrou0EbuRi5JOm20Fq0xV1S47obi4GWAg7Zs0qECfi4T/M4z27hy
lEu3YM+SBz3zVhtszitgacLUDX2c7k9OnXmA5ZNBfKWJz8I2xPOHN0OKkEKZyhv7
uUT5LBtm3uODUYlE4Yp8RRfKOsSwF0GSxBHPwOWZFaU99BkOZiYWsQWsXDIsB4JL
2/VLWW3PCJBk1P/SdJ+c94Zry4t+y80QniTkN2yMDp4IoIurnym6rgA/miDZnghe
XZxeBHZ45lkbbakZqi0RW7SvckupHg1WIWlF/G0mkQKX0GL765lEvQfg/L/zknac
fwukFhe9AyRrn0GXi/RcM9BBqcGrBWIe5qdhxnZO5jlWFi9+XaTXtjUBvHTRI/bJ
Sz7z8spI9dFB4i2IcPRHjqxj/9EWDAssTge6a2QJlV91QfP+qmpSlKUZwxVMYNJj
pJ8KR9u5ir9nMtR0kJUDLowh30j6JM5xWDuuI+/L+3Fe5PnaOsFBTwp0ySpxqfiE
Rls5hy3bm6AKBhH5bgl6OhPJzWc0V2B0V1IkuGHJyPulFw+lGZexRAza+5l+QLZE
bBYPUlB4qxhyuwCkJugBkhCZIOreDkJPPRY95afi4LXR+rjigfKoVT5uFt9XBl2K
J7ubJ82GpNMIKgnk2uB5i9dBlTYN22GnZPJybL3yFH/YENLsBZfYc6cfoI+ahaDR
SPR+PtgFF/ZPUFPg4ZBLQM5Qh6BD5X6dyym/CY4LXOmMeGR5frbPyBwCw/7BgqD7
o3C6S4VPK0oGCHOLgcvqJaRNEf/NkhjaAU8fr0cIy1e2klYypHOQZEynRhCoE+tf
a3FTzIR+DBBfeuEd5Qpo5iyTWSzKgRN7j3t41e2tv/QvN9AaCbnjyu5gUJzjKQsw
hdb/biQfLICjN6hgF77Mua7RR8h+8lm/PWExJ81C/R8KAH2rvuG3F97L8MetPy38
WLGCLwbavDo+89UqQYk6CBcRB0tWA6ZviUG1FQ5N4i6Y2HgmN0CHEWOm2MWMOcsx
16YEifeLnc/AnPQM8C+O7nC4oBYbtRnXeHADiSVJOGntFLz1k2DoOSh/QHnfGOLs
win1z+R75M+C/svH8svqS1e3Iqp9VpPc55fy4AiAvHRbopc1/D0Fvs+5dGx5oAOh
jlpZCYr9heJ+1p1x2qP8Up9ueu+rfsnbz9cNsLA6TD1IlkItKxgT+AV3makNaCts
aYfy3ngGte1cmHQRY7RKTqUHbCuCRwRU0R/Mio3QlHLmwG4uerx7nwyMbtGMaNwS
KZgOi3zj2LCZiG/ZySNCae6HHjBC3tIai/VYMieFHJpOveMrgppDVlf7NBwbJN51
iG+NAJsff3orAdxmVwPA9xaiTPrxLGgT7SuM206ywBDcy7FGamZklDj6YzZPFAOp
aMRJvP2stR/Uwd+rViSJ2Uti02qbIzwGI0qnK4TCNpxGBBEmILjiJN8pJpJWBoOM
p4R5q46WAqDtTLrZiB1/8zLY7hNi3DT0lY9wfyHjVG7MvL3nfvGSVlH7Vn3zzNVR
p3OaEETxqiG9uRm8e/ZGnn8XX7Sla8AAwDvj6cmGkOJ1l8OVLUoMckfhXULixMVX
sfmyO97fprVYt7K/ofyrwqZAN1zoZbHtGfEX6lIvfuM2KiLFAVTlHoGunUsVAygP
auEMgBiVw1FNY4Ln51SwXOCehuIGLdGhvQQEEu/3xmvNrjfIieHeuYLiazhGbL9v
IljM+jaTs+ugn0dWZYzv5DbGtfG0E5mM8qFoSD3CoOczPIafu/wJ/0i66CJ8w62o
IuXyM3WsYmp0e7buQahqUmo45aFWZ2rHg3QZ+xZPU0v5SBp93OX7kxp7oZ+g131V
cNot63puD+z/IdDz83JFfm+8K/r12omeRzgrIFso5JNzDGYlRXqgqglX9sMbenFz
Za0izF/7wg+8duJXwRc7XOZA086xKzFOSS+dY2mYqHamtCfGfOOZXLrz1tnMub/2
q8gVb7Hsv2Gp1oth5SPJlTp2zIkJHfyO/tTJJnpzLs1UCEBeIiJri3ISgJOgC5Zw
9ODG9W0tsMOTWPCWV4cjRSLZgDcZ41vUkZY2xW3WFdLqPp9i8p+DgfXdw/oMQlYa
xzJQAXzpjqw7grJZm9AQy/ZmO/Cg72DI6CGW7JAlQB7eeR588yb9PuY4AGyes2IP
dizzhrkbsrAITl5/ysfK7STcLU25J1hxxzgd6wK4Fs2LGDgC2LNpd7TZwi2JS7BE
hCevOT9AQJ1h0ec73BXS2K0QvYFjhwOyR79q8/9pomcfU0mxrdD6t1b/Eht7WWJF
Iv3WM6em4PD80iG9eYZyUQiv8gsCELd2pgsJuTZ+EWqTduSXttmivipsFEPYo3su
SV3eSMOd9LLU9yxDO6ygBVS/t0kqR60+T3Y4crxRdmwlHJWnvHf3eiIxOEDRzJVv
hNf0MDE273QLoaNkD/75fE/u1XYla0cq1NX/y4qJP0aNvpOznHO0pEduo6plG79K
wfwip8VGKiUiSPLnR813VxYwJgNwH9DJ7itGoPTY+rNnlpyPztUp91VYYejbhY2q
2UJ+imqPgKTTZuh1XR1wFqb4rl7+RAEmTDBbpRxMFbfGMAFh2oJpBaRPHb9NaP+C
mkH2PLse9DYsA1R4kzOW+wAqgWsA9KBo+MSpYqzmgZHhGruBhCr5swiGJdXUXGFY
YAhFHMVsJvZqKjTYyCEc5NvG07eHa+sQMQw1YEYsGk16loOA152+L2Pb5TuiRo9f
lz1rR1qga3MC5wPcMdmgT5jOsIpeV/nRFN9DGYvWeCP/Z0zMGHKBzesL3aTkbB5v
DwrWf7jZVWVtiiC7qzCpZITvJdQGoVGptAP0iJSqXq+PGKaCxQcmBGc2ot1Ytfzd
i2qo7+iwVCy3mbq1pMc0sdbgi/lPlo5tO4tugEjckMx3sOmABbXAuOEZ7dNOmJUM
H8AVthjs7Kl+4ahJr7ics8x0hlnMlgMb+GjSxXd6RG6ZtkDgWJFKn1/5ulTukY9m
1RNurulli2skqxQeXDDgNNI5LoQaF5r8CEnz55xuTVJzyXyZOOmonjl96BBnEQ+h
ZEezJ9QnLB+pEyCszBvi4wc9HC8Lw0T8cv4thvYNtfMq0DlzPbTQ+QD4p5UNFNqx
p3ZKpARe8tGm13gPZiK5l5cIcSNDypABspkIoqMeXAikol8W5sBxFGi1wnlG9Sfa
WuYhRUy5vnFjjVx+6YP4IW4xYkQ8OL/KVPOcA/FyDoLVQnHQdG26/d+3ZNPSaako
w4UBO3rb6l2GZrV02JxYUf8wmVlvmXme+QfVGxuxqrVgg3WKFsZYfWO9D+5YDuug
gd7qndlJJxJjk9nqg427haZud3YMSgitXtFP1fGdV7ZDyKU9ySWVH6KpPJ+7UNO6
G/JZjy2MMRRY7Wmme3Va82H91lK+mbNTujPIpzQF31Ug05MNyrlS2OQtgpRV4J+w
PzVACWloYOE5vvfukbpiu7RCC6rs7f4nUJJUXrExgOeuqBgK4kvxufWdEzYphrWx
I4SNXzm0+kp7yaKZvnqsKee6nhCnmvtI3shWAy0vXR7S81ejHcztQAje+VrpVSAt
Yd25DaCmNn5a7DPQsaJ6AqgNeTKRxe0nHzY0uQ95V0eXWBEcxnjW77boIEQgF9jr
gpHFeWL7d4UuBF3gyvFiubpZ70E56Hke+bgAxqaHbPpyzDI7txrZu0bR4usNG2WY
rJSddLvYeQyhLeLLfnK6D2Ckzg6gfdsNx+v2+o6MfU0aYzsjohQom5y3lWzTU7qp
k+ETOHq0GL5FSOt6jfX7l1f3SnN+TIMjNmgJ9J4v2jeu5EYttKpo6eQPioTxEnRf
2itsNivJz/A12f/HQ862LMaLS0Hdj+viPO3VRKFApdrh2dhOmWSwFRQPjXfjGHia
02WTT9PCCSUGIkM9HsT74S26qETeMsQaU5kUq+aL09nR/9ucti+Hd8OSCf5YdpJu
RMFaN0076Mt2haIYaYXrXlvidg91/TO7ysGhzsz7y327jZ904lEZzXVyOaiIu1XC
B7TJrs8MdVFJmWVRfUqXJsdh2QgbCkvF4VqztzmRbGsW+zJCZG1pFUGLz6kPDMvc
NcEPzVwitszwxQdQvzfdr1yMTzNb0HIjD1nEWdQxRoCtzTFUDpob9WL+zP5DPXeJ
qAmQlVt7xwne5P1yK+NnI+707v+a5n9rZwYaQsSecH2Xx7r4mDn3meriM8osYHQI
R6g+ZVHNr6YYrtNtrIwDOCo9ewsYoDbQU5CSnTPYo2KfIQcgEkQ7fekmB10rm8fe
KHmy3sMKdDGKnmTRNTxxttV0uRzamctxoBRdhUripMw8iByQ9ioM7SUzZGttyUyz
3B6N09xsOHX3iMIL4W1tRvKGc+QX2EuvebOMFXvgqJtIRu7VfxpiyYBhXZ0Finw+
fCGFKj+RCIWdF6ACAeCGfMp8LvKJ1fBDPviD2xh2zBbS87WGXedx6IFTgbWjLiRO
C9PRkebpmmK5TVOmXViSJ21Ejq2Zd+v+r0cUzZ30g1i2sBWtmAU3eXdvdi7su4yk
tKeVBmEkT8xPpDkKYFsBJ8C55yGBjn2vF9UpM6fHO7a66+djpABwccoOxITDe3Fo
rRjy3MwBeB/W3tGkOhg/O4O16mp2pgAUgZfenepZso6795Rvf12WwOzNhBsoSdAZ
tkl4dAmFNvwMLRpSieZoGuSuL00c16xvTtcWazz8OGsL+K5ial2DaNNPb232m+dH
cFReKgibf8piDLs1QKUbndPjqcbUhyxxdF7PQM+kFxiKmIBkChv1qNZhq26O8F9X
jyG0DE7tAUaXN6kXkQVEePTSfdQOQZYwedsNf470zwceR1fz5Y+W29PxdI/3lcMP
a2sQHnlwGjGNSMWZLsojP0xEEdf7fJ7kVfxlIY9/wS5CXVl+3lClxapKIYFYGR8c
tT4nQce9W8JnCRGpIlsM0aLsZ2UjjxsuX+i3+fWjti9+/64LlPBQ+l96SJoL/Fni
o4v/FnO2FKDZ+f+QpJg+Vqr0izhSvmkablxwLJkDFG5aH7efXvPVo61suAHU3ur9
Oy6aCRl4NQHx7XOagMmy+t2KqulyxfVmjASxbNhOOe7R+Eo5i3r1Xu3maToFoIuh
X/ZK3e8XM2yLX7WjvxHnpBoD4a6BLVFQ8OHoGOWPrxKGtWejaaOE6T676JBaOEL1
HGOuS9OSt7hg4Etbp6SxvomAt4Lq2A78AMuVfp8el7jpc58p9y7aOhlytlq9r1Y1
LlbY6TrfPjRvOS2umJxpq/Gv3rZBF9QGuSAU0nkQcNDbtG0lIih6645GkR0P/2gY
61pq4r+qwGo4CAOOP+il0rW+1sL3dBSqUA7HRcw17nhEBj9Gzl40pLAKpjxKMfi+
xexyhvNdJoAPTNBnQ/vENddOmUyJhLv+D4LS3X12TaFk3XN1pxq6Np2Qhej1DN/z
2ESAPDuD3rLiY6vUdkuHjKgYtucuk9hUnFhIlWfeHfstzxy8rl0sL7hVyAP8AJkI
CCAf6uZZGv+zNex5/Jb8k0xJ/fWH1DNf8XdnN0J4N6Tszas8n2wKoG+GtPPTBDGt
teDEiBnCVOkT+8uoyoqYgb/D+TR2sjQUspHS/UmKBLyukcoXinKp6JAlRYcPYWwd
WWdD1mkKXS2gQ/lsAtoy4Rc2YFC8mvIMcELq/SaQfIB2eR4I8tn5PqF2IstNeTS1
0WhucRBjBaUamW0kC+scwIbwNTnRxV3D1ZRUBNp/GmsAFzH2W69T+R3AtVXlxP+3
X6/E28qcFwn8XH69yg54dFYVc5QrWDy+aRLNQebis3he4Mx4E1loxYXskeGh11QT
7HSlIlUw2eNDpsUpS+71luEKGUiTLwCA3kMeqZ5CUwtZgAgk6pHwNg2HYyRONfck
MSsieuga9jBJu9zo7uzTHKqjzqb5RTitxUs40rBtBSDmajV3wBRKQ9xgDnHXZ8vT
yNt0uceYezA6+h5hyDvf/q7h2fz3J21NSGG/xTgcRixGDw4Y2GMfrgRILtTnEfcO
P2BzCS7nE/jNSmhCDjHbKaIDGUY0xrBd4FwkvHvLth4JDyGyUlb7OwEc36/drRJA
qZIeuWl+Q00pOGkTzHvDzGJCK+YdNzHZuYjcF/uNgz8LEs2NLasBn8Z+JDS74cfv
3vsKlWSet500wQeGO7ynwzsllgcfKQbYCWcnjlYfvDjfSqi7aOdOdztyKru/4LU1
tM+q0jUbmX9X/c5Op+ulrJNzqjfbALFQg1pJnzxrpj1us6+uSepYqK8Jdp9G6Iji
qiVfdql8aNfNKgKlYAINhA3UmOBSFVtNTtz9XxhPC3FEGb1tUIFTa/VisTDz/WRi
WY9rWjzJdrCzFwiQKKEMsJQJRLe2svM3sItmHZo6w7Bk1bnsRQvV0YKSP6fYH2fC
8K9Ua1hC7y9eEQt48+LvNbc0yIP9v6aJAU7mMrTezb2cbxH4Q+Mut6tDmXJNkQxn
ZBIN5JF8vBXX5GSDb4ylJrPD5HZrejEyPWzd4O0RaEiWZF8NQbTELZptelLadSMw
CJ3XxjPDYje5h93Qjq9MTBqN+mBp79s24Lm+pflkJ+Bq5DnSCTJWLxp3y3V+G5DN
fJnWRnE813vzMZW3QVkM4jJhbm9yTaFBr2csEM2qz914vfOCIhNe9BGs5W+FzR22
1feeSQJzljIhMkTZJ9uttsRGa08F/jFjK79sOhw212uJCcw0FmVPe3/IELnTs0M9
hNpDqsD2y1Zy5tUGifbNKoCQwEfajl7KyLgCUF+IyrwdwNbGxaWaql++1kh4mvkY
a/n2dDOyYj4jJlonXK/5Lq/LUOVc+da/Spti+HzWEklFDeKzw26L+avvYy5jNWwd
TBMss/6whqQVdpSme+XRaOKSzS09jnmEpWgF2+B7jyxCGkkMtR57IAqc/1mxoYKX
QtpD7DHPaXDjkfIS3rCCKTLkgP3VdyFcifKezRpNQv5nOR2c/qwDgncNT+nFUXkR
EdtmkoF0r6MaR7ko2nzawz7kCwD552BZjqpkNN2aZeeSOJrUW3DKEucbKQVP8Usw
71msmesizHnPgq/JKv2DbHwwCchJF9HlBwq/jBdazvFLp+9FOMQGAjSrx+UHJR/v
u9afaP2Gh2wGH69MCi7RYF/zHf+ii8V0EaB3vzydKYBCeexsHdsPUvudNtFC5P+S
ZneqsvlcPuI4HJ3qgfNTOgh+iOSkS9Hnt9PpOFjxvsgENmSNGIFxvLu2TJ7HAIgn
Nj4say3Zr0SMS16DsKPGbfO297qoVJlQV2bNGlA/VsBIfLrQPgIWQltx0+ADeEQt
yy4BY6Htv7IRZ/KRY4bRcTA/9HMFHbIF9Ebh6C2GJNxlY8TBhRyOc4qYYAhFCXrb
0c2gfZYrc0Z7KZ+mqXVT8a7IImHRGLFl2HKfhyqw7S8JkpPO71mPue/q8RVxHAo1
4YzsfDi8rPfeBJN2sI/i5Zpmgs0IsPqgVADhW7mFbDJzmt8/JINQsz8N0IiMND76
7lXcN5+B5905jj/OjdL6FhU+xMk7sSofNzWShSSb1bjuXuLicRjLw5ltx0IX2kH1
7Ky3YbHzlEldp7FanJFtWLMAEG+NBlQHG96e6oXZtljhADCkvJY3bNwqi13aISva
Gr0G4AyTkvIRFhp4m/vdnvX6ThHHMUzTiNDRvnM3jRXXQA+I2jt7ZRGgxj8qAhy4
9XOXQhNU083l0CCi2P+U/oaMIJqlSH4hpSf0h3airyOp8tr0RERbO3Zo8BuGfVKt
rztpa+clxRtRQ45iI9lY1u7KGFDN/OriPml/vzLr60OTL/RsJvLmIbcTr25J1iuJ
tegweNhiJMjWrq8DyWoddca36WOjh/KeYICx/8/ubhHrM5jk3pJp3H6tjz8pZ0f9
I5rJ2DVBRxDtR8w6dNpG9tQLblYQfUNIKEQmWbIGep7XIIK3bVCmA6ur2a6JjXdj
5JjnBoaEZF0TUvDV36gaTYNfAHeKupdcRn6jqFbQwX0qct8bO0yj7BGH3f2ZLBzV
sor8DU8w3aOKU078bz3u3giAxb2B6rgBAiSv8w2aI7J2R5GpWNZbgFyOleP3Lpu6
7o8k+JhLbr5N7AJac2yX5+QyS550gl/bq0d1swXcmNBurB61A0bWwUCpBAgnZKsk
nkNMx99V5pg5C7kt8hlwP+niVr0gVpTUGcFz7LoUey1psDY+In7/N1mVpncTWukD
CQssVibEhHkz9QoZ3iPEFtlwO7pVkzpWwMljR+iQs4h314d2L/8Fsdd3ihgYd08k
96iuiWbn43BCxldFOEX31gw8XLvTDZJSncJ0ryYv22/u7lkvoIORSWvgL+nORGUH
IrkWcQaB5wsxDSiTmiCA6EZkqp0WSgHezsoy1fRRm1j5R+6apXbPxySktedVtAcE
krob1FxUq52/p7L8S2xQ5G6qa7YmlI4cajbr6lBJH1j0fur356w8L/1fuAC78hA6
VT67ClDzE0GngdmuBSkhhvfCu32KkwHjA6kC8RbUY/Vl6s0bx3ppZZe2n08EcH5O
JGsbQITMCDZhHaPZjjHtGF2snRc541BGvN4oyyw6xc6cCZRzgRgIoXmUuSher7lP
FGWMRDeICW3vDseZ7lZ8CaUKapAAdSSgH36JD/71YM5VKsRoC9xufjGiyzAdfiSQ
oTexdaYdt1ahx1nP3aQoo4f84HnZ8wPcO32D/UK7QRcG08zk9aSNlYw1hogJw0jj
Y2TXDS3YHlRI0afXzLv0nuYmrperaJoRLBYaAPWfJvcF8zPl0mW3nqMIXDmtGMXh
2dpfbt+5lPriISyJZzSoNTdA3S8c06f3Sa5VnXWQuZcTKeJTpyx3fDF+i/6dS3J6
uszM67SdI2gCgRw8/231FQvFnavpMMEU6PcWsuFQ6fyS67SAfJRxpd4GvNv9clWE
D9Cf5p1T5rwSHDe5uXRlaeOp69Z5vRJ/D9ICspuyakCOTqaU3RNPhrksNPRF5DFF
O/a7IwrVPGr4w+BkZk/tWu1PXOnFkM031VHUQGwiR++7eNcVYzEeIASK3591ApMX
YyCwlvFUxz2lv1FeVYrX/6KjwWQz+QjgxcBT5/Eg0eIt/EgyI8jPa5KmCSa+1Gzw
RaCoVGyfGdvnUNNmi8uAbsIuzDpoznC8bDof3VUvA1d/BC8BUNbAopDfhaDskFmk
TCjEgG2922mwR/G+D2T+KmcRmN/UCQIIcT3NzThlph5MVvcETCLzcHEq5AR5QbOy
pXfgA6nbX8Yf/7x1dNY8MS+zmuoYY/XS6Hd2ovbzS5+IX7AvKS+C5XNazlUVXDgG
co1YbxDEMm76bku/YCmFbYMmFFBcOkbubEYaOTcFkfguktApW5fKFcC1ETRiU9gV
iZEkNMd04dxc1qUqgkrky0gIiZ3JO2w42G19oOqKAxVukwQF1xltq92Mc1NGtIIp
nRt3T6fyQwDCrsPLCxIFiNRByoRn5fXkYkZWegj9P9X9a/VewfyqggE0FlAAXxh5
LsnhWmJatw8ml9J8VUrTh6axQsEVm3tNb2pogPSxadqCHGO9u+mQoGXhbn3TSgQY
kVO50JxPmTuenCWXZQifPBfljuX7QnrM4716U2MtH0WhqyBypQbjK572vwqIorl/
v7v0j5LvSa2SO3reET4yqVg7w3B8604i6lyGTVjDPCusjqXGm376CXtNDIhV/J1e
Qdcw+QjguuEqwjJ3WQ8xjKuR9CxEuf6NMbxvU7vtMuwfIR2JENbVMigqgFqnqa1w
uSTt7wW/eOVkI4YV++ufGZQVRtqV+U4P9Ryw/aZSJ7UOa+nFeMWhSeAnUsczcOS4
oqdfjjDN7FdnfmRX8tVckSy43fOL2wE7/8uqp5a887yWDfXgW+7ALN91PJMWElmH
2I/JVyi8aNCcgKHRA+Jz/xg21/gNkyzFnOuUk/L//dprLvYJLNI8xFm44nv01Cff
gCLqvxySdkEG3X0yYkRBqNpEPowcuGtqVYkjJ0jDfM1Kcjy5DER0ArE1g3QTBkNR
ffeONq9Qqo4hpywn7X+6o0pN6fI7VXdqy6+tjgNyoU2Xh6hL8yz+KafJmY5fZaam
BJB8rRY5qqA6m3xu57CBltpRWK6S2bXL1MMTlcYJjT9RlnW7jvputRfUw1+ezThm
M4wbJXKLczG95j7kCbjYyeu4xWRsznKgUtrLrkXCJYX1+oPLFQn4ubOUvdPwumn2
rcehkML91lTeLh6IY3O5ZrsGzY4zHWQaVqhnNskPaLGtAtkhJBnqGOBzQeNXgM5m
ZMnTlHMstJ1JNAyiVADbzhkxsMXRRVFUWZgUjTSd9z+8gs0dJYeI81kpciMaI782
CqW7voIKNFxtXuqiWtxR0B8q5tClTE3ePhfKqbShh5WhFaKpRhMpFASkPyjLyU2y
tpfxEIuokMJJwO4KQuL3398YmpdUDaQYKfrlPstVLSk8bRjGAYgdlsSZOE95xa8q
XT1UeDEU3Ty6dq6DoThPWRKTwiJ/3g/x0gsRIaRTKkg4pTpcBulCtoOyTRZQkSfA
rck89+mpYL5+aqmh5usnsaz4MrUKc8Z8/I6eaSY1QH0YlL1vXJXBVBhsO2/GAgC8
fELJS7p64awLLhhHX03Oom1crGnCKt0YLRb3WFBxLsWkkOfkV8f8dIay6EuAuzG1
oGPIhYidzHgiqK2tznoaRAtTGKx0KX6TMfeK/PO61DqkMh+8rMtanStKxPettoF9
ONC6gUGPpUbPRIKM547TKig0Mz5wYF5A/ynVd18f3V2Xdcd0kZ9T3LoUzB94SF+c
dditfd4Bn6uPxCbRc+egSkIy6H47ALcyPPCXbpUkgcieGocfSNzfB2ZLDCk2+BDA
rn1QfvVZGKU9jpgzeIQ1EAuKBZlJI4oD76l31yRvjZEy4wGep5Mne1peacCxxgLI
ISSz1nXuDlcBlPgzoqCbQ9y9k88mO5h8Z2YFFb2+CH9mmb0+HR7GNvLdkaYyYR7V
Nhi79boSS9+OOxpAkz0OsAcSjq2a5hwF2ETo6/ND1+RgiTFp2YISHiTn4Qbg2Zil
6hYA/JfiaSXMBdkvoeng1B70X4eGiKDNrpPI2wOo0aTBCyBT98WxOaUU2GLj7KpP
EOpa6SUSbjEmVGjdVcHTYFBK2hW/CA16esi/QKC9p7h7jfgVxRpkD2+yxxkgAKP+
Cr/lndKCNg5UE60K0mDIpyCj/g6mHNAU/pzMwJjxNzeswU8grabYqDZ1Hr1fCB73
CTdu1EZM6zq6SCtQU8J+0qX5MJs/mM0AYlyHZluTa6lxh+jva4cDaiAwVviUUz7w
yX8JAlFt4UrgDcpZvA/intULLzZoKl0wzpm3cv3nCnRhjontpz6+kD/tPlusWQX3
quJFBOxitK3tjJwxGg3zS9RiftS+nxuSaYad3bD9hcO4xYUhq4RarPDZO1CxkJyR
TN9boJcJJM5WVB68oA4l0zN/3svtW4DY+n2uTKFDg5+7pDinYSJdXH9qAxY+tD7i
yoXFmon05zcPksxRkPf2t66JPaPGMnQt0bJNY4GCTE4TNEszJjI1oD5jpGrlp2Ej
FmqG31UZXagCuIRK8TC2UFP0l0OzxqikRPSCSwkriEW/mn5ote4rUGjyeNYMW5kE
xVY1fFKOv1SQWldR9cJoRgIn1H1xkVRVpDZJUDMj40bJ3/uj+deenwe8YTMJBZhd
XCEzqx7UfGOXXUAgwu4g+A0vS16uc061XgP22fsF7aAywiGoZBQd6tHOPAHavuW0
E35hxRB3dL9eujKQQCB1esOJ5Yi+rN1wFRJm9g6p+0ChxMi7YRNA4WGaw6KtvBp0
JBzk08oW62grVSyowiaTOxj1Vhss2DEPCCuZa/N20+atUjDS+L/4FtXkSpdPDUsH
inn0ozVLyxNoypPZrcUytIQHNlE5vg0XkaphwmScHPQmM068CiRNTH5/TTBdqsFv
cwopkLxwI+AAOZ+xbTF35tsgaWOov2qPWayOXQ5VJG16d38r/Uwn11e9V8nQpM9Z
U+68L/mLQMBTWQag3kmysudM5zT48MNn9kizJf08A8QCmTaft6FQbzdrYNApdGt/
gSTCRCp+bme6PQM7p9TILRg466JWdgw0BVnFDtKPdLJOhnpvSe3RyVK1gFz4SAps
ebvWxxBR1cARNApuPygcGFF43laHRMsn3ZdRtE5rBNLfAHIglNbl+Ob8kS8xpZHX
apRLYuf8kgVf6zXYXcHVkYdfwA+05WXvRVGAg8wUK4U7jOH9J2RDy60edWT7f8TF
mg+etgaCQ3SBuW35jiI8Cf3EverFQMitf9eC4G66o1S60WPbtWdWx/EZjlATHWM+
BsHakTI/ZkY/5YZUmlaaIaY/7/qnK5VrHqZKVkkyHDNJ8bcECVsgbsCihAg0S+24
19KPqUMMYvZf/gM12XGPICxawDIwtIJA9aCfMvhInqHAdB1J+xXqELqkNkzXynGr
bE0RrZ/KIHGJmpI6b9ZTlQpsii2UT4nBcvq+sN0j4Xd3WwhMLio7J3Rnk+/m5LMh
Vs/8LOHJXfxRT6DA2hByjfMg4tPTVlK3a78c/Xwe6avQygVY8ZfOzvB+usjTqIew
cgLnlsa5fRSJnt0aXFdHU9JhSIWif+/HUK5LHM08Iykd+G5BXjeJf3Sr23v4yL0V
AmnBtlfnzm2PrvjNm2h3UJxRZU7AqT0aWIIV48A4cy45pT6ZScIsEPq81B/Eermr
QnGs6mRdOHWL1Fi/FmqLZ5hKAdNgd32wNFS3cKZO65zD3vL0hAP3KAMKJm2GpN+2
bT/gh/i2F+BR//didT7AKXUgWBfCOrKocgRNG2H8MTqOKg3jB5r+Q5Msj99qbp3s
s83AXDohwnePqA0xxW0HDb+UXmEA6TDHXZcrsrgWJgRGR2NGFLXq5o1x0BJLAMMY
ZlCC2ab3hPREzB0mQDJHtwGSLwScMuhSOgcrTnDVOroAS86yUfzVx8RJRM5t8rjO
Nzi4iVYTZhrTjS07LsDsaoJXbotp6GWi/iUoBQFvu/Epoph3NXHdgraYze5+K7LE
mRR5mrs8jb+B4C/OcA4GmEiEgdktC+C/S3MnDZJgFchDcHTsIbZwtS1ACqA62/Jo
6PSXWlpYejmwWi6ZNK8Z7bCbMVkQMrD6AkPnURFiiiTg1EdQ6dUBVtGK2gaQFd0J
VIGsz0ifZMkpxsJU19z2pQ5MIPpvF6dWcJFH1UIH9axa0acQ9esEoLjJ8NMgkBAa
fmm5ymqtDFUZNi/ABUKee0VLTl0lq9M239iVJ+EqS8g5oSzuT5j1ny7A/5/T9hNO
90osm+gkzbYskZ9K02oYeSmGpL2DicgE/y8nENWw9kBncg5KuEgxEgdeDFjln3J6
7wFf9AeZ4OqeSw5hiqK94SCm1Dzyj2SYwMa42AfNgWC7QPBDjNZZi7cXDR7yY1m8
Fw0Eh6FHuW7y1tsiUkQUkReAJqhoSZ31c33UZ5Z96O4zxrojktsTF4qKkV1OZOZE
`pragma protect end_protected
