// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JgBUnKDO+/Hmau5Bb1wt4QDXUo6mASYx70mFBtUjnS+k5sKJjV3vx02BUo87E07p
3PPitdZnyN7/G/glw1gS8Q1yXOVjdk+XpwoR37azzacvOgCmrVGL5QUm136O0UUc
Os8AGX6BZsuo5zzW4cPTtMM8oqPEXBlgn+TQnurgSrA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 38960)
TzwcSBZNWjtIpqHMslnS9ma+DrqSJeYxju/auimVJq7DU29pUbRevGr9lQKUrbi9
swwerDbAoufuUePrsyOhpPI26NYoRgACtJwwzy5f91uZksFBBTyuytIXHwyxTYJK
sqbC11QrqHrt9gYOLbd/DSN/fEfxfTrzUS44HozZjm7RlxKQH2LUCZeKoRe03Mt0
m7s3G/iEf3Kfuc/pk6aSdT+lYniSVri3oehxQ+H1yjo3V0xYRQHFug1jqU6WeM58
DEpcb12H6X49/AIC/iTWM+79l+PoP3Uynoj6q9+R3rkFY6nysMRfi+2Bz463ka1u
uZURU4+QDVnU/3tFsEITJ9m0hRlXGzjI2R7XpZTSIBjrTfnyPIRttbIlyJobb8mP
iHmGN8ZQttcVFxAsZh5eW7F0n6fU2mMjW7o/0JCVklz5Tw4qboRiuGdGWlshWi4A
B+GmzS4Vi9auQlPdkTyP3DS6GgZS8IH3Uf19qQw4I37swXqaD0/5jxU/CSDP0bv6
3q0Mi41zmrzKMqU8szHUm2TfIhJ9MLIxFK4txGewZZHNDSKG87vvB3gRIjsKi/x7
V5iMZAen3Y88wdCzFQcW16LABg8uAzpjkEb8jrL+msZ7VOlWy8LVnKWNsqppe9wT
aLJx6tftcGKtrWC0Taco1gREwdybDlOZsJh0w+2bFAI6m8ZwHeF/LxZkwfqSsK49
/vln+hayHz8aya6IaSx6a+i6anfipmAIhKGDbNp3p2aJHiwPanue/G42x2POcbSz
xiNlmAfPLffxpen8PmBpQ+OEkM757XIvuqwsrPoQIW813TPRFPsC+T0+BfKktw4M
9uQHQgwZfQp6e2nDHuGdJ2+cPz1iDHo6501EEVTVQJ90/1ojkkoNMfh2b4i/XBWK
TDWq3n8NbkWkVZXrwG/63dhSVb0cRkIYvBgGE661Sdg1z//zGAH3N5wQ33dSqnd3
axNGalav8V9bYuZUhApic1PPjXqXl6xETXvnB0Rv3cnhmH7iqshwHa3Ibw8BSDUL
Jp/EI6af05q1b21pFkk0UlT8gH/DEKlFchkhD/smPSpK/WMAF8ukBIgoZ5czmtQG
BRJzanKy+Dx3I61Z+oj/G1DS4CxzYRTyBjpN9JtAqxFz0vaOW78tdJRiQq+yTwTM
T9dSx+XUg/QyKtCrET0QZBRr5B8vpheBiNvwOxLEqoLeqDiOLDLIl35NQfOwvauD
ICxWEvpQ4Evj3EcMk13Wid4kjl6vAfArKHJipunpAMQz54sGLXyC2XEMcoTrXiku
yEDJ2S4p9imEgZ3HopnAsGL8CitJFsHZJh6iWs15+7tm99ST30epmkP72/PBCvqB
Up8Xhqn4Hu7ILRHXvkb7QlGFFnIXbZURddNVnW28P++9vH8xNQnzfbnVkejLkC87
VQtb2Z7UofPKjbOljSRYc7uH5OvskkCReuekIzeUaA6NGF4TC8/DfS+yNuRx1wdm
SmqyWjatyI9RSVJmz5mB2OPJh0/LFbzVLyt+sf07NSpWY67fznteS8qnzMCY93Lr
RP3lny+aFtnSwUsInHHILYbmwXwtWofx4BAmg1Ev/rYSFhk7agXSKYHVmzKrS+LM
WMaltLO5+U5EnJAw0pv9DQgP74a6yXn1pPXGjuumL/HTH2KmLaxg44SuDZUKqMWj
HRL7WbLuCqvZtr+9aacWKzFX4chVN3ixkWrpPvzpUmg7d+cVBwN4FDFbJZ/wd9k/
9wF+nWRntm/yegac1Jo41ihvjyAod0wKKRmdYu/HGynz5FGQqwy5s1NbXENwA8xl
oucTMu5XGxzCUcXpeSQTZiWa4JRk5Wy0jVvXSwHvR9K0dl48pnxTPGJZWYmhH4eU
yrlU3iQv41BBkSuLM5NOoKYUVGcFKFQS4M/uDW7E9bf8S5Vh55expv+Bis/h9dWU
dJ+rKL9D4RnQFpUCbARwEF21fT77XcNQLnsTebZNxMsDUD8WimXLGglP5BqHQymj
iWTFW8dvrBd9rIBTy9iKdUYn3SKk/E1U3feC4MMOG4Copdg/dHT0XukaQls+kIff
734VpQe5lHys3s4mHXIr4P3Cbo3iPu1flK6sckqO4TuMcJIQVZ1fkMgs8XVYqkbA
BY+YYPjtzt16DSca3+gfjiZPvhrt9R7sM0pmyOpBw8FAog88c06ierotwf03HyPV
LJvgBkf5AIXGd+MWsB21sXVPX0yYBwbLkaG+QVIGX41CDHP0wAiPzpuRa6y3UB8s
lbDUtMqfq2uKmc9pTcYS0YZBzMNks/lO4ce8HBOvA0tlo0FR7z+Qpnp9KLKnLLC2
TaiYn0vwvtHC1QBNMJCb1GfUuvGuJn0hJIfJMkDjqwEyB7/cMnwZb1QjmVTX8Yds
gYQRJdUBgxkEhSE1TOQrQMbKhvDXAJSqCXhzD2Ew1QYnVHK47ZgVcvxzNxJxeFUL
nltWPCR34j/pyOXqPvWIPMJi7Ejdj7WGjR5sNKtvqFrEUGLZNsGbyR42M3WNWv8D
5Nf8J6qNhrN5x1lqNHyDnCjDgHKhLcLk1dbAjs4VF2U39wsLM2rFtnxpi6pYBnHC
2hzOkHKhrjnkcKQ36k+FVxO/Sb1IYqJTDQMtb2sr9MXFmRNa2lhHBFInVYnkbmPN
XXZqqeRGbldWTZWmy0/AI4o1xl0UBKJxhR9nhTYZ+FWID3XRbz1CZIlGgDZtu8Jv
56jGHPDlmZeL8O+D4dGZ8C4XRfqKIHCtZPfT8fN9e51kDyaQg+86LAmlMN/9Nka3
D4a+IL+m97Zh3SHF0r/KVI1+EpgYwndBZc/hac7X6mvisNJb/8OcsqTHfsX61+nQ
Eu1MkiCsU3we/cGIdalzJFAV7BN506bbN8NcWbkR2Xsw7rbMW4zcTJYQg+9jq3Uf
FFBtbSfK/c1uhn2aiMwLvHAnxDSaqxQvNJz59p/Oua0TlLcRDxECxhAbvIOASXLF
o2AX0omRCUr0EUFxm7PYiWNBnrkwPdQPd3G0B9ozuP2FAaZqxIa3kWytEnYpXPB0
Brr4M9JaohJ2i8gDZHzVPIYA7hJY0wEWLkc1kO1Gii5Bzdzm8Z84HUocL2pnOpEM
da8uDL5gHZrBhlCXjJPmWNwrVSFLk48yjcBmpLCphRRnTPdMCBWDT/Xm4t+YDfnf
Clq4PojBqZa55uJlDABtOCMB5ROREHuexn2BV4GySP6nbtzzFC6xabTj/THkr7N0
1J30edO1l9enarjv+hlH4I2Jo2GkXMP+7ilghSY/byoveKQDeOnCIcbfFu/HSrXK
WiiYkpV9KmGa/VdGWmE5h6KbECTWzhejjJ3q/a8/s0rn1O0+R6cPtKGtHtBU/hS9
ssAyso7fk3fRY2Bx877ny4IZQA1oAJow7ggF0eUr8oRO9e9WqJWtKB+ybHxv/jcA
UUBmfLixIOGR7AC6fdK3g6NB5naW7LkJJeMGUQCahMvDVjqCRsPDdiuXmIipXQSa
yFNL9cPZa4lPrJBeKOQKuONPoq5Izxv9p8VBD9iB24idEB/JWPC5gqdK0ohBYnS0
LlsKIzJ8DBgXCnbJwkiu1zyT1JDfBBTzChTMkxjaI1pDBw/SMlDzxDv6jbpbhF82
XvUTbo4KpPQIJ/K9nndhTUJNYCDuJ2teOiMijSknxes/euMvwYkG5zGtKyEwx5ky
CHoF0St+xVCwuXaJdzfJU9tA6p7Bn9Y+cdWirdq90b62digCY9mPVDDJLu1hxaZt
ifp5LF40t5DrbkFmK542ufCtdtUSRth0uWhOhCmrLbdlkNi7BKH78xHpomuC91DK
8LoUZbAw3Nv3ljxux5EjQ0gQ9F7mxeQrq271kYJczvi8HkdaCpQyd+2r7HLqFW7Z
5Tar3NwvpA8RW8wpWQ3awkMTjzOMv39iJvnigDhg4UiOqxUp96emRfWPOrt+E6Aw
kje3PId3zd3y5jl/Om2N3qWfrHkxv4IaBZaqfpZabS08+5O2ablGKqgASRGalIzC
ns49qsq4h2vQ+jeyY1+NsZIM75QNAz7qq88o4StVYPVDd4l+M0hfp7UUx2x4Arjt
d6YlNJWH8+OOK804lkmy71+eKygKaMGYkgDNcRVDq9DmKbMiFY8qOEvNWEP1Oljm
w3iSe23gVc8O6GuFaD5zPPP+Bk8DblWt3wscrl0jZLqibZlCon2o+1DEbHli/drb
kFwnGTUzsvef7mkT0XOZFdAYpyvjoYGQQXJ9xmmEpVccjkR+njiFrB5mseTd6XIA
l8+BBAVmDXFafI0PsWzlszq/tNqwkIfat7nUFvFYEzTEX2Gx2hWCtQ/IdlsU4lNt
/7Q+0Ca00yTjgRLtqbbrB/NSWiZcChykFcs4jyeH8r9qavr1uYfdf+XiRhedpUn0
t6xhqLx0NtDZ4YLxMCkm7Tu1j9fLknM+Yc/7/JCA77FACCbjM45hgmzxaXWQa1RJ
FHmWzRYWL7fDznbBdRir7x/ESEe+77mJD6TY/PwWY0PJjb9+6pNRiUZ8G/7o3x/9
yiGVbY4UlL6yoCHgUJLOyGMDr3JXdcEKVw474vLP7BoSO/Khx6iWzWT54qO0bD8S
6QrxhugiOOyMqDsiBQMkfs6sAGR6+dgY1G4RiJu7R92/pjim37eZolUBbRFD4FTI
1895q3GFAp2+x9cn66xKp4vgH7huunUHhpvtnSzH4vVuXquC3Ek2n2O4CQ1ANhQN
SfXBsZSslvLjCOAI2qZDVyv6j1EBWSRO0vEaep9HOnCSGEJ+4czRhQo+PH853kBo
qID8sHJCz7Z2PuUUJj3xH3aT3amtWMDkM9V4w/xUFFEUvypjTqLDIULcg+wvtNpH
3mrVn3K+WYuktLOvOSpgioUUsi771PkAIse4TMy5jNFFKg13lsbI+wruzWSoS4s3
iaaGHi8NXVBwf+xJ4gAJUudGbG85pXzNplkoKjv0CblXoABJ02CKpGF9wj/vHkwt
Ty7lAgW2KwFlxTyV5YGB89i2kmBHweBRWGI35fnTsS67OotJnyYHEJ/Rojq2Yj3A
nSuGVpFnM011IGizIrJ20vI6P6asSkXdQSmomRing3rQQKJLrRz09cHFEuoSaeMi
GMbBlWv502s4BLWwMxalmhH2PFyaPED0YHs6cDyuppqp//ISz72V5E7wiSOBwbPs
zeaBK4x7YNmPEwNsDh4TLH5fKrukigd8nDvAnIuNfSzz3nvY1fWGG0D7/8IxZyoT
LcSlxsifvVTZ4h/HT/kAH/lLz94m10hzg0bV/jqfJSIC2io/T58kS/5a/sd2cSel
CiItQobU8+MdS2ETY9yOtI4M90XbQVwhnG3q4CQAKr/CTvEtes4DezaIWHeCil1D
Jk4r8cmMFOfIB0OwCKoXzluVZ2SMLuhGKycDUQZeSth/OsADs/KYgq1q4t60mWdC
TMCE2daD4xZH8wlt2IFu354s4uzEW9VQZ5umZTNPXuuRq/fPcKYhkYts/aORzZSq
IQEz040zvWDGrgg/n00h3MxsCwnLFcSdYCrhNAwBx8yg1eFJcQS39WLPYcaqusC9
FzEVhLkM4BynYdDPmKI5r5xrc23zimXYPJ+X9oVl1PVHO2bO0wzMKVI00ciM5ln8
0jgj874JmgiEZtKwJTqmouS0SyefWLuHSuSt+SvMjYqHI6S2JYkraFqeKLgoHNGJ
HOhutPq2+sug1PVP3fZt5IwovMnfT/WsjAsLn4HiNXJK5ES4j6i+8AFR5rojHbrI
flYc63188q60OOZDBb438arD1PQ6dxgfCmLInBaFel/vMlnDUpj7uvvXwyi/6KNg
i9lWWtHY81C+oSWHIQdGbym6AMgIRkVZwjeOCPk2PKWM6bU0LXxMT+uMj639WkFA
hxMJP2SH1wtUB1W37+qhvcxVjJu11puO7RQJtFqOFYpq2ESnJB05NCz31U4UXP6W
nPYVFpO6bhoktmwM2d5L85/DJKumpx2/eXpMcq9fkyEwKXuT5sgaGyN93InQ7iTK
ek45GbBx3VkRW3tajR+pePX7pJhQjcRXRiZQQcpHSq10ecCErCMMrPdyNSt8iWnw
RH9hWcIiha8iLkUeVBaz/NQznKQnDfNhptyjEnSDDKnnKBQHeHz7ufrE0wvL3L5z
z46Dcnpn2706tWlYMdKakuQ9F88frNq/3XLN/yukiCfc/OBg4tlVG5P7O815XmBC
0RanJjYtOBLt5hIh7AG8ByhCOiM4xj0ENcuqzmqVZnQkiJtBLWoFFtPQCKjaAJt8
0SV6/Dgc0sbdDD6e1RI1J7qq973WhZNoxEYKlyx1IxIg5vCGZDveR3XXG0kP6ves
sxSsgB7T70YeajcnHY5AoLkB+Jqa/5qXxHWylSUuTR7UqZ/oVXeveYIFec8fipb5
ut2qTtCEwWuH3zii3A0nlVkL3/ROYv0cVuUaX+L957hNLPoJJtDCcynSYqwNP46m
vOZ7BfTIiXpymrDJgYgOEet0NeiKaKIIkhj0whQSWBb2nQx/dpjEhtOqNJs310X6
Jb0XqRxU6/kZ1+iExHyjBGDhfv4fsLFV8iAretyoHONIVEVAhMvjtAjs523c7w7Y
7OLKLkDAYsoycXi2XgSxtAhoHVVegXYJ2hVShFgo9bKO4oxwbyv4wS5U6RggI9ym
OvQjKoaUIcteezXuxdS0Ktq30mSVYGTYWDY0fuodqHtiv+radvtrOpLa3k/MVHUH
S9NUi/Bg/DvlR9kaiu0KpOaeSNHRYCrLUvaUn90s/NJ2ZVJIc99llR1EplBto6an
hwqLo8Dh0wx/Szx8iUFr8pwxmlfTRU/xd9jOZ2SC2sVuglYWOJn3i577SbrWvrs6
kRY/orxPq0U0/ZBDducsrqRJm/sz26bD7xSWuQZgyOQ4LDkqqryOgQo3KxhEvPbs
3pRDpLG9u1nckDYrLISYcgpZIj11CcZ1Kar0ee+OD6CttUjKF7e5pUzJUu/8pX/A
8Oxwro+ANtVnQOorvSia/zlCCY2ieL4Y9XXkii/xxBlCObOxjUZU4HHPo4mDZmBn
L2ribSAcoVpB9w7RGzgXOapAQUiuawj4S5fZrpGYlWtzr137qxHs51ibRlfHvB4t
GVpOxUMoh9U9ZwPDWn5gEakx5eh5ITYdsbsEQ3dUSp+hZaezMByWrzV+PcpJCh5f
7XEVdfDHgspPmxfyBPMYpYzrt6xE/A0wJeTWO6IixGOrSmB+Tsl6xR8lPGgITYLH
eM9wioXNYQ70SK0SjsqHcNUKS3xmjThfnsFXN/RI1lTNIWxHj5efiZD736FV1Isg
VRwlGUcdkEfLA5bo9mWA+v+0wT/FvlEzSR5pCJCCkxYrZPm9tqxIxOKlRyHu0Erg
vD07PqCRDlEgZ8bivFTnci7nDJuYj8MW7VhLRji9qvCIajZR44IP/HMruOoKHydr
44bnmaSNeOGEfejm9KUmKOlpdpEVFznW31SdMKf+gGRmbsBA8wXPOFpDNxMUoFOU
eeicJlor/RVMqcQNSYJcE2xbb+5bgr8BIdiu16ljfgT+OvTYVji1fxd1pFcxLROC
qWVfbVYRarhOy/bTvbUW7ZTP01aMSOwtll5VqGv2BEnjLxfvBdRMlXim6Kkr4pnV
eZ5Xc1JLrgwSUQ7M7d+KoXzlDtEvuTS1Anzxk76S18c2PNZxO4BpTJ+e0ClktJi4
gbAGWys0a21lW+MLGneXKfXkCh+9h/uJcbl2BUP/hQGF566j4HU63kZTGvfQds6f
+OO1dBTo6YF6+vP+bnwfj2vztQyeloZ1ij9m58bWooju5ZBsJiA0IIUJ5Ogyy57J
5jXq5chXc9qPUhZEJQYMmJrOI9DlKvWvRI2/lsBLH7gZgK35P0jZui0d5YtTfu8V
HRBcmYdDS0z28L731sKG6DRHnaxg9/wuyizZ9/CuzGiQ9tze0wKV5/ILb3g0nwWa
sjWFoTOrRf+a8tUHHpzTQTSXbr78uaZ3LQoROSYpxa2l6PNSIIltNo5O1k7a8pv1
egLBY5ePBsBF1iVCJPP8CIL6+lg16/l4DYLYb0ZcT5jxMygbJc2zsoGnWLe1mWRl
HVAjbTXXPYxMMZc8kRyTk0eIA/LEmPEMBtNiEFfYLyTvkzKOWvwuHDqgsV+cwYVA
WXumbK+jjKY3R971cEKhRjAaX6VoSusdWpJbG0ySXm2y1QAzjX+g8ojPcs5W8E+d
OYBYtFULSqKWrV/dUrd2ViZdP4UzDqbxETKLBjGkCAbmGUUre/J6CLlr4CzKQ8o/
ptbd9Ksg8RV8Ay0iZ2DBop9sxQdrlNnuxXdTR9LEL7xjXow8fLtmVGvWP8h9XACU
Rvs0yxhP5uEYHYgNyC+PB3wtQ4lz6ej+Itsh+Im0maVXDjiMPSDk2KB40csqrDG/
WekeSid9fjYO0+iAhKu7ejt1maYF3SSN9TTf8e5fMdHA78VwhbkjPQpt8h7RxcLb
94bp6LCPLehWC8q9yimgoKMeqMzy1x0+HLAVJlgNdmHVyPhLqZhl447awRPSvT0W
l6ngYwrbj6Shc6N/TQkHkp/oVmY7ltJigdefP9UE4jqBTujawzMvS8obnMhDwWok
SDCSYm+7WWJW8vc5TtVBo9wN0eq5Eah56HjtEEL89u9Kgv/ZHYTMiljGF21nRSwr
O+yLoE64ssQpIauPImBsgyPh/3Lfgko8hlA4NZZOWY84Gd6Yg/h1zKXI7GkwGA+J
xKNBi6rQpclznJPoi9kHb7FQPgW6lkxdvNrc3Aa+LDvb9GWsC6hVr3b4ZMeYrmFt
lgZDAD51x0YnnqdocFCA2zKOp3HNGNK6DLyOmCPkJnjnGqDL0H/+rXd8EbiNt5eN
sQXNVFzNGbToG53acsKm3eSA6MhRNioxTqi6ipPJJxJy6BUpZrzBSKcNnv6r3aBj
V5aLM9+BU7DNeTb6GLwbesNjYRANFVcx1uJgCsR+duSXIQ4rzjJOKZ85ZtDEEwLC
5yeBtdI1GK9lqmu9rBmHSkfsctbjKVcaw+JiAXRZTggJBYFLtmNd9H0SlAPSwi5C
pagL0RsZkoyiN3MSBU64olS0xH6L3y+S2UQesi9mBWSwboXi434cO6JJl6s+1cSq
gNlHpqcHdmaQrB3wXq9BPWCqsP7cp2x1hEO0wKW3gv84Yuf2Z0zuEd/eiwsxOlTV
m7dhKs7o4ROVmm8Nq0lahK/DK/1Lm5m1i5E7ABIYITBfmkW/MCIXZydQq0LOrPys
DT167CfQaPPkPluOyVrAQj00KvZ/cO8xQUVbY5KGMDZ26CSOxUj78XuoHwtm4gZK
J6EsqqjFR834p5LwVpncMbb33h++JvvL4e2HXYRa7qyrqxDQMcydOykfiBL47Vm3
KNybnWU6pRpb88Q0PsTY/TjjozU5PkM/92wP3LOXYjPJgtj4MlAnficXlC/Za95j
vZjlComtxF8zpN+sfb0YLFA435j2rg8E+m04Cf9rxpQyq4lap9p+GFjLdMh/Vwoc
u0YEGBzGmPRD6aEOsxz2yGCk3kglVAcld93ZPcjavtCY3ADQE7o2Ot3TUnvpF+qn
qQvHR2P7xGolwWPvLPtjgjSl4Eogv/FAogp5MZtO+DvtvVdXlLHgCCpDi9IK5XaU
ebkpDPQbBow2I7STqqhsPKip5q0fmrjYQZw7s2/VZiTmZQFwUH+aUTAsRl4GUmhp
FUC4xvq4623tPDrPlQWSpWcPkK3EvHlnN2ERlrvYn1NAB6pjygbdlBs6U7GE6bwD
TPsYCMUyjNrniWnvod9OD75WPTp+voUI8hwFhT9uhEFR7XYZCZPMtVX2uFjXjYDJ
AtMas4QjbZ5y44mJNI/yhxImWn4J273LbqyllrWk176VUCdyPtol8Rr5cnB4+TMP
CkDV99+CO4M3bXhx6h14taQv0Zs0RJMfny7Ba+PDfQYMPAUO7wFCHxZb1Xma61pG
55mP5Bbb2+nbB3uFoMwNQCAg5cefGQ56rjr50C6FNR3/KLpJKlm6AebkJMF6PCHV
Ci7ksm+IGaNuX0HUd1O1zWlGmHum2JpT0KKgaqy5nkCMgkqi38WZ+6deT41qLkr4
yNGFBFwQWhsbxDlhJv0YoxvWQrJML7MG5RePXCluzmLwpIrzCF+KV1ShiV81uoUm
Hrs9Xa91jxHumgdYKSySbO32nLpG3j3TPHjgfUdFtjg31uKb8XhCttJqXivRyaVl
aeEFjxqK9OfqkURuAVr5oMz1A7pefDmNNPe1pBEUFOq1rRuuYdwpmNTqgH5Tmt/s
taj/Bo5lE1BW8RL+mJKjmlMZE0ltmiBX7Jmyl2kmnWG0AY0ZAKGG/XH2ApnxdkoD
lgSBRhJdb+tGYyNaA5xxMp+gYZNOPOTO92cI2AvEfWDuEi4LLGJxE5YxhXbAhbfK
uRGcr6eZEkXc+UsILLqjbEHQ7U4ywfpYFr8nPU42NcmAc1Y32cj7WVp4HRkUYkne
owXTuFdxqmAbZiMLF1sBUJ5W0ipT3j/SRF9m97VAeuXDe+euPvh8dWQ9eNFVE3F8
7/e/vOeu49KOoP8wSP/5BWadPVOno4spDS1pPqZp2Cp0pMPJ40oFmMJRvKR/7Sfp
0gi0e/ggGPXONH8or3N6aIEIQZ8nW7wO5uwaRXnfS0eZmSplydgJN50MUkmdKMmV
kyJ+GE4cZ8EcoCRwvQombcLJAYwGp/j5U4Iq2gXb0ctm4QvvrzTYDxMbI0zFo+n7
jJ990raOu+517QGvz6Cvjh92N1HqZ/KbcmopkfSY80fmLolY0tqQy8125TAN/4Vu
mxjCSg7PaH+8E27m2wTo0ClE7PJssYr6VuyWOps+ee9zzNvDzoBiC557WP3O8FHq
qostCPPjay/xE/nG3KWM39SM3CiBM20wU6WejzBxvO2nq0fOTIENR6Dvoc49Q0/m
w91On1tG3mH0lvdlJk6IqfC5silBIKMe97h/7pbjqvajRpRASov/MCZQIxSIoLHi
kN3bVHISumVaMbzqahYom8S9RUMZfco2WLWaH6hJs7efDX3WBXyEyDEa2ZbxENT8
T5zJWmITvaYD7gM0XO5J0S+rFwXHUZQ6Vnwugp1JKvYGG6Hr2o91+1nAg3WoCyM+
5tABQZ8gp6DtPFaccjzWjTvk3erotSBqrvET6aifrCrEbRuTndHKB+RICLGaWgp5
fwY34kSSzRvHtU+9uXEBKFuyxb4Owl/elUF8We1tWA/w9HAGFpHx8gZt6z30YEth
oijVtDZzCyybxgJs8BIH10j115+s3GbOBQUM5MF7uo1IBdKDra5/ZkmnsFtD686X
COroXXQEljnxywS4SWbZLu8xGcEZ70iZP4Q+8dVO6tIdi295ck66gjAY+Qs76LKt
CvCl/U7NTsiEZkhYZ61YN/JlarTlhWLZ9VP3480vWsVTWdIGx/xP3KbBmJxQlwUO
y7P7au+ayaqa5kUIiI2W7BRzp3Cn3DcQZHeIGhxkL+BIGxUYm1wM6Gxqa2LxmjrW
sRKhCc5GXA97tRs3BDslMcNRHzHrmeVjTdDoqHL9K7rPd9APR6uDba5dSK5LNyN7
zFqx8kXq2ph3d9GbjEJZ2yGFoI4VMyY0sxisE9gGVO7liedYuoBlUqFgY+NUIok2
g1hM6L49PfFZNGnJgYmU8vH75TR/rJ25ybE/W5VTAaCFT01i5LbqUgXu7hAW0CAi
CErg+2LKz59PE3PSP+jZb8UPSVs93aSlQv+LM4A0/or3IJSWO+q8VmvEFo4bkfXE
XqaOG8xQ6n70I9scWcs/0d1QwlSBA3Jnalmq9q+64yMfPWgzu8gFV9GWbS1fei21
6Pq/p9zqFnJTwwqT4TdhN51Aw7LC5/GMHHC3oujm2cGylzWqyq/1t63cAf88QbHB
kZOfbF/xlgawhquZAshbti530yZjB1gJglqRijGpdPpzIViKvGgirKO6UkaUZsBD
CDo19EDxtGuijtFLWu28Wta723ZUY39jR7lxANeHDqaRfWMXRD7mkXsabplpue6z
WXBF7HMQHOhzSJ7EUxvqpgFsQ4dsOBZpQvhSOeSul1QOGQBZlSjML6ooe+e4Bu64
+boPAYeBZ46VZwiNdrExifyvdmc0k+nW15MzdQlbLQWAlvZIFIlAPcaHskexSE3I
/xT+5JwxNGjJym174ysEoCMGurGbvZTFHWHGl/tvS/DdJPVHtkA1p1pTLLY1fVQS
YZ5C/5pfXAY1EY52TKj11vRz/AbhPxTiafPE3zTNgbxL1A8NlwTz5igG6hzJ6sFa
clZFXeHwvLG7jXe2DQbk1Xmnf1yQdYUNPj1pDLYP7SkAHqjaY/FLv0VTcPIs8V1T
hL3Hf88LtPU3s/LtvNVIOnWxeQueNhP6SRGGBuZ0yFZzciPMQ002iwbrn+Hr0Zwr
Ib86WOul63aNvITfkYp0RzZH/qaZ29wz5Me+BsW48vCkVJbYwSVPnOZVCwsLhRXN
6LI/w6WDmc+jhfT1WACdVeJ7xDRnh/FjA8JbJE2KM+CV+Tc/pAyOb4NRGlKarDbY
37zJDuoXNQJ2PPcYQVoInHQvrtinp/PAl4SNrs3bi6vXmP6RAK6OT2TWhlQNB/hi
nqnLG+2TloeQO112OWOX/+2zqgYZQAxr5IOnVahA8Rl7cSjKLAuDbyt/qGdKVYRI
/7ckGo1G2KxmGWFBew1RVOJfm83bwnWPhXrw7LobGRPgLo+B3JRxPbH/EzB0hw72
Hkg2SbtvnRvAsvDGx5q7xZ4DtTon93AN8+dbthyE6nZKoblALqU32GHZoMijb3MX
08RBFgcrKivR0R1XZaYeXDYnuyLFLHjyPx998c9kr9ad7V+UDeN5C9DmV8Cpqy+2
TmSBGuPZXbu2bxBRAaVxRjoZK+vLFin6RmylEj7FPRH3IuOAcTG5lvpXtXyVFpaT
BozikrDnzbPUZKm+rmeL00MlJUbq6EkM1MQASyfgJ9bu0ymGbyKbFiozBw2D0zAB
03zdOnJhEy6ZKjXVwszHZqTMmKIHfBxKAkRQxRdCuhCjZGxs9yc2lfo9S6N6Y6nS
uMz7Gocav6OqQRAvAsg8z584S4xiiS71q7LWMdGlWXE8xT5uzuOp8sjBKnlz6sTv
kJWNJmTSSS99tm7l13/LUzNKwanI3u2/1q90g/z7hB4fLh92HiLXkaEB5bqRWdrZ
K7Pj33sXZi/t32i9oH11ffRBiv7QGFz9M9RelzeCmU+wleazcVMcsXWvYkNK2XjS
dheO9uOout952sSvJ/QHcoxaHSMTMahWGk/gLTSWwwSiqtY3oA7/XmJKwmR401tu
pk97IcNAy+zRG04Kces/LqX/58djIm/iz4y4rkNKq2KtLLbi7l4Ir1E40656dvuS
9divfGwYpDrAHwVyttTtkwJkrYnCcDkOG1uwiPM3HWfM5FosA0wxlXIiQuiKveq2
A63+BmfUe+XYXWwu9+urFsDai1ijUKnBl7Kf+CKF6m6UD8DvCUp3WZ5HFszTx0iJ
1qId7+E7RjgzKocyQ/pSQAyxaNP6qDvyONCvy2k3+1YTCmKeGz03BMZmwrsHlnp0
AhAHrQ18MqyYtOcFhYMc3Vlv28svGpbr9kKdIgPdRG4S+EucXriirOJS5uB4A+o5
kBsmfKH3ishQcxGr6b7GDS8XJMkdSbNAb7bmqJTtF506LXMbasO47u2ss+c5JbU/
ck/pWvSuJO2/d1QZLLF8G6IB3HIS9HLUggLm1eYETRyfYHVTA5yMf1KC43RT1ECZ
fYRlAaaIdB2Rh9ltwjyxMlM/fvoF5wAFzVn+7h/MW6rENSwbNhA49GfpqhrpE6qn
rZUmQfpysnBS6D2d+xdXLqpHaTXqiAo1xiN8TbdM/JO/G9RuAgY/+clXezCL+rHc
oiOB1Mp1PxV567vsgcJ1ZKQnpRF9fXiaM4KIYt2BgGiTis53SqtrQkiDuNhGWrm5
Jh6wlYY6vJVzMG6yF5bBuEK3T8IsADgNUmdmr6S/prjRTbsf722howxJz4CEKXcN
EYqe8fKD+mkPKExAq4n7SlqZGtkloOrHZPx6/qDhO+OxtQWgQDfs1JneCeyojhIr
Nedukfv5HVpsweAxZaGh/UuByHc6H/qbatZMzORylhq/EQi/2qHVZAzTm6jmmZXW
S9wlVdYNUsQ2/yJfKotLpGKEl+1YboPomycbmtJj8KCr20HjPHBqnoPLbzxoOm7R
hzEIh//yLDHEisy1qg4Gmp0bVMTsI1D/NlYT2/IH03CwR1jLZ+e1ZO3N091pqW1K
pOohAb4HQfD20MIDI4ehtxk1SgXULlkc2cwfkbDcEGQwEqA4WKOFyOCJUXGXxZ31
gE8zHi6ROviqsAFifKe4hAHjvcZN51R8ne4k3qrE00WihkwQ19nWZXepTT5kDxPN
Y9JQe3VnJhm91ClpNNdEsZrBMm2airW+FdHFzRXA+fkPGnlC5NYYHZAg7gmaFisL
QNkGqHc44RK0ZVsRaLOwQuWRZV7dizv5JXOLkcnpCcBEL1E6awFlZvQyS/Cry1a5
bX3axTNnu9j/EXyxbTgJpHvRqOIxd0srz4zBX6ezV2D40JjjaeXS6HI69HsEnsKU
8/y2M/R8pMXFf6AteOIy89azCbk31ztaB0mVk9w5J8x7y03KiS6AmKPFuKhGWpyq
mKfRiUEsPTXMCa6CKW9wG0WLQf3uIyHIBQMib+y3g+rM1li8W7tntnKjNA4Sorgt
ea9HnGSNLKcbMHiZ+hC0P53X8wkmYDWz9Mmqc7xcHwM9J9DaAYgGUlDApHt4/cc2
8t8pJD0rUH92EJqkWOShQfu94xSPDATVFSTCTrqQvQmGY5qLRCwlCkCxM+GrFriv
Qzi9DOPFJeKtxtXM88XDCtEdJhlNjifRfSLAN1mNtv+eKN5o0jUXwD4AqA41JWtp
ANdwALBCMRhlDgudQmUraAf3dxjSC4HWArpBeXFSbHfo0XOEv9ULDlCr/lhLa10C
n9emR+37HkUUP+xSqX3l1furn7HeGhOx2lUzPkTT82awSOv/L2/EdUgAa+Z3lrIk
cOOThe9Y8cT2Ytvu6eiI7uuVS7b1oEycLQncRYQY2ONEGOaAD3cB39khs/6gHSsF
IjRaq62kUZNRr7H2VYvciCfsNNfd7nLce71FM6OCWqecZihwYjH0BCCDMElEJsmp
ybl8QVfpSz+cLuQAbLx2UvtZi6YZYODgvR31vi452wL23NzLjIbaNQ1y8SvH1gBg
6Bb1zUGKGPlT+0cetct8Uo2kUikCbjqjGarkIcpXKSF6HChG6KJ24K0wRK3K1UJ7
+YnIKB2DVaO/M0hxktaMyNr5r1Wd9W1uGGmTgPkfCcpUzlcxPCT1bU4UQmgnCGS5
cUePuFq9vxklT4p+d5gyW5X1WB8qbWdZwN0KiUjzhEG5MA0AYEhjOu3nEg8XAca0
wVLQ4ULvefnJETog10/kIM8MeCY0HR5GdF03/25h/mQSru0++QYlSk0cNWV0//v4
6O7WwXFJ9oFiyxv1MdBXrz+HsVwRLCtT1FdJfHOgRf0AmrnNmQJn9YtLqSakX0cI
M1FRczmdUzZB0F6sHQ/KLY/F6yAGaUFxNzghLtu9W/J/BweGO4wRCU30l4+UjqYe
p+B1/J+yQrNRFmZkIO/CrBJeBqIGflqun9CPoyOJhh8fik3KkKEdaeq2MLkZEWlN
9V+4gsYGNwV0F3ux5aZ1wE8oVSFahWhq5lYEpyKWaayR1cuD1ECMo4gUfvWCjVel
BgDV4+XiNTP6IXOyB1s2QzaGizhlVGpv//7mH+omK2eb31Fid1GXY88lmB6Crqrp
8m4fXEHLR4kP34JseYY8XUC5PysNhmEB4YvVson7+/T7AChRm7+Ns+U9nqICxhJR
GsIGAGY5G7E+LHpzVZ7E7B+igo6shfwF7TLZ38UQs3Pszlkp+s40G6bV6F3cxYry
5T8E9SvoUs3GSBi4SAYj9tuwLpuTexYSYcBQYNcMOpNcRRBtmCnkkdFafXQ8iAKc
XD6QXwaDUfoRgZcF8kI7SNkBHWuTQCgaFR+/gXpg6mz4QSUz6usJ3Gh/6DpfpR+u
AWY05/mZ69VuaK0wYER8b1iEpfB7+geBD7N//FdemDzB7mDFFGAAggIDEXeWBFdU
L4DLdL4ZoVfGIqdV+JhAcMsSGdzntChDC9zZI9uBLiQqHKeuRrmjOUTq9nKunu9i
04dKe+AMrC/SSDCNyDHacqvJSgePxltEy5fphcLUJM7U3ZpLEwS7N7HrBEMPPg+Z
5VHykzDCxH8f+AgeBvVDyu4QzdN9LskSiio413tV9U5/G3CKHaBM2D5IilFtep4z
/CMF7afINf1ybkL79Kg6vYeiYi+koZcUkZZmMzzUpwPOQsq8hBfjUJbau0Rl2FAH
31aAOtx2AITj0RVmnAyBIwj7qE4NEpbb6lTttjzEzcGT609qUAjd/SgPa09UIGcn
AX+oQgndAmVQ1KWPGrZpWLWcrCgeKuBJ/Qf5t15/7vIiWnA/v4m4Uj8rfO1NbmLw
Bk2RUD64Pc5J+dep7QCIvrxtEoMDmderyTHbZHHbNUYfkk8QYnL2WB/AGcrZsdDw
DFe4X1oLhRodbzwmBnVC8ePsk7vnIaRw5ZeeGi300Bwp0Z3QJE37NNFj0PJqLxHG
TzsyvocdNvnIKczVtRsU5q5u2Bfw5b+0sity8gUa8Te2+f9lZju40zazCAk9uA+L
SnTPZp/yPGFv3XpFv4u+kHKaTXOooyPhn5xRadMWQpTzgm2Iw0bA4UxbjDHgsBNY
QW00aIkqO6QqYghzeuL+UHj9X9LCG6AIDNZ58v5D3oSWTWwdvrLndQyRU6W0D1Dv
O7JA/Xhp/4TGSLUesTlgXDoQ0hf9eXZcyEi8YWL+QIblri6tE6Qy84M/Y7QPZx1e
Lq6HUkNbhzsguhojnndhUikZ7CiLig6Ph4mL+05k5u3pikIOK3NDX8+Sg2Lv+/5c
ofxdLaUDNKtNxPN3dAlC+0lpxn6K80VocUy0HsMW69h8wEXcQ+wOGY4NbhpeEqmv
6LH6jBJ9uIPyGHzkKYDm++5+cEMonLTgPYvDsjyfFLfyAr/kXNJOAvqCzxrHQKx+
op4Cms4X7scIaiB0b0h8/MqIBopqTRVoX8UN/VUSpZJfN5yoRp3GqvP4D+98g7D+
eY2mjtYkrvXhGlWe0kEW2mVew8Dohvwq9ss8ut0cSYFomEZ4/coEyDZdsDBzK/8D
ajUD3XI2dcZuGCE59+51d5nTMbyTSasheahxZmn9M6JA96ULuFB0qHR3jQhFGwpz
ns6w0cWMLkg9AS8evAg3PIN5l86+Lt6YmvVBKtT17j24jkZFLYv1/TBc+yZpu0jp
BhoG6EBWJz3qHiR6xmiX6SwGrwQdsvqty/vsil91jVNJo7e+UtXbp7W4jqih5OU1
90KQUlKd+ayM4rObqcLzhce7hqhgzT3EihmK7DPexfupbvh4DHel6unuR9ckYefj
Nh6TVUjTjbRQDwmf0xA3YSjseODcB+JPwO/HKtSFZD9fUudKvEAJO+IyjW1oP40u
4ScFrj8N6FkV2aIuwDpmbIjIEhyv0PjRH6PxO/So7AHW4yFUwsGyt8jtRQbFbOoE
ZDBbnwXXrio0SXNZZws/JmRG/r5a3IUqTvYrBL2ntuzX3+FMFKCkn5d9iL948GgF
YSXIUnlly6RginJQGQbWpdAlY17zjfFnEyv5RMSS4K6gF0rdIBKNTcHO3vXlLpwa
ZFIxocsfqkGCWlbr79nY7p0m9Wa8pN6pIsMj5sJ0x86QLwajC1kl8axSMSaZkh7H
/BQv+B+hpadhUN1iBu42L1Mr2n7JL14bK7hBqJLioOiN9EsmgssNYfI6chD+aHZ7
HZ97wPjoop588t+NNYiv2H93s7stNara8rrYeo/R4sXJzwAT3Xy88+Fat7MWKWUG
6lpxulL4+1U8mXLvfPeCBnGWu5QEsTTouebPfjqDDR5vcQLKoOj1bHibL/VASTjy
UUv+FbAj3Va21uuU3juxMV9jSfCYjWjuqIqp6st3Z01ftJ8Yc4MsyOBgzm26lcGr
TWxX/gFuMZ4JBWADLNF/h/f7SpdRyi0t1BTz3dfpci0tpBDMZk4Ed4gBBgtrBSzj
0csJX+Rq8ZpbAl8bOhtBnfofuAv53gsxIIfgRfFveJJ7hfSQ7W7YmHbSYuCfvW2C
eH1HazmfiEZ7cIF3tzJQUEPp3UlyALtZ8vYCNNSDnkqMPPTjNDI5soKIqVmMMzz7
x/czPDj4Ru89g1ng+p3FnKA7r1e92mOB5X2rAMVNFp2IPx0Er3MTLPeLEYS2fb/G
Fmn5QD6QL8iELFUcoIXtjW5AXo8Bw2NMcQvKjGkT1x9YZMKBC+TAG/7fN8vEO1Zk
V6f+3h0GXM+MQ6sBBgk1UE/4nw6ZmO0SgNYGBkgO87y4xi1ec43Yb8iLjL7fEo2d
1wQQiDx7P3qK4q7g3rK8rZan8qTGAA1iaAKWSHfOzwOPP6eeCRDlPEf06fpJpX97
jUOIAooVMQkBIpYIKZt1RTkDr29s8e8tgByhp5g4wrhRwP+qbhGgiqqu5t7XUF57
WWTgJgXfco8OsPxrq9KVMKkuAZLUTDrEUpjluhGxx0nGcxo5Vyrh4BCuL4WgKDjl
WUqeiHxgODvpc8M/2PJvC25nPfME9GQEyZN3PGhteRf6tPw/iCexqUn1nn23u391
pNzzMI7o6z4ihIPsTaPS568FbuRWAUn1XpcTZ9aT4GlLikLu2LjDJmKs0xqvhEgU
RbBcPTPYmw3siL4WlADRT7PY/hvjFKPiwb0ugJjaCj3MEtywyLyTcl/mG3oA1CvB
gSb9KaelyeicLKMgezgeyF02nH08gVkTFUQP0tSeR8Om2iZz1jVUBQv4/yJrhts6
RhmoAbmQfk65NoVYIoaeQqUzx6+IU6JTHahnb9rZmTrWHBMuKT/F3okiRKbSNNIy
S9abhQ/MMJWqtxEqV8oDyOocvrgt2S3X3JS5OeNximx7HUapCol9QCiuursxbsIu
0EAadYJgOYkOdawx9u4s/ZddLTrzwpJiri2dPYCmgmV56Jghzq/QwvtRT0kZ0svr
BznRLWIZ7wV2O//jCaQN8U+g67AMxUHZeOfznU9MFyWt4K81z6pImfeFR1E1DuKs
/q4hqAWtVYNdo+I+ZrYm+eRwEn/OiRTnbp9TSlBTeBLA4Uz+N8kEm4NsLX5vQ/Qv
CvCf15Q5y7fZjrOymZH/4sjiB7X3gXtAur8ovpn0lQGggdSaG8MpjVEDzAG8QlMa
J73hY0gR3Np/1DmEv20FJCQ8j4TEmwbyvVM/TKlhGjVpbxlNE6Ndje1+kFt+f51A
o43JUNzTlvroG7+TLzTFSycA0MWD0QZ8Yg2TnNqWAGhLKCqwiXyIHOiBZfaopCSf
wElMa7iMPdL9K7fPU8WD9BOi5QwTngheB2Hw63mO/s0pXqG6QUTii3J32fj2heL3
Lei1sVSJeB335WHmOOEwyoEKIxoFrMb13DYRLCbAGAsiqlBh1lzesJBzdCXsD564
/eTkGSBJNb8ZSSkFakrfOif1H5LAFf3yGSniK9v3HaONADERMvIfYi/PHN/+yG6r
RHA/O17jog6Sn7D/ovIL8NO1e7tJpvz7IfYJRqqyb7EuAWgWPq0xVd+Wh8PkPBBo
NPSY+y3EMs+mznTkKzkA+u8wHgfh/ILv7ckpeifHBy10dQ9KU1Yq3fJ8nH5zfnyC
orUqvH5WeGCx9OaDsSSYw7dIrBLnx0S1YqJR37f1EeJDixRPig4vqFfFLh/x4LfB
u1SC2GGnj15s9D17swit3qh65ecURlSv3kWBLoCIEzGhWn7aXk6wOiwZKAUd7Ta9
lTV4olNSO1IcYTJN2BWC4EFhSI2HV+m9pbiyVFuQozGoht9PRZTj7Nsks93zH/th
g8Omx9ohLlQRC63/F+dZAQhdObESbSs1eYTb0wjZh/HurD7ERCrdmzwj11k29tOe
RL4CigDC3n8GvSC7LCC1LcfOeQUTQ5X1G2gHiySDAJW4Wv14HqiLHMNEHD9qFf7a
msRtYXnDTgesvFwHhwSzsEvQp1j0exJNuKhxS+2M8UZvKKqPm+FEl31dFynRb67a
+JbUHQTNluvhD0PBw+U49yXGfn4rjZLIUrlrBesRTa9uWo8ZdB8ZtMo/Q+SV6UW3
RdsgVW5/yz0N6pgKQmyu1RgfKxFzU6/TO2n/DA0bbIl7rgD/eeiU+yj36Rsis9Xh
KV2QL1ut0yqqoU8FL1XfhBksooM+H8HGUwp3pnriYKTGghRbT8awY6+j+rMo59j8
yBUP5G4EmuEOffQfkhq3zKscPqZ+v9KQluaGXCFITI8TsDASAwBT15JX7Vi6fBpT
TD4NsefJWC1o9DELaNiOLMhpnJkluChjggvTfpndOaJEk8u7fAxcKoGOWGs7otFd
D+ZavHpZsoHqZOK8m6JUBYYoFA9LPBQNv2Jt6exD8rdVLlvBKO9ElBaT9MGCmmiD
ihMmSGrvKj+1itjVHUJ2K6wbG+S30hoNijqA8N+VZWgqnn144kE1DOGC+RVi//Mq
/v4spp6f0IGSTQ/9BADCeNXbQAFMP7aoBpZ+ZlvjdkEjJgaGvt1t3SsgGBxwmuEJ
pxSniKVEi4quoNRmugP0xeslkhdtoPq7ezbpc8feFYqb0s7NMKXR5xcIje5qZltp
dlUefF/CGAmltIf8GrfRpTMIMFM/VDuiMctXjGMZsscksI020AtF//saUvkxPL9O
e9HEoeI2bd7lQVN0FeHTgLhFYl0XqYfh/W4BtNWVS4/0/mbEV1t4kz1hhlelEWxp
zCfxjUwiP2vz0ri8iITPdxpo1kp+lqrVAdCYhrPQlPH/Avgnkh2Af8Y0elnEwoAN
PpL3z0TBcqcqssIVZUY5y+J907+UODsr656Czy6Eus73DIryrb2oRJKqaKZ5q4dS
RTF9/aD/wPoFG/a9h0UgtSlFYAqY6YkUVgxLsCWAL6XwPKXId9pTY+iuSN09IpBU
sZ2gs7hcqdgtPfUxN8Fq60SfzmS2S9kSskV4mgBEweMsRgQ/PA4lVU3twS5xfEar
Ae1PFBfa7SIAFC2m1po37PnLMNTC+Sr6FexHreJO+8MH2WpzFBJoe3zuWwyn4Jku
5K65ypVCLmdjB83tNUJMra9aQCdlY9we2Ig0qrHXZURql54IYx3O39IdBzaT4VBQ
7kWYRRLS8hlDknDA9LdY3TrSErZx6/7CQqt1KHpRYbhssUsSOC14dBII/iseyKA6
3fS9vm07pB+/xQWd4M9Du0n8+Yg2eqDWjDUWOeaIcd/4P+7F/jfxYImhRHt+h746
loBggO6OnZARiJZ8NkrWtMXVWGvWDaxcjhj/iJSgd5SYmmCVsb2pSNBVRDF27QFR
40etBnohwNM8J+tGQzhUa7qynSZFIYhUR17aqX6XrNvjj2mvh8aF+8teOLYQ+zX7
wtv16fEYX5sjN8i5OeMEP7hjNFuB/wOC45sGAC802i13M0wXDKXoaVwFARoRd/Zd
iYAb9DsYhry2jZIXewdlSHk2UoaUP4CmWcvKrhpNH4LRqBMQ06FsK6O92VwIhKxI
FFdEo2hb/uYSGBiRC4oGXr9gJyDgAVdCyDURkJQ1CYA+Dou5Ni9p4Yc21e704/Wk
WMBoH+QV+PSGw9WoZkl+kNX0juC69svMbxKOnoZd/iFpON+AxxKyXUCt6yRcRBiC
rlg+jws8cmgj1yIg3+LIxtzOgrh8mIaqfahkIwDSzNQ+zbtiOynyFRZ2lxnofZWC
vNHCOReT4dvNhGQUU18azH7dfzQgJ+DZSiICM3nDL3FrZ3PflkkgHj24THaxHgej
qi8r0ZcXFiMjlDL0gJpGHkM+FryR7NFZUmrhlXxcpu+S7o+23ZdMczYAVDNNGOEK
GE58K7S2nQpIuX5mHfI0OaqjTYaDHcLPDMYPhBF5f2rRP/VZ4zJYwGNgDey1Hdgt
ibn5/cicH0VkrrRCloT/9Igsg2LHq568bSX7D29x1femxEZtnySpnVzZYI+WrNv2
3AidR/4Xxr9fdLQaKSv4LhgANfK3Ud6b1YlXT5jbYuvo0Yu4M6nVlm6rTdizXaHq
XqMJH8CHI9eYcWKn9zKqIq6a7KYXVQvxAYKzLlJb8cnhFmMWYtLoLYlZZgQVErpI
a4juhLD77vnilG/mNwKR5Zz2Vh3M9A4KATvz3NldjmS3O5gQNo8DGSqfsxYJS63y
IMr85OOdLdxvS5DUNG1wEGiYgm/vGz5ez1uZnjsNpUZvnjgx4B+oy32UfhpZEZ2B
xJk4x3Wc8zXYkjrtLSQyk3kCru+Fndn+//lx6LPN4lytYZjrNXr8puSjPodyHPR8
MBdiJaq01DGJb9fqS7bh62iHsM5HWqv8NAnBcnObNNpOyEck3YD3goRE9DSqLmkv
F4Lgjsusbe3mdZWrimE1PcEiXotOzJmiFok030GxAHjhoRECDJ41Mf3Tb8nCPbFn
YUbAjozTlRPt3npWH0mjoLTdtO41JXyRGrkR1e7b4WL2SiJx2JyRSNtei2DEpNJQ
jsBtfArZsSTqDOtegvagfTEOW1XKNBdOdXuKxyalEqTc0XUgBkNpLmpkZhjsltBb
iv2Etj5Jz4hIkrZSjzRuZ2/wHRQWMHMc1aFafRWiid8ZZgWDLC/TM7S0nTQV2N/F
UP72IDbxRKPPtsOIfVHIUPHRfs1+L4cVSsyZu87JP/4tcAl+QsR6Os4xwdFsxs8Z
gYYSY9CFVT+8PrZhYSl1yDSUPffxyKX424DhTyF+30LQgYjoloqGDqpGw2ivPy66
DFox/mf8y/B/86Dkji7xBSca3ARjdw0f8Lmt2qIZ5exWFvyh4IS0pAgW8X7izG5U
F5PvO5rqhdqlQJt4nqYOTYEAOnwiDiVW5P4oZOMyJ7vF6pPuCx8/B0eBxYCvAO5h
dglt0IQJgYLUcFDLY1K/abJLzBWAaR0jz/wEbF+825wJEENgkosMO8NUbvEfrSSh
BXunEoRnDREmGm7uddJJQaOLARlZXjJD8SIOhHobzrJmY5F8d7tkjlXzIaYMXy5G
y0wEx6X76jJUpGJU72zQAvuj6rrOwCnfMd7srWhHLlhTMQf5APjp/1ILJPPTi/zK
iHmtU192U++GkcifTYJMR7rjFy3s6XR/AJDE334aRzSBCh7Aegk3lHY3JHpK7nf7
8P6uUU2pIoiMnMd95Z7h0GBhlP2x0RSe3dXDewi8Y4Xsgrtb9gALGZGp1/pCVcXl
MTLhfgxLaLLyeEpZ6P4dTCBInVEPaTF+shh2XeM2yW92U9ve3aATWhZ2X8Bb5XO0
diL+9gO+PTBx5vvgvoUxNC+3AffmZDo7eDfuS2ackIzGX7La6GtGpZp3j7nB42i0
U9VTbQZIr29XP043py42CfFPwK9Z7Yy/nkOKTgPP1n1f629aFKvsRLOsABvtXKLC
44y7NaKzTMYlrb69f+WKfM18V7liLje1Mv+NMuFrdhfzaMx3BbkPyHLx2j21JqAr
l+hNfEoi45yaTh+lUAInj1sr5F+u15mFqN9mvQ5C7rR+1dZ09l2VELTaQj3GbUMo
BLXJzRYTkNOI3KuW7uvY/6m0ij1OsudYI52J9GyFVR+wwMHevDDScWbbY0csy+8D
LmlKOsWs69yLclUnMb+LmUdPneivF1ZxbA/iA2GaCkPjaFzYYDPHkwpHLMYqoHjt
0x2nSTEtUSsoMHz8ktykH0y7nAhl0dkzcnpGQ39zimODn0oBJK8YaYyiMFed3Aca
xfbzndGZC/qA5rM2ADeK6r8mBvNbmZqcjClhhANTQxgTQulsE2QXSjBghTorcoJj
xl0VYqiMFPY7xX+tqDk9CY7cjiiSqJFzeMv0CdYRrvsC88CBTIq9iPQTaXR+SBAU
4f0YMmx+AtbMMmq2iP/Hdqg+s/SE9f0LUxkikU5JMYm87xJtB0YprNtO9gQYG/Us
yO1nBhm/j2AhsMf0GEm3xh7E+wzhuzjhKi2W4q0Fru9KdCs27UUakKTXwFcK2fC2
elHkMFLFiRj9mEgAy0UppmgpgVJP/YtEI6opb3lYMBNgOnc77w8Bz+u9mrcEm0Sp
Muo/FlHuHBAZ+c/5qBtDOetxPi1tfcA+rhEBu6FnuWzTryUKqUyMPM+eZE3fcplr
CsccoBDDokiFexnjQTiJ78prRtNGdYcO/emnmKqowlUbpdgt1sowMvHl64CPkWha
flYhTg3LpvCnERCrKEfCDllBUf+3AMe5eFRiFC6iZw5RuMjKq3PbDGZUdk5IUtYG
hJLpcjG9rKdrv48OxNMMPwK9D5/ywlDGBrcrmm4CERG6nwVQp510IJ893pYBO1oL
rhC8Mglz+3VC+QmfyhbteZ9ZtN5caAPRHmllYAgjhHCiE/nZTtueNgMc0Gccq+Gs
o5gQgZvmFCcIQaRdd2I3cG+RINp/4s5NBJLcw+J0na7VPHlS+VJ2nmaFbwTBP4ZI
hb5tBlFTp1+sxO7VbPBc1zjbltZF6rZUUHkRwp9BCWNC7ikH4+gyDjsb57Vm9b1E
pepIBXmI3qmmJHjtRZpLzynPBoaHiuNRr6NRxYFl234QNJZKqI+NMbLDYZ2cxa+H
qBpDRxl56AYYrQWgKzhxcfnNKWssc6LIZSVFKGyoec8HLUMluWt7WY7gx2tpi0YQ
m/XWC7Y1GhK9J9MK+olKLmWy4Wtb4FAKpUNCyGB72zXcoyzxQk2AiqaMSXhgpCoe
Zp7xr0HJgUDIvEzWFp9TY6EznL0OJUVXfkjsqm8t99hs3nyYhmiY+dC8eL+3w66p
0kQuA0IAxmBFvt6215ssjEyM0Axn0BK8YtRD+TDJ/FSWL90Blf5k6V9TmhiTSm4O
tl9eNjlJE7IvEk46wPu+cEu3hPwn67QPifmuCGQMjfpqAm6+8ZYsD5hZOxbUjE+G
ds+PMuSXI3f9uJ/VpMj4AQtvdFxNnbDUKmfll8dhl/ewyTrdxUJsEeOmLYaSzZ1A
gxyt4juwvXAH0+3roJ+yDg1GQS8oGe6cwRoxoj9Bry2tCNgPkhUBqXLuzLv+mDLY
L31LU1t/K29JA1v2xsvrIOn+76jst2sZi84gA1SSMcDNzPVkfFNVUITI0gQBL2XI
h2uTz6PzXRDKml/1F5VsBDhIhckKAHiGkYvQewJE447mejkmGD6YNLduzRQA9mOC
Dd40uPAATZFLZHTrGKx6jM76LrXQuGkhF88b/t8Et3vB5oaqvSX6u7WsXqoNxO0x
v/izu1wb1jdGnX8spOoFzMWsN19bI1xMycopg9evk3WzhD6dS22WJi1zGJpwNy+q
ChhuhvIg9b+LJ9cJQXox49eBE6SSaMyEfadqn6739/AvhxjhMHr8jiUX+2UxnL6T
NUCtOec9XlZUmnSbG4MFDcTKV1mrTISnIIHfPIq9WdOOY9XNtAeHGX2qZGA43neA
KLrGPkZ3L9DmG2hiaCKkJXoK7492GfY9om7IhM8f480WBB9cFl7qEg6twPUBkq9p
8jAVSr5R5NOPKPFSGt+xQNeU+/CK6A+uPfYUoWnqz54CrS4cNYls+m+Ys2DHt7xd
nrMt957GFp/8RsqkJeAUZ2Pjd5wvXvQt1M6JuMOt5VZjRoIYv+R1hF2Wkie4LWw+
J7SMoDt6b8K/s6CZ3bnrT1ZIDCPHUuxZBWtHYg2u+hy3ysroUuceJB+UbXn+loCg
oXcaW1ZsgTHEAbswaqKaY933ejERvOp19TneWTTyZn+qsV8z6SNoED7Af2FbCRj9
HbOmck5WOfFAKT0vPvBtSpFXXM1R0zwLMik80KLQijadLm5IRcc3+3RHw4Y+Jh/W
ScIWZu1QwAzgLURwy+mQ1/KbVvKqaMGOowNC//orNmEpoTaLnnKoYddUt0SBxsWs
YTMB8O0A93epZp7S8NM3c0mJ8UGqfkHtrZvtw/WWQ43u68v7PbCZYn/GiF8JbOIc
mm/oIv85y/WpYB4YdzERofvCiRvaOtK82mXGdnBzeiW9+XWVUm+fyjWHakYCWdth
IJ4Y1yzSUKfC+M7r8EhYOV/r2vRUUPfquWMoMAwq8U0BEv75Hq6iTpf6k8aIjFZw
ZWzVuHgpqTsYE5Z7d7qctmzGnqZgXq/bAhZUsAvyEzsjSSTOxkFPygVIbFPclNMN
qGfVeAjR8HAXMiRuXGq51LTpHhKsMSCzED3dJ4RT+YCNAGPjPtLTwgPU9+n8vf7x
adaKak1qqWPmwq/YXggerMKkexEyLOt+ciSN7ey8hhjeIqGft8P1l/7cKZKsPcsW
LRAiBwMN57bIZKwAG56sH6yuYnSt+Reri6Cf0TBewlX1MmD4YBnIWjBwEVZSHg1y
h4EixsukQ/HfXIBiasYF4BIHkh7n9sX2oOwuTddK+dkwzio2mg9CYygBej1UH9II
HpkIcWtZ2SU7+d2SdpthgIDPaLJMbX2qlGq33sco7gyjTHfEGPeN2IU5vkCSYRdi
uaIv76qMhhzDuNr5vx6TtkgWZK6ITmcbnteROwYLODuAricJpAKxDTfBoWzw92DN
WmaRa1SC+8CUfxf5kljQA21D7iXngFgR1CMhqyKpVYvtSSF/egGM3S8hhtgEmniL
IxRbGNT5MkYeoS5kYe7h70b0UiJBNXJI6++75N1xYw/mhk9hlk2GTR4xEJNw2jJo
4SLA+Ya2RJEA4QUO3ft27KQeqnR5S8u1QKI96sD4im0iiICfl8oJfPt8oFsQHsvl
adRN52VOtJksErKhc+ZbCsYYrI9O/IdxSQEObMbNviPOaOPftqhnwPyL2CdPRgtV
2agE3a4XCVjOgqo3yFIVEYGDC1lWsMFN01e0lrOWtQvvRZB6972fWvwv2zkvFUsX
z2NE9ClagFsdRu0Jaq2CKQ4kqs8Kdmm54omLDcCOF3OYNmwbCfaxSyG/mbuY9gZv
dhx0MGb1AV3w0Ch4/zY6XbqTZPnpDa6hwcr7FnJBMsjAz6FbtddQeg+X2RImc7/B
fy5TsKg6Yz2f2Hr+nDAK9FMLkSHYqHNQAXdxwyhXeuDXSqPLtQ4VT0YYDs+D4+DZ
rx//YWkAkoZVkPnMAWASkkc6dDqNZo7WXgMt5oHxkV+Nc26vrBrZ+XPY40GFTT5c
Z0vdJvJl3E7ncuOpjfFj/3bmqmCsJVkdwcoiFS8yfRtZD4/aMTj40+SyPm7Ek7we
C5QlpOgSqsz/dx0Vt9Qi0MACsu5c0IVf93mZmOR1g6XMAmilZtd1oFChHyAhPxvH
kNSa/pyY5JLFHDtRpXm4agvE3kizmigXSzG7k/CFbvxqokSpmROKT2WpMk/a0EY6
tISN2LEElEjnhMVUNvcbcrwutiAaFBo3Fukqk7DlADSIb630+35C/LBCE5lm6t5B
wq3tscWRyQKUEZkzgGLkkjOVvaYn1du2efAL1x0iBMkQMae5ozJIIkahHf4hVAt6
NpN+hERVmDQNOTm+bUZL04EVL9GK/Q7WeC3SF8lm5xGI3WKcHpdGKj1fL3a/nVk5
dWA12eetKhrvRJuS31cJ54m7FOTkxseJHkGEwaWzENLTA+abbMxYhtXX4TPsMFF3
jmIO3EnprLQc/4aTq/I7tXWfQ7i3kjQh+bvT2V/52BpbnrYzZlmqSVSUmnRw/c71
uzX7//8bYwUyz2su9rTG4WZUuY4rjTpr6f+xOp25BOBwmespOi/JjO49rXgqRb6E
yDKpq8OVJurYVV/iT2d1z8yCI8kvWrmiGAf8BAtByfRhk3rJfvu5lrpGArac9bM9
U3ZgpLtOkS/4LYYQQZFh6yCNbiWnKDBR+ORjrdGgObcr4VusbZdxWg4vzeoVEcMQ
TuKllMfWYPRnn9u4ZriSCaHgNgs2Kia7UcX7tuzsnRB20o9oeOM5mb4Sirk+lUDN
KUdZ5mRcvP+Cwb4eMpsA6MlyZaZQMTf5WuLkj0NwFZ1Jrumb+HV4uosOfQ80lvp7
DspqPOcv1dkI0KewUONXTabUyNGyrrHPN4eXQDRptEss/nzbwdBYO33LyhjXMFtA
UJkehs+sVUyLVQgZEiXaw+sm2tTlrDxR0gnWxjqDJ4kEX9k1HbYAmxqf9Tw6R2q8
CusnYUdxPSKctJ5q/22M28C9uERR8qxe0fttUbGJs+Yb7S6R7VIsYPJF7kVwqmoc
Pn/2RnyH6fZRZPy02x0yX8O2daTp3Gs1JCHLN5Xg6xBByLvE+lv9ngSNp5adMH3f
65HYU2eiHfkNKIuM8MfZzb+bOkULMivfuJXhqeKzINTWYlkLRmcG76mw/l6VzIuE
7+rk2QTJsAFMo28Xo5S1TxxX52x2Dm+UIt/kDSJ0ac9ta/gi7rSUcObeUqty/4uk
0EoLd1PlnWJsUySv4qeJ235jN6k1ARNhQ5Kf9u7WgDYlpAflNO4Ss14x+h7azyIE
5f9cwMphYNgnQG74dKBhuPXFr20UYKPAxIDySYaK8mBAekZkA5VZDK21P4qNz3jy
MYzOl+AwFe/lhTo4CEgWZPbgQPzKf7mcvtEhhpIy5fVR/wlIFCwAk790talKcRqc
dBiHw/FpEe6IHwYSXN13wV8KKlS+JbD/ytD7TYmC/ApZMSwA2AkRqL+b+9lZU/tT
QeLCqWo3wn+RTi76wYDF4cu/0oy177O3xnImidKsMBtvv3SbRAz06K16Cdnev2oN
tpW71PbzIXcLdwftH//lhwqqn90g3DB52UIP78nEJ/MXwpC3tAvMHE0ycxsD6iYL
Eeq99Ibz8aTruqbirgvIMr1qpYZwJOvu78/TDslNHtxk7QuEiCFrIjl3ZO/ZlM65
o9ie4dYgGeBypmTNu6E4gdBmO5H+lVvKdO9/ipTfc9ZLqYeRlj5Z+psySxGfTAzV
FzwEU0+6+6QWew5gE1FJme7q1LgC/S0oQav3J6poO0bn8SAuXZmlPzqNC5wLGfGr
BHQA1ALutDsBIg6v23jY6JET8g5kH3ZnQV/OmtPVG1FeDgRKbDusFkw1QNwGh12D
mAvkWUYoHRW4Nshg/ugQ47TbhDzn2umyLdG0/4sjZffyu2yM3d9Ib8Y/Ef8xxESK
6MJeiw0oOz/UJwDyI/kHuS6GITY0CY+Un6UpyerN573yWMMMKTTE0vv+u1jRWszV
KZX9ZCVxQVgicqiWUxP26r0SGYYtozXdbvdt0Va8knhoLbvymAeX9b2qEjnTkJA3
nsjVV3cCBhAIFAfqFZf7hOdxd/PH5WCp5/vIOo23zRpeGh336qVJelKn4CPtneRt
JgeIhWp3VpPxT74wfB9X3djUpAGm2fr1g6c5XewPHOmd/fQVzrh+VUCT1LZSmnj/
g1Tf6m3zqsL1S4e9JWCB/efTo7uZ/O6LPSk/n/WOh33Q6Fbd2Pfm8G5SIJxqnNPJ
rgWgrc5dxxW9VYokad+6RUHed9BqQLh4+SfVVPgfs7593cfA4XIKSHUE75QleDFy
SfhpKKFscIAieAlKHwPkFgO3uqIXg3EPs4bJU/p2o8BySPrxLaE6aCffU0B7nJio
hp8ebWc+MW00EUYe/N+dscyHUubYoZ5pN4KdgF5EgeSAne99/Abf3YxmFNYmVElo
CjSH6mOpWrbC83VuqGB0CcGsr5599agVttnJ74OwK7z/Br492c2zioq2CiRy2Arp
DiVWyyQ+Jq3WNlOjWSoiQbgBbgihc1Jt+mvpuClKxQz9PRk8D9Hkg7aiVKDAompZ
RqCCG91/cs584EETq49ws7kNQKUYv0hkuFJa0PJnDOfVXX5jTA4R35VYXXjrw9+r
1ju+qsfoiZf4SVuWN347LjOUAsz9CV7U9hp4/0sDrTAmHj3Y+y6esvkbD8X6LsxV
P0Ry0+XII5dHetgqRE+bidEiy8hkmvbdxBmopnQIToPclQKX6/JAwieWcDh0N1ZC
HF88p/r6siT6TcB0eZgbUAgE9YkcKPUgi7Va8Q+EvMRvfp/YqNCcVBOFkYKKn6RB
WB8U4hnaLcm3i2CP407XM85IPqdMwOnu6+2T7xj77vz0xkk8QGd1bsX80y7/TtWW
inT9z8PvZegPO/9pVjp3BG1OzpWqzDoWUlXV8P9sVFN/MnRfXZjGMjK3owizHjin
qeu9cRoVApr4F7tXt7T0nigDq+u5JHq3HsTQMLaw1GdIE7KMt24HxE9US+GTMeE6
lj2W37ycM2r4RSvfdd26Y0FGr4SPkKavoNxb6F623tDCHCesF1m1IE/bn/6v/rhh
xfYOPcSa+bzeQK2nCs0MYI8NoD8hn2PSNPO1mG8+KLLKsgorwNi3Z0URxzgdgWaX
vlUdtXiEHcTnOndKhC68iMS8oMFw4AeRZpEgNrHz0V2zXC65iubyaKZ5xvQ97Eta
metZcCJUGm35R2OJU+c9Cqvlu7eTOVCrbN/tNKV7uy+gD0QQaZeTWqwzynKwUoBn
UAxY4DaeJToah7/vYRimpEagxL4DDOx9pMCeliqc1GPeFzh8dx1lFc6MqX89oqz/
SPx6rRGVw6j3h0heRAVc/HHJFRS4gLaAYMPIE/W0HNcV4VNfKSuYLp4OIxrfE0aQ
ilYjIoLGcX1nzT4Mfh+4F5E3WhYYiQ4bmGhJ7aDam6V/PTERx4FgTCvztnU3emkU
26HlArmK0RWCSPbqwCi6YuGNgk875uT3oI9q+ZXkvX4Bf3dh7UUj1INFo/VZVjC2
S/A2iR1tPqZ9q1CG241th12a8fO0HkH/VHn9rZzZiAlkvSFc6APUIq5xaUBAQUX5
H3675+FBQB49sHWCJXKQ06SvlHt77ZRBnqJ5pF/SBwP2E/7aodUz5HVx02g/Te8t
hY/7PvyCIhS9/F8B/njQrTCCwIkLQ43/Y4FnElylsyf4Mz4vOV9rOnugLlzh+s7o
MgKS8U6ynJdcIbCSko+NYnkWdgcDEysL+oYiei5eIXYtjUiHRSDL+eYSQmDbnQFh
VexNgGZ6HjjtWlwNSMU0+/QIqyPd+/OPThkqwz+czDt/Z6AYt/acNzRU1DuCRi47
rSPPeBrRbQkz8Z3tfBIrCW2Wz1zH2mqTeHQUys+fRObKa5XoAoSGgIsN6n+DOqZ9
8QDgP09duQRibZ/tbGN8r0FbP3LgEDJ26yqEcuhs/EfwogeQDx3rCk4JeZaBHr8q
MgBliJ3BcsieV9FXshz7UdhFArD9byQyxdTZRq4kPvvemjyIfArOLer47qGV6hyR
ipqLq//FGwyoZ757vB7UoahrQ2tBVVJLNyOVg996KRoLFCTRqIdIyoPTGz0BTC8O
/7M75TYiW3DsrKAwF8PWZREzmLwPOlLtaUjgmLa6Roy/GVtdqxRGvf2rbMJzAjJ/
kMbTK+gj+tmLZlEaMSUH5HVOt5QBDNl8OKxpP4GoLMYnqKRKerxlCGGaa7gR/WcZ
9eOrV8x/oMWyuqdBi2cGAAsZufydHQWyHUsO5GLhG+amiNuZhC4HQ/D+HusGOtax
0+rtaY17HL/PMcC1MABY7y1kqkirdVrzo3ad1/rJvjaBDzHJCbwxZ2MIp6yCtKN5
ucEQr+f6ZMypSw93fcskzH2/PSOTQgZVyevg2ABFalj0EEkTER7oXdhJc6WhHRIO
8YQjZMpy0tNTEEQdRgFj8bezzDs1ev8FVZslEt+DYYzUqTVoJlggY663ef3+xR3p
b5/w6ZgQZvEMUbeA8F8A3EWJs3SipNFND0ON5+pNKAKJ21S/PgvG55oLw/B3ZPHF
oL4ZJCeFzIfpPUsOAJM6oDgtFPsePCLkB+xdb6SaOsLxPZPcuD6/zVa5VUYKGYls
0cHJbHW5Gwt56848mwONJ7YNDDcQ5TH1gJQS2NOsrJFuqQYhdM48EMCofnEyxeG2
bxKftG3xiuwSOW45/vS9a4Dj70/D1pDVruPlkKfuvGHyqQPko74YlKMVEw63ZMtl
sLmBIx60t+YcDf9M/ddfMnZLUc/vuxV3Zi5vJ102exRnkQTl8ADUGuJL9IcvLy9G
cyP0NQFRq12yvXLsGYC1oGCvWdcfOAZ92AtkQVm9uEiC3+DTddImrnACVNtnuBIj
oy/rrHhYSY6jO4IVCTB50WcAbbM8lez4fnFGmYJ1FlQwjZzUq8ZiN9Hbr8l+7Vm6
cvve7167j0mFL4XMJunLlvAkNr8N0j3c5A0tlcT4fLTdTtwIitUPIbRRjzyBqetz
p7RQhaX6C8irNEvCkfO+cDUX75Eu2me3nz5n2qAA6iHs3wh4QnTa6CMrx453AxN1
VL4Fhmd9KeU6MhhfVhq68Pcd5t3PjWgHye4TNk1X6NCAT1pzP2Wt/7U9D1YLYzFd
9dAEjiE6MtSQEW2BVOfsAqUdbq7rXFTCtHPWW57hNbWky3O3B+XGJmXTBzgUW/ic
lZl4cVwjBd1ih/KSRVorHF1p3E1w5X9eN544wgXwqqSbIEJ+diMeOynfaFVyyvyw
EEM8Qs/J7t/7LjUmia2D0UVyU02zDrsa+pwv1dgxXsA5sd03KjW3vHcZLVvmMh/K
qZn2mNtGvW+D2toTY3fvBiGvFRmiZg8+CZxzoxz5XQq1X9Agc+JYrRBs+ZSvZ5Cq
O6Zb/fzUVVjMj7vTe5AkRVU6ByqkA8gGrUISk/Ov67uSV18UVFAPiDH7tzxikznh
yMHoOaNllGtgJFZMyR1lpHWFFzmt7gcvXmU77ZadQ/CWZ0jF/i9F9zMfdXnx1y1J
Ft3j48/NEkriILE5dKGzPydzbQTCQU8a5cBYcUSaGyGk6Bpt17t/Q9+GdxcybeOs
SuOahYRyfop3Hm6sAU8o0oLwrGfFuZc4J8PJ3AT9VlS/Eh5OHCfcvGmnJ9D2NTe2
D0aE5sn1bLdc2dWmaCexOUvbC3XSUesE1K/W77n8UMWHa/7sB/XWaD8QrbXI1GDE
b8xvB5MxSxQ6Hk8brkodSiaeaZEPifFDjrGuuQeDqpyNlTBeV8r16GuRZibo5ZDy
TtL4C7G3hR3NzV7PQ7+oKAuMSsUJPsSN19y34PnVjkn0Z9OeLvJElf4Jc6ulhCL3
ROJMhWRWiE4fLHQ5Uik7qKKEMZempEuxA1TrekXGS9Ew7ONB9G3uo8pgt3U0T2XQ
mDanzT+PCbug3AjY5PZpoygwERLyuAHKP57ZIZv5/FHfXQCABPMZkkX1vEccOTyi
u+BaFtQJ7LgsfAQ8in4FtwMkpio5QCc06n9nsYreK7BooT9HQ3OjX4OtrdSKUyPG
o+Cjjup95aXoRx+KDdPfnNnTpmOyVDfgKT1jo5Ljbzull7IeVnMLhlhnuQpPwzRy
VY/zy3moQ2/YVlZv0Ox8xYVE9gKMbdEj4MJgadZeobOi7El2mtMu1fW5mpAk9t3d
FMbFRmfTxiD89eTSca+XtdJNXQe9Emi+TV9vGVDJgQW23Z0su9ytJ4+nDpn3DoaI
JvDV/Qn1IHjmz0FAZ8fZ53ChVIF2nLgkUQbGPFsd5ZjdZwjeGwM9n6hSWl7R5r1a
mzpkIC0FTqUh1GXUx99AhY1OCBxzviPxqH545tY8cte97l1UeNRLrWVTG7lBvV9q
E/V1RerJUXhaEnok0lM1UhbX/Lk4xkyjE7dNqBtCyHtVr3YQy7E4TUea9NL4lTMt
B7y/Dm665VWtqGAtwaSoaKowfkmkBJRvMVDHXmu9gs/XBYAlGy7eKSoL+pmESy36
cFt/b+e6GVVT6W6oPdV54xxdqexn3GNXRfayn7OZOwa0ZgOiWVi0n70vPpLDefNu
9HK4YEnDUaKDImwwjWr1s0sjFUytT/YkKCZSo/Wiar8+nIDM5UMa8O7gj/tvHXYr
GcAyYHKJCebxCTlcRmax+KDtDx0OLXTMxTFZ+LqaNbsc4RD3vJbG+3fAhLB6kBwe
sIPKn4UYRsuqtZqldIBTkEo4Vh1iUI5Z5XKkBnWAp9a1Pep35zw3zr6weNrVgdEd
VgtxFtdSMdUWvF5Fjc6hynEy9TGuQhTsfoW3/NkbhHDk059GVZh1cr05sTmhGmtX
EK9GMzwMKYUabvQ4MQN/tulwe4ZEkkRU1uMZLB2VSXV1wRI7jasS6+4y6Jwk+kmL
V9J1DSkJPJDqELgL0SMwh/IZMi5HApsQRo4ZlBedN4Ro+p7D6cZRPHhYKZfwuAne
zkNXyulIhiAyuKdhCWFh+C+ywW8FILfCfGSFBIuWHOQruzQQL3NU6lOY6o5onaAc
C1lTKGdWnTvGy8nGq+jyCzO5d2UeF3nO31UMrL5oIA8/0DFabBjAWNU99QH++d32
n2aCaEalkBLN5hwFq76GDsmnK+MnTaCX4um/sgWl7A33PxcUNhNmyW8Cz+teoExp
TYM6S9Ybnaou6lQjOYU/qMqmg6LV5CNmDXFzu09JtXZ0hQNKkM5MjSRhlsLVOC4W
vCLrM0BeslilfK8VyHLHu8e0iePVY2usSJfrSEALXEelV3+fKaLAgo7NIj00348i
ueSGOjrqPLUzGthu/HIUTI5EX2JjeLN1hHO7t9zZ4glT7NnM2HAqxOtnDsWKoo5V
8C7TLHftm6KVTDsEomJkaLl82S+b2QHw7KldxdKFhfsdNTW2r+hpGE4zJj4NuPxm
/b4BBhwPgLui5KDaVlf6UebhOfz9KBsrZ3jRXTMg8G1lEDHNnq1nSzIIgX5kfPWi
XCnXKvYc1nkTPVXGBKQqPLMh0y9GkKpnCE3hLa5QL22X/0tH5iIUY/nX+kblLB5a
krAUdloHSNuNbxdVOU9FP1GTkJyNQOODmH1vK5GkR0U1vYdL3jizbf085KUFXhNB
X8ht6XC71tcS7h2XcXVBPr/XDF3OHHaSwEVCZX0n+e+HEBO85wx8sfT9w7T1V1R+
kymZ1olLdA80obHv30AalTpHiMpXP8CIQJibaRGbFZ9YFSr9kaG71wiqQ+VmC5al
KqeWm8JAjd3z6KOopLSIX2mCVLl8QwzMIHRAzwGVqX7w4xQfEAq1RsCQitITdeVu
px3/ixdNsrwJjCvWlMNR4DrcXH1qHKklj7QR3GrPzhU0WZgyTc14iHNc6/wRfGmR
5CqGedV8+95KDDU6sKbIVCpxP/b3gql9y5YL4y9s300lIh1hFZKES8sRgRT8WbTE
z4Pbd0Z31IG8/UQVkL5/5ooKwQbdJlkbqc/TK5TuqB1/qb1N6NamtUZwDcTVfjce
ie4d+psuXHBjmkiyQ5NOVujomAK3MD/eFiwrb5XV9Ln3vBbAiiiVHkTy8XWWJnxG
0724zPKexys5uImmd3o14MEp/50MHY2qEMJEQeu+9jYk5ZnEYXwShA8hUF7x2k/e
IxAPA6qkeZfPtoEZG25MAMTFI6VofSl5VbaidvkZfcQS6xSXVGAJKy1GltRbMvrQ
tqWkPEMQAugb/ILi+SLnEjuryUqWH4evCu2NGtWAneGCYNcVH/+xU2rIM+qXFpb/
WA19Qi5TUAJHadvQ8oWS2v+hs3RPyHLjuOjZ0tFItLlxiDQ/YcDOcBFslKNH0B/0
+midW3hAHHhAkYV7/IIUAoTQm2G1Xl14oaWC0uc//NQJL0U3Pg1FzyXi84OiUluK
1mM2MfP3092mhekQn4vx/dUp+F5+YzgfdQdGHuyY9mersDoZxu/WskMr+mrGBdV8
Ify9vfyKZYhvSJbPYOo/dA6SFKE5jlpqtTg3p4XgCRaqj6MDfcFyj4uDRoUBAbVl
DaZFebn9xgtOaaAaiEMIp+rTl6zL0UvUym9NY2PyBTw07s2GOlrRa3unuSmzgkCs
6Vh5Y3NqpLw7yvy+tptXOc5vhNOuIUE8YHgnl+L8nYk49kU9mdhkpOgwe+prQs5x
egSWgZ3FN9B6hJ/jCP2+iXi4l1roKZo0t5V7mjabQHqmbJSFn0Vrj3+zGQUp6oKs
YojxxRXngH7Jzlk8zzD9UOBmbSfsZ9Cdk8JCVX8SPpimxkJpQrxYLZQKTZfylJPQ
Fetx6nry3MSFDVpjvHrCpOZlTOzjFiCJ7z2bncSuF8Idzsu/rqp2FmLPFHPH+oLI
rO12uGUkRgGzeZDmduORy4znj3bgIK5mfCe2Emt6tGUYz5xf1c4pgVW8xfnOYuv9
9soH9z5ogQYRKgYXwx28ggEFbdZSuoZZNwRc6f2yEOQmhHOoiXlKqy0ovTL4/afH
61AU1RBIbNUkmXQ7Ivl15lTpbF9d0FulVqFkAj9rtVZIvsdDlPukxF1Otk8qmg8V
t6HkYEqpQ+P5b08FQ2Sv/JH5gZTtXZCTA491rgl11ykdWwh/7GrucbXjXK5Udse5
uSnBjaMuL7sF/HtiP3MlGeQCEMtvx9mZF9gIBB98LjBklzH01Tj2ZlJr9yHXJPHm
7uID9Dkcd0ZiGl60dmq5lsi8QsjDlb/98WMtIy54muNxYD+qpzGyvj9jkxgizKPX
7q8/u6PuhANIAveba61vvXQ3b9iCpygvrvRSLqTgkkpIEq3uG1QQNaJO26daxKX/
+zDaCiC7+1sZ+sVNQ+LpyLTpwLijILDKeYUOg99wkeKUY/TELdd5HYF/3+s+LCWN
OCuVnPX3sTmQi5ycMqqMotPs3+OlECIirRydkkEcxXpeojf0kdfEHO9ZPWmmCRDu
iNSR5ndIbwlTFWPC7eNYGDs6IrVIT5lnK5gV7xmLPUkRsiGY4tD7SRL2WwdZkkEd
rXaQ8ZXUY5mgvMntfwClMseF+YTjfmXni5UHpYOEIbhwVqF8I1ufhvgfOrqLbKnO
RXzlC4webkLQfgLgVvjM7ZSSUwQ0wuZMM6xzKuQ6Ijjq3UWr4EFrtt0HS2l0pwIb
vnj2VVXoQi8Du5HuXfLccx99tZOmGK1HH01VuBHBAnYfeijNaD2Cyknl8Y8ZfBdg
fdMIGcdjqsf4OQ8rqcig6HjCEAxJirWpXVQLEGeejnFZbf+qOw9mzOcOw74whNjl
3ruGs3FXi10Zu1jfP+R9aQ9xhQLE4hGw4L+e1lOcbbbkHeLSxpc/drcSGz1fT9o4
5lthZP3idklfegXv8yJgztP/LwZ9rUZjv6S9o5lTQtBf5bKw5aNElol2T964+c38
z2oLA6B9cPL6tb5B+QXim8tvD9IAfUXPLqxhivfdIWr2KrixHjYTIF7tcJnQpJP5
t4uN/kgKaFowAMjzRWjnAnbO8xoVPRDG2Ci3vbMetqVNkwQv5/UP6L9yAT1SGrLU
3ed7Std49pbQ9InbQuD0kW5DA8oF4KSDDXydo23DboS+9ytJB6UyYRQuVGAj9Ipc
EjsK5B5hFa1eBZ9nB5UGdDI4rO4hoYAXlaEcW2RbWBM3/TiYYDpu0Lc3qpf24u+B
nWonfjsff4JeCQExN5CcD2N04cwwfBzGjJF8/vWxlioaWAHUAvueMquuLLNkrN/g
d3q6MmwMK90+PvG0ilpymIPZ+fv9tlI+xb517Pt4tyQpYZNyKLqdTE5N0C8TCW2p
ZA0+mZgSacWRPAZTTM8a+wHxgZGnvqZxd+GqTqzygntsR7oXONXYHlgB6BLMdT+r
8hGkEuj1vL9mAmi6LFjxQO2iqsnEDFQvFX/XqwbqyR/N5QnbX4X2DydUKwTNHO89
cqhYRogrn26iGyomhlyH6mLr7UgUlf2cwpiX+rOyDQbg4765WXbnoPU9MiQSxIcc
+NdRkOj8qtakb/9U7u6HovFnDX/mwfy1TnqSqUrNEfUsoLfxi35hGXOO8ZsltoAX
kMf3RTvXlMphmJEAsdhzbKvyh5vKGaoJSpO2awRwm2TeXhXC21jqU6WuMgv2c9RU
mJD/k0GJ5fcc4hq9KkIYHhv6ho8FBh0O2raC0BW2mWaP54WWPi+TPoYMO9QT8Wwf
zCJKJ52w7BCNTsMb4rHT5ck22vT0gUNEraiTuH01IEa2iqF9HzTegePzX4uZxJn/
GuuebXcj/MzfnoB9SORy0rcFeUfCfiZpnoRQtBlcXPxXWQAdanntfA+ZLE7K+wsK
gGGUluUxBb1mCO4Dwtu50MGNZvZvhOgfe0WvCkC0aC9nUa9Dz2uMwAgaT+0ZYdjg
c8kVmIEpytfA6znzBm/qN1VgkTurs56fviqWcP9A/M7gbtzq2EIqv3dK92sC543c
Yj7KapQDHkOJ7Dv7IdSDjGmX6NO5tzZie/0KmF6kIut4VMrmpd6Z+lMiAwPJdLPQ
U68UroENZ3bwDtASnaYHoVVY+EUPNssexN9CmkP6FopvZc7XXLVt1++IA6IgmUZb
PNEYe2JF5EXADtjIXG5TokNGi+5EdxLP/IaWwLsAaVGY7VHxDVh+2DsgUgU5imNh
8U2jtOlRrMHyuOFr4IoWYFCD0fSxUz9M/2hiqy8i5jrwfKP8buAF8sarbwV8w8P9
nXN0snYJIyQKnTvq9NWiWDKV0KPxfXbJeqoWUnAUCO2LkX94XmfWEiN/vA4xFXwJ
Brnte+d6u109z4OPkgruq7yJ7Wyxw2COdd/zYYf/QVtnW0sbgzUFG6LlnqXYZTA0
0oXKivOXkR8raILLf9zkonrRXcvlY8sUumIbgH4NBE3OjYWF88Kcyh834oEg4ojY
uX7V7WGo6xXXroCC1i/pT2vXF7LjqcVot+8NyJ0Mfs1JN/0uKEg3X3QD4GlR2/bR
UmlLAofsLzYHrfcvHJqlZJZYv/4rKK6gi22CIJx03dc9QyXUMkQJuFbEmgQ7A3Lr
4D65owNb1BfJ4gxM2dBUllSJS2VIBG9eO8kY0H5Ayx7fYQO7KF9aNngHegDvIlGo
Dl8Lq8A6zoyLDiw5Z9/EboobJu7OaFGWgT+OfWIRUvWITTneBlBlE9shYq7XzYql
Abf2rTZmOUF6G9obXPyNbxurnfahATBaiXKYMloWROhoWO6Tjy1gjhVhsM+7eFmA
gv5dVcddyP8vI8e92RDIx0aL+hLZ00Cue/UNjB+atE+eWQ/pBnp9AeT96PJWbbJO
Pa9K3igxVIDhYCLpujg/VKHTwcXEABTfIzdmw6usyVBQyFch+6wBP3jcDTevvzuE
Buk+u8G+sprGLVPjfC9gxiK8kZNw3S+U/GuwYw3dnlzSUtNXrH5s4tNMaDU4NgMY
kWRpBssW+5xlOjd99rySI51Ij/v7F5Y1fTLbOSWQjy/icrn+zdp6UO6Lhn8slfZ6
Tw9bGvJ4KSYPeBl+D/ev377RIqoAPkgjW3+4WTVKKVEfD3jkZvzXJXk11da0Nm43
DwhAhopYNNtzXdv7vrxEb9o34PNnoMmezLGiYU+SHQXnOhYDEzA9qaptDVQC1f6o
PfcTdTpd7gHrCG+o9IX7A3+qneYDYJD7phG1X1hqPUxgZYorbwpW9QVbiSt0rW2S
42M262rxze3n9B4gx/WPaSq6ScU7HxcpLuwJe5VI4EXSyVrtlECu3sfR28Iu3Td3
rDx1Sun/b7uDvOn57QarDc1AZ/JWz92qxH/G+Jm2HdZwC2llnRaMggU9jeN5CLxd
X6DA2OAe3yzUtKAbRVdjehrlGGRThBCv1EDxRNWLT3ssEveBHknD6L0HUEPo6wwC
Ugv/J47RCGKQbUg2F6XgBH30AR0hezRDCVBhB5OjXAiacmnxspxrtMztuqhyBfcs
xdv/4JPmmBYxv4ayN6gdtB42UJGOPiAb3CudwlTsHJpEaA8SERmzQEr3Zij5gI/b
cMjefajxSUutI0ZPuw3DT3sbpW0r0mEKIQxKQ9xXk8GjXVvhstjWixncXlysoinw
55AduSLjzXk3vfC7HI7cSmlzmjYx++w7ofCv/YmeiLZssfbUTyKAyYV5S6nfMAMA
VVqGCT9MU34uDJez8z3c4GxBdwvbomGIfnt7MWgE19oB+VTVw/Ux7ek9Jpf+HclS
jCp5iKMWgp33RMNMTcXW9QMDYB2YA2RYNk7IXbKz7B67pmVPz1JgXO1MJzrhctoJ
BUYyF6Lv5t8tpK1xegJJfoYNDAndnvd9PUl4LlRXit8grkxeKT/eb1s5a/K7spIx
o/jqk1+ufKkWsU8rmGshH5YbCSaBK3hTB6Y3l02502g/8BbZLWiwxyaXlXXEYiut
jnwtLlaARmzpypEJpNwzYyjUyuQeLSgvgMpC6Hnibg8TCJy0PtE+VeZ4/+IJbkgx
wIdqweOgi1F07BcSf+t/UdInzTpeUhqa075TQrWMCG+wiW+VWi7Aveg59/IcMTrC
tIJmVFdKKkc3PIUqBu9x0nHlgcr0AQJ+ODNSqRsrcDcspGIoifu02j6aPt2tCPLM
VDX3xgsPiaKKfZeM+iZvHlyN6UjzPi7eWg7JxSpNmg0rQ2BjxKluuzqd4CnPBK9E
psmKPePj7k133ZXS0waJqXCZ9mq8Pjq28+Y7NBRgRysXS8reVIIy+hXB04dD9OIR
ppgUdDqxogb3T5CAN9cacJcXaR6Z8wCYCSNQMx17K8jH5ICq3tIUGIT1q7sDhmjo
P7CWQ273LsauD6pQNEqmbg1Hv3IG1NX8UW6tMbdmd0TpvTDw1hxyxHHltsYcPVvE
l5O51l1dLXxa8QMdSI53tKNBZWv8HPd0udEAtGGxkDXwF1viY+A6liMgWXaWoseP
Zp4C6J32PtBcEzkHuYFnGxH2mJ8HcWJF1PVJPECrXfU8E378yRDIM7LvImCOUsEA
MLGtm+bqt7WsZ7dtyjFCKhiwvcyKO1p6D6hFRGV58Rgh1L2+QjN1JvEYCjVLVn2m
T3X1itHanTRNHxsxDJ3mlmX4rt+wgz/3JynYbZYyVeT2uxqz1pXEWMnqY8mQMjEU
EBfm/AJrXD8mF48D7NmfTYDVpxjTSmttvnC1TiDEXN4u1lll4FJbsbRgp7Fz7OA6
5v7IsRX21OAQSXZd8zLQ+VCYm7g2i8QSjBrjgDuHFYUsMImFfHcv4PC7+oo5OqPM
TvGF58VaVKgdu7tqJv7BccXsYN8wFYe0N7d9YR/u0SpvbZSfrUrHBWK1a6rPQma/
W7WpTrjPbvblryrgbtergIC6JyMTgY1i0T292Fbd02fkO1/q+/pH+PGiU3hxFnXX
ujWyghmVIBu4cLjIoijiG772s0PRlCqXivCKo2aFya9J3bX+wrVOjp4VCRmO+p8U
nfuIJA8gBiIOePimDA9sf+LWuiNbI9HtNm0ybpnAWLPQoP0Wp60SxAsrlibC507n
QcA4ewUieJFBIdbiO1zezSPmaL+y1PJXYhKkwLhE/qLigMliGv4ckzvDuEUzeCEh
Q5SmHOR4qKXsi2Pbxf3mDPANSKlzeQ9mLWMiV98ANM0Uy+Q3+Rolwui5598U/ljq
JZD0VK7K2jNjXMGxsfOM9uDBolCRolRWSx59L9AzpZqfS1eLRyp6tqhmQqEC+jtS
7gVImVeZe3OhDuLIN0bHrc1WE97f6oZtEpLS6DjTid5lYXnLeDZCkUEIsdVdkC0M
scbqp5rBTDJsaqORGOczQ0Y1JJ8Ho+bqGQuTYc3Szeahbmm0mxQE8SLWNASRyu9N
xzXG3i7lUvEr3wobGbRc8quWSaEn7nc2j8C7jRVdwiJd84su0ZX5GqlQzCBSQrJi
darGleuqOuWKK8roD1LUWWe4lDvF/dnq0/DDaTN2ztjOW+M4GFcxSCThYeQovyuY
QpUMDMtB5teIyXjS2jh9Dqb66ukFGcQ7l/xjbAmzJ6QnyvomjtoPrUK8bw4W3kxD
oYJOMzG4nnCw6R82RAcrOpixzfpkvD71V06U3as3PfDRq5vy2EKr8srLztgy9Xja
AtX/9jVBjrlCWrzbVF8p9z0xyke+oTKn1f/Dv+J0C7sQLeQJuhMIfQQmL/TE8Jev
s0abUvB57iYP/J88YXos3fN/x/Kua/2kNp9EXdnAjoDS9BTjAaVTHqmoaEiNqHTi
WtnnAtKPlO1WKfhksk13EMDFDUI3ikpNob2RAc4J8fWvXEqO8zEW7LbyEKkVZgQt
whQW1P9HGZsiMJLXBi8R91h+9UKKSzzrJUYhVweslwqsoX2Bv93k4OK3fyBeO3t0
BR94/ElLpsmOBFkT/qNp5Go7EjP2mobi5c7sgliCZIbv6Q2thqQ3erLTm3Lzp6Fh
EXVwsUKjHm3zaldk7VD9hoyvyyBHGVa+kBvysNFABjndnBp3HsoeuxBIr266D/WO
6D7oF2HiAQDss5PDvgXc5FHgGrdx0RmxMsnYdDwXTVRiNkvNkOofYIq+nnoZCtO5
wfAJWI2zZK4UlDE5oC28AbDLuqzo2eMHMW+64/Hzurfq8HLh2V8mqmH7JS0knGzt
NixfBmrky8LK/08veoo3w3XgLihbVAA+3AQBJ2AgcnRfjEiOGnWA724nJkoPiFew
k2Cysq4v107D9V1+iGRhJ0iYSMNoLf/o4FvreC42zYdFf9ZrJEG8NXLguml+R74d
NgC1HVoIo3Ou5gaJKkavZY/mZdKZ8CwlgoAc192Te7nBmD5bQn+Vm0lfHHUAigA6
E2vLPMaAYHhmyh/bxBRRKR3XKrMWaNakpR0ojTIfyfOXrG4gFP+Il97u38q7jUZ1
8FuH3ZZdEAv58Pm11RAdKpEZgjPRxIlvvV6knd03wi5bLkQ+k/LEudN4UV2qxIwf
hA2Jr/ctZdNc2QOy4gJ/XNjTbxii2oeDgls/H4D5Gs9d52L14uBrP17n1blJ8m+U
au0Lgpgfmff2LZhNM05/FIkhpyi947G0cekSLTAwwCXQIBv9XlStl5JedDZFC3kd
9/0GIVzC7mA9FsW/rd4laC2c18lKmvQtzJCFsY1OyvtpmfhMrohke7XamN9cDmHp
dMNZ76EgEd/Ye5sa/oRZs1oEnn46NyjjVMPhVALR4H7MkZ4W6stCER2FHZ48JwUD
tGnly0d8AuMe1w5zjwcMHrFSt348jF+/+2IPX8ys6I5LsQgBniKB9eeQxOb5NqhW
r4Dha2sPLc9S8V6Y1ns8If7yFezoPVqLyZLGZ846t5DUNvVdH6ZH0yjE8vBoPtgH
fZvZAtCzwq2b8lCYVNwszl5enBwgE0dcD6cfE9eSfVv9JipFLr+ueDdf8AOGzPkB
HnUb7Fx99h/pXLg1C9eP1uhc4EtPgDO6sfwPGr++q3U1lH7MbpcsK3xoi3lV+cJa
nEXkM+fJ9epNLgC5U4CIaWYJSfihTMOimC3UaoE07ejv1gadZW8vOXVDaUm1ka+g
WJuahBNcnq/RdUG3uTYePTaWjjAe5mF8PUJHJIA60p02Mr29OfvqHR6DQIrd5wH2
1f7G/WXDd+cNNopE3mDP9umrp5NNy/3oefiYIK67y61Q+oizSEmY7ZwLqwdMkniO
hwaUtYsLmgALIvXYaicUNhIGtbQTspSKauhsMF+GnYjEh88ayqTSfuv7KGuNdDvk
47vWhogy4yl2YUkCc8eRAZOlPA74T+herYuHddRuiVDzm/iFjIeu+R7C0EGQRBoZ
RlKQEvI6Hver55HR6OTjZ8PM62JVFPn+NoZyyZOocUX5M4DcgRhiO27cZDW4qUmZ
WBbFpBcliTLvE9hTqusTWOpUX60biSllFSYdjPr/Lx5limKaGkyUptljrVy5Q2VT
xBKaWEwjiTaNttFSedlw0ZVjeuPSs67OhS5vFZkoH9/0nLS5NcM9tHjos0G2qkwJ
C9/UbZ4OVOM9JqZHQ9TADDhUnwYPk+Fb9IzTHgodixMf6SN9fqlt64G9hxx3yIz0
JhgsBz7dxUctkdsC+zy9OfQ7s68mdp7wp9MYf82MCu1WLDKWrq4+JI6ZlppfUZVn
i/P+uW+kr9dYuf1WBdu10GhMY9KegD/eqAoEmSnPauyhp3b/aDdyKV7jeCaKLjtj
8QLzsPgTrCU9cd23RnuLnyGx+jwu00p+sbBVFovaieqDTs4IzOlUPJRFWtz7ICYT
SAFS5ZcoB2/nW6XAZ7Jg6fPN+nUpkEViYsy4LZoFINhyE9vigfRychlp5hErTokt
ZMF3sh0Zz1+OqK5Ia763qif9Nz+/8vE8NXNftqw7mu9cdEp2pxvL+hJBJqq8JyJC
kLySKO5rmvW/UYEfRKsnngPPtteuKCd1eGtbekQmFR4HmxtdYpqsUFpU2IRlrGyJ
R0vKlOqHKK8EUdwTFoFQRx5sxorJ4yQKsCDCEBgACXLX/L7nlLN6iSH5Mz0/CSnf
M0x/wMPrzr8vOGe3E4XxhOnko4M3FMUDMhq4ujFHcIeLbyng+6f0MJVhgny5RkEH
R+B2JShkQEKCIhVRE9WviiWNsOgYQpnWh/DR6/S4jxAGLzTY3gJ0HXWPXkRxnzbr
wbyCTgqZLBkXD2z/Lc5JMvyOSQcT9ky1muizLjRW8fQo8Eo5VTBSagRON0hgjq0B
zK1qao5AVCqUjfG1F9ZZ7az+d/A53YLPYcqiw7t03dmsQxYdciOhJhHo3grYaZDu
emKCi9/+X5TmZd1dTg1eWe8pgibPeEq/OeYx/jENbntWRJ3nQcZRBBeKo3C941M2
HGefuHRUElC23D8yrEeknk1A/vtE++IuCl14zgq5ji97JFl+EdNSzgv53BgWrW6Z
P/Cg02vsRK09sYLj9f1FUDULs2jYIeRxcsR5jc59YDV82gas0706qyVNCYgEGkLq
Dc99lgjdbBfPcwJG5zFBYe1VX2KIHVTvPHCznZzOBvjSCr3YwfSvztz58V06qvoJ
VhgT/kHgb1nkUVVsIR322UCUfimxHhIvJxtX2Zy8C17T1NjGl4hWmXQ87zI2BTBX
2RtY/BxWAQJ8rWRZwsxySTw7NXbSFqL+r1GHCqKlwwnDXDzCbIt0fBfSAQwh3SuN
UNy0oaXIp81qCn4BXVMHOt1tSUaakhQEly9MQkP7gePvD8vuzcVZfKWbgQSBIWnv
qZzXE5q91YOIK8PI/a4KZg+BaCniGWHujd0tJwAvezB1WYTeIWV1EdXOO7sRwJhn
q6xI5n0vIpth77PyMQOJsSXBLpgRIqBvhdG27jdxNkxcloFkqpGtFogr1hY8uOyY
ZEELo2RYrrimu2OHzDUB2gYR7C9T3cn9Ejc1DtQ/25GQu4eeZcBWwfzynvd4n7eD
zCbGDOM0Y2omS5s1oiDgXn1WnC8KV2/R7qP/evfRrXtD1n0L4FtyNKctEu4YxWqb
FBG8nwC/x0hDQuC/JGXVPbZO/7aXtwNmjNbYGB4/7rE81fxpltwyxvaUdZs1MTwB
7KORfWxqk4c71Sk5eaUnHGGn5fIgjYLWBbK7ZCHoa80JmY5xwVh5diFVZUqkSuYA
WOTt2ySIr/yVrIqBeBUwQBPDaWMYrOyWEraX1YwxFLChlR9/xPGkYGA3aRmGLJsI
+hmQWzvfprRf4k+Ne0HOHd34LP2CosmGDYrq4EnLKVX65KRR9jabzYcdFCiPRRmV
FHUva9ZdIxvlVcIZl51ZJL7Fh6yKxKUgDF75WHHa7VbMN95fHpAm22ZwtfcOavZs
5WFfzfHgAmYriAugzmeH+c8RPckMeIYSzFCRKEsY5xOOLlup9K3MR+5RF79Ifn3V
pAbKQq04pIFeC8b75IH3rOruUe8gSCQRiKfpzYpQK5zDxTXupHFC9UeRsa0dW5BV
37mG50NTE5po3h5IUOcLnQHpvk9BIuSbfhz4gfxXVg2if+/pCOgs2z59luGw60Xk
8w/Jjy88N00/ZL/OWS1ieNWXD6auCDdEiqasUUq1u8RkYg1XBdN4WIAq98k8FihT
ljTREohzs4BmLb2f6FlOXUOegR42e+SgK1RvXLqBw072WJKYxG4TbJzARwjrcynl
xpKcw/BnpC38rNMq16li+WiY1YXKxAqWpZb7nq+m6ghoKA4/c58eKc0Zazv5fZph
hGU/mIUogCFkEPU6WphDL5dg94J6oaKVDVeIPb8Tl2RloEpj1DcjkZCZogd9sV5a
QoioHDJr+AsPnrzdKBQ1e5AeCd1Rr155X5HaEEl1phftUiqU2pUV4PIwSrqZRb9I
X9mv9PxcqwKz6ksLAsYQvfiM1gtFSaXIGl+nW8WMvJc5ZXZTLPbJhO9DRfRZbXyf
nX1JnuyYgwmVlqaLXBWhPsf8sbOE4q+aFG6HNL0TojDOlZlo7Y9o8wkMa+udGARB
CqdQl6i/aiMzflDFBf2+fuqyD2Bf1hwI72sS2uBoP0Ni8Dio9l7ITipQoqAscx1f
QPCFdnkOismHyiburPrnV1igahpODw4uaWtXwAFLxqPRRmNfcxIBn7shVxSl5X2x
0mCiTqOPOAjF59GL2xr72YhxFg7ZFDGehf5M6ZBaDkOI7MVpVTiaV5bPaU47nM+z
Timu5rzYuvssjzG0m+e8Mx3NC9RQBL6w3BxU6o4TborS6TpcbU3oOKok7/44hrxC
rnDJbkj9I9UpTvTTvqGpWi2OQlkJLUodUPLF16aEjr2STvQD/6qm0RRutJsj6PhL
iFkmd1xM+xh+/ETyaiJUbwT76dHAj+fTtS5MtXiKw8eeX1gvlihUlVxPd5fIDGGj
smZEj4gAXiDZ8lTxCzGPSCNMuHVXY1X94WMm0HzXVNcATJr+mtujbXnlElzGLQSj
X3k1tQNO+RkSlT0s3mVTOvakJgq9gNh9BAGYMBejG1+h8ko+Ghb69lPdO71TE68s
J3gt+DEgC6b6fMUJUpGAqd9MSNAMnbJaF5Te5Hq68c39dTin8RjDgkDEipEZxgxD
BfU1BO6I77ockUWz70NZrHTTSOPP363HzWXbxPIXUMsv3PQ64FykmftNT0sMbEJC
ZCNJpRuHPjxU+qtI/28iA9rW492jB+Ldr7iPKSF97OMuH0GUiyC2GANLIPkAqZJc
MhDgCfO+iHw9D0SjF4fF8M9NPOdH4lO46B7wpkgMZKtotAKPgKgfsoUfXImLgnyK
ZlGUP2WNxPsV6vxBVS0Ch7x6Y2YoRHkIIQ2lkRS0wK4EmZEl1itrlLkEjer7294k
u4q0gVcO6Xr+SgUQJvywXnjOQJMoYf13YwwMjXY7l8w63HTGgggwcb3JmDS7+xOh
0KOemjaLMfH0WPnqK/Trc6eGcoJFBldLXGD/VuI0MaKWA1UOhsBbANCPa7iNqWmf
sVlG6HDWsq9Kby/iHbXMOTTnI+RrZGZS1OWC55AVtkZXfu/9YulZD+FUFggWvMEs
pQ4yPgIJT7xN/xPgEISp5HmaNTMDeHesfodOehcJ2eJ1P2z74QX5Y6VC6I2P+Qye
0B37h66p0gvGlaXwI1lar875jkAnlaKHqCXHl8wj+M0Sb+VYg1npy36F7jjZqJNf
SBkJe7u5cK2EqhZ1axj7/5uWMCb0ymYjO4EwTGjU5Bwj+whFQ6RlRPLb4R5FgwH2
qrezKK/76fSIHoDxmLvrGosau1PxvAxVj87+U67f4q3sEdCdEIVYV0RjJQ+BmxJC
yJd0LpkO+oPzqrkbPv8lkT1C1t61m5bqgf/PW++fRWWdv1t2k4AUl+B/k0VVyJZD
EMuuL4mIVBAYZaF3rZBifRJ8t7AK/onUd0kvi5Tjk8FB5rlRrWIxnRVjFRPnCIbZ
dkwbx9poimiYg3vlL+HUNAMgrCoUVQjVJGNQAxhx+X41PgKVTBmzEEtbeCSgyuKD
eBGuUKHPl6WtQ2ICdibycuF8ietvq2675zDKl0AB21tgXU6zzQW0nry3TdLZxI+A
y+JwyeA11hpsuQF3eJdGHTaYgL1i4miMUhY18DqNK/QKtEScjtWKo372YFLhXHo2
dAGQh54usJ1fTvxfSuc9WK2d7iATK+/1GTuWMFSFQd/uwBmg1E4E8OREMQc0hhRE
xd/lCTrBSkZs9RehZfB6kktMblXvDO9D4ftIxKL2woJOI14MfGnzgljTm5e+8++H
V8u00+gNn7IoIV9aoew0KaHZh4sunhdhE4JBd44pKCYkOyaRvs8rFPSaoGn5m+Ge
Ev9FI7xNe7/Ngj2/WGYopkj6BLSkc9L934uML4AIDiM9KdHnM0t01dJlcOKnURRX
nOdB/1gRlV6CS5Ww7ii7EQKg50WWr5SzYOe1xKVBPJ1SOxC+gRe+UvxukLcFIhKi
J9Eq308Lz/CTEA4nARlyuQpTVcYkuuGnEO2/5ZZageE7WEq9PszbcZIZ8UwAdGRj
lm5Lq/7DCP0Yit5tShu07O3dFhmexNSi2JZGRzSKCq4tApfgpyw6NqOAQ3whj/z6
Iy8mLyktJIurdwzBdwU4ftNd0nGtmvr6+eb4dg0tvF/xelh8jo3exBjNEpDBr9kP
su61dpV3lkGklnzCInrMuIq0vyn3F5lNLsT65jkELUprSZNavPegxbRHw1voEh8D
oOT1pd7Dwi67Aeypll7vgsHIDTNrFAvn95hIytptCB9PuoqJ61IyKUXeFnjN2Zmo
KofQejdKIiHfXERqbbXUO2SQdDJscsZJEZBqAPGOXomikyJNK6CBzP7vZSnwDBB0
rEn25ceXbBUAw3bqlRejnH1Dm+F2Yw956PRPvXfzmUKtZWfUS4WeObWxLqrldCbX
DiYd7KSmIydCwHsgglnce9rUH1YhJWPQky7DxdGktb/Ie+9yRp78plErlXsafE5D
tTeYBc0iTJ/A0cLGDEe4yZL92DKPvY2zIhbQQAdrdDgfpk/KLwbs1KpTqjMI8ztV
hJlaOeFDW8HCl18STPCPbzM8ygzL8Dbp4134hdC1kL7ZWZ/jxLEwXrFKkjhRWol7
zFugO2TxTBVXcnrFNmPZ5dcx/j7EFnPCYBXr7SFXP3mQiBe7IbZZOiIMvm+07TdQ
OBZMSBM4BcX0R4IEReXSThlH0SbAc2X0t05JvcZElv+uIGZtreuDjbkoS3zyZzmx
nRxKoYWhLFd/fF87vPM1WHqN8dN21wyRQUDqG9yv7BckFTELPzXNsqWFayEVc000
dglmEUMcD+liS69UMjdPdkj6PskPb+oyBgUq6htMDzviIrsUmWBW9jYuxusP1wpf
/5MG4p6eMyogYqTLUVirZLrkzeVfpnuNrUfa+kEPMrCpqIOUkHMFQNnNaLFbjn0P
bi09SSLTAYaLvceSqbXxiTBT6PJa/UB+6ps4jfACSYUtCQQZvx1rEyza5uikSUVg
5k8R2W73pCEq5BJ7ekFkOl0vgkKnUvvsV9+dq59CQ1UsBdQ75TZ+duZU0rpsqUGL
avSFxRqAsTFvrB4S6ajXmCyY1xYO1x3auFPrI4YfUUfrtomLie2jfpW7cPuDb6Sw
fSpNdfNGFcGOeTFl35244wN8D/CcvRzXq5D2qNt7/TEXxJ9ALM5pvJJjKw4bEj/+
MLZPpLu7gTjtwO/lC67QA3AM2U3Z9M6BdEzByNAGwEU9Yneizfik6JMJgMhIHz5x
zht0Z5sWJlZ83iKdTuDhcLaQ2EufIg5+op6018GM6xdrWxKk4GaLeauN28dJPISA
CAmMSqR4ZDg4GZn+pZoog9ALEpIMlNz1IHcaXZ/VHnMI+S5rQEtfWJwb7nwPLbDn
uNghJJvZnqo34GiJTwWoN5IRNvY1wC+0RVm3w8EvZp3tGUHOgWxX1Bj8apNt2t/a
KtxPElf11IBLqoDKAohFSZ8IirckuvEi3B3yZD3DQyX2ina4Sxvjhq5F7KrQt5E1
Ylup0/fKJzQWxuU2wmR3SFVdZkYiUmDU2NmImy4caN9yxPRQshPXZfeb3beWemt/
UduspgPFfFS5yeav1G346js56yvGvWsuEkdE4Zt6lHUBx6BRYGoN8gLgH9GfHxVB
bPCISKMuwv0xMikaBoL2gyLmeJIQOuVipkH0fahEs737KlgpcNGxApBhKQBjQ11r
ZjOgiiTxXlpNxpZ96E/axQ8/k+pTeDpbYHPIpRhNx4gRhQ9KQ5Od9dAIgSJhXiRt
q+eJklpPLxGFnBnoYArUNxO1DVu6/CgbZaryn5SxKjS2PUISN2JHsm/fhqCHxwmf
Dj0l1P6dVwa1ZQU1ilqJ1+GGDvcMWiScMOst4VeqvdHX4A0uKTKsD28b1YsMvuqo
H36LPQxWENHiV2oZJfn1U/Ar90dRhyw5mfrGaZG/n81fQrKaGItNcmr1xLnnPsRf
O2c7nUvWmaZ50rL/8n9oWBAEfXv4XlHPeSI0JPXy1w6b4iBX6FovhkJqIim8em2F
I2lHj9ApwlpJ3r42bz7pyUSdulbpV+l62lIvRvzcP3faFuePIoaShrfU/2S8rZ0V
amB0lo2FY+m+SHe2lx8MP/T5Rk4W+nxCPg9LqHH9yTi1f/M19aqF0gPH3Ws92i4W
9zvBJvMB7GcQGMFBDs/b2Klm6qjznRRcePxllLRHp4VNcsOLu+a9z/wEqTutiIxw
pM/jN2HxnatMaBfSiLRQXRz5KubINY1I8NtdCw32zuAydX9OnesP4DigfBZA+n/Q
OvYqWhRCG5X/zp2sr1bDFylE4Jz4erJpjVeN6inbMBuxq6hLaec9mFo9TpcnRp87
CwaI1MppjPpiGblhmXnWCls4QEeDAYtuCAw1PGq6UyqgspR5eltbMT33Da3mX0lu
QTqPMJqh+Cz2LoCBTdNe3febGYAkAYzVrwIhoVatHdtJj2Cfw/t7tK2sxW4UEeLo
fV1TnBYP1OfQmMsSkkPPQ1B4329L+AAFrlw8k5OZkxxSqrXAKPqSJ71k4/zlYMST
v4JqZslqgEnfAaBiZvYLUn0iPA+AowJebyFwdyjXjvJx15l5rcu5oM1FtbxQQR0J
u/e9vpA/yo+vp+mBxsedylmwKCIS+FEhp5N2pt4HOM3yPp6FU5r23A5WkMZvbpFw
FvV0E2cDkQCDEkeukjbdS8MhIAmJLOTXuMKYxrEm1DNCVZlu9dp5OSxYM89RrrZv
ERRnODSkeiQNM6UMQ/d8ixVq1chAYN4R4IRWS5Dmo+hEs/J2BGxG88M/cZeYa22E
jJu20fdciTKaL5kB09L41W/ZcFtPUhUGnwF588OlMcmmF+nqJOBLeDPV7Ga2PJ9l
GQyD0CL9MkDGY320jkeU9UOqj20hvOzqk5mcYe77pXokYH2yErog++IYrZqkHgx4
SbZLgVAQBWwgLrGGvkq49vjWbjFlpw34ik07DnzsvWosQHpbGjrXAgkCTZtOPATR
lSgVsJXgGD+6gNWWUChpOH9eOYItDIPPeemnotWmdPWtvLslSbtew5YTfRmDWZH5
CM9uzkUsuRYc6duRkuy2nI67DGAVcLJKj7kEyN6wO0JW2mKs4DMkEoKY0lgVWJ1t
FBDj2heXgqGqt21RdmLLk4nSM+aR7BROsywDlTFXLoCrdzqzlgPxF5AQ3UX7b/VF
64opXw/TGLyYW8lgjCFG1qjTFqKTsBUoG3kAZFMs+rlI7bVzS0+ZHpjG7YDaipFf
36/HOgl6dLTZqO2PVvuo2+Yv6EdfGse5OOmkDxwwpol/J9DMYxorGg9FPA+BiEBf
m7luwKSweBdXoODY5PnJrEtzlzIQppD1kZ1fA4hR554QsURHgqJXe4paglfvcuFO
p3WvvAHrNEtMRBHjp6wuB5aWMf6JILq9sLv+zXWRvE/A2yany0k0avdp6vMGPf/5
XUfE3r2b7lz1yYg1pZzCKGN+FSpqW+MJYlYNzE/t/N5cBjlsdfcJC9BsvrxUYN16
k3KzsT4wHcTXLoJMApnBFfW9kGDB4PRAZUUHWUgWsjP5BYB7ita6t1zL12RrFLZR
/81BZW4oPaE38gQ3atjeLoYDEumdxBVkxBFo+vbNiOSEevIxhfP9E8smH6Mq4qsI
sWhVVeftCUvx81aTpayXCtYLOIivOIS0M3hxO33I5mUj8M2j6YmRzRgknTgKGoKn
ge1oU3TjJ7ilw6iSM0LQS+O/b5fUfYqp4mZcW5ZFxiLdXR/c+N27ZI0OB3GsfNPr
1GqUgNKKpT8O5Vh2+7/nT20KvJvvrrNDloPCdWegtpn1seylhaKSvHp4M2uY+BvC
LNqAh8djFqWHP1VLjXyJlq/uXfgACY8JKsyp6BsKVllo1fPcxzq4C+aUPtewrq3H
82OeRVRKBQwSBp63yGxt6yKnEixJt3phTULjALRhrRCg9QYyVmDJIKpuf8d4kEJ+
Ltr8+PzWG144j8fGcPNn0HHee4Fvv0ZwTx95PhiEQKtlaKugCeGRJItpRtjKrg3j
W1zHdcLx7ElMqfXU8AkMeK1/D67C+urkWq34KAGghR0EUJpGCVFH/9YP0GE9/uqJ
5qJvKePYDqyJaJFKkypFpzO1qaNDnrcnbJsrEk16Kz6Ku2MCGJaICopTmdF7/4WJ
ehq2YgxkQQ/suycG98LFvW0n670letbWREgyxvXoKaKjM6WtTFGwxSNPq3BJlKVR
qO8yI4ofLlJsp0hCOQaqfyGmAt4mm47aMUtnUNT3kyIwKiO0Jd7Mn30/EdC4uM+B
qpC09oQQp9ECul1lvMz5gr/Wm2QHwOkBfF8iLft+uhXbHZG8+DRC9rba+ZMWHB8c
dgdBWCgokfpKVQuOrliv+YupoD/9TaCYOjOgxG/SemQ=
`pragma protect end_protected
