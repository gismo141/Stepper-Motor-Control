// (C) 2001-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip, Riviera-PRO 2011.10.82"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC08_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64")
SULBB4yIHzMYvO5D1oUHcYOSgnoJW8tMlhMI9Dw0HCg0sYYFMRFh32hYNjZPvgXyxMrqUhf5o/Km
7s481yhaKGlfeMGcdDHT8JbLv+t9ghKEzjwc8pWtNeP6BiPosok2eVqJSKR6etAhrOCJXXP+AaFQ
Km+NBOP7bPKg9Yk7zuWDoKQUnEA0++HNlLlLl3x3J8aZO0s37hKsA4JzC976e/ng9s1PixJh4qtX
nBASAf0/5fkVPvIVizT/trvTX/wFdJE1O6hweQ5FmmbiL0uV0UV3oHDv+WgUwaGjhhXvi/abBXV9
bHcPkhMYQB+ciluwtPnUUzHUWH60RBanKRFA3Q==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_method= "aes128-cbc"
`pragma protect data_block encoding= (enctype="base64")
Y6ztvdvli9nBiBtgwfdKv925hfaqopb73Z6hlxOFder+8A5YUvc5tyZFrXHTmS+sSeabL30M14J1
t3uZb/77iZ8yxL9GH0df0WU8GWZdbotVgViKGzKFxD3A6HCo6Ww4K0Jn5NxRiqbv2A9LQBwj/qDL
pX+BRv+e4knCMEahQb5OkcQyEhCkiTIcVRSe7/tAHfFzt1hLYfX9LINigHhfxYb2FvhuD1qoAV4H
sHj7PU7krP6CgsHzSG7yRs7Wdln9p6CbdHelbYNuv6htqC3gnQ2vQfnr/B+WV2qJicgxaQ1Ht9Z0
9Oquirllc1fRxumlshajGzX/wGDJpCUzM1yTWBrRCrDIlBgguCq1ztpZe6Th3N/klLxGbvPK1nYu
pVFg7bFwAKjoYZG0Ji+FrtX+iO2Ww3O6qJWahDadn6IZoA7Ydg5NXhPTVWl6N0MEdwf8eBCV9iFH
8MwmPxxERdgNON/b3kJOJSnVYoeU/GLbJpsZNo7u7+lcE1ERd8xorLo7PBnd9lZVvyozS/3IehXB
YqYl0H26D9u0VbKxnGyaZmsZFS0RBwxz8/wGVfAcS2NGBNfKvUF+qxTT1MkexniL7roLvOv15+1W
28i/+/yxQuMmJitbCXbFkT4XHg4sXSZt2rmVHsnTHsafyG+LLM0Qee1QWuJPdL8YcG/hLgbdNcs3
42KOF3CJcMXdljBs6GezAy4vgI6RaUdqEBZMmbprv2RLlufqrmlwa/ZYVkFGdugZEvpvARtqwLsD
fdfZzwvXHCZe9plh/szmClPvNnwrES3w7SoFlFoAJK9h/t5ETMGcEPy0tufcW/65Hx0KEU4OCeYF
gYMwBJYn1XZ+HNcoeyD4FaifThxzAvpY6W/V3J/2ABenUf0Vl1tCv3kthsoTWwb9sM0BABgwEGSb
tnSQBoTd7MDLRsbfSFGQl4ztFb0wLlvjHJNbA/fHqzK7P+x20XsWEcvRDiGb9DVwk9cP3cRriBE9
YTFfIud4O776Ra7gc5mU10Bbh6wBjh8/7LSF+PCg65wwFnoYr4IZd6OyITCbcGjLcGlFVXx4ucOF
Ikfho/OGdmm0Sf+xtgvj/z0qPuF43QltSB6BqMgvbCgrTajUwYr4d8RRMCsMIulT8KjkineWwQCT
fjTkTx27HM2sueV5Ba6Lr2QF3bAv1+ca1RX4YWoHxc6k9qYBfb3Ki+6U4W5xrN8yYvlY5lnaIvl+
TmLGBqhQCBsvNZ5GJIpcgnO9zWd/f7ZGJAUtqajTiyoEqv162Rp4uZK+UUkBKtnK06UI995huVhk
41VAmMa7UrvGwq7J3Sn8r0OjSXi2MoYtk9CnT0v70DIHgV3nUiIyj6qrJDkhac+0pvIKA3Yy8os8
D08RhoOI7u3mqaVJdcNLR/1FiJrVcl2faNzbcejtICQnmcQJx6mRdJwUk9G1SA2LuTcY9SkzIZ3k
6YjkffCWtJdqpYq2Lc3Lv19Gd7ZPk1iIs1ELos8f/FH1GxtdPleQMv3MKtF8u4omI5gu1ilRlJ7s
0pEc/Rl4NJqLIiBiCiyEAqO87sbD6CSsBLVDFfpIV2ES4pjUBwCeXSV5HdlwugHUNpqvxx6j5VUd
MYZglgKHwLkCDkX9fUeQzEGMRywbkYV4QU5cig+1ooNL0dA/ZP7nmCEQZY5VlpOqufs2Ici2viYz
H9UpVhzcStp94CRL34ww4bOiGW7Gyv9+sfzoaeA1fxzmi2YS9WLHVGeb/AZiDcK4HBBR7yGYcQ0Y
r6MmzeqfwXYrwwtr0uT1MK1MRW4RbOJ2rlNG8EJLmfr69ey8//3MH1D4k6+rqn3vocuciCr26YLT
pnTMoftSC6DFIJR5exkB5Xc6KrQzgdE74PEKG3QfJFwt4iKXIYE61eegehCMShJmPqiEApkcjX3X
1G15bBUOx2ukbK2js7sn+TgWzxUDGcpPejXioM2yP5+46cEs4l894aiakqSzl7Bms0OlJvCgQZb8
SMj5xkbs3CO5ADJ4J1Ovu4jCLYjY3iUXP5XRcASqmdsjGMGskdy1o3yF2kjw1r3gMge52jze7Gzw
mQSsSGWVTR6PRA3JvkKrUpXfeu/GT4gBuxWqAl5frwAz+OKdKJSGOu2qnSpyS/2Ng/BYtXReP0GM
LkJs3jIV3PqtUNkTTMzX8Gt74mIDkQbsbZBo4cqiyWVLvAuyQEi6JmGPvtnKZ1AyGF+MkE+/3oQy
YIrUOXfu5Vgu0e5t1BPcXcoDVt3Xvwefa/pkbXlnan3ACjLINf/hETivRdTr8+8RdjOI5nW4qgVR
DnNm9qvCGvQz0z+Rx07GI7a6w5d4m6e4ost/p9iUjfqKBY7lJQLbmADLxaZBq/WWFPHcxIxmeZls
quW25kzhKsSW1mgj3IKU/jq3+vDIuvtzceI/p+CcCZN++GihdphQMr/uHBgnkstU1iER7tQYAJJv
IvBb1RRTBGEWBjtYY6w7WTtQls11WpKau7kHjQ5NW4+f8F5MNQVEOegjQn4cPu34ImlsEkfu5V6v
qgcWNd+MDlQEJEudUQsudKspKzdccEkslUIAklXgAFeQYn4hv0twQ9RxKTAC0wr5BQ69SZzVq1tP
cDTMRpW6FBYiKIRm/VIzTchOctxMM1S9vSjzBD/3JQHmYUZvPVbs1QZc/MFs/99nF7z3Hn31NvfX
2ILmPkncKUn9WooD8Ca53C5M5KcYYIFql/+8v9H/Zsce0wacw61Vucd54ZlZrONlvvkgr1pgZM+m
bd5CeRDsb5TB1z8BQvXv/0st2ms5TKq3CFE2TMff892gNrgmE/AhVyUPskhLYmMAPiVY0sIqBjZK
NMMfABboSoDJVMwDLYcqdrW99CSDhyCl+Bv3wP+sihNhxDmD4JX6CJO1SRVSn93fG7o61uhbSaR1
pQMwNX/5LgM1mPwu3wUZAIdNCE4fkeJ1HZ2YkKAbCv9ZJs8mtGcFSEwLGje/b+N189QwxtBTQGqt
8+Fxcce0qZm6/wD5hSOpddmfDI+sdIojQ8lfPQMjWIaJiTADuccmPa3PHy7/9mmsfzj3xMMZzJv3
8CE9stqKdQoDy4p1zVUlGMju67u8Ql06LYfrd+/sFXJkgYjf5Xf5tsEhkd+X+oBCS1stT2+Nt9qi
q78NOCR3KrWxK2na67wSrBwj5TH8uDkpDkkPOLb0C+MN40GMABGfESukLKf5ilwASl2jSsHK1qJf
hpNzQHlqmj60/E98L+2gRFWjHPJg+PtyMyhoOii73XSwK5oM128sHLhdFC+P299vCs3zsjJdsoqK
PwHuTM3fuf4ZaT/flQm1uR9aK/sn+E+/PBGzYyNcsOOuRxIuc779acEk5JxhMrYOZbwz0YMcaF2s
GJ8777qES5cyIX1y+Jf18i0OCT4CwkkMtwgqO0llzeE09QaJ5p7RiLhDzj3t5QOtHPvjy7XLisZx
gsECOM90ccyiVKYp71QDg2wRxOx1M6tgIEZDrz8kJ/3320A76qToQtjIibmZBnNYLKG3oyd/yAzq
dLqiIDfpPw0bUJq6g8SfQtQkGR4qPPky+cZCo5sKkh15aXDeasLItVJbjOHkRe475Ce/rqED+Biu
smPg1aC7nSkHX96ristqrpXtDs+NeWUKsy/HrPEiLWoRCzhDmqd+zZwKpIT7UpoJ0ePRhNvZzKjn
EQZSq4rAZ3lCI6xezwnZwkBj8sPzWxS8QdrnqnIyIyPQ7MFPetO+4hFmksFB6oc726socJdQAQkJ
gWPFtmSjVjD3x/P6ASi+MFcskwr7+/vijSSQyWRRsk/BxxEWZgY4ouV8aMvvPRDWRbI0kl/QyBgK
DTG/b4DKQWiST+15Ar5Dkx43rXQnSRKh2XNo2jOAa40qlykWOAMW+bC+9KcYHfr0pfe6eOUhC52U
wTDYJ7aeiAdYfBLzvbCxHKV339lWZoqb9CiVYno+Hf9ailwesGA9+ls9OE+iiQeXCeXvXAmXNR9A
GguF4hZVRs1j1fNtzf0lFmXVNE79I0/cJGHnrW5kZ7JwcC341OeeSTL394onUjHKMNQbPXkZ92EK
qEclcDXg0kqFCUY56742V030WFvq6z1QC9ZnI2ZbqhOCT39w5JQf/zEPjvP76W69l0+rI3yq6O/h
iJyFDJXOQTedjL8TrKB8ctLlNvExAtlGIGkSv5XS6hd7LgOfZpnj+0EXubm57mD4mvhahrDVLZLp
+Rl3IgLhojl8/xWmnF6wZwGnFM0khGJggToxc+mVsTIUkuhEtL9DE6cvp0ugKHG8qgB4ZKOg0TZW
LzdCM0d18r2y23aCd+G34hcqlet+OBwQr4r3DsJR9j7QA7iXJAQXUKxcooTBk2zcF9WPXbG+alHI
aksoTu0ZbZ0kMAXe9+n3GCMvU+Dwz9wcbbQfas+7Dedcrb4bI6ZoUvu7LIhFDEvIR1LTgRxmxy4H
OQA/Rkv5MXYeYcGJ4hLj0yNImjaSyTqAdllPyAQLrBTffMs3LMjvc6lPD6IqXJKMZcck9/g516kb
W9lQtc171/bQGRaJCekGbe4z/EY9OUXc04GsfeBNSl7YA0hXvPv+pF5NxVTQu7H0c5NMgD+YpSps
KH1VKkdrpESeohPRBykSgVE0Rv5fVV/pJiX5YpwKI+q5iNwn8Hb6fYWtHI3+vzgliSjo/yUPdDjw
97yQrZO0yA0alnI3p4mOirY1KMrJHF22+iUuv5OzzqVZZEorZNWYZGoDNUaJgEbx8Fiz8k/LcmeY
TDBCap1UMXQkGwK3ygln/vEEFiMIw90RLGrUlpMte476rkxxD9WOwO/LJcnx2hfVZL23YXIJDpBz
YmTm0eP1ZWW7cfje77RxFrZ4vDjXM0zPMuNLAr7du1QrQ3UN1jg4RWKwg7PEqcF1eRCpSPxwiWTg
HhigeFYC91lMA2cd/36f3COVtiqgMW+mLJLZRiCiU3qL9p2a+UeEjxZ7cqN/f4Qi12mynvmLXQRP
XwUqj2JB+sGaapDKUSDA37BV+csOSFHlja1W9BlEmMtyqZOVha7Rje2g2TX/Ra772bsO8IO8tcan
g2xsIgESWokj+4gHiBx90aYyNiR2xAR6/yEJc2OqSfP0NvFZQ3vlho2/TT3yA/Lg8F30NqkxQd2o
wxyek2SfwylpT8hvtqk+IdPkzXfQcZcUFra0oiLeC4Ez1mwx/7Vd7Aok/J+XGTMillr42QgMTeGe
j1I3xMTInGaExFezvSlC6JT+wILczv58vcMqfYUJPXbcqO8IgzoqrA+g5l4pkQz1OalaXvRiOwb/
ml/GJJzBjWZinkl9lDUayajT1H7LMpif/eg72Sy5UOnYOEHjvc5Hjpy13lO9vI6D6LBrPu+6PdFP
Q8lEJfQHf0hNLppNXuzoWQ9agLE2FwTb22U9rEaqzanx3mjzhm35ah3HnzzdhstIlgnx4ZBSPqZs
T5goR4yOv0YCKZN4PdtZhdlY2LlBhqQzorvibMRjypvlSSVVamWoRe5QWA6zAkd6yYwFvoDyJDPH
ZBtGphBUtwWtRQr4cpZB2fE5vEinuXQleqppJMHMvyTmHiVArh6xykt2p7G3OmVOE+eq0MJXD3N+
dkRcw6uvADe4AEtGOM3/zbUkXW8qxlDtxTLYBUaWOfk9oTv3ejuivlep82quEIWIggeYQBvz4c8F
VWx56fko1Jso6bGt/3qrKxengwMMFgZ48GRdDURQtUEOPyAVyBce0YA7enrj2WQX4e7WPJa/xEmt
+ULJGpmR9Ii8Yo3YNQvYvXVM5CMoQQCcUstpE5VLIqQme+Yu+2iL3uVkq4zIGOVcp9PNHOL3aU9O
e/p5YpJXcRYfPzubqqrGmGZsmc1eJI/bbLqMASu15nQVGdoLTnxKHuv7aCiEf3QR4VpBBGg2B6JF
Hqx2DtcpMYDl3LhHft4gqjVwyXMnsW89bE6Nu5o2NfeejE5YbSWdXi/gSiZkzGcGqZYNRIlIoySq
Yes54TAwPGDFdn+vGZ9/FGwjvuWNIOqe39dRFwGZCuLEiST+OB4qcRDGqP9SYkBL0E5HuKOABcOj
m1uRj7qmrcKxs3tj545rqEMtZHBDTpHiWoK6wC5D/BGAijtV/RMhWrx3nHia/Rw789bxrEonQQ4d
a1Yro9q4C/S3yQIYHrPh47uT4ZT8EKNhBbq50l+KqiWfPJYiKWqALDocoq4gsEhWpUrExDXqhGBt
lOgmQ7srRl8cowzAVV5kyBE3g8vT1nSF4KNYztrG2Zk/MyGcSBSPE1+zGAUsGfwP6dBT0Jn6H9vK
1Aq7a4spCnIm7APGCjFchvL/lGX/QSxAmavMVollWcc1WyrLBkoDEjhrpzxdJQ67ldsddhlbpN5w
Me4YwWgf7OGz6dCpqnyYoMKoVxRk8/YBJjd/ffBiEg8wY74o8vh7ynmLd4eDzleMqN99Qq55Gc94
wprhSDSDI/is3XVe80LJbgZYf2qAPyuLfwW8nztTfgxc7k5jE+jbNlBnvwCOghor4/d5RxkImTur
asepiDgOdr9+PjkkIILIcuBZoPZLTv7gKhEoR2oCl7F7KT3Rvp3XiqMyOgwSAO44s2m6G8PMynHA
4Mu9pHUza7T6AnxWOOPFir2dwtMcFrrJkyTzB+9ubsS/Jo2WijkxpirPaaPzgEsPurgyWCy6zBKX
3EutLJNbSlHpQv2RgWM0+Rm5l0Jk4tYyXVYErvpaDUgZhOu4W7B/R3WizWAmeBByIZzQ4yckgyFe
r6FjIJuvRLhkq6Be/Fn0oJ2DVThxvSxvKh9oHC3op76S+f9X0x8P1JnKXiktOYT+Pe2bWj9EmCYp
NwnL12aKkBhaS0ZHMTOOh2+iYUfOtNnsESJjHIHaM+NvDBpl9oY/KdJAm5yTVMuUgxXss7+KJkmf
jF6CA5FfaDHC6dFXYo8IFVuYJlmu6RBC4YWkIKO+LVfH2rO7fqrBB2ZbapiyCbYtC/hGXtryL+wM
ekoSfao6UEtNh8Pax3fSTjXHTdHMasvA09gLkR0SOnH9jatPV4/w0sBNTV2C/0/pC3/RNETNnn11
CQ2yzVmFM1T9MvdSTrn9zyhsiRYzUJCBOMgIk0zB9ebebMs9RqLzalNJtrfjv0YwQzdeOVRrDF/6
z5U4dV/d2EkgJ0p9coaGgPnR9W925pzYeEzIoBuUdR3jOA+6DJTa5kQjc0H6VElCarH7VpIUbEnn
2CUl3KqCJytbZcd9VyPjXf/szr3dsn5cr1Fuu3bNr0/ClxvkMewX0Bbn2BKBpYVoTH/uCxjgBiuf
0eXTYWysStmINHZNTvSxVCPkdJ2TYdRdCgTzcBgJMBL2tWIzEdO48cyOmIZLR3Z2XquEgBxgUkmC
kX+QQsO2ab0o0sL8T4R6Ovhp10/Q7muujh1z+pNClaFuPX/PHUc9MH+KDR6XodSHV4CUIaBMvNDC
UW2w5HW9Osxujfb0AIYTQW5HbjfjDIZRRocd2unkQBhK4c3lIybp9mGX2YL1pPvWCUcuH5NwjVWG
dfovf0gAPrNWxEoVN8hQNrVVg1nRNttNYmz9E/mHaZ2uFwm2uyacbXvaoLAElqwCvWSQMG6QRaoK
k11g+5IP1gBQzCTzPm4Nib2Uiyntt5armFb+LF1GtIJ3BjHhGSHo1Y+/UH4ptsr3x5ThIKKNh3Zg
8msOgokmQrWBldbsHb0Gk90STeWrevUTHdlqSWZQ0fLTfMG5Op/DN1sD8GZi749Cd2Avk4AmiSaG
OjzQk+vkMV1DBGJOxhOSqm2bmWGdzhWMS3kLieVcetIHa30GgyRnAfpGJ5GbYBPs5ozi28uIqj0z
3LatP9Abr3RJrwygz70cIo8xDPWbcRbC7uRVb/6b07b8CFJRFf6eGv1uJpWR/uPAAW07Ict5/sWm
hEfqeag8MKYwuKMF8TnOGwOcgtX76x5tT7dioHT6IJkty7ZUK/ANQzgG9tb6Ba4Q8TPqO4AgNNKv
D0Fi886WPbYavGc4zltXfdvcrO3J5lqmNG/iouV/yjIskpsXRf08vo6DMW5M3XthECgM0gxHUGMf
ntjo9v5jhUumZShiX7JGTY3MXyPjhrn6hWjNRNPyUyc57dexm2ul1GmvJUadUS9xaojREHKdu4m4
4VOEqW71AI17Ln1YRpexA6RPcf4vhIhIJpt/Fu49ovFQxQkrg0mOZtpv6othG7PyZn9XMUhIcFdS
zMqLSFyT5gy6dsuw+K1079RCDaMFw/SsyF5uEJ6P/XdMDbRUQGtRywHDS/fkkuKwYbAf+Vl/KTX2
sFb7aNI4h/TezdhyQByi6efX+gWDL+LCabFFMoB+sZVYOdIvMLi4OfjePN9jrSV1Ewt0exkcTZxl
JG5NjcAR47OZsSo3ri23Y5eHyq07O+CwQArqvQFofU3i1WxyStp9zWTbHQO6EXr4sVmjjiEHeGB3
QPBNAPlHbqGK4gxCGWZZO1pHR3Sf5utQo28v4IKvGlYImwkzTfqimuAOhuTB0MEqIeKpMmN0Rcl+
DUdXbc5kc8ShJeP5pBj/DJLxrl6fIrwtWOgJeUODVPnZRsujKSUM5E14hctBSNdegW0CHqzHGQU1
0YlBt1wx8LK37WcYl3gz10IIxl1IVxpvCeIC4uG0t00ngLPScgLsLc1rs4kUfH6LOOnpxIYC8Z4G
NITCsAukUBLXV70x6kwlP5jvW2icHBOE1jIqDdTAkQFnMpE/PrtUKxS3azlgHrNIIsYWzz1Tfjbf
0oO+kflD5k9QNjUDp6iuyJjg9vsjq/9LpolY9O/6gRmErWsk0IicAEfu0Uq+kRfcZbfYdd9J5u2P
Qo93wKprukl2HqPAQUQa5MrlXlRaipZ0XFHFkzOq+4OstTDJSO1Rxvl8/APEbbOEkpex06Fe4TFh
XUa9B2wtwy38b5Id13XJg074XXyIsQ9lbbpb0pRYm7J45KmkjKKUt57VL+HfpIBFEPNO0de7veTH
yJe3sz+Iy9x6XFi36I01fUwZkQiYCUpYjKmm2DOKi00hfwpGdEL0yo2qbFORhReExripC6g80LtQ
t1Od9Is7hM/BetARkg5nX8oKNu/liZ9xV3tXkiTZVXilUWqqk8q6//vhNt7/V7l2Hx3ue3+Y8f0Y
nRn5YqN6jb/zTlQurJqusmyfUqIOs1nluYGLO8kFVwZ4T6lvRYL7ck831qwlS3IlSnE4eQ/6gDfj
BQqgfHJNjwaVnnPymCCHg690KXRuHzwYBxYFrpQ5g9wGsak88IQjJAAWyATV0THd66ODrRyIt2FT
MBXleH5xUAKVcY4MYzsb+U+F0XI1+xhEpEElhrpT2Th+kBLnEBcDta7I7t40IJHGT2lBWo+hTt/T
Jq8dEg8YJVBdKQFUS77xSFJVgPJhRoTcIDlebqyP4HD9R1BMttyiMb+QEpRktmDUiTRal5AURRdQ
1DRCdSLii5GAIFkX4t8fu+1PM93Jdh4ffbFF/awRpt6CdqYz4u6TxZjSRSOqCs2HAFvkMuQXaoKz
c3zzM3M6AbraxvrBY+gk/owxqDoqzjudU5n578xEedPfGHavcED0AzwqbgluEhShp9ZtX3AwFcNU
uD0wY7g+cY1ACpyk2TR4J8Ru/7CQfHf5jTHMBPBH0cy+I04My7vN05xsTLpzYS9Gc5nDMn0zcTbh
Yx1RE4TTTq5Oq/zUZrlin/BD9VgnWY9MSqkWbC23g1ktsDKeGsaEm4nfc7WLk6Uc/kaQRqEzCtWd
VDGDaW4dAJrSH2NQ0ttqfOqheN+cyH0/Lv1EDdIXE2CcikfW1JhXlxBGs5I0bsZCQopRrLbcj+V7
rk3fKdR8spv/l2KYwWt+VvrHa491y1Lqbm43+Bghzsf7HBaLp1Mcsdc8Pxr2ivsPNmEVTJzPSlW9
/qug2edU3KRalhYXyjWtDKO8e+SwQOQFbfiylM34nwdwv0jISVE0C+mrt3uynr92J1umGSNhoDcX
LtlnWX0i+H/7Z7DDov1rjMv2eLis964oMC7tIzdqQAuiD3G3bsrgeZmTwublmKMinTVb1iVkZnmT
4b6DeLdUfZ9Hc6FuY/h725rvTQEsY+wj+pFJbdj4XR6fshk9N3rlAQRJU63bFd8rved8v98rD4Ey
IaLTaKeEEtC8R0dyZH1sbt6Kx/UZAHECruX9n2WEsRAhPVdryzDUmaqApYorYEzhwkiogA32HmbR
RFx1MrsYFNv0+MgKOqorxaNLOS7Lx9VL9IVyme802zJltMBTxmvDlVe1u9On3CB7LCzb3w49BlbU
RqOnKUZEgYw8Rv/1UvNSbX8WrjzBV2h2NwPPdc62MzUklVD9wQ7qE1U1OT8AvJ7d0gv9LFO4jx/U
tX3rw01oGv8KWQlxMbXzNqBh5q5WQBl2VPSNq0n00H/znoXgk/YAv+IjejRabIAbAXGuUn5ZR9Y9
HlVDnXgE7zxl3aAUGgwYYQUqhXnSRjGWiPjlAUj25HCY3rRoAJ14xYoykiyKGK94tysAbuc+PsUI
d+5snfeQoRnBrSr27wz5RZUDM3/ucT+3chbZT/l4DfFdadl/Tg2YvXjxb01vAASHgwvrlvq8ntPZ
JgwLm6wYWSiMBD6jdnDeMpBB6zGCEozBqfwGoi4unHkjDSUZ9EgUScLgJF/MLNEVlx77uRbbZW4A
4/NlQDuGMXW+5pqfkeECJc+2ZFI6BE8ObhEapY93DID2YA1+U3dlHW0ECMS3jes8QsxN4WG1BihE
0Xj1msvytNTQO+ELDGZJv3N9gByDFiZl3CadUA1ini77Mkz5DpiXH03sw2+bxYT49JJs0Icwfzjs
iUXbv94Fa7GZLD0HxdTvKDbdWHCkma+brA0dzxK7ZwlM6NYGXNb5ClBi/Xvbx6LdxyDBO7XMYndo
HRX4RJ7l1i5fImW4f6qr3NSq70Fh2lmuCd/QDNd/7FbYJ2kPYjqyCwTsx8w1HQoSlPqQiH9EUwY8
quXdWHdXm2HEYs5UeHCFS8iLcvHYMo/u8/C1hFd1c97VYz1NTH+jH4EgajO5Lhg0+qflmd6a4hLT
pTZEIZR0kG0O8pySZ+4xPQk7TM30TVA1YFijTwoy0DykCe6Tg3uq8sPDAZ5FVmGhW/JRPWo/n+OE
1yTfXusFIqfygl4KJDjFQIHG4nIq900q0yRMV9heDJyKRLYFROsGKhSfVHemhIPqLhL3gonoJruE
mN5JoNrs0I4lZ83JNwN40kaMkx0dQc27quhjSrlJRRCztfttUBjKn0M0GXpwF7RdsuhMdL8uzPkt
5GEeh6rfZSnM8pqLoBZozxBXOPhMRII1purazznobWHyGtEHwzu73mDSZHHSCZnE9bdzA+RBQm4n
5RyZUPh+mhjfvTHB6eCyirNzsXP4roWcU49D3scwU0fUseHgRgtePD8Go/g1QSxfxCupPvykiI+V
l2tIkzb7Yj5Xk59G0lbw3hf6tcLRMt60HbxtRhJhMMWyxYfQvYzLNaOcJZ31UJc3FTL+J37urkCs
AHL5SJrTSJsTEZdYJrt76v/7WqFJFQHix/x9QDQsLKUb4r+fbN0LLO+UZeX7Uj8Z2Gu7tk4b6IUk
2bgTX9jTP3UPIeAYy/mmt4beM4ok/Zn7eHOnAHCivXcgYXo+0S/phqiWK9zW7u737xJo6s1wcdY5
hgcv28HiRl+SIuQcZBLxIFl1YcVII3mBKzP7Dgg/fq+2Od8Iq9aRVludb/a2s26ifvGASB1ICv8M
9WB9QMIjFs8SQtkAyr3NROWx/AJkHWTi53ulJ0JrqodNDezWCjWS2zZsGsfrGEAARROfYXt6/ok8
bOAubR6BQXrl17xZk5My7zmkRExAu+nsMhi7zi0mzb08q8NS2wBKiiQ2VDjOhgePkusur8vIefCH
emJ/FXVgdkZiaWZWnd9KtYPCyl4KPGSl+W+a4eR8FHkbmzz4cADm0mN1TuUJ03MAbcRjGxXVT4YI
nTDvx6ZGW91eOj+Jeba2sOCHqvgoQzH2y8739B/Ox6e3a8g419LPs6tr/2G8ZWUxpV9ClQul5YmJ
mm4fxXK3sazKj8X7H+QbzXwIUfVpJGa5ozHWlCVfSn7NRsGPIhK2nnmqkrIxA7kPIyVP27AwsMJu
cGzDGXzAiQKrx0CK+SP1v+9l23zmkxZoZiWkDlvpK9MdmocTaMLe6zMbhF4oF5ivh8GdObd5JRQ6
SGr5IZs/DQRg8Y6kM/fi39vge074R6/HKYPzwl5YMtAPlwuqs5aciAx8KFtFsKy9/brOP5m+gwTD
PCL1NGr7tgCCbe8Gv3FO//WGLZ+GlJWV80cXA1x/v3ArO6M+9Bmvy/qOF0ZHzobFYqFP+yLKEmIn
X2VhSN8DWw1SUJZgG2X4EVH4w2UJPp3tOewtaBKGWGSN9xSf0XZDk5u4nR2j5KjkR13mVuL3MHq0
fZWE0/gKaZRj+6v/xf3gT9cscYrLDdYbEgvydTcc7tnQLF3WllVBSt/DMYCKwOoq8rTjsq3sfi9o
4ARA8eqG2Bhi5pvG6YhNi7gE9wYvL38txsVnZ0t3Z71MvLpOx9zk5ql/li3YRl9VTpwwBV2cQjBT
eEC457WX0X1FxdTeGS5h07GntI5wC7qd7G4++VLX1zlT6+nSBp40h9Q6O2Os2GJdFl1FoYy78qJo
EREq20cBqvc3wmD+4oJq4XQ5zE4qPziN2XcPa2xLCjHMAmgL5ifad8h3h0jQ7fuA2sSCBfzKb46x
dMnNo3vMAHUtX/wRFMVmrTER04tMc7qEqMRNhyuxJYr1T4/bGMuWfdiBpyQQKbovi63R6HATu+Pn
6zHwByX25QLtvAE7lcH3GIMxU1qfui6X+IjxgsjNAvxLYLBqQcc217ynwjJHkGFvlFABf8l+Y1Ur
K9HQCvui77dTeXtmRBl6c7tjE0nM4k8Yd8kcU+JX7dOmK94U9/rS4PidB2lgvuuAttEL035Job2l
zpBbjp5qu7fjrlz6969U0aQgiRF1pEt4jKQFHGXmgxycLUQXW8M9I+k9c/zEvRFUayaXCgnDH3Bz
F79MnGDjC9idg9G/vNVewMwfs/T8c21bJH8Dy/rgSgFWqXWVlPTeEXrjp1edeu73W69k2ryyb3XA
itH0r0zRjgba4JcK+CXSylqudIE23ax2B1S5em73MMWCl38dI98anbbEQrb3N7BSFlJO3v6BjLtF
OUKRh7EkLCfDlsiYIhPDr1HXo5/VN2DFFsD5nOPaQGIW38sfAw2IkymyK1U0ELqissYKnbnbjK8R
QOFnT2VYK/PJcnHZF68NuuEQJc86TbMvmEif9nCFeyNIqaPYBDsR4EwLakCk7AF+sYLjM1u02BQt
mtI2SzizLV+RXjAIW3jt2as7ytxaqWOkECTL1zro5btc/xcsYvchRkhX2ReWmeV1V5RdIMm77/XQ
sPHpu7QiqIjnEOroDhAluEgDxbSLoE7J25WnglWMBFtS2hEcuDn1zT+PR9Nvn6qr3jaHxYHcvWyj
xHTF87agGgbg936XVqKYjx5ACCkXUoP1YX9BE14Q0sJ6jsLkW1hrIAkk1anu1uVHYY83gE3KICQA
pZ0Vt6c6HsEASqhp3JB8Td4D73STnT2i5mbopJXe+LIgUsLrMdkuXJ2j2Pkjgj6Iv4yyWEE2fzkB
2DccepxBH4xxUUOrp+u+E/hZ5vXawecCJndoNjK7o2z8EutEdmmLjhha33LO6KaB9F84MJLzlyLg
FjWu9rQ8l7ZmTFZps4007w+KHUUJLZt1Ea7UzNpZwurc/+sHdIdjxa9C/myqSaMZVhasuBQEdrq6
1MFMtX1WASIUDsrtcWz0CgIOVJFrFeW8RvtCnuR8wuCvc6LWQ3kR/imJT+haKpvW3NgTNyw3gH8Z
fUX69Cb11TsoxSBG4tof0hcl3OGa+hdvg0M1g5dVkfheSl4Ylxegi8Hggxa2zTsomzl9slTZChy9
Sq9vor+PLuzPcPkNlC9GlFgnd/FaaQiy5usupuklStPfZQ/Vc9x2EXQjOGzmNS0AJWyDB/jENikL
DCERnsRndZdBqNWRX02sKOjAs01/zcQbt54ImkpqGRG5GqTTV7FluiLEeUvBrxP16wNQlGsPthO6
myBBSIx33REvCk5Bbg6xSt69PSHOhud9HVJ/vGA+Knted6+xIFhZbr5zMw9J/8ECvRGiEsurlj/M
aud4BJO62WgwhLILqWre5Wx5uFvPaEwHzigzkJPjb9R8Wh1YvXXR8kGMtjYtTH9cs3gcFsYmfTBt
PQ6xztsAolBvlzEUjZ7o9sPTjcl+joZ7QgzjTK1WzPNd97ZOBwuZH6GbdZPXn7dzBKns0YWDdOPg
3tIi18rrrxvBxP9h5Za3MU/B4WqXF+qWhwX1wbEEUN25HAxvJkyzyLvAglGL5W365AoRnCDriopD
cTzTn1W8K4Ho6Dha/tCq3Q1tMmHcf0PklgiZ4Tv29xBUKyhbmWKIUwvpaoT5h+cXNNiJSfxsRldC
PIvseYTDUrFvzZEMazPPL7oJWeieRjveVMPq+1n87hsgFCQehvJ/mXyF6uR/7rsbt8pM4Al3AOOx
EPgWNP/okAZe1I35QtdgYLSuoiLvadghw934PmbCF8h+vLWsPT1kh/48YwX0LDohUonmerj6Bfrf
sYi1lMYEGEQK68bYlMIF3OV3nDvLw4xcHvIAqIUrLUp7or54LDo0EkH67sMRlTlEMU9GMowbfSVE
4fup1peA9yxgpSjpqLGV8aHx4awdWLv4rker0v+9RpuLciGLnZ1scWRR/e4Mg9aEz0CO1hHyOKeQ
nfGIgDDEjuAtMzx2h7b17ujoSiMUU5Qz6h40G4JLdJHs/MBQD9Cluf7svlyrbbvRFD348vdLnodp
UIfpxfGd+Xsc5WA+wkK0UZRIsbuUkibDWwGQ2h9aaiByHNNgCKayrEZjUa2plAdv5pMo8MlqPCSl
b8rSlfTcmsUDYVKfGx7QWCYSqDWz1FPJ5+C2nGY5KpQAXoHZWQd+DH38DaZHIXFxuMT7E259aIyU
ogXVxDIp6ODmx3R4Oj2/68TkMTE0HUWITU+r7ntFcb2W7u2iw/nfTzlnmWhdTYvpF/dV4OMoGLRp
Wn887SPAkMvBOxpo/gd1E21tBSilVtjRb2Qua2I60+whASj5r01jW/9TF3bHYp1n6yP2zgrnXH7V
o5KVFxkKhg73+jTNhDX2Fk/Kk2aIohRlvarXQlN7SI8ZUmSRZJpt4MMwOQqs/rKwcGI9lJPYGqxJ
nTRJ4vgxfKHa0ffmlZkQ7/imhpHyf8rdoVbBzE3e1yf5zPDKi4PKz1YJaGw2xuf9pk53vuk2Dhrr
T9r7xP4JcYjsMwK5+XqtCzuPcU+KltcBjjrfG+pwyVvvDRvIgA0qu/58SVxM+UsBZrK55NXu0lwI
hjQncJNLkiXe0EOTXN4A1Wl5cf/H1MJQ3EpzxGUo3HHXkMn6uHPcd4NcjMdV63/dFPWE9PTfTPD3
Jz3uBBbYPRgFVH+mzqsj1gjnjLU0rsDJjpelhrWgwuCNk3uZpVcEpJF2GL0/1xXzbsY1nINu9uFN
8il3i7v+EBcd/+8KokdgXmmx5/c7mxcPZ9N6uVe7t08J72TtM87BLv872RkJHHDRsDmxtvtjnc9s
8dKYu+78yb7rLWNmzrayPZfGGvjHgUGzKlYQxMya1MX2UQ4l92cwQ7rGFX5mThYyKKEeefN1PSde
d2P+ekLfk533ybopuiL13JB+9aptfT4D9DFp2BdKZ3x92o87OI2MSnDrx25e4Zp4GioaADOeEtrk
wF1cio+QEK4Abn8xgIg82893QooQwY7EgeB2ilwpYkGDWJ97rTc225D0zYf3USBVr+Z+heMYY3i+
SUKvdW98hskb+pndBe9tOkB8o7CEgMjxaZOYDGZ/w7bd1bVLYeZO8Id3nNhT/2zlN97b2+8K7Tsu
WqrSrmbUIUOhlr+pjl0pmXQnQNCVnvxqT7stJwqdCcGOqYYOO9P8AydcAOZ8DeWQ2uJ0mDq03eSH
gUIwddsvx/9NYziMsx+G9IQgzwzajuc1WKn4KWIisIDByDuwldq3RcaJOh2hkJm2PYnVWFDaagcZ
u6qt5Lsrx/DqR31kSNFMMta5JHHG3Hm5t04JXsi0mhtA9G7UelGfLNiFKpWqNsK3vsIH1o1jmlJU
7CYGJnWl4YZ8STvIhY/8J/ub2Bl6LZ7x7jd2Fd032kKiKkbmgyfIrjvow9MLMF3u6S4ENkRBPRBo
bpqrLhMcNZWs5yFnThol5aB8hfD6yG2DfvgiaEZaFeEvz0Ncf76AfMdnHh4s2lwwpUdpJ4uyaf6m
gAopdGktcJXQYzexKQ8+VyEq12EUp0YsQSV46cAaDLduUmz/fnP4genltDNq0honwkOallfYuHFi
i6a9tZa5WNNHf1MRR4Cjr4q+MO55fAMtsUxcem9L2yqoUzzKDYgYIePjmuu9Wn8ZVEI+2NC8bxQs
ZsdgaapzCM3eG1PUWlOpARVRgbQpGowA3R7U6iTPnu0ooOrllX9H9EQWEAAy16UQ5UNWRIm5RlqZ
YhtjRoK7UYuYogfUj583x4yuRXDvZq0m7fcbXu95zFUOCHLux4nJ3kTKBq8cBVvMLaTbmA6e/UKv
HfPNedz+1jxAXkrNph6m5l4J6vRnF1uv+L8AGEVV+jpHBLQQpmM3oEO/l6mRl575ddp+HQqiVo2I
V7MPv98x5maCziNwP/lXNGvNbFa7cKykPFyAvaphLAuoyLhLsSNndGTHvbe4psf4U913lrZ5KVZa
ub6eh0WbtYnw7SOpY7HdAR9VZKXSPZy/ROrP8wlhFSy2zzk5uUq5exOSdMUSJ0EdS0oW2s0kUVmx
mbLwosy5unkVvcS3J+rL21+52Z0=
`pragma protect end_protected
