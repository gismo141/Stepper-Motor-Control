// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0
// ALTERA_TIMESTAMP:Thu Jun 19 02:53:49 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
STvdwBQp27NqYznpdz/OU5imSxOc3UTUAL68xi616zaWaePe+uSW+fPckSk7LBGN
My+dZy0/f47G/EmFxWgseeZbY6LBlIsEn4Pq7m0ZHWm7UH6VNvfYEBji/Xdgg2nu
ZerupL3+mKik5nwWPnasl/5Ze55CgGDxRFy3ipl/Cnw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13968)
gYbVA491yNpszHT4SPjwT74yT1QHCDqP9mouXLI40a4OMjfrOI1T+VZVYw7sSM56
KntQwfl1KZRABTebFnLzk2pSFOryJcrztq6BkNul4m2mf7HRw9J7XBgZd3UwFKc4
nmLyaR6g4nAum8eZNurAqekBKNOPUWydMSrjslyOi5OsuLv4bHGLI1ZzpPHCe4mk
DzY0jmumt5uXOAeAEzFJk9Uhif64x/eOpnOLzKmKxR3Feanc3fNvdWf7Ao7/O2pi
W2hTMXdpAD9Ha1f+0WevWT/5yUVwobvEq/QQrhZLn3B9GNOJqY+NWUbzKWGQYx7q
A4nvHtEIUSn9RcpSS2RFzkcCJZiFdNO8k7IYDP8ktZMz4XWxMNXY/faq2pnf73CK
JvWPMrPH4VBv0nEAMpRSlPD3h29QYZUFw0gx7byU/Xqt3izdcwKLqBwaDd/F3hCH
8x4B54P7E9QAFVW0ZnDDMc7k5/ltJ6hOVtdzag6bZfN3Gr8XFdONLeNy83x4w5rG
WseJQKftJV6y4BIkPg9uqQoC1IlZwOri6zYvDqg4Npq6tDLOa7cQjSnouPrQtnSz
lUWYmFN/CRdgGa84GF42Qclp5xdZedAYXHH8tk+ogyHJMRO4O3KdyEnaPgm6Efuz
QCirnpAQ5M45xye5HJC+ACarFl0u7SyedxgQhHoF5AtAZ5p2YbyWKgkStdGbUEQe
BRKcZwb6IBi+dPGCRhKMBpquFEtbkmGl7nfQB9qJ7k0ZVPeYRB1zMWOYPIiRRk3l
ZA9z88Z3o9FL6jGy6NH03/fC3G+DtbFBrX4MCloDEfp/hF9/zlu0W9l8PIIyJ8lu
WtZVCcxzCUKcI5BXfPxSevrIhBELS06LBR7yHBR4mDJ/hTVGWMRmA4aF8kNe8k9v
hJEdy1/lpVVJWu9fMHfbzj5EXRARYAnO0VudY8q/v3b/9cXnKRuVm929r7FEyCHd
KQr4oV7Ia7tINxMi9+itWUy77hbeOoznSIAG7FsARR9d0to9y2WQ4TmTHSs7xJQI
y2ZXReMirg6s+OS+G77Lg8lB/OsZfEMmXGDaTLs/ZloxYPcjKVO2YuohzsNI1THd
OETxIQZqx6Orf8pnMIEOolITTFNBGt2rZk5wsf5nr7CBq5S6IAme0HdkXSHNkHbZ
lwowD2tzr+ZTBnmJcfKoTU20gIwu4kyZ0uqK+xsr7Ims79N9I6pkO69YVMPSOi0u
cIIJaIrTCGRS4nMnQ9Omm58UkPQXMpYxB7ECgxrNClnLMUDJw0DNb3onfIzMF8wE
wux6giGdVt/IYTHBHuPlrM26hIrXDLa5gcrDCAsQC5W5m/TgTFRs2bx3ceFe2GTW
3BT3tkPqi3nydJnu1rxRD+nJZGOw5WYItMniyskUaLF2NIR5+T/dIn6okrCkje7t
2rM4cseFpYLbvNPKZKJTHU6rkc1g4FI1ILePR/lJW8VPWdvfX4AAHg5BNqIIpMsS
FVGFlkevM6oaOKuu2avrncCydaCFGzYE0XTYXOL5bHwKPCDkOAKaNbP9Ik3wNScw
JwrHurHCe87VdiV5ZjvLaxJHBhCjQCh3iAlXJofEQ9FrdDnVUp0ofPIugZbXIWPM
GHBnC1lQQyqGQ0UqybaBicctiphu1xZ+DMUZbo/13yC7BM/yQZUzCqlKAUhhrwPG
WLX2OcQSOPbZz+iGm5qw4EuHLoOOcr7vufXwtS6gSeV5uv+Q3SmLZq/lgbzMvegN
J0r+3QSDKa0ISEfXaS9PG3YvDgwOM7XmfK9G2sHpPU/HEzzbVC8aOHcdAo0KDAuL
+HdB/F+rNpbNaCuzZ6KDKdc/IYlpQ82QH+SaRmbgsSNquTUWjiMsVqgoaX3V1QPu
QRa9Xja31/C4af+blJnp5mWD3SfW8vKQ6+yyTB+4F5pYjwGkAuFD3SZxZ3xJn0Fp
up3IjqEBxDZ5oFTLaYv1MGvcoYlj1+IEpIpe65PzDJVndBcoZGi5Sc3+038VJxNd
9CNjmTxvpc/EDOeDTWZpykp0+rFtGJiANmTrjHQ8/K4mBEQt8ac1e41WBoHtR67r
Ihau8t5dokYEDBTb1D/Z5dLwMBKgTeqSD0sLo15IZV9x/Zv3k2NHSwTPdWEtLdLc
UHlawgcLJuJyodfhLeBCEQuJlugbz9lvl9pyHDC1Hfm9dDU/tOl+4X1+G0psxL7A
Ic7gcSKxGLlI8OHlW6NLfHiJrHrz7tEpdrW038WGG0VKg1oxRsIU6eC6Rl5vIES8
hZeNexbXgBtJoDHFW9bnRkEQwV/KlsJ6ewsy2SxVHnEwqNKRulRLmDoNVcf67v0Z
NZqiDj/QTx9TZ+AQ2nj9n6XxhrBeNoPJizccb92wlPzb30CgqshvueRlveUtIzwx
2MfDSrjXS6cMeRbkKtiQe2SjL2PEGD71KX7lD0ebompnu2CYmapFJOb5Zj8njvBG
CfE1TcHMnWxMHq/q7xypyS30ZBEcb4Pc2K1mZBsezgbDe0QpN9yCYPqMPfJOpwk9
6Pdwzx/6ZB6FZaUvgDyrhfU9Z44QrTFUPNptR5CA5FUKD+o948thJ6NZYRCnatlI
y768ifGwM3mzvv5AgSsPYmgNxFpGK2j80sgZqld3lKaOtw5hiupSicewcAdiCN9C
sKU76taNI+5ccmfTRGbOHKBcTMQLEPzxEgVzIMiIlUn/sbKApCtaonaKEkm+1tz6
lBY5xlSnOw2axQAgOHZjM/D5Qp5mPCcPKuaxqtlmonC8tlS+BHkDXDzw5Nd2ou3J
9H1Xop1tlFt4C3qngf6FQhrBHMBKB+GoRCqJP/+EEjLj/V+TZj+MPQf9ZUtTqNrO
AyvVOip6p+XEhfzpyT7BTA8HpjI2+csTEkr2pIE/6NIGjNfmAb2ruijbppVAa6WB
gPXQlzvJSia/MUtvS2wQjZA3UeX71xXFUYlEXNCBZV/ZhTdiIn8Gq3Hcz3eFynzZ
s/Ig1heZWlvLvRTwBjGCGsCCRlz2sCiiWloT3lgyDcxQfcQ4WUrt36MAwcbOtd4J
n5cwtoYCRYoZqIwAaqwON0Z4/hnrKjTqn7hqwgStHe5oiRzHrasxxwyPhmHe1Rfy
b5XCz7GxSWDry4qMPkehbusDwIRlrOV3HjNw7zGWFkkhgP6zZbWbc/4hAEChNKPs
PsXC9jKWmfS9Oj0AwR6CnHGt0DLA4JGT3Qlm3aoV7tejk4n6q8hDrpS4N4lqrBca
JcwCWjyd4BUi0jJj5cbh74r4x8oeSH3E0EeXL7v+h/8HNSfnfkVqFJlHrdbis86u
bMdI0O2Kep1ztD275sfMFG6dCueQ1UInKXUNAStBqvlhL0iJTf9pq01XNDJM0YrX
RiE3eJhjtCIOTGfOBRCkhD+Nt9GILRrxgI3CjVr7nthF1RneUPDeYwDbzfbyY18s
BefUTKTHTgFzSAEKzF6FgPGtQ5SnmRULpkm0uL0/rKF8IhLq3W4uramrrgNVDHdM
zEx/BpJHlMTGe3/uyXi41BTImPzrUrXamUvKf5nCvX2M/qcSfN2bCknCWvvWMdJ+
5QtyU9jKA8WnVhMVaJKH3o+gSBOUVtS75RlfYWSCh8VNw0G4KJvrnMSk9Uu59ENP
DALg4GaxMr7J4NcwFeTKBlsXGYjoR9PsdtfAV7BP3X//CGdvWp/8YGCoRV/mumtv
D/Ap1HlUEAZbjZKBe036dNGdlM36y7+g2kvCturc69ocvJYyePd481qMBRMW21zp
0O5lc/68NaUYsgUXR/JiAFz82NjtLu4mNI/rvo6HJN5R6QDAn4+6crIuGs/k6njf
ROI3MfyWOB0yikNOIEnZk/n1W7/QtXVHDl0+NNDxUvOeNv6diybTcxFAsmRuPT6/
BF+AP4MutIP6V2no7Rdw/8Enp0+BsUF3VYlg6uCyRK5q2OTVT8wKLBQWqoJUb08T
a+GuYKStFhw9ea7Zzw5J7DDCSd7xX9wBcaTmUxGuaW+bXhpQMN7PwaFozkBFf9f5
2r3rqVyehg/CLVzKdEqsfF09zm58rECiNfZbTjarx8Zt4XhnhS2J/X1y4Y1+xwgl
tmt+EzFimCGsQQZGDMa14w0H3mzjkvHHe6EOTGhFw4kfjW/M2qPDUpEFBSyQL6N+
7hyj1mI8YIbk+zpiGj3JBkYWQeimRTHhptTiP1AAgwuji08gfiNHYMgCK7AlM/22
kb3jPMGGy1iHPxQ2SCDAtf654EoxRhDRjsHCTesryhE8QrqXzxWRcIVGK4GorHr1
lwmhhtBE4r/yIVHVrhA58tq2H0loF8ADwP69RTOGeMbX0a21d2rRu3wQaYdyB1hV
5OT6kGCjoxE4vxr3fx2+IZpjoO5kyxGIKl2xdiFJyu2mveblGOTM6Il8Tjv2G1XL
cTD5EGAC5tLahev34bHB2mbLh+aT7NlItcphGVur+Yq5frRxrAHKcTWSCxzJFt0Z
JzAbuW2DqT+CH+YVQ4Jg+x1A+XQpJ6+yMWEusQ2O2PGOFJAWXm+1fveLKpICrwst
9mpzl3S3dcMJlp7T/miBSfKOOkUHk2xhjJlwTdBYTKSf1vkvQZv5PYvB/CoQdbnP
93GY6lxSDcZgmuYoDtoCbnUVJ2KX7016sZhXxcFbJZKRcbfmgNY147n9ujqRjz7f
FZWH1mQV9qzAjsqBpKPMS99seuk/uPzi/VGOtT+QnJPJ+sTKuhxzF51k3arExpwO
5LvyO7ke+wsJPin0GGZH5nd4ugudY0oJeMGM9tlQwcZfGcI+sb8SVWUFEfFJRIAc
p1fHFhfnFwcMrVWxUFtlFmE+OlxIfC01PJf2A7XPK6/Vn50XZAODz/kH23lG6zw8
XFAugrsNa7yndW5l5xgvqcygekEEkPtZgrPgtAS530fVAqpskPj4hlu57jlKKpGO
0AC66effxZbsAAEJWR8hm8jEqHxxtYQ87ytT6NswUUiz0RZ11VXYwx4/YqqURhUe
AD3YrkT1J1thPrTDsMPf7CnGLdxQjTlANJ7kxE+Jan27RByi8MFTiXLOihrzVhiM
ZxzD3zNnJB6Pcl8AVvM08QTpQ9YLlfyYTQPdPDqt10SGSL/blYwSr/pK6+pDdH5P
3/Mvdzgga9y22/8lZ7ndn7aJVvjhviWY1F42glSTg/Ez0oVY1UQc7kUw+vPMnc67
ugqpBtfrDu1eeoJstsX0H1TFl4HAHA0nqj6RzerTubLTaSpFzQftUfXc9s6XfcSp
o5vid5YLXQtiHRKOWZkBdNsdxSgO+i9py97kal73HUY73CxF8ppjNLfC8x5+AR0s
EZmeI5VPe7FAk2GuPT7PfDLKsUzFhVyUi/TXjHQteQINkfbKGQRyx/KlRiEyxnBC
6eDTC6eCBWxnaQOJS4LNgq3tnYknM0+jdtio1YipkYY6nN4AXrDwl4GbTtssoPRa
kAFu3MyLeqo4sDmz1/2Nk42RnpK8Z4pZt6YVZbJQyPBeGFJRUZagE5973FiuEfg7
JVkaKgUXhUw1jEvfX0KQgIdXYLnHm30oHIPpPJXbPBxfYgXJAjG7pDOm86iGhcWs
HTsSY0pdgWQzap0QZV+lZ4UJZUUPMopWQwW34ZefbLMiL6b6ebRZudwE/pQYsg90
KGlhXLYCL4lp/d9Ftj5iE+urCQRoROYMIp9L4WkZrT8Lhbxjpz4UVlBecxSflMI/
DUf87r+kLL06xkpCVzdLNeEvzN8nJu520l2gxrRUA9zalKmnQtUgDOuElXAnbiMJ
23X/3W9PPMyGDDBb6poP8bP3Fq3hoiCfCFgGTImf/wwlvD3nOK7OPd3Q8ODbywpk
04N36cDdNBU8552U457ZaesgtPakzwL47srM7QTyi+QG8baLv97T/RqdhOa9a+JV
0IxoHv7WrUC5xoPCYxYB+jekoxw/ok+WEzoQldqp5pcIEKLnjfSfs+3KJLrtluXu
fCwPy9IBGeNrid21nI73kljSaB4PRVoGqs+dO/Drl/GR33+s0mk955tbgdIUuWJ1
SPsLgSEoRsMU5Kw3Z+80ZL83Gbtg3+3jTCjMur+lrIKoK8AhqbqXeoEC3sQv0XQ3
s1Iq21ytIfxfH1Au1OfkMkOzTtYpkBiordC3d7KMoA5T/xL9iNTlWpPPNTkpoGdZ
qRY4K0OPsKHKCF8+f9tHjA9lVcGWZNmqLr1dkPv3hOIUi3opxjdRmWlDqeGtX4cI
0UT2JRnfXZAsyywqOP1Krqe1O+1Z2F6si3LUDuli3Urm1JoQZfaxuvu+Q9JulIsw
qt5rZMJOJxOflKp+T8BHNrWl4NYMqu5/4BpDjvHUvwMljqEW0H+chy6pvBimqbfI
uwMEsA54Bo858GK/3QqoLdj8Q9b/SFRZcAK86lS2Qt1Do0fMigL5N0vUoLIFTZpf
oM6ckiz4MS71+ZefedT3gLCDqGBmTnVfBiUs0IxmQegsRbkf4XEaXyPSa0qj/KoT
NJUH4DHMgJ4qp2Xz/I7MlloWQGnuBP+CwbWJzpO3Qdc4p/LiDzHyygZ5fG0RnyXX
soPoc4AbgF9fbmH7pVn0hEGvlVdYQERCk2TyRdfhY9QE2ZxHdaDfIJdlmLbIDoTh
NA6ljcp9K4Vl9kK7+QX0JWkgAbip2ZvVfIvqZiCRj018mpYMVpbT59DUshBEL33y
pGdqsIqhpvUaDQCFrSHKSVIViVMY+7QmCkcLe1bSnRlYT7ZnWQBAezjX4KJWBUHp
z07vM5jIcSNdZ2q8a7NSaZBAolLbrxfKDnCyk4VzbXOh1fvMCJb8TkIQI5aqD3Ng
y7frSOK8pHoNlB2zQwHW3Ab4Xllz1cT+ioj3wDKA+KR9fudxC/YSSqmRrRbQhbJz
1VJwH9XAP4anXmdAaGmb8jD/ntUA4LJUD/HCetxlbMLL3fY+eVH6W1FF64FBZFB2
h+dgA0ilyuXFE1BVcNnLWTtJ5lY3PS7mlSvAqHkqaNoW1w2G4NyDP47lfDxWG9GY
JeZgE4R2lkThLuzlszrdDHoyMMzkKxEsdccXeam+CYlOFjUW6jcbe0c4Ypc+ALO1
gtTPugKPAh7FEgbIC6OHlIlPLb7YbtGxt0DuVba+D28Y88z5arBaYPbK2sLYbMYR
f9XeDZ6FXjBVf1vJtluhzDI4VXCEG7I8arusdned6ZGeB/QFssI5XEqXtYkYqPLo
6dWEsJE34yHx2e8SQEkgpgAyXD6HrZoLL6QEbnm2vp2sn/ZkTFGtRQKsPlWp5/BI
OtuU1b29If7gd9HTTElDVkXp2aQ7/lVMMccIevBibM3Fe8wAjtLn82Ig+gO+ohLY
FUEM/arLdKrrmk7XOmw4XEGBDLIws75yB5mneN/YUYo+7kTml+HF80jvPdiO2Xl7
TupcIlHI30/zSXltIThRBmv4ex5iVbHnXi2/QLazK2UDgYwA23WPcrcCNkgj/7/S
yrs77s2Tm2a0Q0z07odUY17NMTzeqa631GNg1vlLRLwx8QFtn2f2P8stW/uLSoyN
1Iqnpl+69f/+SLRh81NAu037EpOGnwbPWTOWk/CMkUv02/E3taeNf61OCVK/e2xg
2xQsq/FrOOqhn0uCWp93lF1E0BB/qmXVBLiYVLwsMmnUT3IQaJc08zs5KB47Vngf
ovTDjclLehbpHxvRUTUSLNANloiBwAkcPjAPaDPrym8edV/WVS73B6UY0dInzldN
qsXIxrUNICLWLxqUZDdgmtGZJ0LT21P6xhoX6s+gCAIwmT/55wd9cuJ3oKblslpy
23W3nN7qwc7VSK7C69eIjb6MISu+zIgSQTTW2zdEk6HOIlyv8jSmg8lvPJLKpzaM
jNKf7QDnGPFEZ4gv4kppTE3i+xVoHAX+o6TDMqcj4BkbmiKSUrzVkdF9rS8NsjAC
EHW6jMKwo424PWGp7XHv8LkRMjkNMWUgWyh0VSCAfA8MuIIWnY9XYPZ3otisarou
NaZK7taIYudnN/ggA4TVuPx1JopoTjjPGvAF7yxnBShun/8sMy4IvbWSNCRfIT1j
nmpEkxjQ26NZ7lYNYHQZQqGra9Ald65Zy6LhQanZQMpgJsHhrT0bNat1oYEQThaD
s+1WTRV5QLAOyn8u4fSVYIczp/aEf2h3mkxAjxrTl2Wyxuz3/73/aJ6gqaRXiKOD
N93T4ENd4gvuVD/Kmnkubv92CncIzeMZEYtobpR3Y4ec7rmAiq0bhVBInwqUJIQF
EjjbtKrhrTQEQc7wktNqhYHBPXJ3BvwOXq6CmLorIRlsk6sUkUmeOcGyBWnr9CeP
Ue2gSXwY9oOEzuBIWrO/rXlGhQvxQlmqb58l4U58IBUsThIUql6dE3d5yVfM/vFJ
Hi31W+w2wjf6FJgVC8xmFQ/YNK5ELEVHRJFzX+u/JpTPsXYnVyxufEjArWRvaTST
hMPfgNVvQaNRwHLqliI8AK/7qiw4Y5OEFLpNynerPjKqGme2NoLOLlwA/41dX92q
8GJJqUSEMu+FXZiR44/E2KhOLVhRyuIJJvFs8aVFxgPbMZMM51sdCUtbKTRGnkK5
5UjB1MZ7jSU6Nrq5t+hixcBrTdO6DR2K40suaz+eMu9zP0FqlKke5ntF0HcDOqsj
B27lLun4iLGnuKCaVjWOdkfStmAahinHBxwAXREWsA13tztUBK6BzIzzr2KAzncy
E/ngHGWuZiIDiPuWMREDdmV6n/3BfNjSof0Nck7wmIn/A4VG0h1247kysmqcSJe/
Ai31UuaavdPsjr0FvoGz8RFKqRr0kOuXmxF2VBqz6tQZX/F4fD2+aqNR5WJSoatV
EMkG3B65Y785j4QgaLMO4S40NjJqKDKj3Dg5GOhjuFbuTglzxm9nRvHX3eXzDFNR
3EYoBPxrAUu+CX7w9/UuyJS04hKdqcy19ioy5PdaB3h3eRnnPIHvD8f1XXdd/aYx
qWfUs7Fu8US68nJf5OyJEeASv4jAh0XnNi0vxtY+bYqb5Mi0hLe+2u2GyLHEGEb/
jG0l9HKGXdWpRWUaSWDC7R1tihlSDRh+fwTEJ+T+Xt4Xe73Wgk7udeiQI0Wb8Grz
XML71n63wLOaREApS5kfL3pw6Lx53xjTVHAVPg/qt6QZoElFqN4JNc9sT0gU+BYN
cdGiE4c9C496chumFbP8GtIYQuBAp+JiQPebDBXHTKg7pO89GYN7rLaMuCqllhPy
nqYbNR9KruGPX54vujyasirgpl/MLQQ1h5O4ScImZ4vzc1pi+3/uz2sWE6dCJDZq
BvXvDFiJ7qj0luSldrJxpJioSmFc6s/1aNAgkF3/p/Qxtf/AiVkDzuVDFLvd87Kq
Zm69It0SiHoEhGxD4ICRKXsPsuYDB+ke5xtzRi1AHLOZlxOOkhMY7+8VHjQSMuu7
zyufIZAaZlcJG8nInVsptkyw9rHMiOhmzlfsCGCDgKs8B5xoypNjjp9BimegSiey
a71OJKVlr65+I7hNtr596h9nkNLM0JaZmlKlid65fWUBhdooBY0TCa2P5pDcjkbI
WD1nAUT4kUo8CUAyS6a/XDG2JEOm7SeIK0wqUt0Pi32Q9CgaN4JGC+DFlaGIYV6O
GyNFGQBtDADhuAPWatng+gSFhYuYfTth24d7hrBZNxFyOMqfA+bnL0zV+nkCvnbB
upmooEBgsISy5E3gv0vF8i2i5gd7CrUl5IuT43eCauwkwJKPk3XCBg8XsF7EfdiZ
7S4GkaduoPfyuCfxQvL7hqBHXkQvoEOVHSKvYOd/5iz1jAkH4AoBoxk3oL2Fv0SI
1jiRZYgZcjNOqiyuVsxyd+q3jSM44uklcucKIQpyWWDcme531HMJSjIf1TFiWXhb
TaNc3dymetDvRe1mkJRWWJvcppliPIt9wTEimflHzb1TYQtgYUm4m/FkNnM2V3mg
HIDYZbk9ZDsqtu9vw/PB3LF+wVkrAeBsegOT/APlDVvowjCIvnoV2VorS0HTbOpF
e9XkcMwnddGqGZsXJuB16Ny8NulBaBBQ+5aqbWWQtWsdf6mVhkrgXiZNi1mEufFI
sCfJ5wDgjaX4G0Yyb8X1mtgUL3QbxMwLuxpT7HVh35BwCzK/WayE1n11OVuF8DED
NP5cf7u0zVU4hfqYWMfiosAGFlbBNmcdFUYQv2ekRbLJpYXgjSdyBPZISpBrkdh7
pLQOOivN7vxX8PNs2uQb3Tl47URmIrYYRvjM0k3Ik3p0l0Bi2ANC49p4GjM9ry18
kb7mgoQFyKTI/DxAmlURJBOVT9kU8IH2jANY56ZGmg04eeAHjXc68vnmmXVOBXPa
fa9kzIDbpvcgoQj9whV2rVtXd1iXAfneS45E0bYQ9fmEML+7we8Euxy96kV69O/5
lmePWhClE2lXk+P5pvVhapfQU6uAcIsQ7yKv+4+JMTfD2so5Ue6zoViI/j4olBoT
34Es9VV1Pt3tfUXZUmiisv8HEm0ItCdeDX3fVyJQdbk2RQLrbGaco/BjriLk6OT7
rsXsIJz2av/CqbPT+uD56/OWDQ9pXa6JezkZA9KwIWGCTTW3pRkYBRc56dM4Movb
OrY+YrIGFdjhEILnKKMrJb/nAla2GhsMy42qkY/tPfEvLaaEorwM8VHt20kFgfEs
6FoiPx0Ao6FJkpacIPuDoYHZuA8arBWEnRxP7qVEqRd62sukSH54ut10xWCIvIqS
F5mRZXIcI9FQTkowE61wL3vOCfubVnHJnGKiz5yu4B5KbJ89sGYid08/t2Np08eY
D5SRaTkwgqIaJk12uwsyzDPL9V6chEp3qG4Nhi9Qd4wm2++8E6jn+Vlwy44xOJ9+
KTrlS8yrsGh9J/uAFfg6/NrqOxqJJYUMzDCfmoBzqcHGVNVUAPm04ftgNurffOip
lxLGrYCmE9o9+skkffLsCdPwUahDfbPmLW+lmvAjjhO95P4L5uIMSWBcQPOpNVLD
m3iF5VBZcisl1Kl1iRDZ2Nvco1RumOYwT93V/S31o2lNk0AV8J+FSgxfBpRvDr4s
43iIY1S8psBk6iCTKK9YXIq6690tgCs8lnLDCgpqiUU5LBg3Ubzp7MPVaiWVo66d
WgZUfwNnMccbqBes6kn7u3LmHgh27XIC0FZA1r48ibpEdeC/GUlnc3qPm/yydsEk
qynfvXnaeEI332gnPVo+A0MuJo2VqLYwjqOVVzRkOIu7N7kkmQ+kt9r654ck2nW+
nlbq/JzU2zNxPHCF6xv8gnH99X54KMoyzM/nvg4N8ESq9alXjRgY/kao6Gfhx5PL
QcTT8QED26uOgsquWYwOW9Wj1q2joZ1ESEvJys70ZtTLUn96ovGHGT8ESUvDrGpx
e4jqqcnzz+iON52SPFsBw4uwXAemC+VuW4U0HlRxkICpVYW09Ym+T5jLKZPgJysc
nbgAPQEL49/UOzEvmLsh6ucZGXrRTneMIt8hX0u/kv4pdiSN5PkjvyAUq4yArtD/
bwlZG2P4UhY/jr1IFQmHX0b9oN+pfbLHbxqZtKSvbDvruPVKuBNAXKEJlsKV3A91
8LE95u5yGcwfCwu/jylERCDmaTSRu06KPQoZLsJvQxNeevHCbsXmXW9AH1m8yReQ
yM9q0w+1Q5X9tEe+AKQJYhKTmb3/B7QRIVR6c5SAIqNvcntpqBlzkdaYkVuq/S9r
2fMmp2wyh1ylECAhsWfdRvJy/p7KUdOr2Ljyn2DtuPsjPiaYU7ckjVDrCILixdcY
Y4Inc2N1vVUFFxNOLnkBzk/ebgsVjzFl9sQng+7dU2KoEpC8iWEpJSDBg6J9NpY2
+ei8ajy+myI+lyhEluIS2sLfIp9dmXEqx302dZbG6DnT5g0RaqpGJMsx4oKQe0Ga
wlNL9d3QP/vnm0MLCtGDYJo8Z/dabOfr6X07ic5W5toZWC/wIikMHsZ7KeiOxjnE
aGZlPMbDSPbAZSkygTEnCXIE4ltvK4KdNouzMxqjqJIqlMLa4va219m3mVprfHoy
A8nQAboevqnY8HvFRG6TfEbclxPZMDBOMn+woW9v1zXNT7xtzuZm59hLfQiU/dDT
AIxgFMpClGMg0UhP3YGFcFdvHupVvjt4roVxKEwouBcsHRqp8KV+qlJt6vcYzpHt
x0k0ftH+CRIbIVXbUPq+g6HWgmGWsnVRrB+KJmL7DnsD5j9r5IlWtICgkdQXAsiA
CSW1QiFjUJV+eVHFdgEKDqyH914uLn1Z2rCqOdEXHEWv7djAuFghLSrsEclaUHc5
gTvHO6cqfZrfLXi+8mIPk5cAUXaZMQnXJjECtVtUUkOdik/p7FNnopmqw36yJm8b
4xSuzJlOpSuoYpxrJy6IDmAtYLK5kswv1FpISOc1IQdSZe7tDX/mPxtW4fZUMFb9
2qarXKfdvka0DlzC/139x49b2tPI9Ry/+bVsEVvlftA2e0zFzmMx9bZcn3zEOPpO
89RT7xs752QYIUTUdbnIaeB3sR+DGpBS844wxEkVAi6Ll7zfvXP4FjpFnQpypERk
Hn60lCyffXjqHguCfz3ucZ6lkHiFzgLyNgCCOMlNzew9qP2LteEc+NEnt/jk1Lk6
RpTMCXn0oo5qKxyAd+9RBS3eSwS3iWWgzdUwjUPtxpFBV4Sfeha+JIWtgtmDgKy6
blJiMlEA6hVTxrsq7BsVo5VAHgTT6mCdGEUbnrYZ0A4vgdxeTXcpRfZGY0hNOZUn
UaAEAEVWPqxDCHFquixFW9dhUyMoa5BMms/ODrkj7/7aVuVGG0JwnKz7FHPe/ZTR
oM7LpNi3rzt7Y+Vq5R72scGfXvKF/MVOY1S0KkoEox6iZnsYP4MJuX67iYyp6eOv
Cil1UPoZx0F50QBUBc2roQEWwcx74lJv72cR4IxqNjGpAedX35rFxQeIRwVIEAru
f+tplUl9SwSswcLV+oOHCwCgzE6YYuJjQmpJhQZV6r6WNJ2uUse+wVRNjz+5SKuF
AlcFRtKXXrikLvjbC6klMfSB38kaltFnXeAxwVaXfILr4ek0nHXsEz3oeMxCDim4
STtIEWuprcoSE+luozusavWqU9AhIIYRsv4QR+zx+LJj1OXLqzetsIx11/otDvBE
x+wVJQnndv/bDC+/g14I1CY4i7zop303qPKXflzUKXVSOurR1rmSA4FgfBNKzvcm
tdOy8uDXqtFU+U6KcKmqrqTNYGNolrtr6qAe+5wtFBBvOsnvb0Pl9bkgfs4eS3W8
prnhP+eMKhRXdv+VvVQExzsVwKgwCIMGT0wdi0WWn5kc3C5WZDGerAKdT95+4VpF
C8DAvI9yRoiwhmqSDwTb1d2B6EXoU+rb0iyWGqtjiYXSLSXQ4RrDO82/XzCPPSHj
M7CsFtIGdP2dHmdnlHEIZdZTjkPY3R1oQEU5AQ5YgXd+aqCde6pGLbEe2IogJOZV
AYABLO2IXY+Z8d8TDUv45QAz8cfZIPajJxcTmE1xoSBLPHUt/R/i6UmOhOfwZ90X
wGF44WMVg/PWgxde2fN/ZB6Z20PmveuMKWsaMz5uwGJ+fkHuQeEfs1G0FrvHztNH
H2RJnrUJImTd7ijiJASrzvLyP1pIznV6Hgy2TmYhT3PQ0PTTh7H1H98dWdZAcE96
8zroPICs8zfiedc/NLxaCGb0QcXiJclHK/QycirCpmj1KsBz8Oi+hGXXSkkkkEja
n5cfqqc5lNS8Ik1xohMNBOcWKRKNt73joHM3uMCz+PO5Y6EqqqctecJP+IkeHj98
ib1aivasS8g3jRZ4qRZ8smBNbUTKakF8z+IMwUIQCcte2D2Fl4zrwDxboi8IDWno
eU0udUe7AQ1O29DzY1zwh4F4cBWsK1BWI9GsK3TVtCAOy3tz7Fv38/UKxyZGEwaR
lXGMmvmDE9w5eCcULU+yVxVEo/Me5NogMf8TcmbRas6HKkcyyeNhp7l9ofGsEsKI
ldeVmG6ZJCZddku9dWpF++TAtmxSnUHFcuxre9i9R6TM2O7x7mLm6gALEq6hokGU
zKTyO5eBf76oCwmEtR4LLYrLuQHDB5by6/hgFSnT71FFk+BYoRVYGV+Y0IqByr5Q
7jfU/tK4CQpltEV2MR+Oa2bdZb1zENyWVbFZFDHZ1Q6WuqH2R9GWGXABTA3zavB9
cc5/Pa8laIrifGrkJ0W44CtDByMB3O7VvhEDat4DJVV20XhboWfARtT5FomDKZeV
riz48cgawc2uHDmKIjllVObowiKBcflqZMSOD65+1xPj3Ghru6VRUG71ikviP4kW
sDXcs6NQD9qDOId3coV8qg8/xKLcXn4D+Qik8QEdkhleGyGP13O1WWl2Zmpup/OE
rlJPveeEY1hHFl/1m1cseWFidXaIlwZs2TlBGuE6h+9gMIFXbhuUP4I3E2yLzmi0
psVWZZJjhBkHDD7unsxevsOT1jxw42OVQ5s3tpUeNiNszbElFBO+J6bjBeENgEJ+
R8YTOY1I4sig8Ah0wYPP9glHea9HVHVmGMbcM/U5tESjs6IIOjVVrn0rqWQeVOTR
QobRgm9+lhgOsIpJiHBkNS3ENWTYgUJPtviMbA3RCd4+5kKDVbcjc1Y7j4njWg9n
dwogcb52GiawhaYsSXX8HKfl7G34wjELAUQvSt1FjGRMlBjLKZiQTtQ6Gm4OZtwz
D+jD3FpqP0h9fI3njNpNY5t2v21gW6E4zFu9xR1uZ4ZN8G0bpBmchY248IEbEMYs
BY/0+uY44wz69X87+0cDxfl7dWZXlnN5cn6aqacipPrVyFvIaCP3q6NXKp7+s4zt
Rn6yH4KK8IQCfV6spCVOkzl4LaeGfu5wL90UhA0C68R78gMFD+GFjgU2qTkepxyM
+6l71/sQdHUV85hv1XyNRArzzz526uotLA2sb/HrTAgPwzhDKSDngmfxiVlVWE1Q
mNef9BOCLuv6dYQ/bI7CPb9btenClXHJNFtPo+k/stfmqeES35O3UiyI7kkefi1x
sOMwSCXlO5C97+Lf0ucrQwkXY7s1il1BwKQvY4JtfIseM5WaKSV6ye/IKzFxWbD5
0j4VYy4DHiQOuunO8d+jx7I517jB9PSrzRQzimANVsJWVKpYPCsV7lZqlPoyRlPG
pVh6/lgHLThpnUryZmW/Hz8qQP10ZuTKxv/HeWSKEugy//OaMlkXYl8wQg5yrTEE
Dwfwi2tMspuhAmj9UsQHOJ9eqDll6lO2/ctMWzcuU/leaAYAkKDOKRqLPmtvIU5N
qyfsYoJ5JHWXIvhzSxq7PxS4PYLzBLHZxSEZToNxMal9JWspTILjuJ2RtoixGf8e
RniN7ND0hJN4VmIDlFdigoDbTyGsZV3Xm+YIqevOoP35S6I1BHeZdzFHRfIAVtnv
1LMhj4aYOGBkihyzPmdohgSB282W4LyD1w07NSzVGpqxoDO/vfminpUVTwPssjnf
Y8DGsZirPpaEEViZvJMtDKGbqujd72Jdjn8HA6XzuOcTq1+bdxQWC7UGCq8izIOZ
7Yx6TOhCq1Ed+jxVAlp/Ls30sextD74GXHZSQIrMcNN2x4XRE2w2n5q2xxpKyAyZ
H6pjE8v+g9HYg65vO27ITB3LrRDHAb3WaIlRKnBM8jnFrcULagPm/4Vg06iOP/Rr
B5J42dolBM1ZnVAfvejKvOXFDmZe6NtP8wFEcHQXYyJOTfccLUM8f0K3krck3a/3
odEFY9zSypMETknkSjt0tfAUJ3FuYK/V/zOnjJ4qvOTzuhK4HqykC0Ujt2gWA40G
eKujJ8p7QvdN1rLoQww1AOJLrlcFAkT7XPZWWbVPj78zb2bxTTa86v6f81RKHr/P
PcXFGFHNOxXCbb1tbihBZCYdbS/IWVoMg6OMO/0g0cY/IckUv2zXdclq+JXz9Gga
mwAtbktXLdV1nSVCZGnSkOnjuxc2F3AWOkWPUbzeNwTqrqhRbUYmmybYDvCuYsyS
eMIxV6t4PY0BKSy5v0Er6BASLVUxV5pZ/8jegZx8iGdwc54C2ZnV+dR7ibC8P+PM
7wUCnMvkb0KCBXan1yIycc08hEn/hr+TCHMX/hvAwyVlAvpXUugsgLM+S5XfPfWk
XcAidPvgPpvvcECEwVJV6/65F2r0JXlKsAzn4f8MR8FqCQY05z5iPTpF9RaAii6H
m5h/f84TUCvysF3XjVJ9+XsevuOzNddUzJi0QQII1Hr6qqECt25stEjgDhEadHUo
+y//fRR2J6kgz+9hFjmmv+Y51/W9eCXZpEDPJOxhUh2FiMjSEveEpZf3epGAn5sf
UDsn/J26WaIo0d0+FYhIgkdLWOays7n7huVN/Tx/ptABACEOTrlccbj+CtcslyGB
MCpg2apXvb8OzwqtFlIlK4zBSX54uDA/YWlklJ0uWsrFYsQiQOy3jF74zbsnwDZn
e6TwXINckeJMIP1XUBM1o23TwddzaDgiQJOQ77AparTDE3lbMsqjqVFCpG5ozBSG
URyPBHUoCIP6M9YM33rlk/PCMzeQRe2t9DD2gMJYvd82+Eb1xce1C0UQezHfpfci
JNXWYEhLKaUxzacPOQAnfCotI9QCtaDcmL5LSU2iMJFqjKQC7G7LUWdRFgyqL0ay
smJhKA4NTbKtW2TqXMOSzBGAD1/VVp2goPD2rcbaQ0+hApA6q53ptRfKuFLlUTEy
SIGL3jH2ZPw5Nw0uZnJXlqqEVQSbHNK7Apnt3riUGz3kySZ/KODIcIfLyh/D1WJo
TofKeRYokFefTsz9jeYz6GjNfVvj80zrF3w1hYuyQ+7LKYDc9P+3YPuPR0+af7SL
91oo5ZnXMOf/tJ1ZbR8stMT1fnJzlep1Dea2Or2Jx7cdvKxCxoF/zAU0K6vrOu7Q
5fmRyqaUaDBCwdVuEi5H7wHGq0m3yrHSK0DcDtwiqnW7BnOqkNjDcrMjvc4n+nkp
13EOkmeldvXsFNGwCBHK7VVerajA6/DsQ8kua/UerUJ4xdJlIIJzch+o41bBOgdd
pt31+neqbb/cIE1wYh7H1bvr3FxAPhg+hWkdOjaqc7RtUlpuuwQ/cShb8QqoHFD/
l1iLAc3KM1xhiVJwmvDw+djxQEZ+pn2DVIptjP3VZ6nKFwndZLN5RaDzJx6fXh7W
NYD6ePLuBihRvFaLYy3LfkpVeCJlXQEJYTJvqv+Rn9pvpKQn8G4a1D9EuI66I/qo
ylsctZ8etsrkvpJ0ed/gB1WE/gKPod/rgngzaCp9+uvCbaUkt5+j629qtxJUp6LI
WP0OCyjI9FcH5hz0PRKvDrJLZB7a26ydBeMYp8LF0vonmqvBGJTAAe4hnxRdUg4p
tXf+x8Lgz2L3qnK+K6H/yvkrziHf3yvX+cNFcAOvttKnwun3jzTCxVahIAfrQfsf
liVnvIRLE08rsE1dxBw1gykdXUjEa4JGDxAa4plx/C3cMdCfeBlsUziEXaqexd5g
PzXIepzCl6nl3lhNtuUYQsWva/pDld0PkOm0KlUpB62rwZm6ZI9KThd5cw5xhKvV
hTl737TNNkU4h2LY/MHmbHgCmEqAJANTLdq6KNV9lsz+R0pjYJbMg5CIk3V03qOx
qbKAqURz+3FtbazEg+sA4Jr64rHG0eKTN44pC8XWZ5TLyiKxp/8PsJmStXE72LEp
1Zs7TMJcY9SgGGIk352nO1TRP80TFKet+xomOyDU9m6tjTYIozZXiP9vPFrvZBgp
TQnTrpgWWNT55Ldm/B4aTbp0VdNmyO4//iInLyUufcoCXADB9CJySMmeNsrJdEOR
Xw40WwAdW6lMXO9atOcuzRyCnfELud4LUftYZIk9JNYSaQ7kyhrvrcc10+rNI0La
jfzdhm1hAJbnHYmWQ3LeNtszhYdeAqAYD+X2UBC/bS7Mmfn932FF4I/nEXjvxG8o
NAnDEx7/PWI1CDuH/3W6u6+sZj3qixE6MYbxV2B5WbS0LMAT18/JZ5g2oye2kNzM
nmhy6j8ta44LZ7Q8ZJ5b0Yx7uWMZM8z0Ya/1Q8WoajxWihTT3661BffVHi/LNGC6
i86ODkg+n9T6y1PfgFzL+RCBaWMoGixhI/q6z6KYkWGJe5VMoyY5LTBEnpfYeLri
pkZXre8ZtsDMx0MspBE+vvFqnaYIClza9ibL0BbWMl2UBhhOOPHPH7aXMPNl3d2M
jxNT1WDlQ8YWER7m5TSzINA110YDcULiHpNWYsykLgN8gezxWgXr+Fs92PXViqlE
x6dBiNZqImjepgoNvRGxEfMrH5segvq3HYczjGrP/uVvYNqa7qEL4neyOfTpWrsW
6YfhPgrpayv+kyv4FJJl2w49DcfGKz43tYxbpjmETNQfDi+fO5+RwYRc7KrOZuYw
JhU643Kk4o9+Psar1YSqaqT7MXmXe4GZRDvRdEE+eWZ19BSI3WgvDh5dpIMUa0hd
JUGKFNaOjzjWV0xjoWEWpZmPlxcto/2XysFi6lriDptci513lgflB4gTcy+CXK7/
Z3oHZfgdtHmK3JAKc/S28oKuvfK/H07Q7onUl5919solGHh8WHWJbSUPdfMB7HXf
74oyHUbjU4RVR4K1oh0T7bovqOU1AO6u/RbfZjRkzIi6RiVDyGO+iQBooWp0X84U
aV8/JpwnKIOrrwduERkrUCPPv6NKa4tXkL4gwI8CF2qZXs+PFFT9O6SvlvcW9mXG
TYI+psk2qBxKFKu5QjmsBvXfbEfjF5FmyCkFiCUkO410yNmktf7qa39RDwBBbzL7
rLsKnaixuOfiNWwpDmq1gIX5uhc3cwteHQKoHMS03BWRX5PnrqN3KUxDNFsS7f5R
WaJYTm/Dx4GEVp/ZF9GJekmNl4yg1RFEYZn+W059YTHaNYQZHpLXkaYQYhpecmSu
`pragma protect end_protected
