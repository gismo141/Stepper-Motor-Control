// Copyright (C) 1991-2014 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus II License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 14.0.2
// ALTERA_TIMESTAMP:Thu Sep 18 10:12:52 PDT 2014
// encrypted_file_type : mentor_tagged
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "DEV-6.6"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MJRq2QScfam5mi3n0yi7A+esk+AvAiSYoUHio25go7NYSQMsdcZvD5s7g0xAZXWq
dphySk3sPffa+0FJen3T7lj+v2NYpgA/nFhEDJvF+8OTfUy5PxYT2b4/8F1JvC76
Z1snD/SbNXnhQrSVsgE4eu5F+mt5joNRug3QYT/NLrw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 12768)
uee+J8P7D8pEytGIPedO4XP7FfiC4yLrbJRtlyL5R7XqeFjWtwdZnXMMgDpZXYeG
sSN7PapooeTLWqbdclKasHqYSf55WOahek2PXITzBuV3JwA4rdDy/fvfTMYwOCZ/
LlCr09/451CLwfpzjgqKgLQ0D9yCJ7ZofP4r1ovYVtNVedMJkCTDLl+D9U4ypGsU
knawajnxEywlEEJ1hCI48EGbenK9CKmyF9eYS3RlIVL9/gLhTE7yKmg6RnTRY/gA
rfg6iI8LJ2Jf6XM+TpOXJ5KaxmBwJU7ruBg7iulmKH/70Videiu/8sNOy0yoYU0B
38VijK6dCNypJ8A73B7k22sGQ+IkGfwdyyi6yVKfLHIoFqnXZ8hHFWHQrIBgazRH
4t5QZ5XDvHnWdLcXDam5aUeXPm61EknO09q0EoI1tQEnj8rRSHYe+dRfbnOpcQ/L
l1KAxIQAcTSRsdVjlUCRb9XHILK9ZSP2ZVo4UaAmY4U9llkcKvxnWtHhR8lVT2zW
qBsPjLLJo+sqSk2hqslp9jHS8PajGxcU402lHlop0Rtj6s9CnhJnTQzua1Lz4IV3
Klb9Kpg73AX/iIcrR3TYcxl3QKvSNwk5X1mgmbYQXAm7JrSR/zGYbhld0ZTLyd3G
S3xzV7A9d+YG27toPahmVL8EvDF86O+9zJTY/tg4CZjvZDlbOD6xQ1m0Y0iRoPSk
OZ4xGsfFz7phhYNpDvpiVUAUPaHj8a+7tlq+niQs1/u3Zgd3Bcoa9dWZDXhhZ/wv
dCeCtNLVFHBnMdrpHHOKLGYHJLMbhm7Ciz9xFNbQeN+F0uHLgbLXRsIVfF8LydIG
Ur6E53EOwBLfQlyN+Sv+sv3pi/F8B+kweuX67NFkdqvoFNUUd8fj1R0cq39LdQdt
VgsxUm9Tb4BwjyRqQ+TWC6cFp7D3vSqWfZtBb6uHiJaob3SO/270coLbyMyu3VC5
grGF/DGajSO6BJjpLOWnQ+zFFlyYh/O72xFtgLRsimBJ1R7qn0N811cnr20rSDUw
E39UhUMPNSpFrRQXIwD2Po1wg0PDWYUvX7f6DMN/iyzk5r6kjgJIzPPZKO3iWjak
FTjqexYCrp6y7l8AymaWGYlzOMAeOdpmgtmAJx3Gkkkk3JghSFTw3kti3UlTt/Pl
xrHFCSH5uCPoxLsf76b5HKB7OHREAzccLKrHGdmjrD6a5+azvP8osKdK5goVlNa8
gDeN0NhoQItsCbRTlntbdE6zA1YULfO/VAHLVP9d6/YfdlwVaOaOjJGlNvA1kxQF
EbO59TxRNWHjEFT44Ln5D2Pa6DCmjXaOgbmn9gjmbrVwY7nWyIu02B37FVogYGLS
R7TppOUGOmPwAx9uofkV4LSDQZZuJHHX3ugr4MVwTjKSl2i9b0HCqaBwnybScniU
/yf9qMSsTYbkZJY/fSmK+QJd2VbzwBCjJBtIsKPwZmBa660hl52Mu1PB+hlmyUx6
WFTlj0A9BVH5pwAxvduOddOteEuNCTaYvGDduXFdFg6xvWs/0G7OioxIF1faiFKd
sLW8tLTdIH30WV+BQMrY0Dfc+7U/Sl26daXsXkZ8vr6C/MVGkccxa7UivV/K4tpZ
2RUn2wlUtBF6SFfBDRKmr/whdkcNEOZ/Xu4DH72yz8s+tdbuujE/WjMy/GREv6r1
lCkY6+imf/zlXbAttlzbvKF0Yk/TvjNGiErJ10NTPTnbfGSCsbYclKDlVeDsLHaj
kj3QdlWvVIWiyLMutopSwGGrUt28Zap6Uh5dBOz8I18k6c4ARy+/7rSfGsnFxp9F
vtdVGQqFRjTL9UPW0+JvOZ/wFPQb7Bm3r6WbbUBLyXsrgqvl2RLP5LB6h6zeBUQw
qjdxDb2nQMyfNez1J7zVVjl2c/sB0dx9sWpMUAsteiMRe1LQEQawU4pwQUAPc6kW
JbZ2pZCOx3N72pLx/UIQG7UlOHEMuGL/w5fmoIeqlZe9cHiDCnYY9m5W7mEPzZmv
WLvwi15SkVYIWYK0csJkMz6og9OMzfx2c2AZ3q9z49Fpfcvmnc7j13rAfGnJGjT4
+DvCDDkl6YIFd6J4lD1R5rwa+OKxOgl3a8fI0iGj2kMkK4jZKPOCvi0MXouIkJ5+
IV6UGmvIa2Okv7aL+FyTrK9Y8ADWvUY5yFaGbbEhMCSk4wQzWp7TObwQeH7W1s5E
ui8P7GKYY8iJviYloc/ENo4pQBefGmqhI6KFB/gJliuIR7VuqVbC0Og/mo8v7cGU
N3nLQ7t1a7a/TNN31zufLGsavmPJ9BXbLttzTVyu/bGrRhY/KeiHms73devgNlvo
Slu6fJHcEGNQHvZ3at3hGXLUjRJhTTQbsz8XmrIWLxi5dWKm3I1CMPleCwl5n5e5
SUDxu4TStwr5TiKFRtx5D/SKv2g7T9ZsltPOjFMnyZ9rStmz1ibkgTOkqBU7Bp/X
OTapaHFl/rVSwCnyr2WxcblViKhlQdPYR98AgRu1lRRWee8cvhHkogdRcRxRiDrE
gkeEj9bJE1WYCG7BlwPqlWAWTGI2/2cZ2JNOvZQAHOFeNBUyz/Jk8/trzKhWvckE
+WQu/tESyOL6JzDjMTE/XukeJbStc3zErx6VUd/LBSSO0JJTCRstswNclwXKONiZ
2D2NERDkYfiK2JEXGwhw7e6EK0zLJ1EdmjnP+7+hFresWzJ0BakdeiZhI1TOiMTj
8GjKBkVRSK0WYTv+Nu+aUAZ51TXoHZk4zhlldlK4lpaOE+N0dDSCC7f2vrl5drf6
VW959FfWLKSwh8luO3FmFEpSwd0zkQgO+bXqTdsVBS3yZY1aMeOzQyEKqwOtnav1
82rIPyxX6Vsf86+G98qE1mRswAU5EeUfvR60bdOHynb8fsWYV+0zXMHdQh1Ig9Ed
zwtmSw2kYiLH6//3hlwGq2FJSatVVa+b19S1JJp2aFYpAVv0Ugcb85trPt3San1S
Vt22iE0g5CF5auqofAnisbISn6/RuomJIx3KSmPFUBukjIePm6IeVHq1mF/kgzcw
ArpaPao4PN503iWsaLiUwxYQlzrmTLbSXqxGsH5I1me0kchI5Y3s6P7oUBVy8gSM
rZLsen5LtFgArS5dgA7ApYwKCieJfQ4XofGTdP/YFJoxQlYZ4eKBFmbXbqz0+XJM
vQdL89sg4AnfZQmGFB+RPubDp6qsoKWc9xrL2/j/4hfqJwCYeWC/ZhBNds5lHvMB
dLVKg15p/t2bz9fNw6p5Pn1EEJx3Xhe8e41KxbaNjAoCW8JrkFpvGAw3HZewuk5n
PEh9fAHjXjx+XiuUApTkDGLkP1W1AUIudVbqMjDJZ31cItZmW3CJ8Y1XalPFl7rz
LCdsyfPCFAuYPu7Md9cRO4GPlP3yuwT1v2nqf1Jd7BgTHEao0fJlxVy9hiysfruE
Y0rhE0SJawx9PT7L7P/Y+HadIc8Nx4j9sWmFz6jHgzp23k9a7U5NTm62t/q1Xf4V
IoQCHK9BUBgPnRyS0NTvm3hTh8i4CPu1RoxtHSgJELOILJ9DhX5F2lOf/jEX4eM7
VkoZP3dceQTf6+krRl6kE0WRQrqbRrXV585LS0tWIgFOGzbQZBUIMYMNNKsqm9jY
+DY7/+Q4WktYGqOMQ0BUL5yspdFusiylW/atkrI2RTKCPQ0Gz6cEsW3kSpiUDZER
prZ4dcM2cbYwMI9BlIFA8hPLallQSik4FCtHB8z549YJ/0LtrawKxn2IKdBBXdIw
L9Klc93mJv08GgInRfP6z/LgXjhhF9mgR2pgu1+B+a4QWkFKl8TTELszbQgfChIz
UPzXlo9rdj/wF6jEby/3S9r8tP3kNejR2TAQzPUucl6+CiHUeou/OdzL66OIgIFw
8XqFJkq8Ug4x7dgNnn1DOlEXqMbLlwMI5YGwmOhOGIz2SLt1jx9evAF+hWa1Hd+7
enw/V9iCcN7bnpeM/ZoMJNza6k792M2bYGVvQwni9nbwWJkjb1LoByv8kP0gKcfk
1SrMaj0/ojVBliqzIfuq10awx3RWEcjY2Mu4J5h7NE45YuriryhdBKmwlStRs8k4
jWULzPGpddm8N1+P7/jU1oGcnJldG4KkaKtgTSATD/2EG6NNrEyXOtb6PuKK0J26
k7a+XGmOP4Ts7vg8NZtCE52UfdcDaWooN6WzHLoYKVdB2g9PC4tqKGB8/y5s0fpw
vCRi6pw9M//+ue1kdmBjtQQ0WxajIxP2Ik4yYbVq9N7dx/QMNU8lqzOu6zcNHhTt
gy3eSbvIbQE8CvyjVA2Vy5ce2dD7/PYF+E1vJQY8pN68QopjEdsllV2UrRDoV2iv
iZe5CawPlzxv2HESlTHLL1yWyYLqjD7N7yoN9GZj814RkNHzJjCRDMwTKNHr6Td/
Y8ND8PrOWW6lYZqL16Luvy+qHMGjV6inyzDScKCWpYhjdcqrqunids0BIwiz/qwo
M9VH7i+K5cO1V8HCaeCBlA3hB9YLvyO+LXMLTygLDiLuLrQzmn7W03iN8OMNFZWn
+BdlgYnq3ZVv3ZCamgM2sDltyoOtbjzxwZvGPdCxd3L4KqOUj1KlKZhH0r1yokz/
FmU+PLCq2O2hZIhNrSpi6mvzHqAN/Ao51/mqTLGhgF/LG2daNJsY+qUC+r6M2Tav
OizyHKA9NBBFgf3V4SK8vFlfozohqiJaUVKigSgdOl9nOKNarznhw/gehHmMWBk6
V8KAmoooUjid+KHnyCYWR63yOjB3/MDICS1P6o+IJT14/XcUKBD1kBtOp3QSOxPs
ggUFd3E9JGXeLRo2njsMTtJeSdZ3dbz1SZBaoArdv0mF/Ww2syNc/G7p3h46Xbw+
PRgpqYdrIydXiVHseElYXZBZUN+j5jDPJDaA7F7132VXvPOAq2m58iOTie8010fH
VD4DXiO4OXco4iltwVJjbbtrTNTWI8eQHlei4Y+eGS/dGPiyCI+U8jIOn/+Sybcr
QVYaNlSaaB993QgF85ChYmW3s1bdnYI9JuP1P628YozMflMSs4Ec6u/7L9Itod00
DRSOaol0z5EVEPPdwD6WqHmGgBL9idW/fxRYJR8atOW23OjMLHPAi2acXxh8Am7s
SmtSNAHg30HPCnhGF1edYXJlcYoJ9QYnHyqq3Ww5MZ6YxeN+IYjWVZOQF+LaDD1Q
AUf9fJzkZh1QjShzTOG/RBOlmQtu6rcPDMg+8lHAm2Pdc0ENWUt9DaGm7OeYWAGl
1G8j521s/s8aWkj7CjQYy8tviT/+bVquo971JLfzy2zcn36TPQO8Mx7tI/MmpTuD
tHZYC+Fcf+Er+akaEQVLZCNXfrETld8+tn7nPkQ7jJE0Pn8ZrZZsVSJB1GSWcTNh
jwJUsYSpUwaS1iqJnopL+QR68NXBTQ/uXZHFacfBzYw258wD+1B0ZLFagEUSAWVq
knMUZikTWFexFutE58p69UUa869m2B2XVMZ5jqDlmhpBzrZT+83pVfKrYIE7dvgw
h1O/oI2ExwFYRNxIy/StHDDJ+fl7EhgBCoKwC4GtunQ7i9lX1IQWtvYk3ejo1YCV
uvFTHTePNSM4eYfrURy8dUGf/l06kE3b6shN5FoSwpM2HKsEMxh3U3iem+f69M8v
nwhjd7oHIb3s0X5nyLnAi/k7XmPVRuL9Tvw9IgyYM0ZAZ669kzRxuETFcpKztXxa
GGLtA5Zr4b64z4jCutTtyy76Y1Mxw7BCi7JgzBtMcSKl4pg6YCfBuxdgM7FQ7MZb
WGKClWokPCsWgtXBGlRAIN07JXlNNGNun4fUqGPlx+OyQ7IagytGNdw9u0Hi8kKu
3R/JasbKJKHSYlgKnceAv9Tstsi8/dAMEf/5E048IF459Wxvp+BUh/xJP1jdMzZZ
jP+wvIpiKeKVd9MRu+n5sf6kwrkp0Ol2a9JRmHFroFDSL7MVAuMuK4lQL2o4P1sD
DdKHYXhY09Yk7uI/BdIAZ+7nJZRLkB0aCeP+vl7qA/vv9Y7UPTyx+/bxovILANpa
I7Ym9W5le9OaHhXE6mtIh5Uo8xNy+LVrvIKhVOS7LXGYBHIUMCBaDf5cMN33oaJT
oaTqXDApRIwXy7Uh1/KavIu/HBKYZ6VBQrwNTGGNNYu2+IAviniE2t8B4dU65eVV
UBcEb7bgrBnrjuN4Tm7s9IbNjfu2TbeCXK8VzJ0frPWg/h86LrvVdpOhp0wVTuos
bdS2XVsf1f97rZyTTZjeB/w1YT8G2GJ5mpj4JJ7w7fkIlbxDJ9wIMfVOprEyRdaU
55vxLH09ALfrUFlXEJck6RkbBVDS7TcdbtDCWbSEF+3YvKo8pWu5GQSgrfsSYBso
fMl4xSiociwpnWQIuQ6ROlh3CtGWiS36rSTpep9MJCcyzTdpMA0LXLwxbcyWRMTO
dunnoDqq7Q9BwKpZ68MlHbSmW4c/7ZGW9GapBEsb7fNnNK/A6Rgpj5afv2AK2SYX
sOuGYgSMgxWz/ddXl675epm5ACZaMaUl4xNXt0LzwXmRXhzqrBYNN2kNkcSFqlSX
ou6iOh/pGJdQmiVSOqXd96qFS30b+5ogRCT3jBx+R9cu3QL6+SB3PH/tqICek4uV
9djz3KD7zaAMnT6P6iFgLrasNVPYgLGQAzaZpEbUo/mhQZf8/hLov4+xtMnn6PJt
8JZFwRdF2PXZ06az4R+3IxwLSp/LNvmj+Bgl6/C6bGwbRXLjtIL0gEUbMhoapxXx
rGUOo5h0yTJBBMt8xiGMNcMx+qV/PYmTazICDyr6V+UGWyThvPG1AjDLsh8n7EMC
ddjWUxSzbXEePfN5ZTKgO/2JT50T85rb61U6X3mNPemfoRIt0RE0BaySZ9bQfj7t
o51n8wnD0GsGLiF8DzLQI2p1x12Sr0MC3liSr1TivA76wRZMZ3d8jbmn+/xbjJJm
FIy2m39KGnprnTsOgslaBazp6dGPY1IYeM5NXeFMrm4l7x6nZcJ5xoMVTb1BstqS
SiFej5eRyN2VcMYPCnc/9dmhcXzpYLv2LYrIpBesICe7chbmq5n1CVYiNbzw4LZy
xZewU0gEy9yw8KUR7gRRfxuBLOxebmAYaYFHzFd+fGnRMv8drGQ2VCkhQZjOR9AK
kSjKzqhCKDHBMvts9g2w+QSbSHEr8ewxH8g3FUOfomVAo62BugbUu6tiI0WTGNJx
WVsNhc9H6YYzHLmuZOZAJ1gqn0pt8VKMxOe505CN6/WJ3US2LohOd6Z2pe6+widw
4toRx0QP7V7fmP/RfTRvh1MS5s2xfLYZjKhaHgnODLbhvludGFv9wy7HZhzg9op5
YCsBEIp8wPQORsGmx0Nu0fDNmHqzp6bGg0PAJTFjKx6pfNI4qpmzWisruqn4v7Bj
ZhKySKRSJiX5+EaMdjcQVgf3mvM19cPENFyDZZFlJN3lUg4/hCxsj4zJogDBN2PF
jCGRWaK8BCBkWXNfO42QK8lKnyp0XJlkVbzp1yKw7GWY5P1nLSAjzuVwDQDJxmjC
bkn1ZGaOZG9yf+N/CivwzuZAk4SEyFQwOzBwp6yys3k1LPL/3ql6DbD+ydLJI/4J
k/IfGcra6pdB4N8EeG/u36SQbC7dGgTVmHdCLjZWqApcZXH1aOaiMyToMwciD0vq
Hwt61I/6ROKTHgIUNkRhHOwlELpsKLlQjjsd39ENxhmuvSki1hyQv8rSx2EbmWk+
RlQ3vZt2wTamoTzlNo+dHSH0Z+A253BnrhfBBXaUAPMHLqqUBGrfu4exwEjPmdkG
9N4bkwtAFPntE3Le02IItGRH3jNQPjmsgPeN2wzmOr4aqrEpxjTwfmBxxtJX882k
1xqy5gQ3fa/DDPrnR256uDtBv7XhPb4BYH37H0nTWxlnXWdghhHIkeqcnDHVXmSS
ce7e+yHq8pHed1AhqXhdMDbFa9dfQ5GRusJAPrlyHx9zoHwt+qeFm22L6a1Ye0qi
bP6oxquQLJEpZInBV1+N+F0nLYYzfOJmIv4aovDZlz5wtQxNhESbLlVbHMfaamB2
oET6B/XluRLB2zgtZcCzJNmk4aD9OXnX6Oz82RE/vbVMCrbrm0Gv7V7SQq2QQzM7
wcMH0+diZ0D7HcDFwfWAiK3IQh0P81EBWsJioR7reWDfPduL2VPSqbOEh9ke+8E6
EqxsJkr6EsoReEU6HnjohtjiXadwxWhMPuq+/3/CxEkhpHL/le4nX1Ish/UYXkJQ
W/xa1XQivuj+fK12MdrWi3kVuZpdFJM2z/q/A1fo9Kqu8fMXqvUmprxsC5amAnIy
QbwdqTO4JglFIelDen9dp7JNifqDQoha5G/OU1KnFwiwbmhIUGKc6f/t1jpKqMih
5z5aOHrcYvohDHHuUOE+y6pokglDTimzQaL90LebfaTrsJT2U/m7SEqv26FJkVYU
/cjomOqmzQXZh2jmwG0xLPDc27uk3+UT3QWy0oTRuE/Tp4Y9QsuZ2/hL2xlfMtUq
V+Hw+vlmGkVqJhPUlJ82KsEtnlfOsw4bBkqlFzO+x0cTDOyS9PElpFcSDiej59Mb
F7tsuvyTJ1WFeNlxvl8SYTvj/BxeNr0i+reAghY3LixDXIgnEux6X0FVoiAMJ96k
pxZuAKkMKcB2BZLz6OmHk+MaLXQQM3nR66FiEoTGsW7WZAK0YcZo//gKDXCLkUmv
9UDY57XrGi2T/pIDjUMr2kitJ06C8dLltzOcZdDXmxlWqmbWrPruMjo7SaFG26Fk
1qeCuzSLETQMwFTadClCaGyf82XQZk7IGhcOnKxd8Zy4IqfwLS0tDEcysuuVcwZz
5wPYZIj64OtTsjHU1iMf5OVCETIKRPQqIncVRQFNQ0T8u0ecifkSZebxN+IUvCME
6vm4ZopQ6lTF+P5I2zGefb5Taza6hOw22/D/80hbOZX8qhudQNI8hPKodhxiKZkC
fKkg5pwOnvcjbjvKWd86UYrW87bkDvk+VPTC6WCsn3jvRqQh1SuYSv82df93GbSb
AIbZvCKhlHqkK8vcAlDFjASyHLon2BUeEoUi5DUHCQiq+QNfduCEddPLyVy5mQny
IsVgfIeXicdkJYFbHqJiN6+VWFQYF/fsW+s8LBe0WkllD85LAFzY0f+hz6wOjyxu
UI7O5NbH1blL5C8qC5dr7gqvcmIl8Yot17HAfNWJ/vLvI08bIXk2Qk9nIBPSIcWh
rC6QrAV+Uu+CVzx5QOhidNVPm95fw8U/YVLra8zlOB6gvM3JLOwr1+KDGHkjHAJR
+WNawbEEvmt/wM5WuBT6Tg8PLXZKgITlgDppz3vUXZCfzOpUHkJ6Wl7/Q3F1VdwA
a0F+MrDpR6LHq74FN4+e3q+KDrfxQnOedVCvRzMKmaZ5jKJlBsI2EuCd8BiYea5H
KWZdnnbPu6ljHPm0xNgVMjiG5/LQYVaoShZgR+4a+rpI2lClH/Z1LkB1dWP3aCOv
i0fCSmXNujFv/iIcbx0mzlfsUWT8hkLiElDIXbriJvF1fj9dNLWXodZ5Ac/b3w0+
Iz0fe4gLbAzod8bymBuHAYYMOECP/6X1eGMUbNKc4QynEHVFeXbgM7SGPbG7To6a
NLMpEKyyt4pFWf2uSSBzhxHf7DjU9nJeV4SjSN19OOrp5eWE6xEKZuagSZS5LuRW
0nfhL+0k3l07h53gabDoqcwBHNmdRIbm+zrt1/S2lUuMcUrTGCK7wH28VwtXmBDm
a1HmNe7q0Faz4jpMa5PfbfG5ASIeOdA+PjtSaaR4flxKuPirAQNG0U3H8aYe0yEY
1OARCSUZKyMxVca6WEvuAmbtYikvS3MLzOUxRbeqt9VrBad6ABF6cLaYzBYnKyCw
xapZBIkSKu0NTFXIoGF3VIHo4NViNK0H3WcbbnQBM+ZUbPvzEgotPArXxJpPfJwK
xMJg/JYRYd9ef3evWIa5zT9exKp05jFiVn1j1KPdu9S17Kb825SKBC+YIEKlfdez
DihBcOtKz4zbEHxDoxzpte/oxC642P/edjxMIbtLOdwJFW/+cKe7EG3k4hi7AJ0j
m6yUJoT+ZTh6NjcuiJBCJ5K1GdejHLMx//u8jPf2l6ZZV78kEoKbYiaIqryG6LdQ
Gjrlt1gasTbavE3rBUu+BxJr43nQNYTtc3PdIaDXndph0IXXYl/CCOeADqxz9q7t
NLGd9MagCbDTs/zGYcT9p3+k1ZLGz+HMSv2oRfT6VnSFN4rePar/NaELIjG09r4n
YWUVFiyRsrhT0Prd1ohe/I3ITKyH+dYmNL6jJs10gdheKPI/mk6xVza+tcLALswW
rF/mhZK/9soeE4WuE2eac6H59ATqdbOXmNNDmUMsRuS0Nc4kwDv9x4BD/6DkKaUP
tDQFGL6odYhyFVViPGekjNi7VH7YWaGJFDpsKGcOqQxVVygnP8iJ6eXJ7Z8Opitk
IybZyVs7ZT2oAAjCyEj0ATUE928sCbgML1QDP7FDua4FrfKxbHlCnsHkgy7oLios
doPeCsAuN6Qde8YOG3lISmGQRUS8g1xxCQUNdmEDSWBHFlDO/XkuoYgCXWK7ILce
8IqL287HCpZCx4ZAM2UDBeHzgavdb431s7O8Q/Ba7GmimXjf7gBAvl1lqkg5WaQh
ptBECipFtoMoTBajLAu05DrmaQNX7jpuPrBtU48eh5RJse2uG+knDuHOcK9WkG3T
9NZ/Hm8p1jHu8rJD9nCGISG0q9CeYGtdMcIoz1UMI5qKPYbVgBGKqJICYc3h4gnG
CPApKPJncJh/mefuaUMIH5YhpHp3Lz5QZ+MuSAxNX5FjYcF55130inEuj6BWkvjN
wZv2M7nr8jqZJpmFGtnAAK6Vzn+vEY2MRkxsE3cDZT44j5DI8b9VoY1CXz7gIuAn
ZWSIQ5tzcf/RU/rlICXdmVmLcXbe8XkKp1EUfzFYemZksFaAQyVXPphDNnutZ1UO
2m3uifDbZajX+k6FhzTe5G7ePlFCRnYIuOS1/frdT4Rxt5SvSMBB0o1YTxajTy0L
smNwyLqp6w+POXd/AQwLwXlXQF5WzpGbOrYI92vhj0iLJeAq5QiwMiR/IMUegtg/
XAx6isLYjmtMZGynm7ulaWmsYGmitwhWALZ2KX/DAh9F1cr0EFlry63vORv800If
XM0Er31nYwfJIivgV93isiY3XAVupVO5jLO97ajUjMkyslEUFWs/BspmHUi+OQMB
2qSlekjBodwGvHNGrnKh4G3bGXSedmgwgE/DZrbp/VQJKkBFlxaoyeUOJtgr8bnX
4m1CZouwrsls7JMchy1tZ1A2FF0+XvcIDxEtMX92R6Zzr75pExU4WjnJbPt1GkXo
KS5S9IUe9WufAi2fwh4tIhmGV5VevTwU5WodpWkDE5srpzUj7RIbUQ/MdXpyjsbZ
2Ge5cmQ+9WZP0VZtmKunwEnselDGcwC1+K0PfrCWep4b2pyElakyj83CcjqUg5pD
dJt0WLEkUAX1m9HlmrrmCIpVgeQPftv3i49GCoAVm/79RrUplLrYkmjRuX+arrDA
zsN3Q0OuwAQLd/8dAjSELClUnHHQDfn1mKkGpheMnaiJ/nIhGNlQqe5dmi4dyFbY
ftHBkda3u6RsCbOmhZeJe1HYsFrZJQtM+ItlbTrkpeo0J3Dz8XlraYs/7NSOsZVl
Z25by8gThi/RWl4TX+E+/hfo5fjCKes56ftduD1o23SvpOBB6zp4AgIgFRLtgNSE
618jTiM4OwzRbrc5kw4GGU5XQ2mOwWrwHUx4Fo049drmiEuLoaBFh65eZXqfe2yD
F2YHmRj7GTn8wSzASl58dFsYYVocxY6cjkJ4c5NPWR1IPb5YeFfePvoFBbh6BVR6
xGvviZFtg4RGXKZgcJo/1gp11rWFtOwgViF4KRZ6WVqxydKnvbHpkZtIrfQrbnzW
xblfSOLZxDZ9OkRC++SxUNAlBG/Kei2IHG0+R/acVKQrPlVs0bQ4d5umdQyOeduG
x6GMLrnWGPuWVFHcUZ82cqjT7qd46A6wgE2JULoUS6plQd58Fk0tkQW64QVYKirj
pwQeACB6c6wynLStigfVg0lCPbwA96qmTpBJCp6d2z7RGac15OQCsg+ysYbEe3rX
AIFA29P9mBLaFXlD8H2VBbaA4SEjBq203UzVarQGENpqAG1du+/Qr13dKEjMgHIB
Jpi+Mrb0roxSdFItmX47RHA+k+VYW5+gViTZjLkIHGQ3LHfjYUBrzPer88fup+dv
X71LQKqyRouv45Ag5Y8PpTyTP1y+K2R9HmP2ejRTqPgfr3AIoeiYf8M/q+0pKin2
DY35HjxomsKsJ2+HOuiPSEVoyse8qcLUmUcLCUMCviRUxs7YwCX8qN9LPwhvWo5F
YKw4gf1zSsRJS1klvGqL78ocgV2t112DitQuubHHF9gH4lwUCH1t/4NpJkYLfNVY
yKf8uTQ+qolYSKeo7CEjXxt9mzLcHRdBUiUEKeGDN8AEjD+QDbJbKBPkHauF9TWO
puiYEjDTjrl50SMvPyxTzBMeZJyqmENpVwdhzyi8aIWpYsTYWkb44rIClHN3c9JJ
8I/Sg9q9TrmX96zBKg+mWM5dHJSlbCKrmmqxzs3zG66dLZspXJb0Cletq9DuKMnc
zbeBWl4vPRkqjVbi1VWo1KC0GVPvslSEKElb/ZXQTQle17FgdvWxzl11eEGh4tT6
1oDEFH94ZKczlksQnnvZHHn/LU2bUaYJggcCSF7qAWpYF/g+kRR6/BbxEsT55nlu
+37mY8m4HtAUIvwcaeqlQuPxx4w4yfwXfhtsK65pT5cwQbwHd+kndUfc+TNVnbzA
zvTH0TtYZY0GjlzEcjzVUT+KRQsdLfTyQA74lB79PaPPL+9jia230+7TQ9PLddI0
7+lzNnB5rckEeQJ71oSxvVMulAzgETQ7pGsBaJgwl0bI5ZXhCBH4UOHxlCsSq4Na
B0vqpXh48NON8++J+oIdfshbvF+DdTob4HAvC1ymi55bIfdN56+v2DoOyhBLKR5f
SGm9+VFWgYT0QpOTgMqSQwxASExkKliuoe91CwekyOqvRbkLAXGP0hTPmNOXQtGB
ENN3E48JRPb+uvEAkcp1I3sDbMScwCowKJKxJUnHHLGt4HO32z8BBc68lCYdssXX
rwYwJ9eGQ7p3dJGC9Iotp1xkh06Ombv7ySTQh4lv8xzyc1TSkz5fFuzOtFJvatiW
2eFVcxTd43MRq7aKRaaxvvmfRGfbOxrcpgPB1mt4xxqGAgQvkkI/hz+KPsGca0yU
t9s5r89d+PIzSxlqsyih3wxl9Hvc2xLyj0eDLZvjVbVxUJsDYHI2oKF5hdZ5ElqW
Byzzhb1kG+kdWKoygH54zEsIxNQmbVbmp4+2bN6NLwGa9waFQ0X0sC1of1dIupWF
ysON8bZNlb51rYInkPYbIdzmFGdlqjGFwgY3Xs2Cc+vCH09mYrXLOYC4n4WpFMpF
wb4Gv8OqdF2fP53CLhVgWD5iccHsUlOINusy2XKPusDO9OdwTpjhFKI5IIBTHSAX
dgrNcm3fxKy0RYUCKac5mM3lujeKOarz+ZZ6tGXjhD71752sJ6A7uklx0DYcfEpj
ZRd42XdIgNR5znMJ6kiY5/8Y8eWjk2dgxZ1qyuTY1RN4vsk986lCKUw91h8AzUZE
d+Zhzs+EcC3+dUqlAexoqDmaRvFtNoM6Ve6WgfJMdWVl76SV+3yus0ShMklrJsCg
Lsg77MQLlQQDLXxJ4jNdGNO+Y5lZtjZhj9S2L2YqeixNxRW79x5mk4piCd9M4iQx
Uvk7XMgYETkIhvr8NHYaXtzX18wkbp3yO8Q/Ja1eELw+mo2uvE++dqpwcJYJ2ZyR
TXWpWVdqDBgy79gUJxI3WjfM7I448g+jORNRhJVHGWP4Kn81iDrr7D+NTCp5V8uO
q6V0aBGQAwJbcZCPaTo9ozXYTDKVBO7wJAG7Nvg7q/FyZuFxsrZD8beB7iRX7bdD
tM12OXlllj12V/ZSwwhDQTSRfrxNA1Xjrt4V8HKUsGV8VoHYfqcvnxMn0FG8GIcx
woa/Ldw9QVhYYgCEobp2QLU/IxBHTcKZmIQpjiywlWfHevVZ0V+St/LgfqWcJqsd
0GNKGexTylup37DWNqIhuJ6hOBxdg4Tu7SzwPdI2hi3YOcwOM3GN1goyhRP/wcay
u+6jYzBL7NoXj+LFxsZlVSgcSge1vq10dM+3uYVTnM5hJk9XDpPcgpOW0qceLKmi
kyBGjXTycwbPIjps67ygYme9h7SWHmiAhrbLMXkZJgAvYjXfUgRx0fQmTj79SOyf
cdRB/ZILDqxr8eNU4EgsywVo00oSvznL15loW24/szYevW7Ii4JXUNoNSyR4jafI
VcNW62V2GvimzX2sOXDDzWvAxrHUng2G9GZY53PqtiRQ6WYA0ZZZN0oHiCOhr7hY
s7b3d2+GsVr4TCXlK5OvJCGmp06njfm92iWwdQFZXGzTPRH694dKs04LGCoENKn+
8ArDwBx/seZgBHo7LOTNzBDQgPfX0A+nGnnT+CKJS8gI2VSU7h1aq4cuKb88692N
kaJ6tLecAWAEP/ffbn03t4wk34egq9Sr6OIykQFO0Vws9wwvWpTvVqRLzIZ2WYK6
F+jmAefBbYdFPQ5dUL7yRli1OqYFMdCZZXG/Rwzue4sucpNMAkyiUJsNj1gnODfu
mOzAMeu4LZaUbMBjAv8wqKCX1cTWY5dqpY8BLiBLQB/gKq4fy3F5m2PASlVQglg0
xbOYrMSiY5gjhUSnaVEQ81VaJCyhBb8G/wV0gOfGfB43xUY/bcZFGbMY0TaOHXJu
twnFvUMo1a0cu36wrh9vYf0R7gnLAKgM4/2FlOPd8pQ0FSsRurVDaRgc4oVOs61Z
s7OcSsJegtrsab5EW9xlX7DQcPgBK6xJC5rQUQIiYRmvwrdLhzmPNfkNZ2qhCKbO
GYC3CdKegkmIgXr/0dUtI0W2+m2ijRoAyn5rZ8nD3/6EMkdZ5D/bztY3qMqlZfgZ
+9V3pKiZ9TAaJxmnD0Lww9NyiySNtjoDbVPdGcYIFP11a5nvrAlCHW35Jv0JKGIw
OqlmIcrSiXwj+InkghLBydQ2XGDwwNz1hNENmWjCdoyyBWR7vNT0ui4MEkSWw+q+
GHLhG2MTEg3BCmVI9BqMt1aM7wl+9fZksvGjrQyJ/db5ls1XRPOO57GMY0c+3K+d
dpInGzUBTQOEiyBW/BJ4WjXwek4POnUTOHydo20cm+AajzvLVsWINoTLuDsjQrN9
ZBMzIjHnb3ruFzC6ea9X+WisKYufz8j/54ghUYN1aXO6BiAu2P5GAqexCHlinWMy
MmZ8Znj4AG+UUoFgELwzjkqRL0gGvKIRxdul0nI6wDTNWc0pD+IvLaLF79FANVv7
55WWDKyw9qIqzm9neeU2wHTCN1WhGEcUICCUFlNqdWkJUeWzEy7n8cxg8Bd4F+uw
QCxf7+GcZD3FNRPptl6QW7CpzLZ6B1Rj1Jb9RTnuW0oBhd6gI5xXnZXZctIqCFUy
WEx52ckzaZ37ffsiGu3SEk3gnOcDci6WVZ0a/Fod7izizuSwJ1vMKCTpdDNPlzU3
bIrHFZBO4RA2ga23h/xnwRUyFhjud0Z1cwARlZCnY+HF58kTBTpsB5wXMLHw2HSI
JPoZho6VmKofUJOFfOSPOx/kChHewKUfGa14sTaAzFY9VwQDky1D3utUaIdajlJ8
l+02toy5uqAO7iFblkWdpMherer4AE2ykCsCaqOzt0UEGJ031FacRMYIonwuehZ6
ApurHO2HgubMxYYPWE4PhHxDJD+KvJl9XS5mKCndfIqtD5ZZzur5Qq7Dh7TdDyRk
b+hm/od1y/LAMpXwEMj4g3r/Djj1qWAHV0XIznj7imemMHP6Acx5KyCI0ZYeZQz3
IY0JshWIUODtwN63GbhOP1y+WWva22muMOfWhvuz6Lw7CFks+nS/mXwNhz5vhXeS
q0V7qgRehvXNCw3HujaI8AUFPRJj4k91wqhmhTXc9NwiqWsWRCfr349vcG82IMcC
scX4bRN+r/9o+/s6Rk4ee+wIUd2yDGuew1UfvIoHD9s4UhXoLVUJdMPIU2+VBueK
TFoKBudKU6DHaDsnHo8nVqH+Bjn5StGtDT60y2LdpZjiHhoCMIqqXgzftzBtaGr/
KVcgJuoAhAPG0j1e+MegwDw5TTPkFuD/WIJp4/r+xjABTB+osJvUMBnOyJV2z0U7
Oz1dZq0IguLt3sg6YHY1zCKU5azWeA8DGYH8nXh8xi/vc/5ANKm/tVMLbo7jhWa+
vhjXH2wZNT8Pv9v3brZ8SVc5LqorfrgU77I1eock1MvSf9Q4SuMCsIuKdlm8D1eA
oCaggsx4bWmkdZyLDHGefNp20ZRU8j+SzlYB4glqTS7O7RN7NhpkEXr0bi9no95M
7mtKv+AHR/WCCh2e+6xYY9hK48wuGl/GW4+tNq+xamV6zZ89PncvS72HDBr3lZFe
8+itM5H5jXSEntGuDnAe/GkO6aZKkBikfGBgXaV5y9JPPxI0E4vrtOZ36K5sMldT
ODEWmldutgYcaKdb+Oet/4vMVeWdsKvbbPluG+INh44yxhXlyM3AJE8DtC2zNAct
D/cOMwwZQgI0itBwHFRE7BFPCapu4+h9BeF7GxbUFu/mWslu3jGmUbZnA+S/IH8i
6u1E5lVauhYhVwZSabnXdcmwLJkpCrrV5sQxTHHMbxhDHuBj6RFhxJYrm3EEIo5M
wc0SkdSymxNSGFMy9TXH854aQz0T+v9176vy+gdTyvJRHbDBZTlkIkgx2KKLTgcm
o2/4QNYX1Rai6VLg9hGoo9eQME7vTGUU+NNB0Jk+LUaC+o7cmWDqTkDC5mRhvczD
homfq9k8ddJ7hyPBi2yH41fKGCRxSPLC+yz0ju+Ky08IeBi0t/gcjs+1ywVhL7O6
O5wHBaSpqPjpJ1PROmMdErEOKoh0eWenM94FfK6LUNU4VntkTVjo2etq4iRmKZ9p
DlBbhmfE9sMnf57qwrlKj7pZXBoL/0vEUaojed5waWy60srEylU5WCyNA9lsdCZm
AAqov713l7J0ym/PCBVRvTrHXZJQaZTaqHrROKxWvlaodCOQC2VXUuXaDkpGQuhv
lv/Dres8b2xqYsTZoA6sSRwGItx4kuif1TgxpbaX+0dtbMp3s1R+2e0DEbbky1Lg
`pragma protect end_protected
